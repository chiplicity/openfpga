magic
tech sky130A
magscale 1 2
timestamp 1605015152
<< locali >>
rect 35173 8959 35207 9129
<< viali >>
rect 5641 36329 5675 36363
rect 6837 36329 6871 36363
rect 5457 36193 5491 36227
rect 6653 36193 6687 36227
rect 22385 36193 22419 36227
rect 14197 35989 14231 36023
rect 21465 35989 21499 36023
rect 22569 35989 22603 36023
rect 4537 35785 4571 35819
rect 6285 35785 6319 35819
rect 7481 35785 7515 35819
rect 8125 35785 8159 35819
rect 11897 35785 11931 35819
rect 22477 35785 22511 35819
rect 24317 35785 24351 35819
rect 35633 35785 35667 35819
rect 5825 35717 5859 35751
rect 6653 35717 6687 35751
rect 14105 35717 14139 35751
rect 15301 35717 15335 35751
rect 23857 35717 23891 35751
rect 13645 35649 13679 35683
rect 14657 35649 14691 35683
rect 20913 35649 20947 35683
rect 21925 35649 21959 35683
rect 4353 35581 4387 35615
rect 5641 35581 5675 35615
rect 6837 35581 6871 35615
rect 7941 35581 7975 35615
rect 11253 35581 11287 35615
rect 13093 35581 13127 35615
rect 14013 35581 14047 35615
rect 14473 35581 14507 35615
rect 21741 35581 21775 35615
rect 23673 35581 23707 35615
rect 25697 35581 25731 35615
rect 35449 35581 35483 35615
rect 36001 35581 36035 35615
rect 8585 35513 8619 35547
rect 21833 35513 21867 35547
rect 25605 35513 25639 35547
rect 25942 35513 25976 35547
rect 4997 35445 5031 35479
rect 5549 35445 5583 35479
rect 7021 35445 7055 35479
rect 11437 35445 11471 35479
rect 14565 35445 14599 35479
rect 16773 35445 16807 35479
rect 21189 35445 21223 35479
rect 21373 35445 21407 35479
rect 27077 35445 27111 35479
rect 1593 35241 1627 35275
rect 10885 35241 10919 35275
rect 15761 35241 15795 35275
rect 35541 35241 35575 35275
rect 8125 35173 8159 35207
rect 13645 35173 13679 35207
rect 21189 35173 21223 35207
rect 1409 35105 1443 35139
rect 4997 35105 5031 35139
rect 6837 35105 6871 35139
rect 8309 35105 8343 35139
rect 11253 35105 11287 35139
rect 13553 35105 13587 35139
rect 15669 35105 15703 35139
rect 16865 35105 16899 35139
rect 21281 35105 21315 35139
rect 22385 35105 22419 35139
rect 22641 35105 22675 35139
rect 27712 35105 27746 35139
rect 35357 35105 35391 35139
rect 5089 35037 5123 35071
rect 5273 35037 5307 35071
rect 9689 35037 9723 35071
rect 11345 35037 11379 35071
rect 11529 35037 11563 35071
rect 12541 35037 12575 35071
rect 13093 35037 13127 35071
rect 13737 35037 13771 35071
rect 14933 35037 14967 35071
rect 15853 35037 15887 35071
rect 17969 35037 18003 35071
rect 27445 35037 27479 35071
rect 4353 34969 4387 35003
rect 7389 34969 7423 35003
rect 13185 34969 13219 35003
rect 4629 34901 4663 34935
rect 7021 34901 7055 34935
rect 8493 34901 8527 34935
rect 10149 34901 10183 34935
rect 12081 34901 12115 34935
rect 14657 34901 14691 34935
rect 15301 34901 15335 34935
rect 17049 34901 17083 34935
rect 18521 34901 18555 34935
rect 21465 34901 21499 34935
rect 21925 34901 21959 34935
rect 23765 34901 23799 34935
rect 24317 34901 24351 34935
rect 25789 34901 25823 34935
rect 26801 34901 26835 34935
rect 28825 34901 28859 34935
rect 1593 34697 1627 34731
rect 2053 34697 2087 34731
rect 3157 34697 3191 34731
rect 4261 34697 4295 34731
rect 5273 34697 5307 34731
rect 6653 34697 6687 34731
rect 8861 34697 8895 34731
rect 11713 34697 11747 34731
rect 14381 34697 14415 34731
rect 16957 34697 16991 34731
rect 17877 34697 17911 34731
rect 18061 34697 18095 34731
rect 20637 34697 20671 34731
rect 21005 34697 21039 34731
rect 22477 34697 22511 34731
rect 23029 34697 23063 34731
rect 25605 34697 25639 34731
rect 28089 34697 28123 34731
rect 35633 34697 35667 34731
rect 36737 34697 36771 34731
rect 2697 34629 2731 34663
rect 8217 34629 8251 34663
rect 17509 34629 17543 34663
rect 3801 34561 3835 34595
rect 4905 34561 4939 34595
rect 12449 34561 12483 34595
rect 18521 34561 18555 34595
rect 18613 34561 18647 34595
rect 24225 34561 24259 34595
rect 26709 34561 26743 34595
rect 1409 34493 1443 34527
rect 2513 34493 2547 34527
rect 4169 34493 4203 34527
rect 4721 34493 4755 34527
rect 6837 34493 6871 34527
rect 9229 34493 9263 34527
rect 9781 34493 9815 34527
rect 14749 34493 14783 34527
rect 14933 34493 14967 34527
rect 15200 34493 15234 34527
rect 18429 34493 18463 34527
rect 19993 34493 20027 34527
rect 21097 34493 21131 34527
rect 21353 34493 21387 34527
rect 26976 34493 27010 34527
rect 35265 34493 35299 34527
rect 35449 34493 35483 34527
rect 36553 34493 36587 34527
rect 37105 34493 37139 34527
rect 7082 34425 7116 34459
rect 9689 34425 9723 34459
rect 10026 34425 10060 34459
rect 12173 34425 12207 34459
rect 12716 34425 12750 34459
rect 24470 34425 24504 34459
rect 26617 34425 26651 34459
rect 4629 34357 4663 34391
rect 6285 34357 6319 34391
rect 11161 34357 11195 34391
rect 13829 34357 13863 34391
rect 16313 34357 16347 34391
rect 20177 34357 20211 34391
rect 24041 34357 24075 34391
rect 28641 34357 28675 34391
rect 36001 34357 36035 34391
rect 1593 34153 1627 34187
rect 4261 34153 4295 34187
rect 6653 34153 6687 34187
rect 7205 34153 7239 34187
rect 9137 34153 9171 34187
rect 11069 34153 11103 34187
rect 11621 34153 11655 34187
rect 13553 34153 13587 34187
rect 14105 34153 14139 34187
rect 16221 34153 16255 34187
rect 22293 34153 22327 34187
rect 22937 34153 22971 34187
rect 23857 34153 23891 34187
rect 27537 34153 27571 34187
rect 35633 34153 35667 34187
rect 4721 34085 4755 34119
rect 12418 34085 12452 34119
rect 17684 34085 17718 34119
rect 28172 34085 28206 34119
rect 4077 34017 4111 34051
rect 5540 34017 5574 34051
rect 8401 34017 8435 34051
rect 8493 34017 8527 34051
rect 9956 34017 9990 34051
rect 14841 34017 14875 34051
rect 16957 34017 16991 34051
rect 17325 34017 17359 34051
rect 17417 34017 17451 34051
rect 20913 34017 20947 34051
rect 21180 34017 21214 34051
rect 23765 34017 23799 34051
rect 25329 34017 25363 34051
rect 26525 34017 26559 34051
rect 27077 34017 27111 34051
rect 27905 34017 27939 34051
rect 35449 34017 35483 34051
rect 5273 33949 5307 33983
rect 8585 33949 8619 33983
rect 9689 33949 9723 33983
rect 12173 33949 12207 33983
rect 16313 33949 16347 33983
rect 16497 33949 16531 33983
rect 23949 33949 23983 33983
rect 25881 33949 25915 33983
rect 7573 33881 7607 33915
rect 15853 33881 15887 33915
rect 26709 33881 26743 33915
rect 5089 33813 5123 33847
rect 8033 33813 8067 33847
rect 9413 33813 9447 33847
rect 14473 33813 14507 33847
rect 14657 33813 14691 33847
rect 15485 33813 15519 33847
rect 18797 33813 18831 33847
rect 23397 33813 23431 33847
rect 24409 33813 24443 33847
rect 25513 33813 25547 33847
rect 29285 33813 29319 33847
rect 4077 33609 4111 33643
rect 5641 33609 5675 33643
rect 6193 33609 6227 33643
rect 6561 33609 6595 33643
rect 6837 33609 6871 33643
rect 8493 33609 8527 33643
rect 10149 33609 10183 33643
rect 10701 33609 10735 33643
rect 12173 33609 12207 33643
rect 14381 33609 14415 33643
rect 14933 33609 14967 33643
rect 15393 33609 15427 33643
rect 19441 33609 19475 33643
rect 22109 33609 22143 33643
rect 23121 33609 23155 33643
rect 23489 33609 23523 33643
rect 23673 33609 23707 33643
rect 25697 33609 25731 33643
rect 28549 33609 28583 33643
rect 35633 33609 35667 33643
rect 11069 33541 11103 33575
rect 11805 33541 11839 33575
rect 22661 33541 22695 33575
rect 24685 33541 24719 33575
rect 25881 33541 25915 33575
rect 3433 33473 3467 33507
rect 4261 33473 4295 33507
rect 7481 33473 7515 33507
rect 8769 33473 8803 33507
rect 11253 33473 11287 33507
rect 20269 33473 20303 33507
rect 20729 33473 20763 33507
rect 24133 33473 24167 33507
rect 24225 33473 24259 33507
rect 26341 33473 26375 33507
rect 26433 33473 26467 33507
rect 27997 33473 28031 33507
rect 7205 33405 7239 33439
rect 8677 33405 8711 33439
rect 9036 33405 9070 33439
rect 13001 33405 13035 33439
rect 13268 33405 13302 33439
rect 15485 33405 15519 33439
rect 15741 33405 15775 33439
rect 18061 33405 18095 33439
rect 18328 33405 18362 33439
rect 24041 33405 24075 33439
rect 26249 33405 26283 33439
rect 27353 33405 27387 33439
rect 27905 33405 27939 33439
rect 35449 33405 35483 33439
rect 3801 33337 3835 33371
rect 4528 33337 4562 33371
rect 7297 33337 7331 33371
rect 12909 33337 12943 33371
rect 20637 33337 20671 33371
rect 20974 33337 21008 33371
rect 26985 33337 27019 33371
rect 27813 33337 27847 33371
rect 8033 33269 8067 33303
rect 16865 33269 16899 33303
rect 17509 33269 17543 33303
rect 17785 33269 17819 33303
rect 25421 33269 25455 33303
rect 27445 33269 27479 33303
rect 28825 33269 28859 33303
rect 35357 33269 35391 33303
rect 36001 33269 36035 33303
rect 5457 33065 5491 33099
rect 6009 33065 6043 33099
rect 8677 33065 8711 33099
rect 9045 33065 9079 33099
rect 10149 33065 10183 33099
rect 11253 33065 11287 33099
rect 11621 33065 11655 33099
rect 13369 33065 13403 33099
rect 15117 33065 15151 33099
rect 17877 33065 17911 33099
rect 19349 33065 19383 33099
rect 20729 33065 20763 33099
rect 21189 33065 21223 33099
rect 21373 33065 21407 33099
rect 23305 33065 23339 33099
rect 23949 33065 23983 33099
rect 24317 33065 24351 33099
rect 25329 33065 25363 33099
rect 25881 33065 25915 33099
rect 26525 33065 26559 33099
rect 26893 33065 26927 33099
rect 27629 33065 27663 33099
rect 27997 33065 28031 33099
rect 4344 32997 4378 33031
rect 9413 32997 9447 33031
rect 10057 32997 10091 33031
rect 21741 32997 21775 33031
rect 22753 32997 22787 33031
rect 25237 32997 25271 33031
rect 26985 32997 27019 33031
rect 4077 32929 4111 32963
rect 6929 32929 6963 32963
rect 8125 32929 8159 32963
rect 13001 32929 13035 32963
rect 13829 32929 13863 32963
rect 15624 32929 15658 32963
rect 18225 32929 18259 32963
rect 21833 32929 21867 32963
rect 24685 32929 24719 32963
rect 28632 32929 28666 32963
rect 7021 32861 7055 32895
rect 7113 32861 7147 32895
rect 10241 32861 10275 32895
rect 11713 32861 11747 32895
rect 11897 32861 11931 32895
rect 13921 32861 13955 32895
rect 14013 32861 14047 32895
rect 15301 32861 15335 32895
rect 15764 32861 15798 32895
rect 16037 32861 16071 32895
rect 17969 32861 18003 32895
rect 21925 32861 21959 32895
rect 23397 32861 23431 32895
rect 23581 32861 23615 32895
rect 25421 32861 25455 32895
rect 27077 32861 27111 32895
rect 28365 32861 28399 32895
rect 3157 32725 3191 32759
rect 6561 32725 6595 32759
rect 7757 32725 7791 32759
rect 8309 32725 8343 32759
rect 9689 32725 9723 32759
rect 12817 32725 12851 32759
rect 13461 32725 13495 32759
rect 14473 32725 14507 32759
rect 17141 32725 17175 32759
rect 17509 32725 17543 32759
rect 22937 32725 22971 32759
rect 24869 32725 24903 32759
rect 26341 32725 26375 32759
rect 29745 32725 29779 32759
rect 4537 32521 4571 32555
rect 5089 32521 5123 32555
rect 5549 32521 5583 32555
rect 6653 32521 6687 32555
rect 9965 32521 9999 32555
rect 10241 32521 10275 32555
rect 11621 32521 11655 32555
rect 12081 32521 12115 32555
rect 13185 32521 13219 32555
rect 13553 32521 13587 32555
rect 17049 32521 17083 32555
rect 20177 32521 20211 32555
rect 23673 32521 23707 32555
rect 24961 32521 24995 32555
rect 26065 32521 26099 32555
rect 27077 32521 27111 32555
rect 28733 32521 28767 32555
rect 30665 32521 30699 32555
rect 5825 32453 5859 32487
rect 7113 32453 7147 32487
rect 9505 32453 9539 32487
rect 13829 32453 13863 32487
rect 16221 32453 16255 32487
rect 22385 32453 22419 32487
rect 22937 32453 22971 32487
rect 25237 32453 25271 32487
rect 27629 32453 27663 32487
rect 29101 32453 29135 32487
rect 3157 32385 3191 32419
rect 8309 32385 8343 32419
rect 8769 32385 8803 32419
rect 14844 32385 14878 32419
rect 16497 32385 16531 32419
rect 18061 32385 18095 32419
rect 21005 32385 21039 32419
rect 24317 32385 24351 32419
rect 26525 32385 26559 32419
rect 26617 32385 26651 32419
rect 27537 32385 27571 32419
rect 28089 32385 28123 32419
rect 28181 32385 28215 32419
rect 5641 32317 5675 32351
rect 6193 32317 6227 32351
rect 8125 32317 8159 32351
rect 9137 32317 9171 32351
rect 9321 32317 9355 32351
rect 10885 32317 10919 32351
rect 11345 32317 11379 32351
rect 14381 32317 14415 32351
rect 15117 32317 15151 32351
rect 17233 32317 17267 32351
rect 18328 32317 18362 32351
rect 20545 32317 20579 32351
rect 20913 32317 20947 32351
rect 21272 32317 21306 32351
rect 24041 32317 24075 32351
rect 25973 32317 26007 32351
rect 27997 32317 28031 32351
rect 29285 32317 29319 32351
rect 29541 32317 29575 32351
rect 3065 32249 3099 32283
rect 3402 32249 3436 32283
rect 8217 32249 8251 32283
rect 12817 32249 12851 32283
rect 17785 32249 17819 32283
rect 23489 32249 23523 32283
rect 24133 32249 24167 32283
rect 26433 32249 26467 32283
rect 2053 32181 2087 32215
rect 2421 32181 2455 32215
rect 7573 32181 7607 32215
rect 7757 32181 7791 32215
rect 10701 32181 10735 32215
rect 14289 32181 14323 32215
rect 14847 32181 14881 32215
rect 16957 32181 16991 32215
rect 19441 32181 19475 32215
rect 1961 31977 1995 32011
rect 3065 31977 3099 32011
rect 4445 31977 4479 32011
rect 5089 31977 5123 32011
rect 5825 31977 5859 32011
rect 6929 31977 6963 32011
rect 8033 31977 8067 32011
rect 8493 31977 8527 32011
rect 9045 31977 9079 32011
rect 9965 31977 9999 32011
rect 10793 31977 10827 32011
rect 14105 31977 14139 32011
rect 14657 31977 14691 32011
rect 15577 31977 15611 32011
rect 17509 31977 17543 32011
rect 17601 31977 17635 32011
rect 18613 31977 18647 32011
rect 19073 31977 19107 32011
rect 22385 31977 22419 32011
rect 23029 31977 23063 32011
rect 23673 31977 23707 32011
rect 24133 31977 24167 32011
rect 25053 31977 25087 32011
rect 26157 31977 26191 32011
rect 29561 31977 29595 32011
rect 35633 31977 35667 32011
rect 4537 31909 4571 31943
rect 17969 31909 18003 31943
rect 20729 31909 20763 31943
rect 23305 31909 23339 31943
rect 25145 31909 25179 31943
rect 26709 31909 26743 31943
rect 27721 31909 27755 31943
rect 2329 31841 2363 31875
rect 6193 31841 6227 31875
rect 7849 31841 7883 31875
rect 9229 31841 9263 31875
rect 16221 31841 16255 31875
rect 16497 31841 16531 31875
rect 17049 31841 17083 31875
rect 21272 31841 21306 31875
rect 23489 31841 23523 31875
rect 25697 31841 25731 31875
rect 26525 31841 26559 31875
rect 27169 31841 27203 31875
rect 28448 31841 28482 31875
rect 35449 31841 35483 31875
rect 2421 31773 2455 31807
rect 2605 31773 2639 31807
rect 4721 31773 4755 31807
rect 6285 31773 6319 31807
rect 6469 31773 6503 31807
rect 18061 31773 18095 31807
rect 18153 31773 18187 31807
rect 21005 31773 21039 31807
rect 24501 31773 24535 31807
rect 25237 31773 25271 31807
rect 26893 31773 26927 31807
rect 28181 31773 28215 31807
rect 1777 31637 1811 31671
rect 4077 31637 4111 31671
rect 5457 31637 5491 31671
rect 14933 31637 14967 31671
rect 15853 31637 15887 31671
rect 16037 31637 16071 31671
rect 24685 31637 24719 31671
rect 28089 31637 28123 31671
rect 30113 31637 30147 31671
rect 3617 31433 3651 31467
rect 4537 31433 4571 31467
rect 6561 31433 6595 31467
rect 7941 31433 7975 31467
rect 8677 31433 8711 31467
rect 13185 31433 13219 31467
rect 14289 31433 14323 31467
rect 17325 31433 17359 31467
rect 21189 31433 21223 31467
rect 23489 31433 23523 31467
rect 24225 31433 24259 31467
rect 26617 31433 26651 31467
rect 27077 31433 27111 31467
rect 27629 31433 27663 31467
rect 4261 31365 4295 31399
rect 17693 31365 17727 31399
rect 22201 31365 22235 31399
rect 5181 31297 5215 31331
rect 5273 31297 5307 31331
rect 9965 31297 9999 31331
rect 21833 31297 21867 31331
rect 22569 31297 22603 31331
rect 24593 31297 24627 31331
rect 28181 31297 28215 31331
rect 2237 31229 2271 31263
rect 5089 31229 5123 31263
rect 7757 31229 7791 31263
rect 8309 31229 8343 31263
rect 12449 31229 12483 31263
rect 13645 31229 13679 31263
rect 14841 31229 14875 31263
rect 15301 31229 15335 31263
rect 21557 31229 21591 31263
rect 24685 31229 24719 31263
rect 24952 31229 24986 31263
rect 2145 31161 2179 31195
rect 2504 31161 2538 31195
rect 9229 31161 9263 31195
rect 9781 31161 9815 31195
rect 12633 31161 12667 31195
rect 15209 31161 15243 31195
rect 15546 31161 15580 31195
rect 20361 31161 20395 31195
rect 20637 31161 20671 31195
rect 21097 31161 21131 31195
rect 21649 31161 21683 31195
rect 27997 31161 28031 31195
rect 1685 31093 1719 31127
rect 4721 31093 4755 31127
rect 5825 31093 5859 31127
rect 6285 31093 6319 31127
rect 9321 31093 9355 31127
rect 9689 31093 9723 31127
rect 10425 31093 10459 31127
rect 12265 31093 12299 31127
rect 12817 31093 12851 31127
rect 13829 31093 13863 31127
rect 16681 31093 16715 31127
rect 18245 31093 18279 31127
rect 26065 31093 26099 31127
rect 27537 31093 27571 31127
rect 28089 31093 28123 31127
rect 28733 31093 28767 31127
rect 29009 31093 29043 31127
rect 35449 31093 35483 31127
rect 2881 30889 2915 30923
rect 4353 30889 4387 30923
rect 5457 30889 5491 30923
rect 6193 30889 6227 30923
rect 9873 30889 9907 30923
rect 14749 30889 14783 30923
rect 15577 30889 15611 30923
rect 18981 30889 19015 30923
rect 22293 30889 22327 30923
rect 24133 30889 24167 30923
rect 25145 30889 25179 30923
rect 26709 30889 26743 30923
rect 28089 30889 28123 30923
rect 29745 30889 29779 30923
rect 35633 30889 35667 30923
rect 13461 30821 13495 30855
rect 21158 30821 21192 30855
rect 25697 30821 25731 30855
rect 27721 30821 27755 30855
rect 1768 30753 1802 30787
rect 4813 30753 4847 30787
rect 6009 30753 6043 30787
rect 8401 30753 8435 30787
rect 9413 30753 9447 30787
rect 10773 30753 10807 30787
rect 13369 30753 13403 30787
rect 15117 30753 15151 30787
rect 15945 30753 15979 30787
rect 17877 30753 17911 30787
rect 20269 30753 20303 30787
rect 20913 30753 20947 30787
rect 23581 30753 23615 30787
rect 24593 30753 24627 30787
rect 25053 30753 25087 30787
rect 26525 30753 26559 30787
rect 28632 30753 28666 30787
rect 35449 30753 35483 30787
rect 1501 30685 1535 30719
rect 4905 30685 4939 30719
rect 4997 30685 5031 30719
rect 8493 30685 8527 30719
rect 8677 30685 8711 30719
rect 10517 30685 10551 30719
rect 13553 30685 13587 30719
rect 16037 30685 16071 30719
rect 16129 30685 16163 30719
rect 17141 30685 17175 30719
rect 17464 30685 17498 30719
rect 17604 30685 17638 30719
rect 25329 30685 25363 30719
rect 28365 30685 28399 30719
rect 7941 30617 7975 30651
rect 4445 30549 4479 30583
rect 8033 30549 8067 30583
rect 11897 30549 11931 30583
rect 12541 30549 12575 30583
rect 12817 30549 12851 30583
rect 13001 30549 13035 30583
rect 17049 30549 17083 30583
rect 23765 30549 23799 30583
rect 24685 30549 24719 30583
rect 4629 30345 4663 30379
rect 6009 30345 6043 30379
rect 9965 30345 9999 30379
rect 14749 30345 14783 30379
rect 15209 30345 15243 30379
rect 21557 30345 21591 30379
rect 23489 30345 23523 30379
rect 24501 30345 24535 30379
rect 26617 30345 26651 30379
rect 28365 30345 28399 30379
rect 3801 30277 3835 30311
rect 7021 30277 7055 30311
rect 8125 30277 8159 30311
rect 24225 30277 24259 30311
rect 35633 30277 35667 30311
rect 5181 30209 5215 30243
rect 5641 30209 5675 30243
rect 8585 30209 8619 30243
rect 11897 30209 11931 30243
rect 13001 30209 13035 30243
rect 15780 30209 15814 30243
rect 16037 30209 16071 30243
rect 17785 30209 17819 30243
rect 18521 30209 18555 30243
rect 18705 30209 18739 30243
rect 20177 30209 20211 30243
rect 1409 30141 1443 30175
rect 6837 30141 6871 30175
rect 7389 30141 7423 30175
rect 11253 30141 11287 30175
rect 14197 30141 14231 30175
rect 15301 30141 15335 30175
rect 18429 30141 18463 30175
rect 19073 30141 19107 30175
rect 24685 30141 24719 30175
rect 24952 30141 24986 30175
rect 35449 30141 35483 30175
rect 36001 30141 36035 30175
rect 1676 30073 1710 30107
rect 4537 30073 4571 30107
rect 5089 30073 5123 30107
rect 8493 30073 8527 30107
rect 8852 30073 8886 30107
rect 10977 30073 11011 30107
rect 12909 30073 12943 30107
rect 13829 30073 13863 30107
rect 17509 30073 17543 30107
rect 20422 30073 20456 30107
rect 2789 30005 2823 30039
rect 3341 30005 3375 30039
rect 4169 30005 4203 30039
rect 4997 30005 5031 30039
rect 10609 30005 10643 30039
rect 11437 30005 11471 30039
rect 12265 30005 12299 30039
rect 12449 30005 12483 30039
rect 12817 30005 12851 30039
rect 13553 30005 13587 30039
rect 14381 30005 14415 30039
rect 15767 30005 15801 30039
rect 17141 30005 17175 30039
rect 18061 30005 18095 30039
rect 19993 30005 20027 30039
rect 26065 30005 26099 30039
rect 28733 30005 28767 30039
rect 35357 30005 35391 30039
rect 2789 29801 2823 29835
rect 4537 29801 4571 29835
rect 6101 29801 6135 29835
rect 7941 29801 7975 29835
rect 9045 29801 9079 29835
rect 11069 29801 11103 29835
rect 13553 29801 13587 29835
rect 14197 29801 14231 29835
rect 14749 29801 14783 29835
rect 15577 29801 15611 29835
rect 17969 29801 18003 29835
rect 18705 29801 18739 29835
rect 21097 29801 21131 29835
rect 23765 29801 23799 29835
rect 24225 29801 24259 29835
rect 24593 29801 24627 29835
rect 25789 29801 25823 29835
rect 35633 29801 35667 29835
rect 4988 29733 5022 29767
rect 8401 29733 8435 29767
rect 9956 29733 9990 29767
rect 17601 29733 17635 29767
rect 21465 29733 21499 29767
rect 32496 29733 32530 29767
rect 1676 29665 1710 29699
rect 3433 29665 3467 29699
rect 3893 29665 3927 29699
rect 4721 29665 4755 29699
rect 7573 29665 7607 29699
rect 9689 29665 9723 29699
rect 12429 29665 12463 29699
rect 15117 29665 15151 29699
rect 15936 29665 15970 29699
rect 19533 29665 19567 29699
rect 23581 29665 23615 29699
rect 25053 29665 25087 29699
rect 27721 29665 27755 29699
rect 35449 29665 35483 29699
rect 1409 29597 1443 29631
rect 8493 29597 8527 29631
rect 8677 29597 8711 29631
rect 12173 29597 12207 29631
rect 15669 29597 15703 29631
rect 18153 29597 18187 29631
rect 19625 29597 19659 29631
rect 19717 29597 19751 29631
rect 25145 29597 25179 29631
rect 25329 29597 25363 29631
rect 26525 29597 26559 29631
rect 31309 29597 31343 29631
rect 32229 29597 32263 29631
rect 7205 29461 7239 29495
rect 8033 29461 8067 29495
rect 17049 29461 17083 29495
rect 19165 29461 19199 29495
rect 20177 29461 20211 29495
rect 24685 29461 24719 29495
rect 27537 29461 27571 29495
rect 33609 29461 33643 29495
rect 34897 29461 34931 29495
rect 1685 29257 1719 29291
rect 2053 29257 2087 29291
rect 3341 29257 3375 29291
rect 5641 29257 5675 29291
rect 6193 29257 6227 29291
rect 7113 29257 7147 29291
rect 7481 29257 7515 29291
rect 9321 29257 9355 29291
rect 9965 29257 9999 29291
rect 10425 29257 10459 29291
rect 12265 29257 12299 29291
rect 14841 29257 14875 29291
rect 15485 29257 15519 29291
rect 19257 29257 19291 29291
rect 21005 29257 21039 29291
rect 23489 29257 23523 29291
rect 27997 29257 28031 29291
rect 11529 29189 11563 29223
rect 12633 29189 12667 29223
rect 15945 29189 15979 29223
rect 17049 29189 17083 29223
rect 18889 29189 18923 29223
rect 32689 29189 32723 29223
rect 33241 29189 33275 29223
rect 2421 29121 2455 29155
rect 2789 29121 2823 29155
rect 7849 29121 7883 29155
rect 10977 29121 11011 29155
rect 13093 29121 13127 29155
rect 16405 29121 16439 29155
rect 16497 29121 16531 29155
rect 24777 29121 24811 29155
rect 31309 29121 31343 29155
rect 3157 29053 3191 29087
rect 3709 29053 3743 29087
rect 4261 29053 4295 29087
rect 7941 29053 7975 29087
rect 8208 29053 8242 29087
rect 13461 29053 13495 29087
rect 13717 29053 13751 29087
rect 17417 29053 17451 29087
rect 19625 29053 19659 29087
rect 23949 29053 23983 29087
rect 25053 29053 25087 29087
rect 27537 29053 27571 29087
rect 34897 29053 34931 29087
rect 4169 28985 4203 29019
rect 4506 28985 4540 29019
rect 10241 28985 10275 29019
rect 10885 28985 10919 29019
rect 15761 28985 15795 29019
rect 16313 28985 16347 29019
rect 18521 28985 18555 29019
rect 19892 28985 19926 29019
rect 25320 28985 25354 29019
rect 31217 28985 31251 29019
rect 31576 28985 31610 29019
rect 34621 28985 34655 29019
rect 35142 28985 35176 29019
rect 10793 28917 10827 28951
rect 24133 28917 24167 28951
rect 26433 28917 26467 28951
rect 30573 28917 30607 28951
rect 33701 28917 33735 28951
rect 34345 28917 34379 28951
rect 36277 28917 36311 28951
rect 1961 28713 1995 28747
rect 2421 28713 2455 28747
rect 5457 28713 5491 28747
rect 8493 28713 8527 28747
rect 9873 28713 9907 28747
rect 10517 28713 10551 28747
rect 10885 28713 10919 28747
rect 11069 28713 11103 28747
rect 12817 28713 12851 28747
rect 13553 28713 13587 28747
rect 13921 28713 13955 28747
rect 14381 28713 14415 28747
rect 15393 28713 15427 28747
rect 15853 28713 15887 28747
rect 16405 28713 16439 28747
rect 18245 28713 18279 28747
rect 18981 28713 19015 28747
rect 19257 28713 19291 28747
rect 20269 28713 20303 28747
rect 20637 28713 20671 28747
rect 24041 28713 24075 28747
rect 24409 28713 24443 28747
rect 24869 28713 24903 28747
rect 25237 28713 25271 28747
rect 30389 28713 30423 28747
rect 30849 28713 30883 28747
rect 33517 28713 33551 28747
rect 7380 28645 7414 28679
rect 15761 28645 15795 28679
rect 19625 28645 19659 28679
rect 24685 28645 24719 28679
rect 26770 28645 26804 28679
rect 34888 28645 34922 28679
rect 2789 28577 2823 28611
rect 3893 28577 3927 28611
rect 4077 28577 4111 28611
rect 4344 28577 4378 28611
rect 7113 28577 7147 28611
rect 9689 28577 9723 28611
rect 11437 28577 11471 28611
rect 12633 28577 12667 28611
rect 13737 28577 13771 28611
rect 20913 28577 20947 28611
rect 21180 28577 21214 28611
rect 32393 28577 32427 28611
rect 2881 28509 2915 28543
rect 2973 28509 3007 28543
rect 11529 28509 11563 28543
rect 11621 28509 11655 28543
rect 16037 28509 16071 28543
rect 19717 28509 19751 28543
rect 19901 28509 19935 28543
rect 25329 28509 25363 28543
rect 25513 28509 25547 28543
rect 26525 28509 26559 28543
rect 30941 28509 30975 28543
rect 31033 28509 31067 28543
rect 32137 28509 32171 28543
rect 34621 28509 34655 28543
rect 2329 28441 2363 28475
rect 22293 28441 22327 28475
rect 25973 28373 26007 28407
rect 26249 28373 26283 28407
rect 27905 28373 27939 28407
rect 30021 28373 30055 28407
rect 30481 28373 30515 28407
rect 31953 28373 31987 28407
rect 34437 28373 34471 28407
rect 36001 28373 36035 28407
rect 1869 28169 1903 28203
rect 4813 28169 4847 28203
rect 6653 28169 6687 28203
rect 9229 28169 9263 28203
rect 9965 28169 9999 28203
rect 11161 28169 11195 28203
rect 11805 28169 11839 28203
rect 13369 28169 13403 28203
rect 13737 28169 13771 28203
rect 15485 28169 15519 28203
rect 15853 28169 15887 28203
rect 21649 28169 21683 28203
rect 23489 28169 23523 28203
rect 24593 28169 24627 28203
rect 25697 28169 25731 28203
rect 28089 28169 28123 28203
rect 29745 28169 29779 28203
rect 31585 28169 31619 28203
rect 32229 28169 32263 28203
rect 34713 28169 34747 28203
rect 12633 28101 12667 28135
rect 24133 28101 24167 28135
rect 33241 28101 33275 28135
rect 2329 28033 2363 28067
rect 5365 28033 5399 28067
rect 6193 28033 6227 28067
rect 8125 28033 8159 28067
rect 14381 28033 14415 28067
rect 16129 28033 16163 28067
rect 18521 28033 18555 28067
rect 19444 28033 19478 28067
rect 19717 28033 19751 28067
rect 21189 28033 21223 28067
rect 22293 28033 22327 28067
rect 22661 28033 22695 28067
rect 25145 28033 25179 28067
rect 26065 28033 26099 28067
rect 30205 28033 30239 28067
rect 33793 28033 33827 28067
rect 5181 27965 5215 27999
rect 5825 27965 5859 27999
rect 9045 27965 9079 27999
rect 9597 27965 9631 27999
rect 12449 27965 12483 27999
rect 13001 27965 13035 27999
rect 18981 27965 19015 27999
rect 26157 27965 26191 27999
rect 26424 27965 26458 27999
rect 33149 27965 33183 27999
rect 33701 27965 33735 27999
rect 34989 27965 35023 27999
rect 35256 27965 35290 27999
rect 2237 27897 2271 27931
rect 2574 27897 2608 27931
rect 4353 27897 4387 27931
rect 4721 27897 4755 27931
rect 7941 27897 7975 27931
rect 22017 27897 22051 27931
rect 22109 27897 22143 27931
rect 23029 27897 23063 27931
rect 24501 27897 24535 27931
rect 25053 27897 25087 27931
rect 30113 27897 30147 27931
rect 30472 27897 30506 27931
rect 33609 27897 33643 27931
rect 3709 27829 3743 27863
rect 5273 27829 5307 27863
rect 7297 27829 7331 27863
rect 7481 27829 7515 27863
rect 7849 27829 7883 27863
rect 11437 27829 11471 27863
rect 18889 27829 18923 27863
rect 19447 27829 19481 27863
rect 20821 27829 20855 27863
rect 21465 27829 21499 27863
rect 24961 27829 24995 27863
rect 27537 27829 27571 27863
rect 32781 27829 32815 27863
rect 34345 27829 34379 27863
rect 36369 27829 36403 27863
rect 2145 27625 2179 27659
rect 3157 27625 3191 27659
rect 5457 27625 5491 27659
rect 11161 27625 11195 27659
rect 19349 27625 19383 27659
rect 22477 27625 22511 27659
rect 29469 27625 29503 27659
rect 33333 27625 33367 27659
rect 35081 27625 35115 27659
rect 3893 27557 3927 27591
rect 4322 27557 4356 27591
rect 7941 27557 7975 27591
rect 8401 27557 8435 27591
rect 13553 27557 13587 27591
rect 15844 27557 15878 27591
rect 18981 27557 19015 27591
rect 19809 27557 19843 27591
rect 20729 27557 20763 27591
rect 24317 27557 24351 27591
rect 32597 27557 32631 27591
rect 1961 27489 1995 27523
rect 2513 27489 2547 27523
rect 8493 27489 8527 27523
rect 10977 27489 11011 27523
rect 21097 27489 21131 27523
rect 21364 27489 21398 27523
rect 25237 27489 25271 27523
rect 25329 27489 25363 27523
rect 26792 27489 26826 27523
rect 29817 27489 29851 27523
rect 32505 27489 32539 27523
rect 34069 27489 34103 27523
rect 35440 27489 35474 27523
rect 2605 27421 2639 27455
rect 2697 27421 2731 27455
rect 4077 27421 4111 27455
rect 8677 27421 8711 27455
rect 15577 27421 15611 27455
rect 25513 27421 25547 27455
rect 26341 27421 26375 27455
rect 26525 27421 26559 27455
rect 29561 27421 29595 27455
rect 32689 27421 32723 27455
rect 34713 27421 34747 27455
rect 35173 27421 35207 27455
rect 8033 27353 8067 27387
rect 18613 27353 18647 27387
rect 24869 27353 24903 27387
rect 27905 27353 27939 27387
rect 7205 27285 7239 27319
rect 7573 27285 7607 27319
rect 16957 27285 16991 27319
rect 19717 27285 19751 27319
rect 24593 27285 24627 27319
rect 25881 27285 25915 27319
rect 30941 27285 30975 27319
rect 31861 27285 31895 27319
rect 32137 27285 32171 27319
rect 34253 27285 34287 27319
rect 36553 27285 36587 27319
rect 1777 27081 1811 27115
rect 3249 27081 3283 27115
rect 4169 27081 4203 27115
rect 5365 27081 5399 27115
rect 5733 27081 5767 27115
rect 6193 27081 6227 27115
rect 8309 27081 8343 27115
rect 9229 27081 9263 27115
rect 10241 27081 10275 27115
rect 15669 27081 15703 27115
rect 18705 27081 18739 27115
rect 21189 27081 21223 27115
rect 24225 27081 24259 27115
rect 29101 27081 29135 27115
rect 33333 27081 33367 27115
rect 34161 27081 34195 27115
rect 34621 27081 34655 27115
rect 36001 27081 36035 27115
rect 36369 27081 36403 27115
rect 4353 27013 4387 27047
rect 9597 27013 9631 27047
rect 27629 27013 27663 27047
rect 32321 27013 32355 27047
rect 33701 27013 33735 27047
rect 4813 26945 4847 26979
rect 4997 26945 5031 26979
rect 6929 26945 6963 26979
rect 13369 26945 13403 26979
rect 16037 26945 16071 26979
rect 21741 26945 21775 26979
rect 24961 26945 24995 26979
rect 29837 26945 29871 26979
rect 32229 26945 32263 26979
rect 32781 26945 32815 26979
rect 32965 26945 32999 26979
rect 35449 26945 35483 26979
rect 37013 26945 37047 26979
rect 1869 26877 1903 26911
rect 2136 26877 2170 26911
rect 3801 26877 3835 26911
rect 4721 26877 4755 26911
rect 10057 26877 10091 26911
rect 10609 26877 10643 26911
rect 13461 26877 13495 26911
rect 13728 26877 13762 26911
rect 18061 26877 18095 26911
rect 25237 26877 25271 26911
rect 27721 26877 27755 26911
rect 35357 26877 35391 26911
rect 36921 26877 36955 26911
rect 6653 26809 6687 26843
rect 7196 26809 7230 26843
rect 21097 26809 21131 26843
rect 21649 26809 21683 26843
rect 24593 26809 24627 26843
rect 25504 26809 25538 26843
rect 29745 26809 29779 26843
rect 30082 26809 30116 26843
rect 31861 26809 31895 26843
rect 32689 26809 32723 26843
rect 35265 26809 35299 26843
rect 8861 26741 8895 26775
rect 11069 26741 11103 26775
rect 14841 26741 14875 26775
rect 18245 26741 18279 26775
rect 19349 26741 19383 26775
rect 20177 26741 20211 26775
rect 20729 26741 20763 26775
rect 21557 26741 21591 26775
rect 22293 26741 22327 26775
rect 22569 26741 22603 26775
rect 26617 26741 26651 26775
rect 27261 26741 27295 26775
rect 31217 26741 31251 26775
rect 34897 26741 34931 26775
rect 36461 26741 36495 26775
rect 36829 26741 36863 26775
rect 37473 26741 37507 26775
rect 37841 26741 37875 26775
rect 2881 26537 2915 26571
rect 4353 26537 4387 26571
rect 4629 26537 4663 26571
rect 6469 26537 6503 26571
rect 7481 26537 7515 26571
rect 11253 26537 11287 26571
rect 11713 26537 11747 26571
rect 12817 26537 12851 26571
rect 13277 26537 13311 26571
rect 19257 26537 19291 26571
rect 19717 26537 19751 26571
rect 22293 26537 22327 26571
rect 25697 26537 25731 26571
rect 29377 26537 29411 26571
rect 29745 26537 29779 26571
rect 30757 26537 30791 26571
rect 33241 26537 33275 26571
rect 34989 26537 35023 26571
rect 37105 26537 37139 26571
rect 1768 26469 1802 26503
rect 15844 26469 15878 26503
rect 19625 26469 19659 26503
rect 24133 26469 24167 26503
rect 31953 26469 31987 26503
rect 32597 26469 32631 26503
rect 1501 26401 1535 26435
rect 6837 26401 6871 26435
rect 8401 26401 8435 26435
rect 11621 26401 11655 26435
rect 13185 26401 13219 26435
rect 15577 26401 15611 26435
rect 18061 26401 18095 26435
rect 20729 26401 20763 26435
rect 21180 26401 21214 26435
rect 25053 26401 25087 26435
rect 27261 26401 27295 26435
rect 29193 26401 29227 26435
rect 30665 26401 30699 26435
rect 32505 26401 32539 26435
rect 34069 26401 34103 26435
rect 35173 26401 35207 26435
rect 35429 26401 35463 26435
rect 6929 26333 6963 26367
rect 7113 26333 7147 26367
rect 8493 26333 8527 26367
rect 8585 26333 8619 26367
rect 11805 26333 11839 26367
rect 13369 26333 13403 26367
rect 19901 26333 19935 26367
rect 20913 26333 20947 26367
rect 25145 26333 25179 26367
rect 25329 26333 25363 26367
rect 26525 26333 26559 26367
rect 26848 26333 26882 26367
rect 26988 26333 27022 26367
rect 30205 26333 30239 26367
rect 30849 26333 30883 26367
rect 32689 26333 32723 26367
rect 33517 26333 33551 26367
rect 8033 26265 8067 26299
rect 9321 26265 9355 26299
rect 12725 26265 12759 26299
rect 16957 26265 16991 26299
rect 19165 26265 19199 26299
rect 20361 26265 20395 26299
rect 24685 26265 24719 26299
rect 26249 26265 26283 26299
rect 28365 26265 28399 26299
rect 32137 26265 32171 26299
rect 36553 26265 36587 26299
rect 12357 26197 12391 26231
rect 18245 26197 18279 26231
rect 24501 26197 24535 26231
rect 30297 26197 30331 26231
rect 31585 26197 31619 26231
rect 34253 26197 34287 26231
rect 2237 25993 2271 26027
rect 5825 25993 5859 26027
rect 8217 25993 8251 26027
rect 8769 25993 8803 26027
rect 9321 25993 9355 26027
rect 11345 25993 11379 26027
rect 16773 25993 16807 26027
rect 18337 25993 18371 26027
rect 19257 25993 19291 26027
rect 22661 25993 22695 26027
rect 22937 25993 22971 26027
rect 27077 25993 27111 26027
rect 28825 25993 28859 26027
rect 31769 25993 31803 26027
rect 32229 25993 32263 26027
rect 34069 25993 34103 26027
rect 34621 25993 34655 26027
rect 36093 25993 36127 26027
rect 17141 25925 17175 25959
rect 23857 25925 23891 25959
rect 26249 25925 26283 25959
rect 28089 25925 28123 25959
rect 33057 25925 33091 25959
rect 6837 25857 6871 25891
rect 9873 25857 9907 25891
rect 10333 25857 10367 25891
rect 10885 25857 10919 25891
rect 15209 25857 15243 25891
rect 15577 25857 15611 25891
rect 16129 25857 16163 25891
rect 16313 25857 16347 25891
rect 19165 25857 19199 25891
rect 19809 25857 19843 25891
rect 20821 25857 20855 25891
rect 21284 25857 21318 25891
rect 24872 25857 24906 25891
rect 27721 25857 27755 25891
rect 32045 25857 32079 25891
rect 33701 25857 33735 25891
rect 9689 25789 9723 25823
rect 12449 25789 12483 25823
rect 12716 25789 12750 25823
rect 14841 25789 14875 25823
rect 16037 25789 16071 25823
rect 18797 25789 18831 25823
rect 19625 25789 19659 25823
rect 21557 25789 21591 25823
rect 23489 25789 23523 25823
rect 24409 25789 24443 25823
rect 25145 25789 25179 25823
rect 27445 25789 27479 25823
rect 29101 25789 29135 25823
rect 29745 25789 29779 25823
rect 32413 25789 32447 25823
rect 35357 25789 35391 25823
rect 35633 25789 35667 25823
rect 35817 25789 35851 25823
rect 36645 25789 36679 25823
rect 37197 25789 37231 25823
rect 1685 25721 1719 25755
rect 6193 25721 6227 25755
rect 7104 25721 7138 25755
rect 12265 25721 12299 25755
rect 19717 25721 19751 25755
rect 26985 25721 27019 25755
rect 27537 25721 27571 25755
rect 29653 25721 29687 25755
rect 30012 25721 30046 25755
rect 33517 25721 33551 25755
rect 35449 25721 35483 25755
rect 2513 25653 2547 25687
rect 6561 25653 6595 25687
rect 9137 25653 9171 25687
rect 9781 25653 9815 25687
rect 11621 25653 11655 25687
rect 13829 25653 13863 25687
rect 14381 25653 14415 25687
rect 15669 25653 15703 25687
rect 20269 25653 20303 25687
rect 20729 25653 20763 25687
rect 21287 25653 21321 25687
rect 24317 25653 24351 25687
rect 24875 25653 24909 25687
rect 26617 25653 26651 25687
rect 28917 25653 28951 25687
rect 31125 25653 31159 25687
rect 32873 25653 32907 25687
rect 33425 25653 33459 25687
rect 36829 25653 36863 25687
rect 6561 25449 6595 25483
rect 8125 25449 8159 25483
rect 8677 25449 8711 25483
rect 10057 25449 10091 25483
rect 13553 25449 13587 25483
rect 14565 25449 14599 25483
rect 18429 25449 18463 25483
rect 19349 25449 19383 25483
rect 20085 25449 20119 25483
rect 20729 25449 20763 25483
rect 22293 25449 22327 25483
rect 24133 25449 24167 25483
rect 24409 25449 24443 25483
rect 24593 25449 24627 25483
rect 26157 25449 26191 25483
rect 26801 25449 26835 25483
rect 27077 25449 27111 25483
rect 27261 25449 27295 25483
rect 27721 25449 27755 25483
rect 29745 25449 29779 25483
rect 30205 25449 30239 25483
rect 31677 25449 31711 25483
rect 31769 25449 31803 25483
rect 33793 25449 33827 25483
rect 34253 25449 34287 25483
rect 34805 25449 34839 25483
rect 35265 25449 35299 25483
rect 15752 25381 15786 25415
rect 21158 25381 21192 25415
rect 30573 25381 30607 25415
rect 31309 25381 31343 25415
rect 6745 25313 6779 25347
rect 7001 25313 7035 25347
rect 10425 25313 10459 25347
rect 11621 25313 11655 25347
rect 11888 25313 11922 25347
rect 14749 25313 14783 25347
rect 18337 25313 18371 25347
rect 24961 25313 24995 25347
rect 26341 25313 26375 25347
rect 27445 25313 27479 25347
rect 29377 25313 29411 25347
rect 30113 25313 30147 25347
rect 30665 25313 30699 25347
rect 31945 25313 31979 25347
rect 32505 25313 32539 25347
rect 34161 25313 34195 25347
rect 35725 25313 35759 25347
rect 10517 25245 10551 25279
rect 10609 25245 10643 25279
rect 15485 25245 15519 25279
rect 18521 25245 18555 25279
rect 19625 25245 19659 25279
rect 20913 25245 20947 25279
rect 25053 25245 25087 25279
rect 25237 25245 25271 25279
rect 30849 25245 30883 25279
rect 32597 25245 32631 25279
rect 32689 25245 32723 25279
rect 34345 25245 34379 25279
rect 35817 25245 35851 25279
rect 36001 25245 36035 25279
rect 33609 25177 33643 25211
rect 35357 25177 35391 25211
rect 1685 25109 1719 25143
rect 9413 25109 9447 25143
rect 9965 25109 9999 25143
rect 13001 25109 13035 25143
rect 16865 25109 16899 25143
rect 17969 25109 18003 25143
rect 29009 25109 29043 25143
rect 32137 25109 32171 25143
rect 33149 25109 33183 25143
rect 5917 24905 5951 24939
rect 6193 24905 6227 24939
rect 8309 24905 8343 24939
rect 8953 24905 8987 24939
rect 9781 24905 9815 24939
rect 11897 24905 11931 24939
rect 15117 24905 15151 24939
rect 18337 24905 18371 24939
rect 19165 24905 19199 24939
rect 21465 24905 21499 24939
rect 22017 24905 22051 24939
rect 27353 24905 27387 24939
rect 31033 24905 31067 24939
rect 32137 24905 32171 24939
rect 33609 24905 33643 24939
rect 33885 24905 33919 24939
rect 34253 24905 34287 24939
rect 37013 24905 37047 24939
rect 6653 24769 6687 24803
rect 9413 24769 9447 24803
rect 23949 24769 23983 24803
rect 24685 24769 24719 24803
rect 32689 24769 32723 24803
rect 35081 24769 35115 24803
rect 6929 24701 6963 24735
rect 7196 24701 7230 24735
rect 9873 24701 9907 24735
rect 10140 24701 10174 24735
rect 12173 24701 12207 24735
rect 12449 24701 12483 24735
rect 12716 24701 12750 24735
rect 15301 24701 15335 24735
rect 18981 24701 19015 24735
rect 19533 24701 19567 24735
rect 20085 24701 20119 24735
rect 24317 24701 24351 24735
rect 25053 24701 25087 24735
rect 25320 24701 25354 24735
rect 29653 24701 29687 24735
rect 32505 24701 32539 24735
rect 33701 24701 33735 24735
rect 14841 24633 14875 24667
rect 15568 24633 15602 24667
rect 17325 24633 17359 24667
rect 19993 24633 20027 24667
rect 20330 24633 20364 24667
rect 29561 24633 29595 24667
rect 29898 24633 29932 24667
rect 31585 24633 31619 24667
rect 32045 24633 32079 24667
rect 32597 24633 32631 24667
rect 34713 24633 34747 24667
rect 35348 24633 35382 24667
rect 11253 24565 11287 24599
rect 13829 24565 13863 24599
rect 14473 24565 14507 24599
rect 16681 24565 16715 24599
rect 17785 24565 17819 24599
rect 18613 24565 18647 24599
rect 22385 24565 22419 24599
rect 26433 24565 26467 24599
rect 29101 24565 29135 24599
rect 33149 24565 33183 24599
rect 36461 24565 36495 24599
rect 6837 24361 6871 24395
rect 8493 24361 8527 24395
rect 11805 24361 11839 24395
rect 15485 24361 15519 24395
rect 15945 24361 15979 24395
rect 20913 24361 20947 24395
rect 24685 24361 24719 24395
rect 25513 24361 25547 24395
rect 26249 24361 26283 24395
rect 30941 24361 30975 24395
rect 31953 24361 31987 24395
rect 32137 24361 32171 24395
rect 33793 24361 33827 24395
rect 34161 24361 34195 24395
rect 36277 24361 36311 24395
rect 10048 24293 10082 24327
rect 14657 24293 14691 24327
rect 15117 24293 15151 24327
rect 21281 24293 21315 24327
rect 25237 24293 25271 24327
rect 33149 24293 33183 24327
rect 35909 24293 35943 24327
rect 7113 24225 7147 24259
rect 7369 24225 7403 24259
rect 9505 24225 9539 24259
rect 9781 24225 9815 24259
rect 15853 24225 15887 24259
rect 17049 24225 17083 24259
rect 18981 24225 19015 24259
rect 22017 24225 22051 24259
rect 29828 24225 29862 24259
rect 32505 24225 32539 24259
rect 34897 24225 34931 24259
rect 36093 24225 36127 24259
rect 16129 24157 16163 24191
rect 19073 24157 19107 24191
rect 19165 24157 19199 24191
rect 21373 24157 21407 24191
rect 21465 24157 21499 24191
rect 29561 24157 29595 24191
rect 32597 24157 32631 24191
rect 32689 24157 32723 24191
rect 34989 24157 35023 24191
rect 35173 24157 35207 24191
rect 12541 24089 12575 24123
rect 18061 24089 18095 24123
rect 19993 24089 20027 24123
rect 31585 24089 31619 24123
rect 35541 24089 35575 24123
rect 11161 24021 11195 24055
rect 17233 24021 17267 24055
rect 18429 24021 18463 24055
rect 18613 24021 18647 24055
rect 19625 24021 19659 24055
rect 20361 24021 20395 24055
rect 29469 24021 29503 24055
rect 34529 24021 34563 24055
rect 7205 23817 7239 23851
rect 9045 23817 9079 23851
rect 10149 23817 10183 23851
rect 14473 23817 14507 23851
rect 16589 23817 16623 23851
rect 17141 23817 17175 23851
rect 19073 23817 19107 23851
rect 20269 23817 20303 23851
rect 20729 23817 20763 23851
rect 22109 23817 22143 23851
rect 29101 23817 29135 23851
rect 31125 23817 31159 23851
rect 32137 23817 32171 23851
rect 32413 23817 32447 23851
rect 34621 23817 34655 23851
rect 36921 23817 36955 23851
rect 33149 23749 33183 23783
rect 33609 23749 33643 23783
rect 7573 23681 7607 23715
rect 9873 23681 9907 23715
rect 10609 23681 10643 23715
rect 10701 23681 10735 23715
rect 19809 23681 19843 23715
rect 7665 23613 7699 23647
rect 7932 23613 7966 23647
rect 10517 23613 10551 23647
rect 11161 23613 11195 23647
rect 14565 23613 14599 23647
rect 14821 23613 14855 23647
rect 18337 23613 18371 23647
rect 18521 23613 18555 23647
rect 19533 23613 19567 23647
rect 29745 23613 29779 23647
rect 31769 23613 31803 23647
rect 32229 23613 32263 23647
rect 33701 23613 33735 23647
rect 34897 23613 34931 23647
rect 20821 23545 20855 23579
rect 29653 23545 29687 23579
rect 30012 23545 30046 23579
rect 32781 23545 32815 23579
rect 35164 23545 35198 23579
rect 11621 23477 11655 23511
rect 15945 23477 15979 23511
rect 17785 23477 17819 23511
rect 18705 23477 18739 23511
rect 19165 23477 19199 23511
rect 19625 23477 19659 23511
rect 28733 23477 28767 23511
rect 33885 23477 33919 23511
rect 36277 23477 36311 23511
rect 7205 23273 7239 23307
rect 7757 23273 7791 23307
rect 10241 23273 10275 23307
rect 10425 23273 10459 23307
rect 10885 23273 10919 23307
rect 14105 23273 14139 23307
rect 15485 23273 15519 23307
rect 16773 23273 16807 23307
rect 16865 23273 16899 23307
rect 18245 23273 18279 23307
rect 18705 23273 18739 23307
rect 20453 23273 20487 23307
rect 21097 23273 21131 23307
rect 25145 23273 25179 23307
rect 30941 23273 30975 23307
rect 32321 23273 32355 23307
rect 33609 23273 33643 23307
rect 34437 23273 34471 23307
rect 34989 23273 35023 23307
rect 35909 23273 35943 23307
rect 15945 23205 15979 23239
rect 16313 23205 16347 23239
rect 19340 23205 19374 23239
rect 26525 23205 26559 23239
rect 34069 23205 34103 23239
rect 10609 23137 10643 23171
rect 14013 23137 14047 23171
rect 15301 23137 15335 23171
rect 18061 23137 18095 23171
rect 19073 23137 19107 23171
rect 26709 23137 26743 23171
rect 29469 23137 29503 23171
rect 29561 23137 29595 23171
rect 29828 23137 29862 23171
rect 32137 23137 32171 23171
rect 33425 23137 33459 23171
rect 34897 23137 34931 23171
rect 36093 23137 36127 23171
rect 13553 23069 13587 23103
rect 14289 23069 14323 23103
rect 17049 23069 17083 23103
rect 35173 23069 35207 23103
rect 16405 23001 16439 23035
rect 13645 22933 13679 22967
rect 21557 22933 21591 22967
rect 26893 22933 26927 22967
rect 34529 22933 34563 22967
rect 35541 22933 35575 22967
rect 36553 22933 36587 22967
rect 7573 22729 7607 22763
rect 8125 22729 8159 22763
rect 10517 22729 10551 22763
rect 13001 22729 13035 22763
rect 15209 22729 15243 22763
rect 16313 22729 16347 22763
rect 18245 22729 18279 22763
rect 20545 22729 20579 22763
rect 27169 22729 27203 22763
rect 31033 22729 31067 22763
rect 32597 22729 32631 22763
rect 32965 22729 32999 22763
rect 33425 22729 33459 22763
rect 34621 22729 34655 22763
rect 35081 22729 35115 22763
rect 36185 22729 36219 22763
rect 16405 22661 16439 22695
rect 18981 22661 19015 22695
rect 26525 22661 26559 22695
rect 27445 22661 27479 22695
rect 17049 22593 17083 22627
rect 17785 22593 17819 22627
rect 18705 22593 18739 22627
rect 25145 22593 25179 22627
rect 35725 22593 35759 22627
rect 36461 22593 36495 22627
rect 7757 22525 7791 22559
rect 13829 22525 13863 22559
rect 18086 22525 18120 22559
rect 19165 22525 19199 22559
rect 19421 22525 19455 22559
rect 28733 22525 28767 22559
rect 29101 22525 29135 22559
rect 29653 22525 29687 22559
rect 32321 22525 32355 22559
rect 33701 22525 33735 22559
rect 35449 22525 35483 22559
rect 13369 22457 13403 22491
rect 13737 22457 13771 22491
rect 14096 22457 14130 22491
rect 15945 22457 15979 22491
rect 16773 22457 16807 22491
rect 17417 22457 17451 22491
rect 25053 22457 25087 22491
rect 25390 22457 25424 22491
rect 29561 22457 29595 22491
rect 29898 22457 29932 22491
rect 16865 22389 16899 22423
rect 22385 22389 22419 22423
rect 32137 22389 32171 22423
rect 33885 22389 33919 22423
rect 35541 22389 35575 22423
rect 36829 22389 36863 22423
rect 13553 22185 13587 22219
rect 14013 22185 14047 22219
rect 14657 22185 14691 22219
rect 15117 22185 15151 22219
rect 15301 22185 15335 22219
rect 16405 22185 16439 22219
rect 17049 22185 17083 22219
rect 17417 22185 17451 22219
rect 18153 22185 18187 22219
rect 29653 22185 29687 22219
rect 33793 22185 33827 22219
rect 34529 22185 34563 22219
rect 26792 22117 26826 22151
rect 34888 22117 34922 22151
rect 13185 22049 13219 22083
rect 14105 22049 14139 22083
rect 15669 22049 15703 22083
rect 16865 22049 16899 22083
rect 18613 22049 18647 22083
rect 19165 22049 19199 22083
rect 22753 22049 22787 22083
rect 22845 22049 22879 22083
rect 24205 22049 24239 22083
rect 12817 21981 12851 22015
rect 14197 21981 14231 22015
rect 15761 21981 15795 22015
rect 15945 21981 15979 22015
rect 23029 21981 23063 22015
rect 23949 21981 23983 22015
rect 26525 21981 26559 22015
rect 34161 21981 34195 22015
rect 34621 21981 34655 22015
rect 13001 21913 13035 21947
rect 13645 21913 13679 21947
rect 18797 21913 18831 21947
rect 19625 21845 19659 21879
rect 19993 21845 20027 21879
rect 22293 21845 22327 21879
rect 22385 21845 22419 21879
rect 23765 21845 23799 21879
rect 25329 21845 25363 21879
rect 27905 21845 27939 21879
rect 30021 21845 30055 21879
rect 36001 21845 36035 21879
rect 8585 21641 8619 21675
rect 13185 21641 13219 21675
rect 14657 21641 14691 21675
rect 15669 21641 15703 21675
rect 15945 21641 15979 21675
rect 16405 21641 16439 21675
rect 17417 21641 17451 21675
rect 19993 21641 20027 21675
rect 22477 21641 22511 21675
rect 23397 21641 23431 21675
rect 26065 21641 26099 21675
rect 26801 21641 26835 21675
rect 27905 21641 27939 21675
rect 31125 21641 31159 21675
rect 34713 21641 34747 21675
rect 36277 21641 36311 21675
rect 27445 21573 27479 21607
rect 17049 21505 17083 21539
rect 8769 21437 8803 21471
rect 13277 21437 13311 21471
rect 13533 21437 13567 21471
rect 17877 21437 17911 21471
rect 18613 21437 18647 21471
rect 21097 21437 21131 21471
rect 23673 21437 23707 21471
rect 23929 21437 23963 21471
rect 26157 21437 26191 21471
rect 27261 21437 27295 21471
rect 29745 21437 29779 21471
rect 33977 21437 34011 21471
rect 34897 21437 34931 21471
rect 35164 21437 35198 21471
rect 12817 21369 12851 21403
rect 18858 21369 18892 21403
rect 21005 21369 21039 21403
rect 21342 21369 21376 21403
rect 25697 21369 25731 21403
rect 27169 21369 27203 21403
rect 29653 21369 29687 21403
rect 29990 21369 30024 21403
rect 34345 21369 34379 21403
rect 9137 21301 9171 21335
rect 12265 21301 12299 21335
rect 15209 21301 15243 21335
rect 16773 21301 16807 21335
rect 16865 21301 16899 21335
rect 18429 21301 18463 21335
rect 23121 21301 23155 21335
rect 25053 21301 25087 21335
rect 26341 21301 26375 21335
rect 14105 21097 14139 21131
rect 15301 21097 15335 21131
rect 16773 21097 16807 21131
rect 17693 21097 17727 21131
rect 18705 21097 18739 21131
rect 19441 21097 19475 21131
rect 21097 21097 21131 21131
rect 23121 21097 23155 21131
rect 24041 21097 24075 21131
rect 25513 21097 25547 21131
rect 26893 21097 26927 21131
rect 28273 21097 28307 21131
rect 30665 21097 30699 21131
rect 33333 21097 33367 21131
rect 36645 21097 36679 21131
rect 12992 21029 13026 21063
rect 17141 21029 17175 21063
rect 12725 20961 12759 20995
rect 15669 20961 15703 20995
rect 18061 20961 18095 20995
rect 18153 20961 18187 20995
rect 19257 20961 19291 20995
rect 21741 20961 21775 20995
rect 22008 20961 22042 20995
rect 24225 20961 24259 20995
rect 28089 20961 28123 20995
rect 29837 20961 29871 20995
rect 29929 20961 29963 20995
rect 15761 20893 15795 20927
rect 15945 20893 15979 20927
rect 18245 20893 18279 20927
rect 26985 20893 27019 20927
rect 27169 20893 27203 20927
rect 29377 20893 29411 20927
rect 30021 20893 30055 20927
rect 33885 20893 33919 20927
rect 33977 20893 34011 20927
rect 34300 20893 34334 20927
rect 34440 20893 34474 20927
rect 34713 20893 34747 20927
rect 14749 20825 14783 20859
rect 15117 20825 15151 20859
rect 16497 20825 16531 20859
rect 26341 20825 26375 20859
rect 17509 20757 17543 20791
rect 21649 20757 21683 20791
rect 26525 20757 26559 20791
rect 27629 20757 27663 20791
rect 29469 20757 29503 20791
rect 35817 20757 35851 20791
rect 36093 20757 36127 20791
rect 10057 20553 10091 20587
rect 12817 20553 12851 20587
rect 15209 20553 15243 20587
rect 15669 20553 15703 20587
rect 16681 20553 16715 20587
rect 17141 20553 17175 20587
rect 19441 20553 19475 20587
rect 19993 20553 20027 20587
rect 26617 20553 26651 20587
rect 28641 20553 28675 20587
rect 29101 20553 29135 20587
rect 30021 20553 30055 20587
rect 33241 20553 33275 20587
rect 34621 20553 34655 20587
rect 9505 20485 9539 20519
rect 25697 20485 25731 20519
rect 34253 20485 34287 20519
rect 16221 20417 16255 20451
rect 22385 20417 22419 20451
rect 24133 20417 24167 20451
rect 24317 20417 24351 20451
rect 24961 20417 24995 20451
rect 25145 20417 25179 20451
rect 26157 20417 26191 20451
rect 29561 20417 29595 20451
rect 30573 20417 30607 20451
rect 33793 20417 33827 20451
rect 9689 20349 9723 20383
rect 11621 20349 11655 20383
rect 11897 20349 11931 20383
rect 13185 20349 13219 20383
rect 13452 20349 13486 20383
rect 18061 20349 18095 20383
rect 20913 20349 20947 20383
rect 21281 20349 21315 20383
rect 23397 20349 23431 20383
rect 24869 20349 24903 20383
rect 25513 20349 25547 20383
rect 26709 20349 26743 20383
rect 33609 20349 33643 20383
rect 34989 20349 35023 20383
rect 35256 20349 35290 20383
rect 15577 20281 15611 20315
rect 16129 20281 16163 20315
rect 17509 20281 17543 20315
rect 17877 20281 17911 20315
rect 18328 20281 18362 20315
rect 22201 20281 22235 20315
rect 23121 20281 23155 20315
rect 24041 20281 24075 20315
rect 26976 20281 27010 20315
rect 30481 20281 30515 20315
rect 30818 20281 30852 20315
rect 33149 20281 33183 20315
rect 33701 20281 33735 20315
rect 11437 20213 11471 20247
rect 14565 20213 14599 20247
rect 16037 20213 16071 20247
rect 21557 20213 21591 20247
rect 21741 20213 21775 20247
rect 22109 20213 22143 20247
rect 23673 20213 23707 20247
rect 24501 20213 24535 20247
rect 28089 20213 28123 20247
rect 31953 20213 31987 20247
rect 36369 20213 36403 20247
rect 2789 20009 2823 20043
rect 12725 20009 12759 20043
rect 13277 20009 13311 20043
rect 13553 20009 13587 20043
rect 14013 20009 14047 20043
rect 15025 20009 15059 20043
rect 15761 20009 15795 20043
rect 18429 20009 18463 20043
rect 21281 20009 21315 20043
rect 22753 20009 22787 20043
rect 23397 20009 23431 20043
rect 23673 20009 23707 20043
rect 24777 20009 24811 20043
rect 25329 20009 25363 20043
rect 26341 20009 26375 20043
rect 27445 20009 27479 20043
rect 29837 20009 29871 20043
rect 30389 20009 30423 20043
rect 33333 20009 33367 20043
rect 33609 20009 33643 20043
rect 35633 20009 35667 20043
rect 36185 20009 36219 20043
rect 1654 19941 1688 19975
rect 27169 19941 27203 19975
rect 28150 19941 28184 19975
rect 31401 19941 31435 19975
rect 33977 19941 34011 19975
rect 35081 19941 35115 19975
rect 1409 19873 1443 19907
rect 13737 19873 13771 19907
rect 15945 19873 15979 19907
rect 16212 19873 16246 19907
rect 18797 19873 18831 19907
rect 21373 19873 21407 19907
rect 21629 19873 21663 19907
rect 25237 19873 25271 19907
rect 26525 19873 26559 19907
rect 27905 19873 27939 19907
rect 30757 19873 30791 19907
rect 35541 19873 35575 19907
rect 18889 19805 18923 19839
rect 18981 19805 19015 19839
rect 23857 19805 23891 19839
rect 25513 19805 25547 19839
rect 30297 19805 30331 19839
rect 30849 19805 30883 19839
rect 31033 19805 31067 19839
rect 34069 19805 34103 19839
rect 34253 19805 34287 19839
rect 35725 19805 35759 19839
rect 17325 19737 17359 19771
rect 34713 19737 34747 19771
rect 17969 19669 18003 19703
rect 18245 19669 18279 19703
rect 24317 19669 24351 19703
rect 24869 19669 24903 19703
rect 25881 19669 25915 19703
rect 26709 19669 26743 19703
rect 29285 19669 29319 19703
rect 32413 19669 32447 19703
rect 35173 19669 35207 19703
rect 1593 19465 1627 19499
rect 1961 19465 1995 19499
rect 14841 19465 14875 19499
rect 17877 19465 17911 19499
rect 19441 19465 19475 19499
rect 25605 19465 25639 19499
rect 26065 19465 26099 19499
rect 26617 19465 26651 19499
rect 28089 19465 28123 19499
rect 34069 19465 34103 19499
rect 13001 19329 13035 19363
rect 13461 19329 13495 19363
rect 16497 19329 16531 19363
rect 25237 19329 25271 19363
rect 27721 19329 27755 19363
rect 30116 19329 30150 19363
rect 32873 19329 32907 19363
rect 35081 19329 35115 19363
rect 13728 19261 13762 19295
rect 15485 19261 15519 19295
rect 16313 19261 16347 19295
rect 16957 19261 16991 19295
rect 17325 19261 17359 19295
rect 18061 19261 18095 19295
rect 20545 19261 20579 19295
rect 21005 19261 21039 19295
rect 22937 19261 22971 19295
rect 23489 19261 23523 19295
rect 27537 19261 27571 19295
rect 29653 19261 29687 19295
rect 30389 19261 30423 19295
rect 31769 19261 31803 19295
rect 35348 19261 35382 19295
rect 13369 19193 13403 19227
rect 15853 19193 15887 19227
rect 16405 19193 16439 19227
rect 18328 19193 18362 19227
rect 20821 19193 20855 19227
rect 21250 19193 21284 19227
rect 25053 19193 25087 19227
rect 26893 19193 26927 19227
rect 27445 19193 27479 19227
rect 29101 19193 29135 19227
rect 32229 19193 32263 19227
rect 32689 19193 32723 19227
rect 37013 19193 37047 19227
rect 15945 19125 15979 19159
rect 19993 19125 20027 19159
rect 22385 19125 22419 19159
rect 24133 19125 24167 19159
rect 24409 19125 24443 19159
rect 24593 19125 24627 19159
rect 24961 19125 24995 19159
rect 27077 19125 27111 19159
rect 28641 19125 28675 19159
rect 29469 19125 29503 19159
rect 30119 19125 30153 19159
rect 31493 19125 31527 19159
rect 32321 19125 32355 19159
rect 32781 19125 32815 19159
rect 33701 19125 33735 19159
rect 34713 19125 34747 19159
rect 36461 19125 36495 19159
rect 13553 18921 13587 18955
rect 16681 18921 16715 18955
rect 18153 18921 18187 18955
rect 20545 18921 20579 18955
rect 21465 18921 21499 18955
rect 23949 18921 23983 18955
rect 24685 18921 24719 18955
rect 24869 18921 24903 18955
rect 25329 18921 25363 18955
rect 27077 18921 27111 18955
rect 27813 18921 27847 18955
rect 28365 18921 28399 18955
rect 30941 18921 30975 18955
rect 32137 18921 32171 18955
rect 33517 18921 33551 18955
rect 35449 18921 35483 18955
rect 36277 18921 36311 18955
rect 15568 18853 15602 18887
rect 25973 18853 26007 18887
rect 29009 18853 29043 18887
rect 29469 18853 29503 18887
rect 29806 18853 29840 18887
rect 36185 18853 36219 18887
rect 18429 18785 18463 18819
rect 21833 18785 21867 18819
rect 22293 18785 22327 18819
rect 23765 18785 23799 18819
rect 25237 18785 25271 18819
rect 26525 18785 26559 18819
rect 26893 18785 26927 18819
rect 27445 18785 27479 18819
rect 33609 18785 33643 18819
rect 33932 18785 33966 18819
rect 15301 18717 15335 18751
rect 20177 18717 20211 18751
rect 22385 18717 22419 18751
rect 22569 18717 22603 18751
rect 25421 18717 25455 18751
rect 28457 18717 28491 18751
rect 28641 18717 28675 18751
rect 29561 18717 29595 18751
rect 34072 18717 34106 18751
rect 34345 18717 34379 18751
rect 26709 18649 26743 18683
rect 31493 18649 31527 18683
rect 17693 18581 17727 18615
rect 21925 18581 21959 18615
rect 27997 18581 28031 18615
rect 32597 18581 32631 18615
rect 35725 18581 35759 18615
rect 15393 18377 15427 18411
rect 15945 18377 15979 18411
rect 17877 18377 17911 18411
rect 19809 18377 19843 18411
rect 22569 18377 22603 18411
rect 22937 18377 22971 18411
rect 23489 18377 23523 18411
rect 24409 18377 24443 18411
rect 25513 18377 25547 18411
rect 25789 18377 25823 18411
rect 28457 18377 28491 18411
rect 28733 18377 28767 18411
rect 30389 18377 30423 18411
rect 36461 18377 36495 18411
rect 19441 18309 19475 18343
rect 24317 18309 24351 18343
rect 27997 18309 28031 18343
rect 30021 18309 30055 18343
rect 34253 18309 34287 18343
rect 13921 18241 13955 18275
rect 20453 18241 20487 18275
rect 20637 18241 20671 18275
rect 24961 18241 24995 18275
rect 27721 18241 27755 18275
rect 31036 18241 31070 18275
rect 32781 18241 32815 18275
rect 33793 18241 33827 18275
rect 14013 18173 14047 18207
rect 14280 18173 14314 18207
rect 18061 18173 18095 18207
rect 18317 18173 18351 18207
rect 25973 18173 26007 18207
rect 27813 18173 27847 18207
rect 30573 18173 30607 18207
rect 30896 18173 30930 18207
rect 31309 18173 31343 18207
rect 33149 18173 33183 18207
rect 33609 18173 33643 18207
rect 35081 18173 35115 18207
rect 20269 18105 20303 18139
rect 20882 18105 20916 18139
rect 23949 18105 23983 18139
rect 24869 18105 24903 18139
rect 33701 18105 33735 18139
rect 34713 18105 34747 18139
rect 35326 18105 35360 18139
rect 16313 18037 16347 18071
rect 20177 18037 20211 18071
rect 22017 18037 22051 18071
rect 24777 18037 24811 18071
rect 29561 18037 29595 18071
rect 32413 18037 32447 18071
rect 33241 18037 33275 18071
rect 14013 17833 14047 17867
rect 15485 17833 15519 17867
rect 18061 17833 18095 17867
rect 20177 17833 20211 17867
rect 21097 17833 21131 17867
rect 23581 17833 23615 17867
rect 24869 17833 24903 17867
rect 25881 17833 25915 17867
rect 26525 17833 26559 17867
rect 27813 17833 27847 17867
rect 31309 17833 31343 17867
rect 32505 17833 32539 17867
rect 32597 17833 32631 17867
rect 33609 17833 33643 17867
rect 34069 17833 34103 17867
rect 34437 17833 34471 17867
rect 35909 17833 35943 17867
rect 19073 17765 19107 17799
rect 24409 17765 24443 17799
rect 28273 17765 28307 17799
rect 29530 17765 29564 17799
rect 33333 17765 33367 17799
rect 22201 17697 22235 17731
rect 22293 17697 22327 17731
rect 23397 17697 23431 17731
rect 24041 17697 24075 17731
rect 25237 17697 25271 17731
rect 26893 17697 26927 17731
rect 34805 17697 34839 17731
rect 36001 17697 36035 17731
rect 21741 17629 21775 17663
rect 22385 17629 22419 17663
rect 25329 17629 25363 17663
rect 25421 17629 25455 17663
rect 26985 17629 27019 17663
rect 27077 17629 27111 17663
rect 29285 17629 29319 17663
rect 32781 17629 32815 17663
rect 34897 17629 34931 17663
rect 35081 17629 35115 17663
rect 19901 17561 19935 17595
rect 32137 17561 32171 17595
rect 18429 17493 18463 17527
rect 20729 17493 20763 17527
rect 21833 17493 21867 17527
rect 24777 17493 24811 17527
rect 29101 17493 29135 17527
rect 30665 17493 30699 17527
rect 35541 17493 35575 17527
rect 18981 17289 19015 17323
rect 21925 17289 21959 17323
rect 22845 17289 22879 17323
rect 23397 17289 23431 17323
rect 23857 17289 23891 17323
rect 27445 17289 27479 17323
rect 27905 17289 27939 17323
rect 29101 17289 29135 17323
rect 29469 17289 29503 17323
rect 31585 17289 31619 17323
rect 32873 17289 32907 17323
rect 34069 17289 34103 17323
rect 35173 17289 35207 17323
rect 32505 17221 32539 17255
rect 33701 17221 33735 17255
rect 19625 17153 19659 17187
rect 32229 17153 32263 17187
rect 35449 17153 35483 17187
rect 20545 17085 20579 17119
rect 22477 17085 22511 17119
rect 23673 17085 23707 17119
rect 24869 17085 24903 17119
rect 25125 17085 25159 17119
rect 26801 17085 26835 17119
rect 27629 17085 27663 17119
rect 28273 17085 28307 17119
rect 30205 17085 30239 17119
rect 30472 17085 30506 17119
rect 19349 17017 19383 17051
rect 20453 17017 20487 17051
rect 20812 17017 20846 17051
rect 24685 17017 24719 17051
rect 30113 17017 30147 17051
rect 35716 17017 35750 17051
rect 18889 16949 18923 16983
rect 19441 16949 19475 16983
rect 24409 16949 24443 16983
rect 26249 16949 26283 16983
rect 27169 16949 27203 16983
rect 34529 16949 34563 16983
rect 36829 16949 36863 16983
rect 19073 16745 19107 16779
rect 19257 16745 19291 16779
rect 22293 16745 22327 16779
rect 23673 16745 23707 16779
rect 25329 16745 25363 16779
rect 27905 16745 27939 16779
rect 29929 16745 29963 16779
rect 30941 16745 30975 16779
rect 35541 16745 35575 16779
rect 21158 16677 21192 16711
rect 24194 16677 24228 16711
rect 30297 16677 30331 16711
rect 19625 16609 19659 16643
rect 20637 16609 20671 16643
rect 20913 16609 20947 16643
rect 23949 16609 23983 16643
rect 26792 16609 26826 16643
rect 19717 16541 19751 16575
rect 19901 16541 19935 16575
rect 25973 16541 26007 16575
rect 26525 16541 26559 16575
rect 30389 16541 30423 16575
rect 30481 16541 30515 16575
rect 18981 16201 19015 16235
rect 20177 16201 20211 16235
rect 22109 16201 22143 16235
rect 24041 16201 24075 16235
rect 26893 16201 26927 16235
rect 27445 16201 27479 16235
rect 29929 16201 29963 16235
rect 30205 16201 30239 16235
rect 30573 16201 30607 16235
rect 24961 16133 24995 16167
rect 19349 16065 19383 16099
rect 28641 16065 28675 16099
rect 20729 15997 20763 16031
rect 22753 15997 22787 16031
rect 24409 15997 24443 16031
rect 25513 15997 25547 16031
rect 27997 15997 28031 16031
rect 29285 15997 29319 16031
rect 19717 15929 19751 15963
rect 20637 15929 20671 15963
rect 20996 15929 21030 15963
rect 25421 15929 25455 15963
rect 25780 15929 25814 15963
rect 28181 15861 28215 15895
rect 29469 15861 29503 15895
rect 32505 15861 32539 15895
rect 35449 15861 35483 15895
rect 22293 15657 22327 15691
rect 30389 15657 30423 15691
rect 36001 15657 36035 15691
rect 21180 15521 21214 15555
rect 27721 15521 27755 15555
rect 29745 15521 29779 15555
rect 32781 15521 32815 15555
rect 32873 15521 32907 15555
rect 35449 15521 35483 15555
rect 20729 15453 20763 15487
rect 20913 15453 20947 15487
rect 27813 15453 27847 15487
rect 27905 15453 27939 15487
rect 32965 15453 32999 15487
rect 26801 15385 26835 15419
rect 25605 15317 25639 15351
rect 27077 15317 27111 15351
rect 27353 15317 27387 15351
rect 29929 15317 29963 15351
rect 32413 15317 32447 15351
rect 35633 15317 35667 15351
rect 20637 15113 20671 15147
rect 22477 15113 22511 15147
rect 27721 15113 27755 15147
rect 27997 15113 28031 15147
rect 29101 15113 29135 15147
rect 30205 15113 30239 15147
rect 31769 15113 31803 15147
rect 32229 15113 32263 15147
rect 33701 15113 33735 15147
rect 35357 15113 35391 15147
rect 21005 14977 21039 15011
rect 27169 14977 27203 15011
rect 30573 14977 30607 15011
rect 20269 14909 20303 14943
rect 21097 14909 21131 14943
rect 21364 14909 21398 14943
rect 26157 14909 26191 14943
rect 26985 14909 27019 14943
rect 29745 14909 29779 14943
rect 30021 14909 30055 14943
rect 30941 14909 30975 14943
rect 31033 14909 31067 14943
rect 32321 14909 32355 14943
rect 35449 14909 35483 14943
rect 26525 14841 26559 14875
rect 27077 14841 27111 14875
rect 29837 14841 29871 14875
rect 32588 14841 32622 14875
rect 34713 14841 34747 14875
rect 35694 14841 35728 14875
rect 26617 14773 26651 14807
rect 31217 14773 31251 14807
rect 36829 14773 36863 14807
rect 24593 14569 24627 14603
rect 26525 14569 26559 14603
rect 27629 14569 27663 14603
rect 30113 14569 30147 14603
rect 32229 14569 32263 14603
rect 33707 14569 33741 14603
rect 35081 14569 35115 14603
rect 35541 14569 35575 14603
rect 36277 14569 36311 14603
rect 26893 14501 26927 14535
rect 28978 14501 29012 14535
rect 36369 14501 36403 14535
rect 23857 14433 23891 14467
rect 33977 14433 34011 14467
rect 23949 14365 23983 14399
rect 24133 14365 24167 14399
rect 26985 14365 27019 14399
rect 27169 14365 27203 14399
rect 28733 14365 28767 14399
rect 33241 14365 33275 14399
rect 33747 14365 33781 14399
rect 36461 14365 36495 14399
rect 21189 14229 21223 14263
rect 23489 14229 23523 14263
rect 31953 14229 31987 14263
rect 32781 14229 32815 14263
rect 33149 14229 33183 14263
rect 35909 14229 35943 14263
rect 22753 14025 22787 14059
rect 25053 14025 25087 14059
rect 26617 14025 26651 14059
rect 28089 14025 28123 14059
rect 28733 14025 28767 14059
rect 29653 14025 29687 14059
rect 31861 14025 31895 14059
rect 34253 14025 34287 14059
rect 35357 14025 35391 14059
rect 37381 14025 37415 14059
rect 36829 13957 36863 13991
rect 34621 13889 34655 13923
rect 23673 13821 23707 13855
rect 23929 13821 23963 13855
rect 25881 13821 25915 13855
rect 26709 13821 26743 13855
rect 29745 13821 29779 13855
rect 30012 13821 30046 13855
rect 32321 13821 32355 13855
rect 35449 13821 35483 13855
rect 35705 13821 35739 13855
rect 26249 13753 26283 13787
rect 26976 13753 27010 13787
rect 32566 13753 32600 13787
rect 23029 13685 23063 13719
rect 23397 13685 23431 13719
rect 31125 13685 31159 13719
rect 32137 13685 32171 13719
rect 33701 13685 33735 13719
rect 23581 13481 23615 13515
rect 25329 13481 25363 13515
rect 27169 13481 27203 13515
rect 29009 13481 29043 13515
rect 29653 13481 29687 13515
rect 30021 13481 30055 13515
rect 30481 13481 30515 13515
rect 31217 13481 31251 13515
rect 31953 13481 31987 13515
rect 32505 13481 32539 13515
rect 33155 13481 33189 13515
rect 34529 13481 34563 13515
rect 34897 13481 34931 13515
rect 35817 13481 35851 13515
rect 36461 13481 36495 13515
rect 24194 13413 24228 13447
rect 27874 13413 27908 13447
rect 36829 13413 36863 13447
rect 22753 13345 22787 13379
rect 23949 13345 23983 13379
rect 26525 13345 26559 13379
rect 27537 13345 27571 13379
rect 27629 13345 27663 13379
rect 22845 13277 22879 13311
rect 23029 13277 23063 13311
rect 30573 13277 30607 13311
rect 30665 13277 30699 13311
rect 32689 13277 32723 13311
rect 33152 13277 33186 13311
rect 33425 13277 33459 13311
rect 35909 13277 35943 13311
rect 36001 13277 36035 13311
rect 22293 13209 22327 13243
rect 22385 13141 22419 13175
rect 26709 13141 26743 13175
rect 30113 13141 30147 13175
rect 35265 13141 35299 13175
rect 35449 13141 35483 13175
rect 22477 12937 22511 12971
rect 24685 12937 24719 12971
rect 25605 12937 25639 12971
rect 27077 12937 27111 12971
rect 27721 12937 27755 12971
rect 28089 12937 28123 12971
rect 30205 12937 30239 12971
rect 32781 12937 32815 12971
rect 33149 12937 33183 12971
rect 34713 12937 34747 12971
rect 37105 12937 37139 12971
rect 23673 12869 23707 12903
rect 29745 12869 29779 12903
rect 30481 12869 30515 12903
rect 36553 12869 36587 12903
rect 24133 12801 24167 12835
rect 24317 12801 24351 12835
rect 30665 12801 30699 12835
rect 33793 12801 33827 12835
rect 35173 12801 35207 12835
rect 21097 12733 21131 12767
rect 24041 12733 24075 12767
rect 25053 12733 25087 12767
rect 25697 12733 25731 12767
rect 25953 12733 25987 12767
rect 29561 12733 29595 12767
rect 30932 12733 30966 12767
rect 35429 12733 35463 12767
rect 21005 12665 21039 12699
rect 21342 12665 21376 12699
rect 23029 12665 23063 12699
rect 33517 12665 33551 12699
rect 23489 12597 23523 12631
rect 32045 12597 32079 12631
rect 33609 12597 33643 12631
rect 34253 12597 34287 12631
rect 23673 12393 23707 12427
rect 24225 12393 24259 12427
rect 26709 12393 26743 12427
rect 27445 12393 27479 12427
rect 29653 12393 29687 12427
rect 30021 12393 30055 12427
rect 30573 12393 30607 12427
rect 32689 12393 32723 12427
rect 34253 12393 34287 12427
rect 36277 12393 36311 12427
rect 22538 12325 22572 12359
rect 33793 12325 33827 12359
rect 25145 12257 25179 12291
rect 27813 12257 27847 12291
rect 29009 12257 29043 12291
rect 30481 12257 30515 12291
rect 33149 12257 33183 12291
rect 34345 12257 34379 12291
rect 34612 12257 34646 12291
rect 21189 12189 21223 12223
rect 22293 12189 22327 12223
rect 27905 12189 27939 12223
rect 28089 12189 28123 12223
rect 30665 12189 30699 12223
rect 31125 12189 31159 12223
rect 33241 12189 33275 12223
rect 33425 12189 33459 12223
rect 25329 12121 25363 12155
rect 27353 12121 27387 12155
rect 30113 12121 30147 12155
rect 31493 12121 31527 12155
rect 24593 12053 24627 12087
rect 25053 12053 25087 12087
rect 25697 12053 25731 12087
rect 29193 12053 29227 12087
rect 31953 12053 31987 12087
rect 32781 12053 32815 12087
rect 35725 12053 35759 12087
rect 25145 11849 25179 11883
rect 26709 11849 26743 11883
rect 28549 11849 28583 11883
rect 29009 11849 29043 11883
rect 30113 11849 30147 11883
rect 30481 11849 30515 11883
rect 31309 11849 31343 11883
rect 32873 11849 32907 11883
rect 33609 11849 33643 11883
rect 33885 11849 33919 11883
rect 34345 11849 34379 11883
rect 22753 11781 22787 11815
rect 26617 11781 26651 11815
rect 27537 11781 27571 11815
rect 29837 11781 29871 11815
rect 34897 11781 34931 11815
rect 23489 11713 23523 11747
rect 24225 11713 24259 11747
rect 24409 11713 24443 11747
rect 24869 11713 24903 11747
rect 28089 11713 28123 11747
rect 31769 11713 31803 11747
rect 31861 11713 31895 11747
rect 33149 11713 33183 11747
rect 35449 11713 35483 11747
rect 26893 11645 26927 11679
rect 35357 11645 35391 11679
rect 35909 11645 35943 11679
rect 23121 11577 23155 11611
rect 24133 11577 24167 11611
rect 27445 11577 27479 11611
rect 27997 11577 28031 11611
rect 31217 11577 31251 11611
rect 31677 11577 31711 11611
rect 34713 11577 34747 11611
rect 35265 11577 35299 11611
rect 22385 11509 22419 11543
rect 23765 11509 23799 11543
rect 26249 11509 26283 11543
rect 27905 11509 27939 11543
rect 23765 11305 23799 11339
rect 26801 11305 26835 11339
rect 28365 11305 28399 11339
rect 28733 11305 28767 11339
rect 31401 11305 31435 11339
rect 32137 11305 32171 11339
rect 35081 11305 35115 11339
rect 27445 11237 27479 11271
rect 34989 11237 35023 11271
rect 22385 11169 22419 11203
rect 22652 11169 22686 11203
rect 25329 11169 25363 11203
rect 27353 11169 27387 11203
rect 28549 11169 28583 11203
rect 35541 11169 35575 11203
rect 27537 11101 27571 11135
rect 25513 11033 25547 11067
rect 27997 11033 28031 11067
rect 29193 11033 29227 11067
rect 22109 10965 22143 10999
rect 24317 10965 24351 10999
rect 26985 10965 27019 10999
rect 29929 10965 29963 10999
rect 23489 10761 23523 10795
rect 28089 10761 28123 10795
rect 29653 10761 29687 10795
rect 23949 10693 23983 10727
rect 25329 10693 25363 10727
rect 26525 10693 26559 10727
rect 28549 10693 28583 10727
rect 22569 10625 22603 10659
rect 24409 10625 24443 10659
rect 24593 10625 24627 10659
rect 26065 10625 26099 10659
rect 26985 10625 27019 10659
rect 27169 10625 27203 10659
rect 29101 10625 29135 10659
rect 30389 10625 30423 10659
rect 35449 10625 35483 10659
rect 21925 10557 21959 10591
rect 22385 10557 22419 10591
rect 25053 10557 25087 10591
rect 28273 10557 28307 10591
rect 24317 10489 24351 10523
rect 27905 10489 27939 10523
rect 30205 10489 30239 10523
rect 35357 10489 35391 10523
rect 35694 10489 35728 10523
rect 22017 10421 22051 10455
rect 22477 10421 22511 10455
rect 23121 10421 23155 10455
rect 26433 10421 26467 10455
rect 26893 10421 26927 10455
rect 27629 10421 27663 10455
rect 29837 10421 29871 10455
rect 30297 10421 30331 10455
rect 33793 10421 33827 10455
rect 36829 10421 36863 10455
rect 22109 10217 22143 10251
rect 24133 10217 24167 10251
rect 28365 10217 28399 10251
rect 30481 10217 30515 10251
rect 32505 10217 32539 10251
rect 32873 10217 32907 10251
rect 35449 10217 35483 10251
rect 35909 10217 35943 10251
rect 23020 10081 23054 10115
rect 27252 10081 27286 10115
rect 29837 10081 29871 10115
rect 33057 10081 33091 10115
rect 33425 10081 33459 10115
rect 33681 10081 33715 10115
rect 36277 10081 36311 10115
rect 22753 10013 22787 10047
rect 26985 10013 27019 10047
rect 29929 10013 29963 10047
rect 30113 10013 30147 10047
rect 36369 10013 36403 10047
rect 36553 10013 36587 10047
rect 29009 9945 29043 9979
rect 22477 9877 22511 9911
rect 26341 9877 26375 9911
rect 26709 9877 26743 9911
rect 29377 9877 29411 9911
rect 29469 9877 29503 9911
rect 34805 9877 34839 9911
rect 22845 9673 22879 9707
rect 29101 9673 29135 9707
rect 23489 9605 23523 9639
rect 25053 9605 25087 9639
rect 28733 9605 28767 9639
rect 33885 9605 33919 9639
rect 36277 9605 36311 9639
rect 30300 9537 30334 9571
rect 30573 9537 30607 9571
rect 32045 9537 32079 9571
rect 33057 9537 33091 9571
rect 33517 9537 33551 9571
rect 23673 9469 23707 9503
rect 23929 9469 23963 9503
rect 25697 9469 25731 9503
rect 26157 9469 26191 9503
rect 29837 9469 29871 9503
rect 32873 9469 32907 9503
rect 34897 9469 34931 9503
rect 37381 9469 37415 9503
rect 22477 9401 22511 9435
rect 26065 9401 26099 9435
rect 26402 9401 26436 9435
rect 32413 9401 32447 9435
rect 34253 9401 34287 9435
rect 34713 9401 34747 9435
rect 35164 9401 35198 9435
rect 27537 9333 27571 9367
rect 28181 9333 28215 9367
rect 29653 9333 29687 9367
rect 30303 9333 30337 9367
rect 31677 9333 31711 9367
rect 32505 9333 32539 9367
rect 32965 9333 32999 9367
rect 36829 9333 36863 9367
rect 24869 9129 24903 9163
rect 29009 9129 29043 9163
rect 30941 9129 30975 9163
rect 33063 9129 33097 9163
rect 34437 9129 34471 9163
rect 35173 9129 35207 9163
rect 35265 9129 35299 9163
rect 36277 9129 36311 9163
rect 36645 9129 36679 9163
rect 29828 9061 29862 9095
rect 23397 8993 23431 9027
rect 23489 8993 23523 9027
rect 23756 8993 23790 9027
rect 26157 8993 26191 9027
rect 26781 8993 26815 9027
rect 29285 8993 29319 9027
rect 35633 8993 35667 9027
rect 26525 8925 26559 8959
rect 28641 8925 28675 8959
rect 29561 8925 29595 8959
rect 32597 8925 32631 8959
rect 33060 8925 33094 8959
rect 33333 8925 33367 8959
rect 35173 8925 35207 8959
rect 35725 8925 35759 8959
rect 35817 8925 35851 8959
rect 25973 8857 26007 8891
rect 34989 8857 35023 8891
rect 27905 8789 27939 8823
rect 29101 8789 29135 8823
rect 31861 8789 31895 8823
rect 32413 8789 32447 8823
rect 23489 8585 23523 8619
rect 25513 8585 25547 8619
rect 26065 8585 26099 8619
rect 26433 8585 26467 8619
rect 26617 8585 26651 8619
rect 28273 8585 28307 8619
rect 29101 8585 29135 8619
rect 30757 8585 30791 8619
rect 31861 8585 31895 8619
rect 34253 8585 34287 8619
rect 34621 8585 34655 8619
rect 36277 8585 36311 8619
rect 37105 8585 37139 8619
rect 33701 8517 33735 8551
rect 34897 8517 34931 8551
rect 35909 8517 35943 8551
rect 27077 8449 27111 8483
rect 27169 8449 27203 8483
rect 29377 8449 29411 8483
rect 32321 8449 32355 8483
rect 35449 8449 35483 8483
rect 23121 8381 23155 8415
rect 24133 8381 24167 8415
rect 24400 8381 24434 8415
rect 26985 8381 27019 8415
rect 32045 8381 32079 8415
rect 35265 8381 35299 8415
rect 36461 8381 36495 8415
rect 24041 8313 24075 8347
rect 28733 8313 28767 8347
rect 29644 8313 29678 8347
rect 31309 8313 31343 8347
rect 32588 8313 32622 8347
rect 35357 8313 35391 8347
rect 27721 8245 27755 8279
rect 31769 8245 31803 8279
rect 36645 8245 36679 8279
rect 24225 8041 24259 8075
rect 26065 8041 26099 8075
rect 26801 8041 26835 8075
rect 27169 8041 27203 8075
rect 29745 8041 29779 8075
rect 30389 8041 30423 8075
rect 32321 8041 32355 8075
rect 33149 8041 33183 8075
rect 35357 8041 35391 8075
rect 28632 7973 28666 8007
rect 31953 7973 31987 8007
rect 32781 7973 32815 8007
rect 35725 7973 35759 8007
rect 32137 7905 32171 7939
rect 33241 7905 33275 7939
rect 33497 7905 33531 7939
rect 35909 7905 35943 7939
rect 28365 7837 28399 7871
rect 31033 7837 31067 7871
rect 34621 7701 34655 7735
rect 36093 7701 36127 7735
rect 28457 7497 28491 7531
rect 32045 7497 32079 7531
rect 32229 7497 32263 7531
rect 33977 7497 34011 7531
rect 35357 7497 35391 7531
rect 29469 7361 29503 7395
rect 31769 7361 31803 7395
rect 32873 7361 32907 7395
rect 31125 7293 31159 7327
rect 32597 7293 32631 7327
rect 33333 7293 33367 7327
rect 35449 7293 35483 7327
rect 31033 7225 31067 7259
rect 32689 7225 32723 7259
rect 33609 7225 33643 7259
rect 34713 7225 34747 7259
rect 35716 7225 35750 7259
rect 28733 7157 28767 7191
rect 31309 7157 31343 7191
rect 36829 7157 36863 7191
rect 32321 6953 32355 6987
rect 32689 6953 32723 6987
rect 36277 6953 36311 6987
rect 33057 6885 33091 6919
rect 26792 6817 26826 6851
rect 30297 6817 30331 6851
rect 31769 6817 31803 6851
rect 34253 6817 34287 6851
rect 35357 6817 35391 6851
rect 36461 6817 36495 6851
rect 26525 6749 26559 6783
rect 33149 6749 33183 6783
rect 33333 6749 33367 6783
rect 34437 6681 34471 6715
rect 27905 6613 27939 6647
rect 29377 6613 29411 6647
rect 30481 6613 30515 6647
rect 31401 6613 31435 6647
rect 33793 6613 33827 6647
rect 35541 6613 35575 6647
rect 36001 6613 36035 6647
rect 36645 6613 36679 6647
rect 26617 6409 26651 6443
rect 30849 6409 30883 6443
rect 32413 6409 32447 6443
rect 32781 6409 32815 6443
rect 36553 6409 36587 6443
rect 37013 6409 37047 6443
rect 27629 6341 27663 6375
rect 29009 6341 29043 6375
rect 29285 6341 29319 6375
rect 30297 6341 30331 6375
rect 32873 6341 32907 6375
rect 34253 6341 34287 6375
rect 37289 6341 37323 6375
rect 27537 6273 27571 6307
rect 28089 6273 28123 6307
rect 28273 6273 28307 6307
rect 29745 6273 29779 6307
rect 29837 6273 29871 6307
rect 31953 6273 31987 6307
rect 33517 6273 33551 6307
rect 31217 6205 31251 6239
rect 33241 6205 33275 6239
rect 33885 6205 33919 6239
rect 34897 6205 34931 6239
rect 36001 6205 36035 6239
rect 37105 6205 37139 6239
rect 37657 6205 37691 6239
rect 31769 6137 31803 6171
rect 26249 6069 26283 6103
rect 27169 6069 27203 6103
rect 27997 6069 28031 6103
rect 28733 6069 28767 6103
rect 29653 6069 29687 6103
rect 31033 6069 31067 6103
rect 31309 6069 31343 6103
rect 31677 6069 31711 6103
rect 33333 6069 33367 6103
rect 34621 6069 34655 6103
rect 35081 6069 35115 6103
rect 35449 6069 35483 6103
rect 36185 6069 36219 6103
rect 28733 5865 28767 5899
rect 31401 5865 31435 5899
rect 33517 5865 33551 5899
rect 27620 5797 27654 5831
rect 31953 5797 31987 5831
rect 32965 5797 32999 5831
rect 33609 5797 33643 5831
rect 30205 5729 30239 5763
rect 35357 5729 35391 5763
rect 27353 5661 27387 5695
rect 30297 5661 30331 5695
rect 30389 5661 30423 5695
rect 33793 5661 33827 5695
rect 34897 5661 34931 5695
rect 35449 5661 35483 5695
rect 35541 5661 35575 5695
rect 29745 5593 29779 5627
rect 33149 5593 33183 5627
rect 34989 5593 35023 5627
rect 29285 5525 29319 5559
rect 29837 5525 29871 5559
rect 32505 5525 32539 5559
rect 36093 5525 36127 5559
rect 27445 5321 27479 5355
rect 27629 5321 27663 5355
rect 31217 5321 31251 5355
rect 32413 5321 32447 5355
rect 33517 5321 33551 5355
rect 33885 5321 33919 5355
rect 34253 5321 34287 5355
rect 36829 5321 36863 5355
rect 28273 5185 28307 5219
rect 31953 5185 31987 5219
rect 33057 5185 33091 5219
rect 35449 5185 35483 5219
rect 29285 5117 29319 5151
rect 29009 5049 29043 5083
rect 29530 5049 29564 5083
rect 32873 5049 32907 5083
rect 35716 5049 35750 5083
rect 26709 4981 26743 5015
rect 27077 4981 27111 5015
rect 27997 4981 28031 5015
rect 28089 4981 28123 5015
rect 28733 4981 28767 5015
rect 30665 4981 30699 5015
rect 32229 4981 32263 5015
rect 32781 4981 32815 5015
rect 34713 4981 34747 5015
rect 35173 4981 35207 5015
rect 27721 4777 27755 4811
rect 29285 4777 29319 4811
rect 30205 4777 30239 4811
rect 30389 4777 30423 4811
rect 32321 4777 32355 4811
rect 33609 4777 33643 4811
rect 34069 4777 34103 4811
rect 34713 4777 34747 4811
rect 28172 4709 28206 4743
rect 27905 4641 27939 4675
rect 30757 4641 30791 4675
rect 30849 4641 30883 4675
rect 32137 4641 32171 4675
rect 32689 4641 32723 4675
rect 33977 4641 34011 4675
rect 35429 4641 35463 4675
rect 31033 4573 31067 4607
rect 33517 4573 33551 4607
rect 34253 4573 34287 4607
rect 34989 4573 35023 4607
rect 35173 4573 35207 4607
rect 29837 4437 29871 4471
rect 36553 4437 36587 4471
rect 28641 4233 28675 4267
rect 33793 4233 33827 4267
rect 34713 4233 34747 4267
rect 27169 4097 27203 4131
rect 28273 4097 28307 4131
rect 29101 4097 29135 4131
rect 27537 4029 27571 4063
rect 28089 4029 28123 4063
rect 29285 4029 29319 4063
rect 29541 4029 29575 4063
rect 31585 4029 31619 4063
rect 31769 4029 31803 4063
rect 35449 4029 35483 4063
rect 31217 3961 31251 3995
rect 32014 3961 32048 3995
rect 35357 3961 35391 3995
rect 35716 3961 35750 3995
rect 26801 3893 26835 3927
rect 27629 3893 27663 3927
rect 27997 3893 28031 3927
rect 30665 3893 30699 3927
rect 33149 3893 33183 3927
rect 34161 3893 34195 3927
rect 36829 3893 36863 3927
rect 27353 3689 27387 3723
rect 28457 3689 28491 3723
rect 28825 3689 28859 3723
rect 30297 3689 30331 3723
rect 31217 3689 31251 3723
rect 35449 3689 35483 3723
rect 35725 3689 35759 3723
rect 35909 3689 35943 3723
rect 29184 3621 29218 3655
rect 36369 3621 36403 3655
rect 27721 3553 27755 3587
rect 28917 3553 28951 3587
rect 32321 3553 32355 3587
rect 33692 3553 33726 3587
rect 36277 3553 36311 3587
rect 27813 3485 27847 3519
rect 27997 3485 28031 3519
rect 31861 3485 31895 3519
rect 32965 3485 32999 3519
rect 33425 3485 33459 3519
rect 36461 3485 36495 3519
rect 32505 3417 32539 3451
rect 30849 3349 30883 3383
rect 34805 3349 34839 3383
rect 27169 3145 27203 3179
rect 29009 3145 29043 3179
rect 31585 3145 31619 3179
rect 37197 3145 37231 3179
rect 26801 3077 26835 3111
rect 36829 3077 36863 3111
rect 27537 3009 27571 3043
rect 28089 3009 28123 3043
rect 28181 3009 28215 3043
rect 31309 3009 31343 3043
rect 31769 3009 31803 3043
rect 33701 3009 33735 3043
rect 37565 3009 37599 3043
rect 29285 2941 29319 2975
rect 32036 2941 32070 2975
rect 34161 2941 34195 2975
rect 34897 2941 34931 2975
rect 29530 2873 29564 2907
rect 35142 2873 35176 2907
rect 27629 2805 27663 2839
rect 27997 2805 28031 2839
rect 30665 2805 30699 2839
rect 33149 2805 33183 2839
rect 34621 2805 34655 2839
rect 36277 2805 36311 2839
rect 27721 2601 27755 2635
rect 28089 2601 28123 2635
rect 29377 2601 29411 2635
rect 31125 2601 31159 2635
rect 31953 2601 31987 2635
rect 32413 2601 32447 2635
rect 33977 2601 34011 2635
rect 34529 2601 34563 2635
rect 35265 2601 35299 2635
rect 36829 2601 36863 2635
rect 27353 2533 27387 2567
rect 29009 2533 29043 2567
rect 29990 2533 30024 2567
rect 32842 2533 32876 2567
rect 35694 2533 35728 2567
rect 26709 2465 26743 2499
rect 28641 2465 28675 2499
rect 29745 2465 29779 2499
rect 32597 2465 32631 2499
rect 35449 2465 35483 2499
rect 37381 2465 37415 2499
rect 8401 2261 8435 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 19606 37562
rect 19658 37510 19670 37562
rect 19722 37510 19734 37562
rect 19786 37510 19798 37562
rect 19850 37510 38824 37562
rect 1104 37488 38824 37510
rect 1104 37018 38824 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 34966 37018
rect 35018 36966 35030 37018
rect 35082 36966 35094 37018
rect 35146 36966 35158 37018
rect 35210 36966 38824 37018
rect 1104 36944 38824 36966
rect 1104 36474 38824 36496
rect 1104 36422 19606 36474
rect 19658 36422 19670 36474
rect 19722 36422 19734 36474
rect 19786 36422 19798 36474
rect 19850 36422 38824 36474
rect 1104 36400 38824 36422
rect 5629 36363 5687 36369
rect 5629 36329 5641 36363
rect 5675 36360 5687 36363
rect 6086 36360 6092 36372
rect 5675 36332 6092 36360
rect 5675 36329 5687 36332
rect 5629 36323 5687 36329
rect 6086 36320 6092 36332
rect 6144 36320 6150 36372
rect 6825 36363 6883 36369
rect 6825 36329 6837 36363
rect 6871 36360 6883 36363
rect 7190 36360 7196 36372
rect 6871 36332 7196 36360
rect 6871 36329 6883 36332
rect 6825 36323 6883 36329
rect 7190 36320 7196 36332
rect 7248 36320 7254 36372
rect 5442 36224 5448 36236
rect 5403 36196 5448 36224
rect 5442 36184 5448 36196
rect 5500 36184 5506 36236
rect 6638 36224 6644 36236
rect 6599 36196 6644 36224
rect 6638 36184 6644 36196
rect 6696 36184 6702 36236
rect 22373 36227 22431 36233
rect 22373 36193 22385 36227
rect 22419 36224 22431 36227
rect 22462 36224 22468 36236
rect 22419 36196 22468 36224
rect 22419 36193 22431 36196
rect 22373 36187 22431 36193
rect 22462 36184 22468 36196
rect 22520 36224 22526 36236
rect 23842 36224 23848 36236
rect 22520 36196 23848 36224
rect 22520 36184 22526 36196
rect 23842 36184 23848 36196
rect 23900 36184 23906 36236
rect 14185 36023 14243 36029
rect 14185 35989 14197 36023
rect 14231 36020 14243 36023
rect 14550 36020 14556 36032
rect 14231 35992 14556 36020
rect 14231 35989 14243 35992
rect 14185 35983 14243 35989
rect 14550 35980 14556 35992
rect 14608 35980 14614 36032
rect 21450 36020 21456 36032
rect 21411 35992 21456 36020
rect 21450 35980 21456 35992
rect 21508 35980 21514 36032
rect 22554 36020 22560 36032
rect 22515 35992 22560 36020
rect 22554 35980 22560 35992
rect 22612 35980 22618 36032
rect 1104 35930 38824 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 34966 35930
rect 35018 35878 35030 35930
rect 35082 35878 35094 35930
rect 35146 35878 35158 35930
rect 35210 35878 38824 35930
rect 1104 35856 38824 35878
rect 4525 35819 4583 35825
rect 4525 35785 4537 35819
rect 4571 35816 4583 35819
rect 4982 35816 4988 35828
rect 4571 35788 4988 35816
rect 4571 35785 4583 35788
rect 4525 35779 4583 35785
rect 4982 35776 4988 35788
rect 5040 35776 5046 35828
rect 6273 35819 6331 35825
rect 6273 35785 6285 35819
rect 6319 35816 6331 35819
rect 6822 35816 6828 35828
rect 6319 35788 6828 35816
rect 6319 35785 6331 35788
rect 6273 35779 6331 35785
rect 5258 35708 5264 35760
rect 5316 35748 5322 35760
rect 5813 35751 5871 35757
rect 5813 35748 5825 35751
rect 5316 35720 5825 35748
rect 5316 35708 5322 35720
rect 5813 35717 5825 35720
rect 5859 35717 5871 35751
rect 5813 35711 5871 35717
rect 4341 35615 4399 35621
rect 4341 35581 4353 35615
rect 4387 35612 4399 35615
rect 5629 35615 5687 35621
rect 4387 35584 5028 35612
rect 4387 35581 4399 35584
rect 4341 35575 4399 35581
rect 5000 35488 5028 35584
rect 5629 35581 5641 35615
rect 5675 35612 5687 35615
rect 6288 35612 6316 35779
rect 6822 35776 6828 35788
rect 6880 35776 6886 35828
rect 7466 35816 7472 35828
rect 7427 35788 7472 35816
rect 7466 35776 7472 35788
rect 7524 35776 7530 35828
rect 8113 35819 8171 35825
rect 8113 35785 8125 35819
rect 8159 35816 8171 35819
rect 8202 35816 8208 35828
rect 8159 35788 8208 35816
rect 8159 35785 8171 35788
rect 8113 35779 8171 35785
rect 8202 35776 8208 35788
rect 8260 35776 8266 35828
rect 11882 35816 11888 35828
rect 11843 35788 11888 35816
rect 11882 35776 11888 35788
rect 11940 35776 11946 35828
rect 22462 35816 22468 35828
rect 22423 35788 22468 35816
rect 22462 35776 22468 35788
rect 22520 35776 22526 35828
rect 24305 35819 24363 35825
rect 24305 35785 24317 35819
rect 24351 35816 24363 35819
rect 24762 35816 24768 35828
rect 24351 35788 24768 35816
rect 24351 35785 24363 35788
rect 24305 35779 24363 35785
rect 6638 35748 6644 35760
rect 6599 35720 6644 35748
rect 6638 35708 6644 35720
rect 6696 35708 6702 35760
rect 14093 35751 14151 35757
rect 14093 35717 14105 35751
rect 14139 35748 14151 35751
rect 15289 35751 15347 35757
rect 15289 35748 15301 35751
rect 14139 35720 15301 35748
rect 14139 35717 14151 35720
rect 14093 35711 14151 35717
rect 15289 35717 15301 35720
rect 15335 35748 15347 35751
rect 15746 35748 15752 35760
rect 15335 35720 15752 35748
rect 15335 35717 15347 35720
rect 15289 35711 15347 35717
rect 15746 35708 15752 35720
rect 15804 35708 15810 35760
rect 23845 35751 23903 35757
rect 23845 35717 23857 35751
rect 23891 35717 23903 35751
rect 23845 35711 23903 35717
rect 13633 35683 13691 35689
rect 13633 35649 13645 35683
rect 13679 35680 13691 35683
rect 14645 35683 14703 35689
rect 14645 35680 14657 35683
rect 13679 35652 14657 35680
rect 13679 35649 13691 35652
rect 13633 35643 13691 35649
rect 14645 35649 14657 35652
rect 14691 35680 14703 35683
rect 14918 35680 14924 35692
rect 14691 35652 14924 35680
rect 14691 35649 14703 35652
rect 14645 35643 14703 35649
rect 14918 35640 14924 35652
rect 14976 35640 14982 35692
rect 20901 35683 20959 35689
rect 20901 35649 20913 35683
rect 20947 35680 20959 35683
rect 21913 35683 21971 35689
rect 21913 35680 21925 35683
rect 20947 35652 21925 35680
rect 20947 35649 20959 35652
rect 20901 35643 20959 35649
rect 21913 35649 21925 35652
rect 21959 35680 21971 35683
rect 22094 35680 22100 35692
rect 21959 35652 22100 35680
rect 21959 35649 21971 35652
rect 21913 35643 21971 35649
rect 22094 35640 22100 35652
rect 22152 35680 22158 35692
rect 23860 35680 23888 35711
rect 22152 35652 23888 35680
rect 22152 35640 22158 35652
rect 5675 35584 6316 35612
rect 6825 35615 6883 35621
rect 5675 35581 5687 35584
rect 5629 35575 5687 35581
rect 6825 35581 6837 35615
rect 6871 35612 6883 35615
rect 7466 35612 7472 35624
rect 6871 35584 7472 35612
rect 6871 35581 6883 35584
rect 6825 35575 6883 35581
rect 7466 35572 7472 35584
rect 7524 35572 7530 35624
rect 7929 35615 7987 35621
rect 7929 35581 7941 35615
rect 7975 35612 7987 35615
rect 11241 35615 11299 35621
rect 7975 35584 8616 35612
rect 7975 35581 7987 35584
rect 7929 35575 7987 35581
rect 8588 35556 8616 35584
rect 11241 35581 11253 35615
rect 11287 35612 11299 35615
rect 11882 35612 11888 35624
rect 11287 35584 11888 35612
rect 11287 35581 11299 35584
rect 11241 35575 11299 35581
rect 11882 35572 11888 35584
rect 11940 35572 11946 35624
rect 13081 35615 13139 35621
rect 13081 35581 13093 35615
rect 13127 35612 13139 35615
rect 13538 35612 13544 35624
rect 13127 35584 13544 35612
rect 13127 35581 13139 35584
rect 13081 35575 13139 35581
rect 13538 35572 13544 35584
rect 13596 35572 13602 35624
rect 14001 35615 14059 35621
rect 14001 35581 14013 35615
rect 14047 35612 14059 35615
rect 14458 35612 14464 35624
rect 14047 35584 14464 35612
rect 14047 35581 14059 35584
rect 14001 35575 14059 35581
rect 14458 35572 14464 35584
rect 14516 35572 14522 35624
rect 20990 35572 20996 35624
rect 21048 35612 21054 35624
rect 21450 35612 21456 35624
rect 21048 35584 21456 35612
rect 21048 35572 21054 35584
rect 21450 35572 21456 35584
rect 21508 35612 21514 35624
rect 21729 35615 21787 35621
rect 21729 35612 21741 35615
rect 21508 35584 21741 35612
rect 21508 35572 21514 35584
rect 21729 35581 21741 35584
rect 21775 35581 21787 35615
rect 21729 35575 21787 35581
rect 23661 35615 23719 35621
rect 23661 35581 23673 35615
rect 23707 35612 23719 35615
rect 24320 35612 24348 35779
rect 24762 35776 24768 35788
rect 24820 35776 24826 35828
rect 35618 35816 35624 35828
rect 35579 35788 35624 35816
rect 35618 35776 35624 35788
rect 35676 35776 35682 35828
rect 25682 35612 25688 35624
rect 23707 35584 24348 35612
rect 25643 35584 25688 35612
rect 23707 35581 23719 35584
rect 23661 35575 23719 35581
rect 25682 35572 25688 35584
rect 25740 35572 25746 35624
rect 35437 35615 35495 35621
rect 35437 35581 35449 35615
rect 35483 35612 35495 35615
rect 35618 35612 35624 35624
rect 35483 35584 35624 35612
rect 35483 35581 35495 35584
rect 35437 35575 35495 35581
rect 35618 35572 35624 35584
rect 35676 35612 35682 35624
rect 35989 35615 36047 35621
rect 35989 35612 36001 35615
rect 35676 35584 36001 35612
rect 35676 35572 35682 35584
rect 35989 35581 36001 35584
rect 36035 35581 36047 35615
rect 35989 35575 36047 35581
rect 8570 35544 8576 35556
rect 8531 35516 8576 35544
rect 8570 35504 8576 35516
rect 8628 35504 8634 35556
rect 21821 35547 21879 35553
rect 21821 35544 21833 35547
rect 21192 35516 21833 35544
rect 21192 35488 21220 35516
rect 21821 35513 21833 35516
rect 21867 35513 21879 35547
rect 25590 35544 25596 35556
rect 25503 35516 25596 35544
rect 21821 35507 21879 35513
rect 25590 35504 25596 35516
rect 25648 35544 25654 35556
rect 25930 35547 25988 35553
rect 25930 35544 25942 35547
rect 25648 35516 25942 35544
rect 25648 35504 25654 35516
rect 25930 35513 25942 35516
rect 25976 35513 25988 35547
rect 25930 35507 25988 35513
rect 4982 35476 4988 35488
rect 4943 35448 4988 35476
rect 4982 35436 4988 35448
rect 5040 35436 5046 35488
rect 5534 35476 5540 35488
rect 5495 35448 5540 35476
rect 5534 35436 5540 35448
rect 5592 35436 5598 35488
rect 7009 35479 7067 35485
rect 7009 35445 7021 35479
rect 7055 35476 7067 35479
rect 7466 35476 7472 35488
rect 7055 35448 7472 35476
rect 7055 35445 7067 35448
rect 7009 35439 7067 35445
rect 7466 35436 7472 35448
rect 7524 35436 7530 35488
rect 11054 35436 11060 35488
rect 11112 35476 11118 35488
rect 11425 35479 11483 35485
rect 11425 35476 11437 35479
rect 11112 35448 11437 35476
rect 11112 35436 11118 35448
rect 11425 35445 11437 35448
rect 11471 35445 11483 35479
rect 14550 35476 14556 35488
rect 14511 35448 14556 35476
rect 11425 35439 11483 35445
rect 14550 35436 14556 35448
rect 14608 35436 14614 35488
rect 16482 35436 16488 35488
rect 16540 35476 16546 35488
rect 16761 35479 16819 35485
rect 16761 35476 16773 35479
rect 16540 35448 16773 35476
rect 16540 35436 16546 35448
rect 16761 35445 16773 35448
rect 16807 35445 16819 35479
rect 21174 35476 21180 35488
rect 21135 35448 21180 35476
rect 16761 35439 16819 35445
rect 21174 35436 21180 35448
rect 21232 35436 21238 35488
rect 21358 35476 21364 35488
rect 21319 35448 21364 35476
rect 21358 35436 21364 35448
rect 21416 35436 21422 35488
rect 26970 35436 26976 35488
rect 27028 35476 27034 35488
rect 27065 35479 27123 35485
rect 27065 35476 27077 35479
rect 27028 35448 27077 35476
rect 27028 35436 27034 35448
rect 27065 35445 27077 35448
rect 27111 35445 27123 35479
rect 27065 35439 27123 35445
rect 1104 35386 38824 35408
rect 1104 35334 19606 35386
rect 19658 35334 19670 35386
rect 19722 35334 19734 35386
rect 19786 35334 19798 35386
rect 19850 35334 38824 35386
rect 1104 35312 38824 35334
rect 1581 35275 1639 35281
rect 1581 35241 1593 35275
rect 1627 35272 1639 35275
rect 1670 35272 1676 35284
rect 1627 35244 1676 35272
rect 1627 35241 1639 35244
rect 1581 35235 1639 35241
rect 1670 35232 1676 35244
rect 1728 35232 1734 35284
rect 10870 35272 10876 35284
rect 10831 35244 10876 35272
rect 10870 35232 10876 35244
rect 10928 35232 10934 35284
rect 15746 35272 15752 35284
rect 15707 35244 15752 35272
rect 15746 35232 15752 35244
rect 15804 35232 15810 35284
rect 35526 35272 35532 35284
rect 35487 35244 35532 35272
rect 35526 35232 35532 35244
rect 35584 35232 35590 35284
rect 8113 35207 8171 35213
rect 8113 35173 8125 35207
rect 8159 35204 8171 35207
rect 8846 35204 8852 35216
rect 8159 35176 8852 35204
rect 8159 35173 8171 35176
rect 8113 35167 8171 35173
rect 8846 35164 8852 35176
rect 8904 35164 8910 35216
rect 13633 35207 13691 35213
rect 13633 35173 13645 35207
rect 13679 35204 13691 35207
rect 13722 35204 13728 35216
rect 13679 35176 13728 35204
rect 13679 35173 13691 35176
rect 13633 35167 13691 35173
rect 13722 35164 13728 35176
rect 13780 35164 13786 35216
rect 21082 35164 21088 35216
rect 21140 35204 21146 35216
rect 21177 35207 21235 35213
rect 21177 35204 21189 35207
rect 21140 35176 21189 35204
rect 21140 35164 21146 35176
rect 21177 35173 21189 35176
rect 21223 35204 21235 35207
rect 22922 35204 22928 35216
rect 21223 35176 22928 35204
rect 21223 35173 21235 35176
rect 21177 35167 21235 35173
rect 1394 35136 1400 35148
rect 1355 35108 1400 35136
rect 1394 35096 1400 35108
rect 1452 35096 1458 35148
rect 4982 35136 4988 35148
rect 4943 35108 4988 35136
rect 4982 35096 4988 35108
rect 5040 35096 5046 35148
rect 6822 35136 6828 35148
rect 6783 35108 6828 35136
rect 6822 35096 6828 35108
rect 6880 35096 6886 35148
rect 8294 35136 8300 35148
rect 8255 35108 8300 35136
rect 8294 35096 8300 35108
rect 8352 35096 8358 35148
rect 11238 35136 11244 35148
rect 11199 35108 11244 35136
rect 11238 35096 11244 35108
rect 11296 35096 11302 35148
rect 13538 35136 13544 35148
rect 13499 35108 13544 35136
rect 13538 35096 13544 35108
rect 13596 35096 13602 35148
rect 14826 35096 14832 35148
rect 14884 35136 14890 35148
rect 15657 35139 15715 35145
rect 15657 35136 15669 35139
rect 14884 35108 15669 35136
rect 14884 35096 14890 35108
rect 15657 35105 15669 35108
rect 15703 35105 15715 35139
rect 15657 35099 15715 35105
rect 16853 35139 16911 35145
rect 16853 35105 16865 35139
rect 16899 35136 16911 35139
rect 16942 35136 16948 35148
rect 16899 35108 16948 35136
rect 16899 35105 16911 35108
rect 16853 35099 16911 35105
rect 16942 35096 16948 35108
rect 17000 35136 17006 35148
rect 18322 35136 18328 35148
rect 17000 35108 18328 35136
rect 17000 35096 17006 35108
rect 18322 35096 18328 35108
rect 18380 35096 18386 35148
rect 21269 35139 21327 35145
rect 21269 35105 21281 35139
rect 21315 35136 21327 35139
rect 21910 35136 21916 35148
rect 21315 35108 21916 35136
rect 21315 35105 21327 35108
rect 21269 35099 21327 35105
rect 21910 35096 21916 35108
rect 21968 35096 21974 35148
rect 22388 35145 22416 35176
rect 22922 35164 22928 35176
rect 22980 35164 22986 35216
rect 22373 35139 22431 35145
rect 22373 35105 22385 35139
rect 22419 35105 22431 35139
rect 22373 35099 22431 35105
rect 22462 35096 22468 35148
rect 22520 35136 22526 35148
rect 22629 35139 22687 35145
rect 22629 35136 22641 35139
rect 22520 35108 22641 35136
rect 22520 35096 22526 35108
rect 22629 35105 22641 35108
rect 22675 35105 22687 35139
rect 22629 35099 22687 35105
rect 27700 35139 27758 35145
rect 27700 35105 27712 35139
rect 27746 35136 27758 35139
rect 28074 35136 28080 35148
rect 27746 35108 28080 35136
rect 27746 35105 27758 35108
rect 27700 35099 27758 35105
rect 28074 35096 28080 35108
rect 28132 35096 28138 35148
rect 35342 35136 35348 35148
rect 35303 35108 35348 35136
rect 35342 35096 35348 35108
rect 35400 35096 35406 35148
rect 5074 35068 5080 35080
rect 5035 35040 5080 35068
rect 5074 35028 5080 35040
rect 5132 35028 5138 35080
rect 5258 35068 5264 35080
rect 5219 35040 5264 35068
rect 5258 35028 5264 35040
rect 5316 35028 5322 35080
rect 9677 35071 9735 35077
rect 9677 35037 9689 35071
rect 9723 35068 9735 35071
rect 10042 35068 10048 35080
rect 9723 35040 10048 35068
rect 9723 35037 9735 35040
rect 9677 35031 9735 35037
rect 10042 35028 10048 35040
rect 10100 35028 10106 35080
rect 11330 35068 11336 35080
rect 11291 35040 11336 35068
rect 11330 35028 11336 35040
rect 11388 35028 11394 35080
rect 11517 35071 11575 35077
rect 11517 35037 11529 35071
rect 11563 35068 11575 35071
rect 12526 35068 12532 35080
rect 11563 35040 12532 35068
rect 11563 35037 11575 35040
rect 11517 35031 11575 35037
rect 12526 35028 12532 35040
rect 12584 35028 12590 35080
rect 13081 35071 13139 35077
rect 13081 35037 13093 35071
rect 13127 35068 13139 35071
rect 13725 35071 13783 35077
rect 13725 35068 13737 35071
rect 13127 35040 13737 35068
rect 13127 35037 13139 35040
rect 13081 35031 13139 35037
rect 13725 35037 13737 35040
rect 13771 35068 13783 35071
rect 14366 35068 14372 35080
rect 13771 35040 14372 35068
rect 13771 35037 13783 35040
rect 13725 35031 13783 35037
rect 14366 35028 14372 35040
rect 14424 35068 14430 35080
rect 14921 35071 14979 35077
rect 14921 35068 14933 35071
rect 14424 35040 14933 35068
rect 14424 35028 14430 35040
rect 14921 35037 14933 35040
rect 14967 35068 14979 35071
rect 15194 35068 15200 35080
rect 14967 35040 15200 35068
rect 14967 35037 14979 35040
rect 14921 35031 14979 35037
rect 15194 35028 15200 35040
rect 15252 35028 15258 35080
rect 15470 35028 15476 35080
rect 15528 35068 15534 35080
rect 15841 35071 15899 35077
rect 15841 35068 15853 35071
rect 15528 35040 15853 35068
rect 15528 35028 15534 35040
rect 15841 35037 15853 35040
rect 15887 35037 15899 35071
rect 15841 35031 15899 35037
rect 17862 35028 17868 35080
rect 17920 35068 17926 35080
rect 17957 35071 18015 35077
rect 17957 35068 17969 35071
rect 17920 35040 17969 35068
rect 17920 35028 17926 35040
rect 17957 35037 17969 35040
rect 18003 35037 18015 35071
rect 17957 35031 18015 35037
rect 27433 35071 27491 35077
rect 27433 35037 27445 35071
rect 27479 35037 27491 35071
rect 27433 35031 27491 35037
rect 4341 35003 4399 35009
rect 4341 34969 4353 35003
rect 4387 35000 4399 35003
rect 4706 35000 4712 35012
rect 4387 34972 4712 35000
rect 4387 34969 4399 34972
rect 4341 34963 4399 34969
rect 4706 34960 4712 34972
rect 4764 34960 4770 35012
rect 6914 34960 6920 35012
rect 6972 35000 6978 35012
rect 7377 35003 7435 35009
rect 7377 35000 7389 35003
rect 6972 34972 7389 35000
rect 6972 34960 6978 34972
rect 7377 34969 7389 34972
rect 7423 34969 7435 35003
rect 7377 34963 7435 34969
rect 13173 35003 13231 35009
rect 13173 34969 13185 35003
rect 13219 35000 13231 35003
rect 13630 35000 13636 35012
rect 13219 34972 13636 35000
rect 13219 34969 13231 34972
rect 13173 34963 13231 34969
rect 13630 34960 13636 34972
rect 13688 34960 13694 35012
rect 4617 34935 4675 34941
rect 4617 34901 4629 34935
rect 4663 34932 4675 34935
rect 5442 34932 5448 34944
rect 4663 34904 5448 34932
rect 4663 34901 4675 34904
rect 4617 34895 4675 34901
rect 5442 34892 5448 34904
rect 5500 34892 5506 34944
rect 7009 34935 7067 34941
rect 7009 34901 7021 34935
rect 7055 34932 7067 34935
rect 7098 34932 7104 34944
rect 7055 34904 7104 34932
rect 7055 34901 7067 34904
rect 7009 34895 7067 34901
rect 7098 34892 7104 34904
rect 7156 34892 7162 34944
rect 8478 34932 8484 34944
rect 8439 34904 8484 34932
rect 8478 34892 8484 34904
rect 8536 34892 8542 34944
rect 9858 34892 9864 34944
rect 9916 34932 9922 34944
rect 10137 34935 10195 34941
rect 10137 34932 10149 34935
rect 9916 34904 10149 34932
rect 9916 34892 9922 34904
rect 10137 34901 10149 34904
rect 10183 34932 10195 34935
rect 12066 34932 12072 34944
rect 10183 34904 12072 34932
rect 10183 34901 10195 34904
rect 10137 34895 10195 34901
rect 12066 34892 12072 34904
rect 12124 34892 12130 34944
rect 14642 34932 14648 34944
rect 14603 34904 14648 34932
rect 14642 34892 14648 34904
rect 14700 34892 14706 34944
rect 15289 34935 15347 34941
rect 15289 34901 15301 34935
rect 15335 34932 15347 34935
rect 15746 34932 15752 34944
rect 15335 34904 15752 34932
rect 15335 34901 15347 34904
rect 15289 34895 15347 34901
rect 15746 34892 15752 34904
rect 15804 34892 15810 34944
rect 17037 34935 17095 34941
rect 17037 34901 17049 34935
rect 17083 34932 17095 34935
rect 17402 34932 17408 34944
rect 17083 34904 17408 34932
rect 17083 34901 17095 34904
rect 17037 34895 17095 34901
rect 17402 34892 17408 34904
rect 17460 34892 17466 34944
rect 18506 34932 18512 34944
rect 18467 34904 18512 34932
rect 18506 34892 18512 34904
rect 18564 34892 18570 34944
rect 21450 34932 21456 34944
rect 21411 34904 21456 34932
rect 21450 34892 21456 34904
rect 21508 34892 21514 34944
rect 21910 34932 21916 34944
rect 21871 34904 21916 34932
rect 21910 34892 21916 34904
rect 21968 34892 21974 34944
rect 23753 34935 23811 34941
rect 23753 34901 23765 34935
rect 23799 34932 23811 34935
rect 24026 34932 24032 34944
rect 23799 34904 24032 34932
rect 23799 34901 23811 34904
rect 23753 34895 23811 34901
rect 24026 34892 24032 34904
rect 24084 34892 24090 34944
rect 24210 34892 24216 34944
rect 24268 34932 24274 34944
rect 24305 34935 24363 34941
rect 24305 34932 24317 34935
rect 24268 34904 24317 34932
rect 24268 34892 24274 34904
rect 24305 34901 24317 34904
rect 24351 34901 24363 34935
rect 24305 34895 24363 34901
rect 25682 34892 25688 34944
rect 25740 34932 25746 34944
rect 25777 34935 25835 34941
rect 25777 34932 25789 34935
rect 25740 34904 25789 34932
rect 25740 34892 25746 34904
rect 25777 34901 25789 34904
rect 25823 34932 25835 34935
rect 26694 34932 26700 34944
rect 25823 34904 26700 34932
rect 25823 34901 25835 34904
rect 25777 34895 25835 34901
rect 26694 34892 26700 34904
rect 26752 34932 26758 34944
rect 26789 34935 26847 34941
rect 26789 34932 26801 34935
rect 26752 34904 26801 34932
rect 26752 34892 26758 34904
rect 26789 34901 26801 34904
rect 26835 34932 26847 34935
rect 27448 34932 27476 35031
rect 28350 34932 28356 34944
rect 26835 34904 28356 34932
rect 26835 34901 26847 34904
rect 26789 34895 26847 34901
rect 28350 34892 28356 34904
rect 28408 34892 28414 34944
rect 28810 34932 28816 34944
rect 28771 34904 28816 34932
rect 28810 34892 28816 34904
rect 28868 34892 28874 34944
rect 1104 34842 38824 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 34966 34842
rect 35018 34790 35030 34842
rect 35082 34790 35094 34842
rect 35146 34790 35158 34842
rect 35210 34790 38824 34842
rect 1104 34768 38824 34790
rect 566 34688 572 34740
rect 624 34728 630 34740
rect 1581 34731 1639 34737
rect 1581 34728 1593 34731
rect 624 34700 1593 34728
rect 624 34688 630 34700
rect 1581 34697 1593 34700
rect 1627 34697 1639 34731
rect 2038 34728 2044 34740
rect 1999 34700 2044 34728
rect 1581 34691 1639 34697
rect 2038 34688 2044 34700
rect 2096 34688 2102 34740
rect 3142 34728 3148 34740
rect 3103 34700 3148 34728
rect 3142 34688 3148 34700
rect 3200 34688 3206 34740
rect 4249 34731 4307 34737
rect 4249 34697 4261 34731
rect 4295 34728 4307 34731
rect 5074 34728 5080 34740
rect 4295 34700 5080 34728
rect 4295 34697 4307 34700
rect 4249 34691 4307 34697
rect 5074 34688 5080 34700
rect 5132 34728 5138 34740
rect 5261 34731 5319 34737
rect 5261 34728 5273 34731
rect 5132 34700 5273 34728
rect 5132 34688 5138 34700
rect 5261 34697 5273 34700
rect 5307 34697 5319 34731
rect 5261 34691 5319 34697
rect 6641 34731 6699 34737
rect 6641 34697 6653 34731
rect 6687 34728 6699 34731
rect 6822 34728 6828 34740
rect 6687 34700 6828 34728
rect 6687 34697 6699 34700
rect 6641 34691 6699 34697
rect 6822 34688 6828 34700
rect 6880 34688 6886 34740
rect 8846 34728 8852 34740
rect 8807 34700 8852 34728
rect 8846 34688 8852 34700
rect 8904 34688 8910 34740
rect 11238 34688 11244 34740
rect 11296 34728 11302 34740
rect 11701 34731 11759 34737
rect 11701 34728 11713 34731
rect 11296 34700 11713 34728
rect 11296 34688 11302 34700
rect 11701 34697 11713 34700
rect 11747 34697 11759 34731
rect 11701 34691 11759 34697
rect 13538 34688 13544 34740
rect 13596 34728 13602 34740
rect 14369 34731 14427 34737
rect 14369 34728 14381 34731
rect 13596 34700 14381 34728
rect 13596 34688 13602 34700
rect 14369 34697 14381 34700
rect 14415 34697 14427 34731
rect 16942 34728 16948 34740
rect 16903 34700 16948 34728
rect 14369 34691 14427 34697
rect 16942 34688 16948 34700
rect 17000 34688 17006 34740
rect 17862 34728 17868 34740
rect 17823 34700 17868 34728
rect 17862 34688 17868 34700
rect 17920 34688 17926 34740
rect 18046 34728 18052 34740
rect 18007 34700 18052 34728
rect 18046 34688 18052 34700
rect 18104 34688 18110 34740
rect 20622 34728 20628 34740
rect 20583 34700 20628 34728
rect 20622 34688 20628 34700
rect 20680 34688 20686 34740
rect 20990 34728 20996 34740
rect 20951 34700 20996 34728
rect 20990 34688 20996 34700
rect 21048 34688 21054 34740
rect 22462 34728 22468 34740
rect 22423 34700 22468 34728
rect 22462 34688 22468 34700
rect 22520 34728 22526 34740
rect 23017 34731 23075 34737
rect 23017 34728 23029 34731
rect 22520 34700 23029 34728
rect 22520 34688 22526 34700
rect 23017 34697 23029 34700
rect 23063 34728 23075 34731
rect 23382 34728 23388 34740
rect 23063 34700 23388 34728
rect 23063 34697 23075 34700
rect 23017 34691 23075 34697
rect 23382 34688 23388 34700
rect 23440 34688 23446 34740
rect 25590 34728 25596 34740
rect 25551 34700 25596 34728
rect 25590 34688 25596 34700
rect 25648 34688 25654 34740
rect 28074 34728 28080 34740
rect 28035 34700 28080 34728
rect 28074 34688 28080 34700
rect 28132 34688 28138 34740
rect 35621 34731 35679 34737
rect 35621 34697 35633 34731
rect 35667 34728 35679 34731
rect 35802 34728 35808 34740
rect 35667 34700 35808 34728
rect 35667 34697 35679 34700
rect 35621 34691 35679 34697
rect 35802 34688 35808 34700
rect 35860 34688 35866 34740
rect 36722 34728 36728 34740
rect 36683 34700 36728 34728
rect 36722 34688 36728 34700
rect 36780 34688 36786 34740
rect 2682 34660 2688 34672
rect 2643 34632 2688 34660
rect 2682 34620 2688 34632
rect 2740 34620 2746 34672
rect 8205 34663 8263 34669
rect 8205 34629 8217 34663
rect 8251 34660 8263 34663
rect 8294 34660 8300 34672
rect 8251 34632 8300 34660
rect 8251 34629 8263 34632
rect 8205 34623 8263 34629
rect 8294 34620 8300 34632
rect 8352 34660 8358 34672
rect 17497 34663 17555 34669
rect 8352 34632 9260 34660
rect 8352 34620 8358 34632
rect 3789 34595 3847 34601
rect 3789 34561 3801 34595
rect 3835 34592 3847 34595
rect 4893 34595 4951 34601
rect 4893 34592 4905 34595
rect 3835 34564 4905 34592
rect 3835 34561 3847 34564
rect 3789 34555 3847 34561
rect 4893 34561 4905 34564
rect 4939 34592 4951 34595
rect 5074 34592 5080 34604
rect 4939 34564 5080 34592
rect 4939 34561 4951 34564
rect 4893 34555 4951 34561
rect 5074 34552 5080 34564
rect 5132 34552 5138 34604
rect 1397 34527 1455 34533
rect 1397 34493 1409 34527
rect 1443 34524 1455 34527
rect 2038 34524 2044 34536
rect 1443 34496 2044 34524
rect 1443 34493 1455 34496
rect 1397 34487 1455 34493
rect 2038 34484 2044 34496
rect 2096 34484 2102 34536
rect 2501 34527 2559 34533
rect 2501 34493 2513 34527
rect 2547 34524 2559 34527
rect 3142 34524 3148 34536
rect 2547 34496 3148 34524
rect 2547 34493 2559 34496
rect 2501 34487 2559 34493
rect 3142 34484 3148 34496
rect 3200 34484 3206 34536
rect 4157 34527 4215 34533
rect 4157 34493 4169 34527
rect 4203 34524 4215 34527
rect 4614 34524 4620 34536
rect 4203 34496 4620 34524
rect 4203 34493 4215 34496
rect 4157 34487 4215 34493
rect 4614 34484 4620 34496
rect 4672 34524 4678 34536
rect 4709 34527 4767 34533
rect 4709 34524 4721 34527
rect 4672 34496 4721 34524
rect 4672 34484 4678 34496
rect 4709 34493 4721 34496
rect 4755 34493 4767 34527
rect 4709 34487 4767 34493
rect 5626 34484 5632 34536
rect 5684 34524 5690 34536
rect 6825 34527 6883 34533
rect 6825 34524 6837 34527
rect 5684 34496 6837 34524
rect 5684 34484 5690 34496
rect 6825 34493 6837 34496
rect 6871 34524 6883 34527
rect 6914 34524 6920 34536
rect 6871 34496 6920 34524
rect 6871 34493 6883 34496
rect 6825 34487 6883 34493
rect 6914 34484 6920 34496
rect 6972 34524 6978 34536
rect 8202 34524 8208 34536
rect 6972 34496 8208 34524
rect 6972 34484 6978 34496
rect 8202 34484 8208 34496
rect 8260 34484 8266 34536
rect 9232 34533 9260 34632
rect 17497 34629 17509 34663
rect 17543 34660 17555 34663
rect 17543 34632 18644 34660
rect 17543 34629 17555 34632
rect 17497 34623 17555 34629
rect 12066 34552 12072 34604
rect 12124 34592 12130 34604
rect 12437 34595 12495 34601
rect 12437 34592 12449 34595
rect 12124 34564 12449 34592
rect 12124 34552 12130 34564
rect 12437 34561 12449 34564
rect 12483 34561 12495 34595
rect 12437 34555 12495 34561
rect 14642 34552 14648 34604
rect 14700 34592 14706 34604
rect 14700 34564 14964 34592
rect 14700 34552 14706 34564
rect 9217 34527 9275 34533
rect 9217 34493 9229 34527
rect 9263 34524 9275 34527
rect 9769 34527 9827 34533
rect 9263 34496 9628 34524
rect 9263 34493 9275 34496
rect 9217 34487 9275 34493
rect 7070 34459 7128 34465
rect 7070 34456 7082 34459
rect 6288 34428 7082 34456
rect 6288 34400 6316 34428
rect 7070 34425 7082 34428
rect 7116 34425 7128 34459
rect 7070 34419 7128 34425
rect 4617 34391 4675 34397
rect 4617 34357 4629 34391
rect 4663 34388 4675 34391
rect 4706 34388 4712 34400
rect 4663 34360 4712 34388
rect 4663 34357 4675 34360
rect 4617 34351 4675 34357
rect 4706 34348 4712 34360
rect 4764 34348 4770 34400
rect 6270 34388 6276 34400
rect 6231 34360 6276 34388
rect 6270 34348 6276 34360
rect 6328 34348 6334 34400
rect 9600 34388 9628 34496
rect 9769 34493 9781 34527
rect 9815 34524 9827 34527
rect 9858 34524 9864 34536
rect 9815 34496 9864 34524
rect 9815 34493 9827 34496
rect 9769 34487 9827 34493
rect 9858 34484 9864 34496
rect 9916 34484 9922 34536
rect 14090 34484 14096 34536
rect 14148 34524 14154 34536
rect 14737 34527 14795 34533
rect 14737 34524 14749 34527
rect 14148 34496 14749 34524
rect 14148 34484 14154 34496
rect 14737 34493 14749 34496
rect 14783 34524 14795 34527
rect 14826 34524 14832 34536
rect 14783 34496 14832 34524
rect 14783 34493 14795 34496
rect 14737 34487 14795 34493
rect 14826 34484 14832 34496
rect 14884 34484 14890 34536
rect 14936 34533 14964 34564
rect 17862 34552 17868 34604
rect 17920 34592 17926 34604
rect 18506 34592 18512 34604
rect 17920 34564 18512 34592
rect 17920 34552 17926 34564
rect 18506 34552 18512 34564
rect 18564 34552 18570 34604
rect 18616 34601 18644 34632
rect 18601 34595 18659 34601
rect 18601 34561 18613 34595
rect 18647 34592 18659 34595
rect 19242 34592 19248 34604
rect 18647 34564 19248 34592
rect 18647 34561 18659 34564
rect 18601 34555 18659 34561
rect 19242 34552 19248 34564
rect 19300 34552 19306 34604
rect 21008 34592 21036 34688
rect 21008 34564 21220 34592
rect 15194 34533 15200 34536
rect 14921 34527 14979 34533
rect 14921 34493 14933 34527
rect 14967 34524 14979 34527
rect 15188 34524 15200 34533
rect 14967 34496 15056 34524
rect 15155 34496 15200 34524
rect 14967 34493 14979 34496
rect 14921 34487 14979 34493
rect 9677 34459 9735 34465
rect 9677 34425 9689 34459
rect 9723 34456 9735 34459
rect 10014 34459 10072 34465
rect 10014 34456 10026 34459
rect 9723 34428 10026 34456
rect 9723 34425 9735 34428
rect 9677 34419 9735 34425
rect 10014 34425 10026 34428
rect 10060 34456 10072 34459
rect 10134 34456 10140 34468
rect 10060 34428 10140 34456
rect 10060 34425 10072 34428
rect 10014 34419 10072 34425
rect 10134 34416 10140 34428
rect 10192 34416 10198 34468
rect 12161 34459 12219 34465
rect 12161 34425 12173 34459
rect 12207 34456 12219 34459
rect 12526 34456 12532 34468
rect 12207 34428 12532 34456
rect 12207 34425 12219 34428
rect 12161 34419 12219 34425
rect 12526 34416 12532 34428
rect 12584 34456 12590 34468
rect 12704 34459 12762 34465
rect 12704 34456 12716 34459
rect 12584 34428 12716 34456
rect 12584 34416 12590 34428
rect 12704 34425 12716 34428
rect 12750 34456 12762 34459
rect 13538 34456 13544 34468
rect 12750 34428 13544 34456
rect 12750 34425 12762 34428
rect 12704 34419 12762 34425
rect 13538 34416 13544 34428
rect 13596 34416 13602 34468
rect 15028 34456 15056 34496
rect 15188 34487 15200 34496
rect 15194 34484 15200 34487
rect 15252 34484 15258 34536
rect 17954 34484 17960 34536
rect 18012 34524 18018 34536
rect 18417 34527 18475 34533
rect 18417 34524 18429 34527
rect 18012 34496 18429 34524
rect 18012 34484 18018 34496
rect 18417 34493 18429 34496
rect 18463 34493 18475 34527
rect 18417 34487 18475 34493
rect 19981 34527 20039 34533
rect 19981 34493 19993 34527
rect 20027 34524 20039 34527
rect 20622 34524 20628 34536
rect 20027 34496 20628 34524
rect 20027 34493 20039 34496
rect 19981 34487 20039 34493
rect 20622 34484 20628 34496
rect 20680 34484 20686 34536
rect 21082 34524 21088 34536
rect 21043 34496 21088 34524
rect 21082 34484 21088 34496
rect 21140 34484 21146 34536
rect 21192 34524 21220 34564
rect 22922 34552 22928 34604
rect 22980 34592 22986 34604
rect 24210 34592 24216 34604
rect 22980 34564 24216 34592
rect 22980 34552 22986 34564
rect 24210 34552 24216 34564
rect 24268 34552 24274 34604
rect 26694 34592 26700 34604
rect 26655 34564 26700 34592
rect 26694 34552 26700 34564
rect 26752 34552 26758 34604
rect 26970 34533 26976 34536
rect 21341 34527 21399 34533
rect 21341 34524 21353 34527
rect 21192 34496 21353 34524
rect 21341 34493 21353 34496
rect 21387 34524 21399 34527
rect 26964 34524 26976 34533
rect 21387 34496 22232 34524
rect 21387 34493 21399 34496
rect 21341 34487 21399 34493
rect 22204 34468 22232 34496
rect 26804 34496 26976 34524
rect 15286 34456 15292 34468
rect 15028 34428 15292 34456
rect 15286 34416 15292 34428
rect 15344 34416 15350 34468
rect 22186 34416 22192 34468
rect 22244 34416 22250 34468
rect 24458 34459 24516 34465
rect 24458 34456 24470 34459
rect 24044 34428 24470 34456
rect 24044 34400 24072 34428
rect 24458 34425 24470 34428
rect 24504 34425 24516 34459
rect 26602 34456 26608 34468
rect 26515 34428 26608 34456
rect 24458 34419 24516 34425
rect 26602 34416 26608 34428
rect 26660 34456 26666 34468
rect 26804 34456 26832 34496
rect 26964 34487 26976 34496
rect 26970 34484 26976 34487
rect 27028 34484 27034 34536
rect 35250 34524 35256 34536
rect 35211 34496 35256 34524
rect 35250 34484 35256 34496
rect 35308 34524 35314 34536
rect 35437 34527 35495 34533
rect 35437 34524 35449 34527
rect 35308 34496 35449 34524
rect 35308 34484 35314 34496
rect 35437 34493 35449 34496
rect 35483 34493 35495 34527
rect 35437 34487 35495 34493
rect 36541 34527 36599 34533
rect 36541 34493 36553 34527
rect 36587 34524 36599 34527
rect 37090 34524 37096 34536
rect 36587 34496 37096 34524
rect 36587 34493 36599 34496
rect 36541 34487 36599 34493
rect 37090 34484 37096 34496
rect 37148 34484 37154 34536
rect 26660 34428 26832 34456
rect 26660 34416 26666 34428
rect 9766 34388 9772 34400
rect 9600 34360 9772 34388
rect 9766 34348 9772 34360
rect 9824 34348 9830 34400
rect 11146 34388 11152 34400
rect 11107 34360 11152 34388
rect 11146 34348 11152 34360
rect 11204 34348 11210 34400
rect 13262 34348 13268 34400
rect 13320 34388 13326 34400
rect 13817 34391 13875 34397
rect 13817 34388 13829 34391
rect 13320 34360 13829 34388
rect 13320 34348 13326 34360
rect 13817 34357 13829 34360
rect 13863 34357 13875 34391
rect 13817 34351 13875 34357
rect 14918 34348 14924 34400
rect 14976 34388 14982 34400
rect 16301 34391 16359 34397
rect 16301 34388 16313 34391
rect 14976 34360 16313 34388
rect 14976 34348 14982 34360
rect 16301 34357 16313 34360
rect 16347 34357 16359 34391
rect 20162 34388 20168 34400
rect 20123 34360 20168 34388
rect 16301 34351 16359 34357
rect 20162 34348 20168 34360
rect 20220 34348 20226 34400
rect 24026 34388 24032 34400
rect 23987 34360 24032 34388
rect 24026 34348 24032 34360
rect 24084 34348 24090 34400
rect 28350 34348 28356 34400
rect 28408 34388 28414 34400
rect 28629 34391 28687 34397
rect 28629 34388 28641 34391
rect 28408 34360 28641 34388
rect 28408 34348 28414 34360
rect 28629 34357 28641 34360
rect 28675 34357 28687 34391
rect 28629 34351 28687 34357
rect 30098 34348 30104 34400
rect 30156 34388 30162 34400
rect 35342 34388 35348 34400
rect 30156 34360 35348 34388
rect 30156 34348 30162 34360
rect 35342 34348 35348 34360
rect 35400 34388 35406 34400
rect 35989 34391 36047 34397
rect 35989 34388 36001 34391
rect 35400 34360 36001 34388
rect 35400 34348 35406 34360
rect 35989 34357 36001 34360
rect 36035 34357 36047 34391
rect 35989 34351 36047 34357
rect 1104 34298 38824 34320
rect 1104 34246 19606 34298
rect 19658 34246 19670 34298
rect 19722 34246 19734 34298
rect 19786 34246 19798 34298
rect 19850 34246 38824 34298
rect 1104 34224 38824 34246
rect 1394 34144 1400 34196
rect 1452 34184 1458 34196
rect 1581 34187 1639 34193
rect 1581 34184 1593 34187
rect 1452 34156 1593 34184
rect 1452 34144 1458 34156
rect 1581 34153 1593 34156
rect 1627 34153 1639 34187
rect 1581 34147 1639 34153
rect 4154 34144 4160 34196
rect 4212 34184 4218 34196
rect 4249 34187 4307 34193
rect 4249 34184 4261 34187
rect 4212 34156 4261 34184
rect 4212 34144 4218 34156
rect 4249 34153 4261 34156
rect 4295 34153 4307 34187
rect 4249 34147 4307 34153
rect 6270 34144 6276 34196
rect 6328 34184 6334 34196
rect 6641 34187 6699 34193
rect 6641 34184 6653 34187
rect 6328 34156 6653 34184
rect 6328 34144 6334 34156
rect 6641 34153 6653 34156
rect 6687 34184 6699 34187
rect 7190 34184 7196 34196
rect 6687 34156 7196 34184
rect 6687 34153 6699 34156
rect 6641 34147 6699 34153
rect 7190 34144 7196 34156
rect 7248 34144 7254 34196
rect 9125 34187 9183 34193
rect 9125 34153 9137 34187
rect 9171 34184 9183 34187
rect 11057 34187 11115 34193
rect 11057 34184 11069 34187
rect 9171 34156 11069 34184
rect 9171 34153 9183 34156
rect 9125 34147 9183 34153
rect 11057 34153 11069 34156
rect 11103 34153 11115 34187
rect 11057 34147 11115 34153
rect 4709 34119 4767 34125
rect 4709 34085 4721 34119
rect 4755 34116 4767 34119
rect 4982 34116 4988 34128
rect 4755 34088 4988 34116
rect 4755 34085 4767 34088
rect 4709 34079 4767 34085
rect 4982 34076 4988 34088
rect 5040 34116 5046 34128
rect 6822 34116 6828 34128
rect 5040 34088 6828 34116
rect 5040 34076 5046 34088
rect 6822 34076 6828 34088
rect 6880 34076 6886 34128
rect 4062 34048 4068 34060
rect 4023 34020 4068 34048
rect 4062 34008 4068 34020
rect 4120 34008 4126 34060
rect 5534 34057 5540 34060
rect 5528 34011 5540 34057
rect 5592 34048 5598 34060
rect 5592 34020 5628 34048
rect 5534 34008 5540 34011
rect 5592 34008 5598 34020
rect 7926 34008 7932 34060
rect 7984 34048 7990 34060
rect 8389 34051 8447 34057
rect 8389 34048 8401 34051
rect 7984 34020 8401 34048
rect 7984 34008 7990 34020
rect 8389 34017 8401 34020
rect 8435 34017 8447 34051
rect 8389 34011 8447 34017
rect 8481 34051 8539 34057
rect 8481 34017 8493 34051
rect 8527 34048 8539 34051
rect 8662 34048 8668 34060
rect 8527 34020 8668 34048
rect 8527 34017 8539 34020
rect 8481 34011 8539 34017
rect 8662 34008 8668 34020
rect 8720 34008 8726 34060
rect 3970 33940 3976 33992
rect 4028 33980 4034 33992
rect 5261 33983 5319 33989
rect 5261 33980 5273 33983
rect 4028 33952 5273 33980
rect 4028 33940 4034 33952
rect 5261 33949 5273 33952
rect 5307 33949 5319 33983
rect 5261 33943 5319 33949
rect 8573 33983 8631 33989
rect 8573 33949 8585 33983
rect 8619 33980 8631 33983
rect 9030 33980 9036 33992
rect 8619 33952 9036 33980
rect 8619 33949 8631 33952
rect 8573 33943 8631 33949
rect 9030 33940 9036 33952
rect 9088 33980 9094 33992
rect 9140 33980 9168 34147
rect 11330 34144 11336 34196
rect 11388 34184 11394 34196
rect 11609 34187 11667 34193
rect 11609 34184 11621 34187
rect 11388 34156 11621 34184
rect 11388 34144 11394 34156
rect 11609 34153 11621 34156
rect 11655 34153 11667 34187
rect 13538 34184 13544 34196
rect 13499 34156 13544 34184
rect 11609 34147 11667 34153
rect 13538 34144 13544 34156
rect 13596 34144 13602 34196
rect 13814 34144 13820 34196
rect 13872 34184 13878 34196
rect 14093 34187 14151 34193
rect 14093 34184 14105 34187
rect 13872 34156 14105 34184
rect 13872 34144 13878 34156
rect 14093 34153 14105 34156
rect 14139 34153 14151 34187
rect 14093 34147 14151 34153
rect 16209 34187 16267 34193
rect 16209 34153 16221 34187
rect 16255 34184 16267 34187
rect 16482 34184 16488 34196
rect 16255 34156 16488 34184
rect 16255 34153 16267 34156
rect 16209 34147 16267 34153
rect 16482 34144 16488 34156
rect 16540 34144 16546 34196
rect 22186 34144 22192 34196
rect 22244 34184 22250 34196
rect 22281 34187 22339 34193
rect 22281 34184 22293 34187
rect 22244 34156 22293 34184
rect 22244 34144 22250 34156
rect 22281 34153 22293 34156
rect 22327 34153 22339 34187
rect 22922 34184 22928 34196
rect 22883 34156 22928 34184
rect 22281 34147 22339 34153
rect 22922 34144 22928 34156
rect 22980 34144 22986 34196
rect 23474 34144 23480 34196
rect 23532 34184 23538 34196
rect 23845 34187 23903 34193
rect 23845 34184 23857 34187
rect 23532 34156 23857 34184
rect 23532 34144 23538 34156
rect 23845 34153 23857 34156
rect 23891 34153 23903 34187
rect 23845 34147 23903 34153
rect 27525 34187 27583 34193
rect 27525 34153 27537 34187
rect 27571 34184 27583 34187
rect 28074 34184 28080 34196
rect 27571 34156 28080 34184
rect 27571 34153 27583 34156
rect 27525 34147 27583 34153
rect 28074 34144 28080 34156
rect 28132 34144 28138 34196
rect 35618 34184 35624 34196
rect 35579 34156 35624 34184
rect 35618 34144 35624 34156
rect 35676 34144 35682 34196
rect 9858 34116 9864 34128
rect 9692 34088 9864 34116
rect 9692 33989 9720 34088
rect 9858 34076 9864 34088
rect 9916 34076 9922 34128
rect 12158 34076 12164 34128
rect 12216 34116 12222 34128
rect 12406 34119 12464 34125
rect 12406 34116 12418 34119
rect 12216 34088 12418 34116
rect 12216 34076 12222 34088
rect 12406 34085 12418 34088
rect 12452 34085 12464 34119
rect 17672 34119 17730 34125
rect 17672 34116 17684 34119
rect 12406 34079 12464 34085
rect 16776 34088 17684 34116
rect 9766 34008 9772 34060
rect 9824 34048 9830 34060
rect 9944 34051 10002 34057
rect 9944 34048 9956 34051
rect 9824 34020 9956 34048
rect 9824 34008 9830 34020
rect 9944 34017 9956 34020
rect 9990 34048 10002 34051
rect 10686 34048 10692 34060
rect 9990 34020 10692 34048
rect 9990 34017 10002 34020
rect 9944 34011 10002 34017
rect 10686 34008 10692 34020
rect 10744 34008 10750 34060
rect 14458 34008 14464 34060
rect 14516 34048 14522 34060
rect 14829 34051 14887 34057
rect 14829 34048 14841 34051
rect 14516 34020 14841 34048
rect 14516 34008 14522 34020
rect 14829 34017 14841 34020
rect 14875 34017 14887 34051
rect 14829 34011 14887 34017
rect 9677 33983 9735 33989
rect 9677 33980 9689 33983
rect 9088 33952 9168 33980
rect 9416 33952 9689 33980
rect 9088 33940 9094 33952
rect 7466 33872 7472 33924
rect 7524 33912 7530 33924
rect 7561 33915 7619 33921
rect 7561 33912 7573 33915
rect 7524 33884 7573 33912
rect 7524 33872 7530 33884
rect 7561 33881 7573 33884
rect 7607 33881 7619 33915
rect 7561 33875 7619 33881
rect 5077 33847 5135 33853
rect 5077 33813 5089 33847
rect 5123 33844 5135 33847
rect 5258 33844 5264 33856
rect 5123 33816 5264 33844
rect 5123 33813 5135 33816
rect 5077 33807 5135 33813
rect 5258 33804 5264 33816
rect 5316 33804 5322 33856
rect 8018 33844 8024 33856
rect 7979 33816 8024 33844
rect 8018 33804 8024 33816
rect 8076 33804 8082 33856
rect 8294 33804 8300 33856
rect 8352 33844 8358 33856
rect 9416 33853 9444 33952
rect 9677 33949 9689 33952
rect 9723 33949 9735 33983
rect 9677 33943 9735 33949
rect 11790 33940 11796 33992
rect 11848 33980 11854 33992
rect 12161 33983 12219 33989
rect 12161 33980 12173 33983
rect 11848 33952 12173 33980
rect 11848 33940 11854 33952
rect 12161 33949 12173 33952
rect 12207 33949 12219 33983
rect 12161 33943 12219 33949
rect 15194 33940 15200 33992
rect 15252 33980 15258 33992
rect 16301 33983 16359 33989
rect 16301 33980 16313 33983
rect 15252 33952 16313 33980
rect 15252 33940 15258 33952
rect 16301 33949 16313 33952
rect 16347 33949 16359 33983
rect 16301 33943 16359 33949
rect 16485 33983 16543 33989
rect 16485 33949 16497 33983
rect 16531 33980 16543 33983
rect 16776 33980 16804 34088
rect 17672 34085 17684 34088
rect 17718 34116 17730 34119
rect 17770 34116 17776 34128
rect 17718 34088 17776 34116
rect 17718 34085 17730 34088
rect 17672 34079 17730 34085
rect 17770 34076 17776 34088
rect 17828 34076 17834 34128
rect 21082 34116 21088 34128
rect 20916 34088 21088 34116
rect 16945 34051 17003 34057
rect 16945 34017 16957 34051
rect 16991 34048 17003 34051
rect 17313 34051 17371 34057
rect 17313 34048 17325 34051
rect 16991 34020 17325 34048
rect 16991 34017 17003 34020
rect 16945 34011 17003 34017
rect 17313 34017 17325 34020
rect 17359 34048 17371 34051
rect 17405 34051 17463 34057
rect 17405 34048 17417 34051
rect 17359 34020 17417 34048
rect 17359 34017 17371 34020
rect 17313 34011 17371 34017
rect 17405 34017 17417 34020
rect 17451 34048 17463 34051
rect 18046 34048 18052 34060
rect 17451 34020 18052 34048
rect 17451 34017 17463 34020
rect 17405 34011 17463 34017
rect 18046 34008 18052 34020
rect 18104 34008 18110 34060
rect 20714 34008 20720 34060
rect 20772 34048 20778 34060
rect 20916 34057 20944 34088
rect 21082 34076 21088 34088
rect 21140 34076 21146 34128
rect 28160 34119 28218 34125
rect 28160 34085 28172 34119
rect 28206 34116 28218 34119
rect 28810 34116 28816 34128
rect 28206 34088 28816 34116
rect 28206 34085 28218 34088
rect 28160 34079 28218 34085
rect 28810 34076 28816 34088
rect 28868 34076 28874 34128
rect 21174 34057 21180 34060
rect 20901 34051 20959 34057
rect 20901 34048 20913 34051
rect 20772 34020 20913 34048
rect 20772 34008 20778 34020
rect 20901 34017 20913 34020
rect 20947 34017 20959 34051
rect 21168 34048 21180 34057
rect 21135 34020 21180 34048
rect 20901 34011 20959 34017
rect 21168 34011 21180 34020
rect 21174 34008 21180 34011
rect 21232 34008 21238 34060
rect 23106 34008 23112 34060
rect 23164 34048 23170 34060
rect 23753 34051 23811 34057
rect 23753 34048 23765 34051
rect 23164 34020 23765 34048
rect 23164 34008 23170 34020
rect 23753 34017 23765 34020
rect 23799 34048 23811 34051
rect 24026 34048 24032 34060
rect 23799 34020 24032 34048
rect 23799 34017 23811 34020
rect 23753 34011 23811 34017
rect 24026 34008 24032 34020
rect 24084 34008 24090 34060
rect 25314 34048 25320 34060
rect 25275 34020 25320 34048
rect 25314 34008 25320 34020
rect 25372 34008 25378 34060
rect 25958 34008 25964 34060
rect 26016 34048 26022 34060
rect 26513 34051 26571 34057
rect 26513 34048 26525 34051
rect 26016 34020 26525 34048
rect 26016 34008 26022 34020
rect 26513 34017 26525 34020
rect 26559 34048 26571 34051
rect 27065 34051 27123 34057
rect 27065 34048 27077 34051
rect 26559 34020 27077 34048
rect 26559 34017 26571 34020
rect 26513 34011 26571 34017
rect 27065 34017 27077 34020
rect 27111 34017 27123 34051
rect 27065 34011 27123 34017
rect 27893 34051 27951 34057
rect 27893 34017 27905 34051
rect 27939 34048 27951 34051
rect 28442 34048 28448 34060
rect 27939 34020 28448 34048
rect 27939 34017 27951 34020
rect 27893 34011 27951 34017
rect 28442 34008 28448 34020
rect 28500 34008 28506 34060
rect 35437 34051 35495 34057
rect 35437 34017 35449 34051
rect 35483 34048 35495 34051
rect 35894 34048 35900 34060
rect 35483 34020 35900 34048
rect 35483 34017 35495 34020
rect 35437 34011 35495 34017
rect 35894 34008 35900 34020
rect 35952 34008 35958 34060
rect 16531 33952 16804 33980
rect 16531 33949 16543 33952
rect 16485 33943 16543 33949
rect 22094 33940 22100 33992
rect 22152 33980 22158 33992
rect 23937 33983 23995 33989
rect 23937 33980 23949 33983
rect 22152 33952 23949 33980
rect 22152 33940 22158 33952
rect 23937 33949 23949 33952
rect 23983 33980 23995 33983
rect 25869 33983 25927 33989
rect 25869 33980 25881 33983
rect 23983 33952 25881 33980
rect 23983 33949 23995 33952
rect 23937 33943 23995 33949
rect 25869 33949 25881 33952
rect 25915 33980 25927 33983
rect 26418 33980 26424 33992
rect 25915 33952 26424 33980
rect 25915 33949 25927 33952
rect 25869 33943 25927 33949
rect 26418 33940 26424 33952
rect 26476 33940 26482 33992
rect 15838 33912 15844 33924
rect 15799 33884 15844 33912
rect 15838 33872 15844 33884
rect 15896 33872 15902 33924
rect 25774 33872 25780 33924
rect 25832 33912 25838 33924
rect 26697 33915 26755 33921
rect 26697 33912 26709 33915
rect 25832 33884 26709 33912
rect 25832 33872 25838 33884
rect 26697 33881 26709 33884
rect 26743 33881 26755 33915
rect 26697 33875 26755 33881
rect 9401 33847 9459 33853
rect 9401 33844 9413 33847
rect 8352 33816 9413 33844
rect 8352 33804 8358 33816
rect 9401 33813 9413 33816
rect 9447 33813 9459 33847
rect 14458 33844 14464 33856
rect 14419 33816 14464 33844
rect 9401 33807 9459 33813
rect 14458 33804 14464 33816
rect 14516 33804 14522 33856
rect 14645 33847 14703 33853
rect 14645 33813 14657 33847
rect 14691 33844 14703 33847
rect 14826 33844 14832 33856
rect 14691 33816 14832 33844
rect 14691 33813 14703 33816
rect 14645 33807 14703 33813
rect 14826 33804 14832 33816
rect 14884 33804 14890 33856
rect 15470 33844 15476 33856
rect 15431 33816 15476 33844
rect 15470 33804 15476 33816
rect 15528 33804 15534 33856
rect 18782 33844 18788 33856
rect 18743 33816 18788 33844
rect 18782 33804 18788 33816
rect 18840 33804 18846 33856
rect 23382 33844 23388 33856
rect 23343 33816 23388 33844
rect 23382 33804 23388 33816
rect 23440 33804 23446 33856
rect 24394 33844 24400 33856
rect 24355 33816 24400 33844
rect 24394 33804 24400 33816
rect 24452 33804 24458 33856
rect 25498 33844 25504 33856
rect 25459 33816 25504 33844
rect 25498 33804 25504 33816
rect 25556 33804 25562 33856
rect 29086 33804 29092 33856
rect 29144 33844 29150 33856
rect 29273 33847 29331 33853
rect 29273 33844 29285 33847
rect 29144 33816 29285 33844
rect 29144 33804 29150 33816
rect 29273 33813 29285 33816
rect 29319 33813 29331 33847
rect 29273 33807 29331 33813
rect 1104 33754 38824 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 34966 33754
rect 35018 33702 35030 33754
rect 35082 33702 35094 33754
rect 35146 33702 35158 33754
rect 35210 33702 38824 33754
rect 1104 33680 38824 33702
rect 4062 33640 4068 33652
rect 4023 33612 4068 33640
rect 4062 33600 4068 33612
rect 4120 33600 4126 33652
rect 5534 33600 5540 33652
rect 5592 33640 5598 33652
rect 5629 33643 5687 33649
rect 5629 33640 5641 33643
rect 5592 33612 5641 33640
rect 5592 33600 5598 33612
rect 5629 33609 5641 33612
rect 5675 33640 5687 33643
rect 6181 33643 6239 33649
rect 6181 33640 6193 33643
rect 5675 33612 6193 33640
rect 5675 33609 5687 33612
rect 5629 33603 5687 33609
rect 6181 33609 6193 33612
rect 6227 33640 6239 33643
rect 6549 33643 6607 33649
rect 6549 33640 6561 33643
rect 6227 33612 6561 33640
rect 6227 33609 6239 33612
rect 6181 33603 6239 33609
rect 6549 33609 6561 33612
rect 6595 33609 6607 33643
rect 6822 33640 6828 33652
rect 6783 33612 6828 33640
rect 6549 33603 6607 33609
rect 3421 33507 3479 33513
rect 3421 33473 3433 33507
rect 3467 33504 3479 33507
rect 4062 33504 4068 33516
rect 3467 33476 4068 33504
rect 3467 33473 3479 33476
rect 3421 33467 3479 33473
rect 4062 33464 4068 33476
rect 4120 33504 4126 33516
rect 4249 33507 4307 33513
rect 4249 33504 4261 33507
rect 4120 33476 4261 33504
rect 4120 33464 4126 33476
rect 4249 33473 4261 33476
rect 4295 33473 4307 33507
rect 4249 33467 4307 33473
rect 4264 33436 4292 33467
rect 5534 33436 5540 33448
rect 4264 33408 5540 33436
rect 5534 33396 5540 33408
rect 5592 33396 5598 33448
rect 4522 33377 4528 33380
rect 3789 33371 3847 33377
rect 3789 33337 3801 33371
rect 3835 33368 3847 33371
rect 4516 33368 4528 33377
rect 3835 33340 4528 33368
rect 3835 33337 3847 33340
rect 3789 33331 3847 33337
rect 4516 33331 4528 33340
rect 4580 33368 4586 33380
rect 4706 33368 4712 33380
rect 4580 33340 4712 33368
rect 4522 33328 4528 33331
rect 4580 33328 4586 33340
rect 4706 33328 4712 33340
rect 4764 33328 4770 33380
rect 6564 33368 6592 33603
rect 6822 33600 6828 33612
rect 6880 33600 6886 33652
rect 8294 33600 8300 33652
rect 8352 33640 8358 33652
rect 8481 33643 8539 33649
rect 8481 33640 8493 33643
rect 8352 33612 8493 33640
rect 8352 33600 8358 33612
rect 8481 33609 8493 33612
rect 8527 33609 8539 33643
rect 10134 33640 10140 33652
rect 10095 33612 10140 33640
rect 8481 33603 8539 33609
rect 7466 33504 7472 33516
rect 7427 33476 7472 33504
rect 7466 33464 7472 33476
rect 7524 33464 7530 33516
rect 8496 33504 8524 33603
rect 10134 33600 10140 33612
rect 10192 33600 10198 33652
rect 10686 33640 10692 33652
rect 10647 33612 10692 33640
rect 10686 33600 10692 33612
rect 10744 33600 10750 33652
rect 11146 33600 11152 33652
rect 11204 33640 11210 33652
rect 12158 33640 12164 33652
rect 11204 33612 12164 33640
rect 11204 33600 11210 33612
rect 12158 33600 12164 33612
rect 12216 33600 12222 33652
rect 14366 33640 14372 33652
rect 14327 33612 14372 33640
rect 14366 33600 14372 33612
rect 14424 33600 14430 33652
rect 14918 33640 14924 33652
rect 14879 33612 14924 33640
rect 14918 33600 14924 33612
rect 14976 33600 14982 33652
rect 15381 33643 15439 33649
rect 15381 33609 15393 33643
rect 15427 33640 15439 33643
rect 16482 33640 16488 33652
rect 15427 33612 16488 33640
rect 15427 33609 15439 33612
rect 15381 33603 15439 33609
rect 16482 33600 16488 33612
rect 16540 33600 16546 33652
rect 19334 33600 19340 33652
rect 19392 33640 19398 33652
rect 19429 33643 19487 33649
rect 19429 33640 19441 33643
rect 19392 33612 19441 33640
rect 19392 33600 19398 33612
rect 19429 33609 19441 33612
rect 19475 33609 19487 33643
rect 19429 33603 19487 33609
rect 21358 33600 21364 33652
rect 21416 33640 21422 33652
rect 22097 33643 22155 33649
rect 22097 33640 22109 33643
rect 21416 33612 22109 33640
rect 21416 33600 21422 33612
rect 22097 33609 22109 33612
rect 22143 33609 22155 33643
rect 23106 33640 23112 33652
rect 23067 33612 23112 33640
rect 22097 33603 22155 33609
rect 23106 33600 23112 33612
rect 23164 33600 23170 33652
rect 23474 33640 23480 33652
rect 23435 33612 23480 33640
rect 23474 33600 23480 33612
rect 23532 33600 23538 33652
rect 23658 33640 23664 33652
rect 23619 33612 23664 33640
rect 23658 33600 23664 33612
rect 23716 33600 23722 33652
rect 25590 33600 25596 33652
rect 25648 33640 25654 33652
rect 25685 33643 25743 33649
rect 25685 33640 25697 33643
rect 25648 33612 25697 33640
rect 25648 33600 25654 33612
rect 25685 33609 25697 33612
rect 25731 33640 25743 33643
rect 28537 33643 28595 33649
rect 25731 33612 26372 33640
rect 25731 33609 25743 33612
rect 25685 33603 25743 33609
rect 9858 33532 9864 33584
rect 9916 33572 9922 33584
rect 11057 33575 11115 33581
rect 11057 33572 11069 33575
rect 9916 33544 11069 33572
rect 9916 33532 9922 33544
rect 11057 33541 11069 33544
rect 11103 33572 11115 33575
rect 11790 33572 11796 33584
rect 11103 33544 11796 33572
rect 11103 33541 11115 33544
rect 11057 33535 11115 33541
rect 11790 33532 11796 33544
rect 11848 33532 11854 33584
rect 8570 33504 8576 33516
rect 8483 33476 8576 33504
rect 8570 33464 8576 33476
rect 8628 33504 8634 33516
rect 8757 33507 8815 33513
rect 8757 33504 8769 33507
rect 8628 33476 8769 33504
rect 8628 33464 8634 33476
rect 8757 33473 8769 33476
rect 8803 33473 8815 33507
rect 11238 33504 11244 33516
rect 11199 33476 11244 33504
rect 8757 33467 8815 33473
rect 11238 33464 11244 33476
rect 11296 33464 11302 33516
rect 14936 33504 14964 33600
rect 21910 33532 21916 33584
rect 21968 33572 21974 33584
rect 22649 33575 22707 33581
rect 22649 33572 22661 33575
rect 21968 33544 22661 33572
rect 21968 33532 21974 33544
rect 22112 33516 22140 33544
rect 22649 33541 22661 33544
rect 22695 33541 22707 33575
rect 24673 33575 24731 33581
rect 24673 33572 24685 33575
rect 22649 33535 22707 33541
rect 24136 33544 24685 33572
rect 24136 33516 24164 33544
rect 24673 33541 24685 33544
rect 24719 33541 24731 33575
rect 24673 33535 24731 33541
rect 25869 33575 25927 33581
rect 25869 33541 25881 33575
rect 25915 33572 25927 33575
rect 26234 33572 26240 33584
rect 25915 33544 26240 33572
rect 25915 33541 25927 33544
rect 25869 33535 25927 33541
rect 26234 33532 26240 33544
rect 26292 33532 26298 33584
rect 20257 33507 20315 33513
rect 14936 33476 15608 33504
rect 7190 33436 7196 33448
rect 7151 33408 7196 33436
rect 7190 33396 7196 33408
rect 7248 33396 7254 33448
rect 8665 33439 8723 33445
rect 8665 33405 8677 33439
rect 8711 33436 8723 33439
rect 8846 33436 8852 33448
rect 8711 33408 8852 33436
rect 8711 33405 8723 33408
rect 8665 33399 8723 33405
rect 8846 33396 8852 33408
rect 8904 33396 8910 33448
rect 9030 33445 9036 33448
rect 9024 33436 9036 33445
rect 8991 33408 9036 33436
rect 9024 33399 9036 33408
rect 9030 33396 9036 33399
rect 9088 33396 9094 33448
rect 12986 33436 12992 33448
rect 12947 33408 12992 33436
rect 12986 33396 12992 33408
rect 13044 33396 13050 33448
rect 13262 33445 13268 33448
rect 13256 33436 13268 33445
rect 13188 33408 13268 33436
rect 7285 33371 7343 33377
rect 7285 33368 7297 33371
rect 6564 33340 7297 33368
rect 7285 33337 7297 33340
rect 7331 33337 7343 33371
rect 7285 33331 7343 33337
rect 12897 33371 12955 33377
rect 12897 33337 12909 33371
rect 12943 33368 12955 33371
rect 13188 33368 13216 33408
rect 13256 33399 13268 33408
rect 13262 33396 13268 33399
rect 13320 33396 13326 33448
rect 15286 33396 15292 33448
rect 15344 33436 15350 33448
rect 15473 33439 15531 33445
rect 15473 33436 15485 33439
rect 15344 33408 15485 33436
rect 15344 33396 15350 33408
rect 15473 33405 15485 33408
rect 15519 33405 15531 33439
rect 15580 33436 15608 33476
rect 20257 33473 20269 33507
rect 20303 33504 20315 33507
rect 20714 33504 20720 33516
rect 20303 33476 20720 33504
rect 20303 33473 20315 33476
rect 20257 33467 20315 33473
rect 20714 33464 20720 33476
rect 20772 33464 20778 33516
rect 22094 33464 22100 33516
rect 22152 33464 22158 33516
rect 24118 33504 24124 33516
rect 24079 33476 24124 33504
rect 24118 33464 24124 33476
rect 24176 33464 24182 33516
rect 24213 33507 24271 33513
rect 24213 33473 24225 33507
rect 24259 33504 24271 33507
rect 24394 33504 24400 33516
rect 24259 33476 24400 33504
rect 24259 33473 24271 33476
rect 24213 33467 24271 33473
rect 24394 33464 24400 33476
rect 24452 33464 24458 33516
rect 26344 33513 26372 33612
rect 28537 33609 28549 33643
rect 28583 33640 28595 33643
rect 28810 33640 28816 33652
rect 28583 33612 28816 33640
rect 28583 33609 28595 33612
rect 28537 33603 28595 33609
rect 26329 33507 26387 33513
rect 26329 33473 26341 33507
rect 26375 33473 26387 33507
rect 26329 33467 26387 33473
rect 26418 33464 26424 33516
rect 26476 33504 26482 33516
rect 27614 33504 27620 33516
rect 26476 33476 27620 33504
rect 26476 33464 26482 33476
rect 27614 33464 27620 33476
rect 27672 33504 27678 33516
rect 27985 33507 28043 33513
rect 27985 33504 27997 33507
rect 27672 33476 27997 33504
rect 27672 33464 27678 33476
rect 27985 33473 27997 33476
rect 28031 33473 28043 33507
rect 27985 33467 28043 33473
rect 15729 33439 15787 33445
rect 15729 33436 15741 33439
rect 15580 33408 15741 33436
rect 15473 33399 15531 33405
rect 15729 33405 15741 33408
rect 15775 33405 15787 33439
rect 18046 33436 18052 33448
rect 15729 33399 15787 33405
rect 15856 33408 18052 33436
rect 12943 33340 13216 33368
rect 15488 33368 15516 33399
rect 15856 33368 15884 33408
rect 18046 33396 18052 33408
rect 18104 33396 18110 33448
rect 18316 33439 18374 33445
rect 18316 33436 18328 33439
rect 18156 33408 18328 33436
rect 15488 33340 15884 33368
rect 12943 33337 12955 33340
rect 12897 33331 12955 33337
rect 17954 33328 17960 33380
rect 18012 33368 18018 33380
rect 18156 33368 18184 33408
rect 18316 33405 18328 33408
rect 18362 33436 18374 33439
rect 18782 33436 18788 33448
rect 18362 33408 18788 33436
rect 18362 33405 18374 33408
rect 18316 33399 18374 33405
rect 18782 33396 18788 33408
rect 18840 33396 18846 33448
rect 23382 33396 23388 33448
rect 23440 33436 23446 33448
rect 24029 33439 24087 33445
rect 24029 33436 24041 33439
rect 23440 33408 24041 33436
rect 23440 33396 23446 33408
rect 24029 33405 24041 33408
rect 24075 33436 24087 33439
rect 24302 33436 24308 33448
rect 24075 33408 24308 33436
rect 24075 33405 24087 33408
rect 24029 33399 24087 33405
rect 24302 33396 24308 33408
rect 24360 33396 24366 33448
rect 18012 33340 18184 33368
rect 20625 33371 20683 33377
rect 18012 33328 18018 33340
rect 20625 33337 20637 33371
rect 20671 33368 20683 33371
rect 20962 33371 21020 33377
rect 20962 33368 20974 33371
rect 20671 33340 20974 33368
rect 20671 33337 20683 33340
rect 20625 33331 20683 33337
rect 20962 33337 20974 33340
rect 21008 33368 21020 33371
rect 21726 33368 21732 33380
rect 21008 33340 21732 33368
rect 21008 33337 21020 33340
rect 20962 33331 21020 33337
rect 21726 33328 21732 33340
rect 21784 33328 21790 33380
rect 23566 33328 23572 33380
rect 23624 33368 23630 33380
rect 24412 33368 24440 33464
rect 25866 33396 25872 33448
rect 25924 33436 25930 33448
rect 26237 33439 26295 33445
rect 26237 33436 26249 33439
rect 25924 33408 26249 33436
rect 25924 33396 25930 33408
rect 26237 33405 26249 33408
rect 26283 33436 26295 33439
rect 26602 33436 26608 33448
rect 26283 33408 26608 33436
rect 26283 33405 26295 33408
rect 26237 33399 26295 33405
rect 26602 33396 26608 33408
rect 26660 33396 26666 33448
rect 27341 33439 27399 33445
rect 27341 33405 27353 33439
rect 27387 33436 27399 33439
rect 27893 33439 27951 33445
rect 27893 33436 27905 33439
rect 27387 33408 27905 33436
rect 27387 33405 27399 33408
rect 27341 33399 27399 33405
rect 27893 33405 27905 33408
rect 27939 33436 27951 33439
rect 28074 33436 28080 33448
rect 27939 33408 28080 33436
rect 27939 33405 27951 33408
rect 27893 33399 27951 33405
rect 28074 33396 28080 33408
rect 28132 33396 28138 33448
rect 24762 33368 24768 33380
rect 23624 33340 24768 33368
rect 23624 33328 23630 33340
rect 24762 33328 24768 33340
rect 24820 33328 24826 33380
rect 26973 33371 27031 33377
rect 26973 33337 26985 33371
rect 27019 33368 27031 33371
rect 27801 33371 27859 33377
rect 27801 33368 27813 33371
rect 27019 33340 27813 33368
rect 27019 33337 27031 33340
rect 26973 33331 27031 33337
rect 27801 33337 27813 33340
rect 27847 33368 27859 33371
rect 28552 33368 28580 33603
rect 28810 33600 28816 33612
rect 28868 33600 28874 33652
rect 35621 33643 35679 33649
rect 35621 33609 35633 33643
rect 35667 33640 35679 33643
rect 35710 33640 35716 33652
rect 35667 33612 35716 33640
rect 35667 33609 35679 33612
rect 35621 33603 35679 33609
rect 35710 33600 35716 33612
rect 35768 33600 35774 33652
rect 35437 33439 35495 33445
rect 35437 33436 35449 33439
rect 27847 33340 28580 33368
rect 35360 33408 35449 33436
rect 27847 33337 27859 33340
rect 27801 33331 27859 33337
rect 35360 33312 35388 33408
rect 35437 33405 35449 33408
rect 35483 33405 35495 33439
rect 35437 33399 35495 33405
rect 7926 33260 7932 33312
rect 7984 33300 7990 33312
rect 8021 33303 8079 33309
rect 8021 33300 8033 33303
rect 7984 33272 8033 33300
rect 7984 33260 7990 33272
rect 8021 33269 8033 33272
rect 8067 33269 8079 33303
rect 8021 33263 8079 33269
rect 15470 33260 15476 33312
rect 15528 33300 15534 33312
rect 16853 33303 16911 33309
rect 16853 33300 16865 33303
rect 15528 33272 16865 33300
rect 15528 33260 15534 33272
rect 16853 33269 16865 33272
rect 16899 33269 16911 33303
rect 16853 33263 16911 33269
rect 17497 33303 17555 33309
rect 17497 33269 17509 33303
rect 17543 33300 17555 33303
rect 17770 33300 17776 33312
rect 17543 33272 17776 33300
rect 17543 33269 17555 33272
rect 17497 33263 17555 33269
rect 17770 33260 17776 33272
rect 17828 33260 17834 33312
rect 25314 33260 25320 33312
rect 25372 33300 25378 33312
rect 25409 33303 25467 33309
rect 25409 33300 25421 33303
rect 25372 33272 25421 33300
rect 25372 33260 25378 33272
rect 25409 33269 25421 33272
rect 25455 33300 25467 33303
rect 26234 33300 26240 33312
rect 25455 33272 26240 33300
rect 25455 33269 25467 33272
rect 25409 33263 25467 33269
rect 26234 33260 26240 33272
rect 26292 33260 26298 33312
rect 26878 33260 26884 33312
rect 26936 33300 26942 33312
rect 27433 33303 27491 33309
rect 27433 33300 27445 33303
rect 26936 33272 27445 33300
rect 26936 33260 26942 33272
rect 27433 33269 27445 33272
rect 27479 33269 27491 33303
rect 27433 33263 27491 33269
rect 28350 33260 28356 33312
rect 28408 33300 28414 33312
rect 28813 33303 28871 33309
rect 28813 33300 28825 33303
rect 28408 33272 28825 33300
rect 28408 33260 28414 33272
rect 28813 33269 28825 33272
rect 28859 33269 28871 33303
rect 35342 33300 35348 33312
rect 35303 33272 35348 33300
rect 28813 33263 28871 33269
rect 35342 33260 35348 33272
rect 35400 33260 35406 33312
rect 35894 33260 35900 33312
rect 35952 33300 35958 33312
rect 35989 33303 36047 33309
rect 35989 33300 36001 33303
rect 35952 33272 36001 33300
rect 35952 33260 35958 33272
rect 35989 33269 36001 33272
rect 36035 33269 36047 33303
rect 35989 33263 36047 33269
rect 1104 33210 38824 33232
rect 1104 33158 19606 33210
rect 19658 33158 19670 33210
rect 19722 33158 19734 33210
rect 19786 33158 19798 33210
rect 19850 33158 38824 33210
rect 1104 33136 38824 33158
rect 4522 33056 4528 33108
rect 4580 33096 4586 33108
rect 5445 33099 5503 33105
rect 5445 33096 5457 33099
rect 4580 33068 5457 33096
rect 4580 33056 4586 33068
rect 5445 33065 5457 33068
rect 5491 33065 5503 33099
rect 5445 33059 5503 33065
rect 5534 33056 5540 33108
rect 5592 33096 5598 33108
rect 5997 33099 6055 33105
rect 5997 33096 6009 33099
rect 5592 33068 6009 33096
rect 5592 33056 5598 33068
rect 5997 33065 6009 33068
rect 6043 33065 6055 33099
rect 8662 33096 8668 33108
rect 8623 33068 8668 33096
rect 5997 33059 6055 33065
rect 8662 33056 8668 33068
rect 8720 33056 8726 33108
rect 9030 33096 9036 33108
rect 8991 33068 9036 33096
rect 9030 33056 9036 33068
rect 9088 33056 9094 33108
rect 10134 33096 10140 33108
rect 10095 33068 10140 33096
rect 10134 33056 10140 33068
rect 10192 33056 10198 33108
rect 11241 33099 11299 33105
rect 11241 33065 11253 33099
rect 11287 33096 11299 33099
rect 11330 33096 11336 33108
rect 11287 33068 11336 33096
rect 11287 33065 11299 33068
rect 11241 33059 11299 33065
rect 11330 33056 11336 33068
rect 11388 33056 11394 33108
rect 11606 33096 11612 33108
rect 11567 33068 11612 33096
rect 11606 33056 11612 33068
rect 11664 33056 11670 33108
rect 13262 33056 13268 33108
rect 13320 33056 13326 33108
rect 13354 33056 13360 33108
rect 13412 33096 13418 33108
rect 15102 33096 15108 33108
rect 13412 33068 13457 33096
rect 15063 33068 15108 33096
rect 13412 33056 13418 33068
rect 15102 33056 15108 33068
rect 15160 33056 15166 33108
rect 17865 33099 17923 33105
rect 17865 33065 17877 33099
rect 17911 33096 17923 33099
rect 17954 33096 17960 33108
rect 17911 33068 17960 33096
rect 17911 33065 17923 33068
rect 17865 33059 17923 33065
rect 17954 33056 17960 33068
rect 18012 33056 18018 33108
rect 19334 33096 19340 33108
rect 19295 33068 19340 33096
rect 19334 33056 19340 33068
rect 19392 33056 19398 33108
rect 20714 33096 20720 33108
rect 20675 33068 20720 33096
rect 20714 33056 20720 33068
rect 20772 33056 20778 33108
rect 21174 33096 21180 33108
rect 21135 33068 21180 33096
rect 21174 33056 21180 33068
rect 21232 33056 21238 33108
rect 21361 33099 21419 33105
rect 21361 33065 21373 33099
rect 21407 33096 21419 33099
rect 23290 33096 23296 33108
rect 21407 33068 23296 33096
rect 21407 33065 21419 33068
rect 21361 33059 21419 33065
rect 23290 33056 23296 33068
rect 23348 33056 23354 33108
rect 23934 33096 23940 33108
rect 23895 33068 23940 33096
rect 23934 33056 23940 33068
rect 23992 33056 23998 33108
rect 24302 33096 24308 33108
rect 24263 33068 24308 33096
rect 24302 33056 24308 33068
rect 24360 33056 24366 33108
rect 25317 33099 25375 33105
rect 25317 33065 25329 33099
rect 25363 33096 25375 33099
rect 25498 33096 25504 33108
rect 25363 33068 25504 33096
rect 25363 33065 25375 33068
rect 25317 33059 25375 33065
rect 25498 33056 25504 33068
rect 25556 33056 25562 33108
rect 25866 33096 25872 33108
rect 25827 33068 25872 33096
rect 25866 33056 25872 33068
rect 25924 33056 25930 33108
rect 26234 33056 26240 33108
rect 26292 33096 26298 33108
rect 26513 33099 26571 33105
rect 26513 33096 26525 33099
rect 26292 33068 26525 33096
rect 26292 33056 26298 33068
rect 26513 33065 26525 33068
rect 26559 33065 26571 33099
rect 26878 33096 26884 33108
rect 26839 33068 26884 33096
rect 26513 33059 26571 33065
rect 26878 33056 26884 33068
rect 26936 33056 26942 33108
rect 27614 33096 27620 33108
rect 27575 33068 27620 33096
rect 27614 33056 27620 33068
rect 27672 33096 27678 33108
rect 27985 33099 28043 33105
rect 27985 33096 27997 33099
rect 27672 33068 27997 33096
rect 27672 33056 27678 33068
rect 27985 33065 27997 33068
rect 28031 33096 28043 33099
rect 28166 33096 28172 33108
rect 28031 33068 28172 33096
rect 28031 33065 28043 33068
rect 27985 33059 28043 33065
rect 28166 33056 28172 33068
rect 28224 33056 28230 33108
rect 4332 33031 4390 33037
rect 4332 32997 4344 33031
rect 4378 33028 4390 33031
rect 4614 33028 4620 33040
rect 4378 33000 4620 33028
rect 4378 32997 4390 33000
rect 4332 32991 4390 32997
rect 4614 32988 4620 33000
rect 4672 32988 4678 33040
rect 8846 32988 8852 33040
rect 8904 33028 8910 33040
rect 9214 33028 9220 33040
rect 8904 33000 9220 33028
rect 8904 32988 8910 33000
rect 9214 32988 9220 33000
rect 9272 33028 9278 33040
rect 9401 33031 9459 33037
rect 9401 33028 9413 33031
rect 9272 33000 9413 33028
rect 9272 32988 9278 33000
rect 9401 32997 9413 33000
rect 9447 32997 9459 33031
rect 10042 33028 10048 33040
rect 10003 33000 10048 33028
rect 9401 32991 9459 32997
rect 10042 32988 10048 33000
rect 10100 32988 10106 33040
rect 13280 33028 13308 33056
rect 21726 33028 21732 33040
rect 13280 33000 13952 33028
rect 21687 33000 21732 33028
rect 4062 32960 4068 32972
rect 4023 32932 4068 32960
rect 4062 32920 4068 32932
rect 4120 32920 4126 32972
rect 6914 32960 6920 32972
rect 6875 32932 6920 32960
rect 6914 32920 6920 32932
rect 6972 32920 6978 32972
rect 8113 32963 8171 32969
rect 8113 32929 8125 32963
rect 8159 32960 8171 32963
rect 8478 32960 8484 32972
rect 8159 32932 8484 32960
rect 8159 32929 8171 32932
rect 8113 32923 8171 32929
rect 8478 32920 8484 32932
rect 8536 32920 8542 32972
rect 12989 32963 13047 32969
rect 12989 32929 13001 32963
rect 13035 32960 13047 32963
rect 13262 32960 13268 32972
rect 13035 32932 13268 32960
rect 13035 32929 13047 32932
rect 12989 32923 13047 32929
rect 13262 32920 13268 32932
rect 13320 32920 13326 32972
rect 13814 32960 13820 32972
rect 13775 32932 13820 32960
rect 13814 32920 13820 32932
rect 13872 32920 13878 32972
rect 13924 32960 13952 33000
rect 21726 32988 21732 33000
rect 21784 32988 21790 33040
rect 22554 32988 22560 33040
rect 22612 33028 22618 33040
rect 22741 33031 22799 33037
rect 22741 33028 22753 33031
rect 22612 33000 22753 33028
rect 22612 32988 22618 33000
rect 22741 32997 22753 33000
rect 22787 33028 22799 33031
rect 23566 33028 23572 33040
rect 22787 33000 23572 33028
rect 22787 32997 22799 33000
rect 22741 32991 22799 32997
rect 23566 32988 23572 33000
rect 23624 32988 23630 33040
rect 25222 33028 25228 33040
rect 25135 33000 25228 33028
rect 25222 32988 25228 33000
rect 25280 33028 25286 33040
rect 25774 33028 25780 33040
rect 25280 33000 25780 33028
rect 25280 32988 25286 33000
rect 25774 32988 25780 33000
rect 25832 32988 25838 33040
rect 26326 32988 26332 33040
rect 26384 33028 26390 33040
rect 26973 33031 27031 33037
rect 26973 33028 26985 33031
rect 26384 33000 26985 33028
rect 26384 32988 26390 33000
rect 26973 32997 26985 33000
rect 27019 33028 27031 33031
rect 27062 33028 27068 33040
rect 27019 33000 27068 33028
rect 27019 32997 27031 33000
rect 26973 32991 27031 32997
rect 27062 32988 27068 33000
rect 27120 32988 27126 33040
rect 15612 32963 15670 32969
rect 13924 32932 14044 32960
rect 7006 32892 7012 32904
rect 6967 32864 7012 32892
rect 7006 32852 7012 32864
rect 7064 32852 7070 32904
rect 7098 32852 7104 32904
rect 7156 32892 7162 32904
rect 7156 32864 7201 32892
rect 7156 32852 7162 32864
rect 10226 32852 10232 32904
rect 10284 32892 10290 32904
rect 10284 32864 10329 32892
rect 10284 32852 10290 32864
rect 11330 32852 11336 32904
rect 11388 32892 11394 32904
rect 11701 32895 11759 32901
rect 11701 32892 11713 32895
rect 11388 32864 11713 32892
rect 11388 32852 11394 32864
rect 11701 32861 11713 32864
rect 11747 32861 11759 32895
rect 11701 32855 11759 32861
rect 11885 32895 11943 32901
rect 11885 32861 11897 32895
rect 11931 32892 11943 32895
rect 12158 32892 12164 32904
rect 11931 32864 12164 32892
rect 11931 32861 11943 32864
rect 11885 32855 11943 32861
rect 12158 32852 12164 32864
rect 12216 32852 12222 32904
rect 13906 32892 13912 32904
rect 13867 32864 13912 32892
rect 13906 32852 13912 32864
rect 13964 32852 13970 32904
rect 14016 32901 14044 32932
rect 15612 32929 15624 32963
rect 15658 32960 15670 32963
rect 15838 32960 15844 32972
rect 15658 32932 15844 32960
rect 15658 32929 15670 32932
rect 15612 32923 15670 32929
rect 15838 32920 15844 32932
rect 15896 32920 15902 32972
rect 17770 32920 17776 32972
rect 17828 32960 17834 32972
rect 18213 32963 18271 32969
rect 18213 32960 18225 32963
rect 17828 32932 18225 32960
rect 17828 32920 17834 32932
rect 18213 32929 18225 32932
rect 18259 32929 18271 32963
rect 21818 32960 21824 32972
rect 21779 32932 21824 32960
rect 18213 32923 18271 32929
rect 21818 32920 21824 32932
rect 21876 32920 21882 32972
rect 14001 32895 14059 32901
rect 14001 32861 14013 32895
rect 14047 32861 14059 32895
rect 14001 32855 14059 32861
rect 14734 32852 14740 32904
rect 14792 32892 14798 32904
rect 15289 32895 15347 32901
rect 15289 32892 15301 32895
rect 14792 32864 15301 32892
rect 14792 32852 14798 32864
rect 15289 32861 15301 32864
rect 15335 32861 15347 32895
rect 15289 32855 15347 32861
rect 15746 32852 15752 32904
rect 15804 32892 15810 32904
rect 16022 32892 16028 32904
rect 15804 32864 15849 32892
rect 15983 32864 16028 32892
rect 15804 32852 15810 32864
rect 16022 32852 16028 32864
rect 16080 32852 16086 32904
rect 17957 32895 18015 32901
rect 17957 32861 17969 32895
rect 18003 32861 18015 32895
rect 21910 32892 21916 32904
rect 21871 32864 21916 32892
rect 17957 32855 18015 32861
rect 3142 32756 3148 32768
rect 3103 32728 3148 32756
rect 3142 32716 3148 32728
rect 3200 32716 3206 32768
rect 6549 32759 6607 32765
rect 6549 32725 6561 32759
rect 6595 32756 6607 32759
rect 7745 32759 7803 32765
rect 7745 32756 7757 32759
rect 6595 32728 7757 32756
rect 6595 32725 6607 32728
rect 6549 32719 6607 32725
rect 7745 32725 7757 32728
rect 7791 32756 7803 32759
rect 8110 32756 8116 32768
rect 7791 32728 8116 32756
rect 7791 32725 7803 32728
rect 7745 32719 7803 32725
rect 8110 32716 8116 32728
rect 8168 32716 8174 32768
rect 8294 32756 8300 32768
rect 8255 32728 8300 32756
rect 8294 32716 8300 32728
rect 8352 32716 8358 32768
rect 9677 32759 9735 32765
rect 9677 32725 9689 32759
rect 9723 32756 9735 32759
rect 11606 32756 11612 32768
rect 9723 32728 11612 32756
rect 9723 32725 9735 32728
rect 9677 32719 9735 32725
rect 11606 32716 11612 32728
rect 11664 32716 11670 32768
rect 12802 32756 12808 32768
rect 12763 32728 12808 32756
rect 12802 32716 12808 32728
rect 12860 32716 12866 32768
rect 13449 32759 13507 32765
rect 13449 32725 13461 32759
rect 13495 32756 13507 32759
rect 13722 32756 13728 32768
rect 13495 32728 13728 32756
rect 13495 32725 13507 32728
rect 13449 32719 13507 32725
rect 13722 32716 13728 32728
rect 13780 32716 13786 32768
rect 13814 32716 13820 32768
rect 13872 32756 13878 32768
rect 14461 32759 14519 32765
rect 14461 32756 14473 32759
rect 13872 32728 14473 32756
rect 13872 32716 13878 32728
rect 14461 32725 14473 32728
rect 14507 32725 14519 32759
rect 17126 32756 17132 32768
rect 17087 32728 17132 32756
rect 14461 32719 14519 32725
rect 17126 32716 17132 32728
rect 17184 32716 17190 32768
rect 17494 32756 17500 32768
rect 17407 32728 17500 32756
rect 17494 32716 17500 32728
rect 17552 32756 17558 32768
rect 17972 32756 18000 32855
rect 21910 32852 21916 32864
rect 21968 32852 21974 32904
rect 23382 32892 23388 32904
rect 23343 32864 23388 32892
rect 23382 32852 23388 32864
rect 23440 32852 23446 32904
rect 23584 32901 23612 32988
rect 24670 32960 24676 32972
rect 24631 32932 24676 32960
rect 24670 32920 24676 32932
rect 24728 32960 24734 32972
rect 28626 32969 28632 32972
rect 28620 32960 28632 32969
rect 24728 32932 25452 32960
rect 28587 32932 28632 32960
rect 24728 32920 24734 32932
rect 25424 32901 25452 32932
rect 28620 32923 28632 32932
rect 28626 32920 28632 32923
rect 28684 32920 28690 32972
rect 23569 32895 23627 32901
rect 23569 32861 23581 32895
rect 23615 32861 23627 32895
rect 23569 32855 23627 32861
rect 25409 32895 25467 32901
rect 25409 32861 25421 32895
rect 25455 32861 25467 32895
rect 25409 32855 25467 32861
rect 26602 32852 26608 32904
rect 26660 32892 26666 32904
rect 27065 32895 27123 32901
rect 27065 32892 27077 32895
rect 26660 32864 27077 32892
rect 26660 32852 26666 32864
rect 27065 32861 27077 32864
rect 27111 32861 27123 32895
rect 28350 32892 28356 32904
rect 28311 32864 28356 32892
rect 27065 32855 27123 32861
rect 28350 32852 28356 32864
rect 28408 32852 28414 32904
rect 18138 32756 18144 32768
rect 17552 32728 18144 32756
rect 17552 32716 17558 32728
rect 18138 32716 18144 32728
rect 18196 32716 18202 32768
rect 22925 32759 22983 32765
rect 22925 32725 22937 32759
rect 22971 32756 22983 32759
rect 23474 32756 23480 32768
rect 22971 32728 23480 32756
rect 22971 32725 22983 32728
rect 22925 32719 22983 32725
rect 23474 32716 23480 32728
rect 23532 32716 23538 32768
rect 24854 32756 24860 32768
rect 24815 32728 24860 32756
rect 24854 32716 24860 32728
rect 24912 32716 24918 32768
rect 26326 32756 26332 32768
rect 26287 32728 26332 32756
rect 26326 32716 26332 32728
rect 26384 32716 26390 32768
rect 28994 32716 29000 32768
rect 29052 32756 29058 32768
rect 29733 32759 29791 32765
rect 29733 32756 29745 32759
rect 29052 32728 29745 32756
rect 29052 32716 29058 32728
rect 29733 32725 29745 32728
rect 29779 32725 29791 32759
rect 29733 32719 29791 32725
rect 1104 32666 38824 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 34966 32666
rect 35018 32614 35030 32666
rect 35082 32614 35094 32666
rect 35146 32614 35158 32666
rect 35210 32614 38824 32666
rect 1104 32592 38824 32614
rect 4525 32555 4583 32561
rect 4525 32521 4537 32555
rect 4571 32552 4583 32555
rect 4614 32552 4620 32564
rect 4571 32524 4620 32552
rect 4571 32521 4583 32524
rect 4525 32515 4583 32521
rect 4614 32512 4620 32524
rect 4672 32552 4678 32564
rect 5077 32555 5135 32561
rect 5077 32552 5089 32555
rect 4672 32524 5089 32552
rect 4672 32512 4678 32524
rect 5077 32521 5089 32524
rect 5123 32521 5135 32555
rect 5534 32552 5540 32564
rect 5495 32524 5540 32552
rect 5077 32515 5135 32521
rect 5534 32512 5540 32524
rect 5592 32512 5598 32564
rect 6454 32512 6460 32564
rect 6512 32552 6518 32564
rect 6641 32555 6699 32561
rect 6641 32552 6653 32555
rect 6512 32524 6653 32552
rect 6512 32512 6518 32524
rect 6641 32521 6653 32524
rect 6687 32552 6699 32555
rect 7006 32552 7012 32564
rect 6687 32524 7012 32552
rect 6687 32521 6699 32524
rect 6641 32515 6699 32521
rect 7006 32512 7012 32524
rect 7064 32512 7070 32564
rect 9953 32555 10011 32561
rect 9953 32521 9965 32555
rect 9999 32552 10011 32555
rect 10042 32552 10048 32564
rect 9999 32524 10048 32552
rect 9999 32521 10011 32524
rect 9953 32515 10011 32521
rect 10042 32512 10048 32524
rect 10100 32512 10106 32564
rect 10226 32552 10232 32564
rect 10187 32524 10232 32552
rect 10226 32512 10232 32524
rect 10284 32512 10290 32564
rect 11606 32552 11612 32564
rect 11567 32524 11612 32552
rect 11606 32512 11612 32524
rect 11664 32512 11670 32564
rect 12069 32555 12127 32561
rect 12069 32521 12081 32555
rect 12115 32552 12127 32555
rect 12158 32552 12164 32564
rect 12115 32524 12164 32552
rect 12115 32521 12127 32524
rect 12069 32515 12127 32521
rect 12158 32512 12164 32524
rect 12216 32512 12222 32564
rect 13170 32552 13176 32564
rect 13131 32524 13176 32552
rect 13170 32512 13176 32524
rect 13228 32512 13234 32564
rect 13541 32555 13599 32561
rect 13541 32521 13553 32555
rect 13587 32552 13599 32555
rect 13906 32552 13912 32564
rect 13587 32524 13912 32552
rect 13587 32521 13599 32524
rect 13541 32515 13599 32521
rect 13906 32512 13912 32524
rect 13964 32552 13970 32564
rect 14642 32552 14648 32564
rect 13964 32524 14648 32552
rect 13964 32512 13970 32524
rect 14642 32512 14648 32524
rect 14700 32552 14706 32564
rect 17037 32555 17095 32561
rect 14700 32524 15772 32552
rect 14700 32512 14706 32524
rect 5813 32487 5871 32493
rect 5813 32453 5825 32487
rect 5859 32484 5871 32487
rect 6914 32484 6920 32496
rect 5859 32456 6920 32484
rect 5859 32453 5871 32456
rect 5813 32447 5871 32453
rect 6914 32444 6920 32456
rect 6972 32484 6978 32496
rect 7101 32487 7159 32493
rect 7101 32484 7113 32487
rect 6972 32456 7113 32484
rect 6972 32444 6978 32456
rect 7101 32453 7113 32456
rect 7147 32453 7159 32487
rect 9490 32484 9496 32496
rect 9451 32456 9496 32484
rect 7101 32447 7159 32453
rect 9490 32444 9496 32456
rect 9548 32444 9554 32496
rect 13814 32484 13820 32496
rect 13775 32456 13820 32484
rect 13814 32444 13820 32456
rect 13872 32444 13878 32496
rect 15744 32484 15772 32524
rect 17037 32521 17049 32555
rect 17083 32552 17095 32555
rect 17494 32552 17500 32564
rect 17083 32524 17500 32552
rect 17083 32521 17095 32524
rect 17037 32515 17095 32521
rect 17494 32512 17500 32524
rect 17552 32512 17558 32564
rect 18046 32552 18052 32564
rect 17959 32524 18052 32552
rect 18046 32512 18052 32524
rect 18104 32552 18110 32564
rect 19058 32552 19064 32564
rect 18104 32524 19064 32552
rect 18104 32512 18110 32524
rect 19058 32512 19064 32524
rect 19116 32552 19122 32564
rect 20165 32555 20223 32561
rect 20165 32552 20177 32555
rect 19116 32524 20177 32552
rect 19116 32512 19122 32524
rect 20165 32521 20177 32524
rect 20211 32552 20223 32555
rect 20714 32552 20720 32564
rect 20211 32524 20720 32552
rect 20211 32521 20223 32524
rect 20165 32515 20223 32521
rect 20714 32512 20720 32524
rect 20772 32512 20778 32564
rect 21726 32512 21732 32564
rect 21784 32552 21790 32564
rect 23661 32555 23719 32561
rect 21784 32524 22416 32552
rect 21784 32512 21790 32524
rect 16209 32487 16267 32493
rect 16209 32484 16221 32487
rect 15744 32456 16221 32484
rect 16209 32453 16221 32456
rect 16255 32453 16267 32487
rect 16209 32447 16267 32453
rect 3142 32416 3148 32428
rect 3103 32388 3148 32416
rect 3142 32376 3148 32388
rect 3200 32376 3206 32428
rect 8294 32416 8300 32428
rect 8255 32388 8300 32416
rect 8294 32376 8300 32388
rect 8352 32416 8358 32428
rect 8757 32419 8815 32425
rect 8757 32416 8769 32419
rect 8352 32388 8769 32416
rect 8352 32376 8358 32388
rect 8757 32385 8769 32388
rect 8803 32385 8815 32419
rect 13832 32416 13860 32444
rect 14832 32419 14890 32425
rect 14832 32416 14844 32419
rect 13832 32388 14844 32416
rect 8757 32379 8815 32385
rect 14832 32385 14844 32388
rect 14878 32385 14890 32419
rect 14832 32379 14890 32385
rect 15746 32376 15752 32428
rect 15804 32416 15810 32428
rect 18064 32425 18092 32512
rect 16485 32419 16543 32425
rect 16485 32416 16497 32419
rect 15804 32388 16497 32416
rect 15804 32376 15810 32388
rect 16485 32385 16497 32388
rect 16531 32385 16543 32419
rect 16485 32379 16543 32385
rect 18049 32419 18107 32425
rect 18049 32385 18061 32419
rect 18095 32385 18107 32419
rect 20732 32416 20760 32512
rect 22388 32493 22416 32524
rect 23661 32521 23673 32555
rect 23707 32552 23719 32555
rect 24210 32552 24216 32564
rect 23707 32524 24216 32552
rect 23707 32521 23719 32524
rect 23661 32515 23719 32521
rect 24210 32512 24216 32524
rect 24268 32512 24274 32564
rect 24949 32555 25007 32561
rect 24949 32521 24961 32555
rect 24995 32552 25007 32555
rect 25498 32552 25504 32564
rect 24995 32524 25504 32552
rect 24995 32521 25007 32524
rect 24949 32515 25007 32521
rect 25498 32512 25504 32524
rect 25556 32512 25562 32564
rect 25958 32512 25964 32564
rect 26016 32552 26022 32564
rect 26053 32555 26111 32561
rect 26053 32552 26065 32555
rect 26016 32524 26065 32552
rect 26016 32512 26022 32524
rect 26053 32521 26065 32524
rect 26099 32521 26111 32555
rect 27062 32552 27068 32564
rect 27023 32524 27068 32552
rect 26053 32515 26111 32521
rect 27062 32512 27068 32524
rect 27120 32512 27126 32564
rect 28626 32512 28632 32564
rect 28684 32552 28690 32564
rect 28721 32555 28779 32561
rect 28721 32552 28733 32555
rect 28684 32524 28733 32552
rect 28684 32512 28690 32524
rect 28721 32521 28733 32524
rect 28767 32552 28779 32555
rect 30653 32555 30711 32561
rect 30653 32552 30665 32555
rect 28767 32524 30665 32552
rect 28767 32521 28779 32524
rect 28721 32515 28779 32521
rect 30653 32521 30665 32524
rect 30699 32521 30711 32555
rect 30653 32515 30711 32521
rect 22373 32487 22431 32493
rect 22373 32453 22385 32487
rect 22419 32484 22431 32487
rect 22925 32487 22983 32493
rect 22925 32484 22937 32487
rect 22419 32456 22937 32484
rect 22419 32453 22431 32456
rect 22373 32447 22431 32453
rect 22925 32453 22937 32456
rect 22971 32453 22983 32487
rect 25222 32484 25228 32496
rect 25183 32456 25228 32484
rect 22925 32447 22983 32453
rect 25222 32444 25228 32456
rect 25280 32444 25286 32496
rect 27617 32487 27675 32493
rect 27617 32484 27629 32487
rect 26528 32456 27629 32484
rect 20993 32419 21051 32425
rect 20993 32416 21005 32419
rect 20732 32388 21005 32416
rect 18049 32379 18107 32385
rect 20993 32385 21005 32388
rect 21039 32385 21051 32419
rect 20993 32379 21051 32385
rect 24118 32376 24124 32428
rect 24176 32416 24182 32428
rect 24305 32419 24363 32425
rect 24305 32416 24317 32419
rect 24176 32388 24317 32416
rect 24176 32376 24182 32388
rect 24305 32385 24317 32388
rect 24351 32416 24363 32419
rect 24670 32416 24676 32428
rect 24351 32388 24676 32416
rect 24351 32385 24363 32388
rect 24305 32379 24363 32385
rect 24670 32376 24676 32388
rect 24728 32376 24734 32428
rect 26142 32376 26148 32428
rect 26200 32416 26206 32428
rect 26528 32425 26556 32456
rect 27617 32453 27629 32456
rect 27663 32453 27675 32487
rect 29086 32484 29092 32496
rect 27617 32447 27675 32453
rect 28092 32456 29092 32484
rect 26513 32419 26571 32425
rect 26513 32416 26525 32419
rect 26200 32388 26525 32416
rect 26200 32376 26206 32388
rect 26513 32385 26525 32388
rect 26559 32385 26571 32419
rect 26513 32379 26571 32385
rect 26602 32376 26608 32428
rect 26660 32416 26666 32428
rect 28092 32425 28120 32456
rect 29086 32444 29092 32456
rect 29144 32444 29150 32496
rect 27525 32419 27583 32425
rect 26660 32388 26705 32416
rect 26660 32376 26666 32388
rect 27525 32385 27537 32419
rect 27571 32416 27583 32419
rect 28077 32419 28135 32425
rect 28077 32416 28089 32419
rect 27571 32388 28089 32416
rect 27571 32385 27583 32388
rect 27525 32379 27583 32385
rect 28077 32385 28089 32388
rect 28123 32385 28135 32419
rect 28077 32379 28135 32385
rect 28166 32376 28172 32428
rect 28224 32416 28230 32428
rect 29104 32416 29132 32444
rect 28224 32388 28269 32416
rect 29104 32388 29408 32416
rect 28224 32376 28230 32388
rect 5534 32308 5540 32360
rect 5592 32348 5598 32360
rect 5629 32351 5687 32357
rect 5629 32348 5641 32351
rect 5592 32320 5641 32348
rect 5592 32308 5598 32320
rect 5629 32317 5641 32320
rect 5675 32348 5687 32351
rect 6181 32351 6239 32357
rect 6181 32348 6193 32351
rect 5675 32320 6193 32348
rect 5675 32317 5687 32320
rect 5629 32311 5687 32317
rect 6181 32317 6193 32320
rect 6227 32317 6239 32351
rect 8110 32348 8116 32360
rect 8071 32320 8116 32348
rect 6181 32311 6239 32317
rect 8110 32308 8116 32320
rect 8168 32348 8174 32360
rect 9125 32351 9183 32357
rect 9125 32348 9137 32351
rect 8168 32320 9137 32348
rect 8168 32308 8174 32320
rect 9125 32317 9137 32320
rect 9171 32348 9183 32351
rect 9309 32351 9367 32357
rect 9309 32348 9321 32351
rect 9171 32320 9321 32348
rect 9171 32317 9183 32320
rect 9125 32311 9183 32317
rect 9309 32317 9321 32320
rect 9355 32317 9367 32351
rect 10870 32348 10876 32360
rect 10831 32320 10876 32348
rect 9309 32311 9367 32317
rect 10870 32308 10876 32320
rect 10928 32308 10934 32360
rect 11330 32348 11336 32360
rect 11291 32320 11336 32348
rect 11330 32308 11336 32320
rect 11388 32308 11394 32360
rect 14369 32351 14427 32357
rect 14369 32317 14381 32351
rect 14415 32348 14427 32351
rect 14734 32348 14740 32360
rect 14415 32320 14740 32348
rect 14415 32317 14427 32320
rect 14369 32311 14427 32317
rect 14734 32308 14740 32320
rect 14792 32308 14798 32360
rect 15102 32348 15108 32360
rect 15063 32320 15108 32348
rect 15102 32308 15108 32320
rect 15160 32308 15166 32360
rect 17034 32308 17040 32360
rect 17092 32348 17098 32360
rect 17221 32351 17279 32357
rect 17221 32348 17233 32351
rect 17092 32320 17233 32348
rect 17092 32308 17098 32320
rect 17221 32317 17233 32320
rect 17267 32317 17279 32351
rect 17221 32311 17279 32317
rect 18316 32351 18374 32357
rect 18316 32317 18328 32351
rect 18362 32348 18374 32351
rect 18598 32348 18604 32360
rect 18362 32320 18604 32348
rect 18362 32317 18374 32320
rect 18316 32311 18374 32317
rect 18598 32308 18604 32320
rect 18656 32348 18662 32360
rect 19242 32348 19248 32360
rect 18656 32320 19248 32348
rect 18656 32308 18662 32320
rect 19242 32308 19248 32320
rect 19300 32308 19306 32360
rect 20533 32351 20591 32357
rect 20533 32317 20545 32351
rect 20579 32348 20591 32351
rect 20901 32351 20959 32357
rect 20901 32348 20913 32351
rect 20579 32320 20913 32348
rect 20579 32317 20591 32320
rect 20533 32311 20591 32317
rect 20901 32317 20913 32320
rect 20947 32348 20959 32351
rect 21260 32351 21318 32357
rect 21260 32348 21272 32351
rect 20947 32320 21272 32348
rect 20947 32317 20959 32320
rect 20901 32311 20959 32317
rect 21260 32317 21272 32320
rect 21306 32348 21318 32351
rect 21818 32348 21824 32360
rect 21306 32320 21824 32348
rect 21306 32317 21318 32320
rect 21260 32311 21318 32317
rect 21818 32308 21824 32320
rect 21876 32308 21882 32360
rect 23934 32308 23940 32360
rect 23992 32348 23998 32360
rect 24029 32351 24087 32357
rect 24029 32348 24041 32351
rect 23992 32320 24041 32348
rect 23992 32308 23998 32320
rect 24029 32317 24041 32320
rect 24075 32317 24087 32351
rect 24029 32311 24087 32317
rect 25961 32351 26019 32357
rect 25961 32317 25973 32351
rect 26007 32348 26019 32351
rect 26878 32348 26884 32360
rect 26007 32320 26884 32348
rect 26007 32317 26019 32320
rect 25961 32311 26019 32317
rect 26878 32308 26884 32320
rect 26936 32308 26942 32360
rect 27706 32308 27712 32360
rect 27764 32348 27770 32360
rect 27985 32351 28043 32357
rect 27985 32348 27997 32351
rect 27764 32320 27997 32348
rect 27764 32308 27770 32320
rect 27985 32317 27997 32320
rect 28031 32348 28043 32351
rect 28626 32348 28632 32360
rect 28031 32320 28632 32348
rect 28031 32317 28043 32320
rect 27985 32311 28043 32317
rect 28626 32308 28632 32320
rect 28684 32308 28690 32360
rect 29270 32348 29276 32360
rect 29231 32320 29276 32348
rect 29270 32308 29276 32320
rect 29328 32308 29334 32360
rect 29380 32348 29408 32388
rect 29529 32351 29587 32357
rect 29529 32348 29541 32351
rect 29380 32320 29541 32348
rect 29529 32317 29541 32320
rect 29575 32317 29587 32351
rect 29529 32311 29587 32317
rect 3053 32283 3111 32289
rect 3053 32249 3065 32283
rect 3099 32280 3111 32283
rect 3390 32283 3448 32289
rect 3390 32280 3402 32283
rect 3099 32252 3402 32280
rect 3099 32249 3111 32252
rect 3053 32243 3111 32249
rect 3390 32249 3402 32252
rect 3436 32280 3448 32283
rect 3602 32280 3608 32292
rect 3436 32252 3608 32280
rect 3436 32249 3448 32252
rect 3390 32243 3448 32249
rect 3602 32240 3608 32252
rect 3660 32240 3666 32292
rect 8018 32280 8024 32292
rect 7576 32252 8024 32280
rect 2038 32212 2044 32224
rect 1999 32184 2044 32212
rect 2038 32172 2044 32184
rect 2096 32172 2102 32224
rect 2409 32215 2467 32221
rect 2409 32181 2421 32215
rect 2455 32212 2467 32215
rect 2590 32212 2596 32224
rect 2455 32184 2596 32212
rect 2455 32181 2467 32184
rect 2409 32175 2467 32181
rect 2590 32172 2596 32184
rect 2648 32172 2654 32224
rect 5810 32172 5816 32224
rect 5868 32212 5874 32224
rect 7576 32221 7604 32252
rect 8018 32240 8024 32252
rect 8076 32280 8082 32292
rect 8205 32283 8263 32289
rect 8205 32280 8217 32283
rect 8076 32252 8217 32280
rect 8076 32240 8082 32252
rect 8205 32249 8217 32252
rect 8251 32249 8263 32283
rect 8205 32243 8263 32249
rect 12805 32283 12863 32289
rect 12805 32249 12817 32283
rect 12851 32280 12863 32283
rect 13262 32280 13268 32292
rect 12851 32252 13268 32280
rect 12851 32249 12863 32252
rect 12805 32243 12863 32249
rect 13262 32240 13268 32252
rect 13320 32240 13326 32292
rect 16666 32240 16672 32292
rect 16724 32280 16730 32292
rect 17770 32280 17776 32292
rect 16724 32252 17776 32280
rect 16724 32240 16730 32252
rect 17770 32240 17776 32252
rect 17828 32240 17834 32292
rect 23477 32283 23535 32289
rect 23477 32249 23489 32283
rect 23523 32280 23535 32283
rect 23566 32280 23572 32292
rect 23523 32252 23572 32280
rect 23523 32249 23535 32252
rect 23477 32243 23535 32249
rect 23566 32240 23572 32252
rect 23624 32280 23630 32292
rect 24121 32283 24179 32289
rect 24121 32280 24133 32283
rect 23624 32252 24133 32280
rect 23624 32240 23630 32252
rect 24121 32249 24133 32252
rect 24167 32249 24179 32283
rect 24121 32243 24179 32249
rect 26326 32240 26332 32292
rect 26384 32280 26390 32292
rect 26421 32283 26479 32289
rect 26421 32280 26433 32283
rect 26384 32252 26433 32280
rect 26384 32240 26390 32252
rect 26421 32249 26433 32252
rect 26467 32280 26479 32283
rect 27522 32280 27528 32292
rect 26467 32252 27528 32280
rect 26467 32249 26479 32252
rect 26421 32243 26479 32249
rect 27522 32240 27528 32252
rect 27580 32240 27586 32292
rect 7561 32215 7619 32221
rect 7561 32212 7573 32215
rect 5868 32184 7573 32212
rect 5868 32172 5874 32184
rect 7561 32181 7573 32184
rect 7607 32181 7619 32215
rect 7742 32212 7748 32224
rect 7703 32184 7748 32212
rect 7561 32175 7619 32181
rect 7742 32172 7748 32184
rect 7800 32172 7806 32224
rect 9858 32172 9864 32224
rect 9916 32212 9922 32224
rect 10689 32215 10747 32221
rect 10689 32212 10701 32215
rect 9916 32184 10701 32212
rect 9916 32172 9922 32184
rect 10689 32181 10701 32184
rect 10735 32181 10747 32215
rect 10689 32175 10747 32181
rect 14277 32215 14335 32221
rect 14277 32181 14289 32215
rect 14323 32212 14335 32215
rect 14835 32215 14893 32221
rect 14835 32212 14847 32215
rect 14323 32184 14847 32212
rect 14323 32181 14335 32184
rect 14277 32175 14335 32181
rect 14835 32181 14847 32184
rect 14881 32212 14893 32215
rect 15838 32212 15844 32224
rect 14881 32184 15844 32212
rect 14881 32181 14893 32184
rect 14835 32175 14893 32181
rect 15838 32172 15844 32184
rect 15896 32172 15902 32224
rect 16942 32212 16948 32224
rect 16903 32184 16948 32212
rect 16942 32172 16948 32184
rect 17000 32172 17006 32224
rect 19334 32172 19340 32224
rect 19392 32212 19398 32224
rect 19429 32215 19487 32221
rect 19429 32212 19441 32215
rect 19392 32184 19441 32212
rect 19392 32172 19398 32184
rect 19429 32181 19441 32184
rect 19475 32181 19487 32215
rect 19429 32175 19487 32181
rect 1104 32122 38824 32144
rect 1104 32070 19606 32122
rect 19658 32070 19670 32122
rect 19722 32070 19734 32122
rect 19786 32070 19798 32122
rect 19850 32070 38824 32122
rect 1104 32048 38824 32070
rect 1949 32011 2007 32017
rect 1949 31977 1961 32011
rect 1995 32008 2007 32011
rect 2866 32008 2872 32020
rect 1995 31980 2872 32008
rect 1995 31977 2007 31980
rect 1949 31971 2007 31977
rect 2866 31968 2872 31980
rect 2924 31968 2930 32020
rect 3053 32011 3111 32017
rect 3053 31977 3065 32011
rect 3099 32008 3111 32011
rect 3142 32008 3148 32020
rect 3099 31980 3148 32008
rect 3099 31977 3111 31980
rect 3053 31971 3111 31977
rect 2774 31900 2780 31952
rect 2832 31940 2838 31952
rect 3068 31940 3096 31971
rect 3142 31968 3148 31980
rect 3200 31968 3206 32020
rect 3602 31968 3608 32020
rect 3660 32008 3666 32020
rect 4433 32011 4491 32017
rect 4433 32008 4445 32011
rect 3660 31980 4445 32008
rect 3660 31968 3666 31980
rect 4433 31977 4445 31980
rect 4479 31977 4491 32011
rect 4433 31971 4491 31977
rect 4982 31968 4988 32020
rect 5040 32008 5046 32020
rect 5077 32011 5135 32017
rect 5077 32008 5089 32011
rect 5040 31980 5089 32008
rect 5040 31968 5046 31980
rect 5077 31977 5089 31980
rect 5123 32008 5135 32011
rect 5166 32008 5172 32020
rect 5123 31980 5172 32008
rect 5123 31977 5135 31980
rect 5077 31971 5135 31977
rect 5166 31968 5172 31980
rect 5224 31968 5230 32020
rect 5810 32008 5816 32020
rect 5771 31980 5816 32008
rect 5810 31968 5816 31980
rect 5868 31968 5874 32020
rect 6546 31968 6552 32020
rect 6604 32008 6610 32020
rect 6917 32011 6975 32017
rect 6917 32008 6929 32011
rect 6604 31980 6929 32008
rect 6604 31968 6610 31980
rect 6917 31977 6929 31980
rect 6963 32008 6975 32011
rect 7098 32008 7104 32020
rect 6963 31980 7104 32008
rect 6963 31977 6975 31980
rect 6917 31971 6975 31977
rect 7098 31968 7104 31980
rect 7156 31968 7162 32020
rect 8021 32011 8079 32017
rect 8021 31977 8033 32011
rect 8067 31977 8079 32011
rect 8478 32008 8484 32020
rect 8439 31980 8484 32008
rect 8021 31971 8079 31977
rect 2832 31912 3096 31940
rect 4525 31943 4583 31949
rect 2832 31900 2838 31912
rect 4525 31909 4537 31943
rect 4571 31940 4583 31943
rect 4614 31940 4620 31952
rect 4571 31912 4620 31940
rect 4571 31909 4583 31912
rect 4525 31903 4583 31909
rect 4614 31900 4620 31912
rect 4672 31900 4678 31952
rect 8036 31940 8064 31971
rect 8478 31968 8484 31980
rect 8536 31968 8542 32020
rect 9033 32011 9091 32017
rect 9033 31977 9045 32011
rect 9079 32008 9091 32011
rect 9582 32008 9588 32020
rect 9079 31980 9588 32008
rect 9079 31977 9091 31980
rect 9033 31971 9091 31977
rect 9582 31968 9588 31980
rect 9640 31968 9646 32020
rect 9953 32011 10011 32017
rect 9953 31977 9965 32011
rect 9999 32008 10011 32011
rect 10134 32008 10140 32020
rect 9999 31980 10140 32008
rect 9999 31977 10011 31980
rect 9953 31971 10011 31977
rect 10134 31968 10140 31980
rect 10192 31968 10198 32020
rect 10781 32011 10839 32017
rect 10781 31977 10793 32011
rect 10827 32008 10839 32011
rect 10870 32008 10876 32020
rect 10827 31980 10876 32008
rect 10827 31977 10839 31980
rect 10781 31971 10839 31977
rect 10870 31968 10876 31980
rect 10928 31968 10934 32020
rect 14090 32008 14096 32020
rect 14051 31980 14096 32008
rect 14090 31968 14096 31980
rect 14148 31968 14154 32020
rect 14645 32011 14703 32017
rect 14645 31977 14657 32011
rect 14691 32008 14703 32011
rect 15102 32008 15108 32020
rect 14691 31980 15108 32008
rect 14691 31977 14703 31980
rect 14645 31971 14703 31977
rect 15102 31968 15108 31980
rect 15160 31968 15166 32020
rect 15565 32011 15623 32017
rect 15565 31977 15577 32011
rect 15611 32008 15623 32011
rect 16022 32008 16028 32020
rect 15611 31980 16028 32008
rect 15611 31977 15623 31980
rect 15565 31971 15623 31977
rect 16022 31968 16028 31980
rect 16080 31968 16086 32020
rect 17494 32008 17500 32020
rect 17455 31980 17500 32008
rect 17494 31968 17500 31980
rect 17552 31968 17558 32020
rect 17589 32011 17647 32017
rect 17589 31977 17601 32011
rect 17635 32008 17647 32011
rect 17862 32008 17868 32020
rect 17635 31980 17868 32008
rect 17635 31977 17647 31980
rect 17589 31971 17647 31977
rect 17862 31968 17868 31980
rect 17920 31968 17926 32020
rect 18598 32008 18604 32020
rect 18559 31980 18604 32008
rect 18598 31968 18604 31980
rect 18656 31968 18662 32020
rect 19058 32008 19064 32020
rect 19019 31980 19064 32008
rect 19058 31968 19064 31980
rect 19116 31968 19122 32020
rect 21818 31968 21824 32020
rect 21876 32008 21882 32020
rect 22373 32011 22431 32017
rect 22373 32008 22385 32011
rect 21876 31980 22385 32008
rect 21876 31968 21882 31980
rect 22373 31977 22385 31980
rect 22419 31977 22431 32011
rect 22373 31971 22431 31977
rect 23017 32011 23075 32017
rect 23017 31977 23029 32011
rect 23063 32008 23075 32011
rect 23382 32008 23388 32020
rect 23063 31980 23388 32008
rect 23063 31977 23075 31980
rect 23017 31971 23075 31977
rect 8662 31940 8668 31952
rect 8036 31912 8668 31940
rect 8662 31900 8668 31912
rect 8720 31900 8726 31952
rect 14734 31900 14740 31952
rect 14792 31940 14798 31952
rect 16942 31940 16948 31952
rect 14792 31912 16948 31940
rect 14792 31900 14798 31912
rect 16942 31900 16948 31912
rect 17000 31900 17006 31952
rect 17957 31943 18015 31949
rect 17957 31909 17969 31943
rect 18003 31940 18015 31943
rect 18046 31940 18052 31952
rect 18003 31912 18052 31940
rect 18003 31909 18015 31912
rect 17957 31903 18015 31909
rect 18046 31900 18052 31912
rect 18104 31900 18110 31952
rect 20717 31943 20775 31949
rect 20717 31909 20729 31943
rect 20763 31940 20775 31943
rect 21910 31940 21916 31952
rect 20763 31912 21916 31940
rect 20763 31909 20775 31912
rect 20717 31903 20775 31909
rect 21910 31900 21916 31912
rect 21968 31900 21974 31952
rect 22002 31900 22008 31952
rect 22060 31940 22066 31952
rect 23032 31940 23060 31971
rect 23382 31968 23388 31980
rect 23440 31968 23446 32020
rect 23566 31968 23572 32020
rect 23624 32008 23630 32020
rect 23661 32011 23719 32017
rect 23661 32008 23673 32011
rect 23624 31980 23673 32008
rect 23624 31968 23630 31980
rect 23661 31977 23673 31980
rect 23707 31977 23719 32011
rect 24118 32008 24124 32020
rect 24079 31980 24124 32008
rect 23661 31971 23719 31977
rect 24118 31968 24124 31980
rect 24176 31968 24182 32020
rect 24854 31968 24860 32020
rect 24912 32008 24918 32020
rect 25041 32011 25099 32017
rect 25041 32008 25053 32011
rect 24912 31980 25053 32008
rect 24912 31968 24918 31980
rect 25041 31977 25053 31980
rect 25087 31977 25099 32011
rect 26142 32008 26148 32020
rect 26103 31980 26148 32008
rect 25041 31971 25099 31977
rect 26142 31968 26148 31980
rect 26200 31968 26206 32020
rect 27062 32008 27068 32020
rect 26712 31980 27068 32008
rect 23290 31940 23296 31952
rect 22060 31912 23060 31940
rect 23251 31912 23296 31940
rect 22060 31900 22066 31912
rect 23290 31900 23296 31912
rect 23348 31900 23354 31952
rect 24210 31900 24216 31952
rect 24268 31940 24274 31952
rect 25133 31943 25191 31949
rect 25133 31940 25145 31943
rect 24268 31912 25145 31940
rect 24268 31900 24274 31912
rect 25133 31909 25145 31912
rect 25179 31909 25191 31943
rect 26602 31940 26608 31952
rect 25133 31903 25191 31909
rect 25700 31912 26608 31940
rect 2038 31832 2044 31884
rect 2096 31872 2102 31884
rect 2317 31875 2375 31881
rect 2317 31872 2329 31875
rect 2096 31844 2329 31872
rect 2096 31832 2102 31844
rect 2317 31841 2329 31844
rect 2363 31841 2375 31875
rect 6178 31872 6184 31884
rect 6139 31844 6184 31872
rect 2317 31835 2375 31841
rect 6178 31832 6184 31844
rect 6236 31832 6242 31884
rect 7742 31832 7748 31884
rect 7800 31872 7806 31884
rect 7837 31875 7895 31881
rect 7837 31872 7849 31875
rect 7800 31844 7849 31872
rect 7800 31832 7806 31844
rect 7837 31841 7849 31844
rect 7883 31872 7895 31875
rect 8294 31872 8300 31884
rect 7883 31844 8300 31872
rect 7883 31841 7895 31844
rect 7837 31835 7895 31841
rect 8294 31832 8300 31844
rect 8352 31832 8358 31884
rect 9214 31872 9220 31884
rect 9175 31844 9220 31872
rect 9214 31832 9220 31844
rect 9272 31872 9278 31884
rect 9858 31872 9864 31884
rect 9272 31844 9864 31872
rect 9272 31832 9278 31844
rect 9858 31832 9864 31844
rect 9916 31832 9922 31884
rect 14826 31832 14832 31884
rect 14884 31872 14890 31884
rect 16209 31875 16267 31881
rect 16209 31872 16221 31875
rect 14884 31844 16221 31872
rect 14884 31832 14890 31844
rect 16209 31841 16221 31844
rect 16255 31872 16267 31875
rect 16485 31875 16543 31881
rect 16485 31872 16497 31875
rect 16255 31844 16497 31872
rect 16255 31841 16267 31844
rect 16209 31835 16267 31841
rect 16485 31841 16497 31844
rect 16531 31872 16543 31875
rect 17034 31872 17040 31884
rect 16531 31844 17040 31872
rect 16531 31841 16543 31844
rect 16485 31835 16543 31841
rect 17034 31832 17040 31844
rect 17092 31832 17098 31884
rect 21260 31875 21318 31881
rect 21260 31841 21272 31875
rect 21306 31872 21318 31875
rect 21542 31872 21548 31884
rect 21306 31844 21548 31872
rect 21306 31841 21318 31844
rect 21260 31835 21318 31841
rect 21542 31832 21548 31844
rect 21600 31832 21606 31884
rect 23474 31872 23480 31884
rect 23435 31844 23480 31872
rect 23474 31832 23480 31844
rect 23532 31832 23538 31884
rect 24762 31832 24768 31884
rect 24820 31872 24826 31884
rect 25700 31881 25728 31912
rect 26602 31900 26608 31912
rect 26660 31900 26666 31952
rect 26712 31949 26740 31980
rect 27062 31968 27068 31980
rect 27120 32008 27126 32020
rect 29549 32011 29607 32017
rect 29549 32008 29561 32011
rect 27120 31980 29561 32008
rect 27120 31968 27126 31980
rect 29549 31977 29561 31980
rect 29595 31977 29607 32011
rect 29549 31971 29607 31977
rect 35621 32011 35679 32017
rect 35621 31977 35633 32011
rect 35667 32008 35679 32011
rect 35802 32008 35808 32020
rect 35667 31980 35808 32008
rect 35667 31977 35679 31980
rect 35621 31971 35679 31977
rect 35802 31968 35808 31980
rect 35860 31968 35866 32020
rect 26697 31943 26755 31949
rect 26697 31909 26709 31943
rect 26743 31909 26755 31943
rect 27706 31940 27712 31952
rect 27667 31912 27712 31940
rect 26697 31903 26755 31909
rect 27706 31900 27712 31912
rect 27764 31900 27770 31952
rect 25685 31875 25743 31881
rect 25685 31872 25697 31875
rect 24820 31844 25697 31872
rect 24820 31832 24826 31844
rect 25685 31841 25697 31844
rect 25731 31841 25743 31875
rect 25685 31835 25743 31841
rect 26234 31832 26240 31884
rect 26292 31872 26298 31884
rect 26513 31875 26571 31881
rect 26513 31872 26525 31875
rect 26292 31844 26525 31872
rect 26292 31832 26298 31844
rect 26513 31841 26525 31844
rect 26559 31841 26571 31875
rect 26620 31872 26648 31900
rect 27157 31875 27215 31881
rect 27157 31872 27169 31875
rect 26620 31844 27169 31872
rect 26513 31835 26571 31841
rect 27157 31841 27169 31844
rect 27203 31841 27215 31875
rect 27157 31835 27215 31841
rect 28436 31875 28494 31881
rect 28436 31841 28448 31875
rect 28482 31872 28494 31875
rect 28718 31872 28724 31884
rect 28482 31844 28724 31872
rect 28482 31841 28494 31844
rect 28436 31835 28494 31841
rect 28718 31832 28724 31844
rect 28776 31832 28782 31884
rect 35434 31872 35440 31884
rect 35395 31844 35440 31872
rect 35434 31832 35440 31844
rect 35492 31832 35498 31884
rect 2409 31807 2467 31813
rect 2409 31773 2421 31807
rect 2455 31773 2467 31807
rect 2590 31804 2596 31816
rect 2503 31776 2596 31804
rect 2409 31767 2467 31773
rect 1670 31628 1676 31680
rect 1728 31668 1734 31680
rect 1765 31671 1823 31677
rect 1765 31668 1777 31671
rect 1728 31640 1777 31668
rect 1728 31628 1734 31640
rect 1765 31637 1777 31640
rect 1811 31668 1823 31671
rect 2424 31668 2452 31767
rect 2590 31764 2596 31776
rect 2648 31764 2654 31816
rect 4709 31807 4767 31813
rect 4709 31773 4721 31807
rect 4755 31804 4767 31807
rect 4755 31776 4789 31804
rect 4755 31773 4767 31776
rect 4709 31767 4767 31773
rect 2608 31736 2636 31764
rect 4724 31736 4752 31767
rect 5810 31764 5816 31816
rect 5868 31804 5874 31816
rect 6273 31807 6331 31813
rect 6273 31804 6285 31807
rect 5868 31776 6285 31804
rect 5868 31764 5874 31776
rect 6273 31773 6285 31776
rect 6319 31773 6331 31807
rect 6273 31767 6331 31773
rect 6457 31807 6515 31813
rect 6457 31773 6469 31807
rect 6503 31804 6515 31807
rect 6546 31804 6552 31816
rect 6503 31776 6552 31804
rect 6503 31773 6515 31776
rect 6457 31767 6515 31773
rect 6546 31764 6552 31776
rect 6604 31764 6610 31816
rect 18049 31807 18107 31813
rect 18049 31804 18061 31807
rect 17880 31776 18061 31804
rect 4982 31736 4988 31748
rect 2608 31708 4988 31736
rect 4982 31696 4988 31708
rect 5040 31696 5046 31748
rect 17678 31696 17684 31748
rect 17736 31736 17742 31748
rect 17880 31736 17908 31776
rect 18049 31773 18061 31776
rect 18095 31773 18107 31807
rect 18049 31767 18107 31773
rect 18141 31807 18199 31813
rect 18141 31773 18153 31807
rect 18187 31804 18199 31807
rect 20990 31804 20996 31816
rect 18187 31776 18221 31804
rect 20951 31776 20996 31804
rect 18187 31773 18199 31776
rect 18141 31767 18199 31773
rect 17736 31708 17908 31736
rect 17736 31696 17742 31708
rect 17954 31696 17960 31748
rect 18012 31736 18018 31748
rect 18156 31736 18184 31767
rect 20990 31764 20996 31776
rect 21048 31764 21054 31816
rect 24118 31764 24124 31816
rect 24176 31804 24182 31816
rect 24489 31807 24547 31813
rect 24489 31804 24501 31807
rect 24176 31776 24501 31804
rect 24176 31764 24182 31776
rect 24489 31773 24501 31776
rect 24535 31804 24547 31807
rect 25225 31807 25283 31813
rect 24535 31776 24808 31804
rect 24535 31773 24547 31776
rect 24489 31767 24547 31773
rect 18012 31708 18184 31736
rect 24780 31736 24808 31776
rect 25225 31773 25237 31807
rect 25271 31804 25283 31807
rect 26878 31804 26884 31816
rect 25271 31776 25305 31804
rect 26839 31776 26884 31804
rect 25271 31773 25283 31776
rect 25225 31767 25283 31773
rect 25240 31736 25268 31767
rect 26878 31764 26884 31776
rect 26936 31764 26942 31816
rect 28169 31807 28227 31813
rect 28169 31773 28181 31807
rect 28215 31773 28227 31807
rect 28169 31767 28227 31773
rect 24780 31708 25268 31736
rect 18012 31696 18018 31708
rect 1811 31640 2452 31668
rect 4065 31671 4123 31677
rect 1811 31637 1823 31640
rect 1765 31631 1823 31637
rect 4065 31637 4077 31671
rect 4111 31668 4123 31671
rect 5074 31668 5080 31680
rect 4111 31640 5080 31668
rect 4111 31637 4123 31640
rect 4065 31631 4123 31637
rect 5074 31628 5080 31640
rect 5132 31628 5138 31680
rect 5258 31628 5264 31680
rect 5316 31668 5322 31680
rect 5445 31671 5503 31677
rect 5445 31668 5457 31671
rect 5316 31640 5457 31668
rect 5316 31628 5322 31640
rect 5445 31637 5457 31640
rect 5491 31637 5503 31671
rect 5445 31631 5503 31637
rect 14734 31628 14740 31680
rect 14792 31668 14798 31680
rect 14921 31671 14979 31677
rect 14921 31668 14933 31671
rect 14792 31640 14933 31668
rect 14792 31628 14798 31640
rect 14921 31637 14933 31640
rect 14967 31637 14979 31671
rect 15838 31668 15844 31680
rect 15799 31640 15844 31668
rect 14921 31631 14979 31637
rect 15838 31628 15844 31640
rect 15896 31628 15902 31680
rect 16025 31671 16083 31677
rect 16025 31637 16037 31671
rect 16071 31668 16083 31671
rect 16206 31668 16212 31680
rect 16071 31640 16212 31668
rect 16071 31637 16083 31640
rect 16025 31631 16083 31637
rect 16206 31628 16212 31640
rect 16264 31628 16270 31680
rect 24670 31668 24676 31680
rect 24631 31640 24676 31668
rect 24670 31628 24676 31640
rect 24728 31628 24734 31680
rect 28077 31671 28135 31677
rect 28077 31637 28089 31671
rect 28123 31668 28135 31671
rect 28184 31668 28212 31767
rect 28350 31668 28356 31680
rect 28123 31640 28356 31668
rect 28123 31637 28135 31640
rect 28077 31631 28135 31637
rect 28350 31628 28356 31640
rect 28408 31668 28414 31680
rect 28810 31668 28816 31680
rect 28408 31640 28816 31668
rect 28408 31628 28414 31640
rect 28810 31628 28816 31640
rect 28868 31668 28874 31680
rect 29270 31668 29276 31680
rect 28868 31640 29276 31668
rect 28868 31628 28874 31640
rect 29270 31628 29276 31640
rect 29328 31668 29334 31680
rect 30101 31671 30159 31677
rect 30101 31668 30113 31671
rect 29328 31640 30113 31668
rect 29328 31628 29334 31640
rect 30101 31637 30113 31640
rect 30147 31637 30159 31671
rect 30101 31631 30159 31637
rect 1104 31578 38824 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 34966 31578
rect 35018 31526 35030 31578
rect 35082 31526 35094 31578
rect 35146 31526 35158 31578
rect 35210 31526 38824 31578
rect 1104 31504 38824 31526
rect 3602 31464 3608 31476
rect 3563 31436 3608 31464
rect 3602 31424 3608 31436
rect 3660 31464 3666 31476
rect 4525 31467 4583 31473
rect 4525 31464 4537 31467
rect 3660 31436 4537 31464
rect 3660 31424 3666 31436
rect 4525 31433 4537 31436
rect 4571 31433 4583 31467
rect 6546 31464 6552 31476
rect 6507 31436 6552 31464
rect 4525 31427 4583 31433
rect 6546 31424 6552 31436
rect 6604 31424 6610 31476
rect 7926 31464 7932 31476
rect 7887 31436 7932 31464
rect 7926 31424 7932 31436
rect 7984 31424 7990 31476
rect 8294 31424 8300 31476
rect 8352 31464 8358 31476
rect 8665 31467 8723 31473
rect 8665 31464 8677 31467
rect 8352 31436 8677 31464
rect 8352 31424 8358 31436
rect 8665 31433 8677 31436
rect 8711 31433 8723 31467
rect 13170 31464 13176 31476
rect 13131 31436 13176 31464
rect 8665 31427 8723 31433
rect 13170 31424 13176 31436
rect 13228 31424 13234 31476
rect 14274 31464 14280 31476
rect 14235 31436 14280 31464
rect 14274 31424 14280 31436
rect 14332 31424 14338 31476
rect 17313 31467 17371 31473
rect 17313 31433 17325 31467
rect 17359 31464 17371 31467
rect 17954 31464 17960 31476
rect 17359 31436 17960 31464
rect 17359 31433 17371 31436
rect 17313 31427 17371 31433
rect 17954 31424 17960 31436
rect 18012 31424 18018 31476
rect 21177 31467 21235 31473
rect 21177 31433 21189 31467
rect 21223 31464 21235 31467
rect 22002 31464 22008 31476
rect 21223 31436 22008 31464
rect 21223 31433 21235 31436
rect 21177 31427 21235 31433
rect 22002 31424 22008 31436
rect 22060 31424 22066 31476
rect 23474 31464 23480 31476
rect 23435 31436 23480 31464
rect 23474 31424 23480 31436
rect 23532 31424 23538 31476
rect 24210 31464 24216 31476
rect 24171 31436 24216 31464
rect 24210 31424 24216 31436
rect 24268 31424 24274 31476
rect 26234 31424 26240 31476
rect 26292 31464 26298 31476
rect 26605 31467 26663 31473
rect 26605 31464 26617 31467
rect 26292 31436 26617 31464
rect 26292 31424 26298 31436
rect 26605 31433 26617 31436
rect 26651 31433 26663 31467
rect 27062 31464 27068 31476
rect 27023 31436 27068 31464
rect 26605 31427 26663 31433
rect 27062 31424 27068 31436
rect 27120 31424 27126 31476
rect 27614 31464 27620 31476
rect 27575 31436 27620 31464
rect 27614 31424 27620 31436
rect 27672 31424 27678 31476
rect 4249 31399 4307 31405
rect 4249 31365 4261 31399
rect 4295 31396 4307 31399
rect 4614 31396 4620 31408
rect 4295 31368 4620 31396
rect 4295 31365 4307 31368
rect 4249 31359 4307 31365
rect 1394 31220 1400 31272
rect 1452 31260 1458 31272
rect 2225 31263 2283 31269
rect 2225 31260 2237 31263
rect 1452 31232 2237 31260
rect 1452 31220 1458 31232
rect 2225 31229 2237 31232
rect 2271 31260 2283 31263
rect 2774 31260 2780 31272
rect 2271 31232 2780 31260
rect 2271 31229 2283 31232
rect 2225 31223 2283 31229
rect 2774 31220 2780 31232
rect 2832 31220 2838 31272
rect 2133 31195 2191 31201
rect 2133 31161 2145 31195
rect 2179 31192 2191 31195
rect 2492 31195 2550 31201
rect 2492 31192 2504 31195
rect 2179 31164 2504 31192
rect 2179 31161 2191 31164
rect 2133 31155 2191 31161
rect 2492 31161 2504 31164
rect 2538 31192 2550 31195
rect 2866 31192 2872 31204
rect 2538 31164 2872 31192
rect 2538 31161 2550 31164
rect 2492 31155 2550 31161
rect 2866 31152 2872 31164
rect 2924 31192 2930 31204
rect 4264 31192 4292 31359
rect 4614 31356 4620 31368
rect 4672 31356 4678 31408
rect 17678 31396 17684 31408
rect 17639 31368 17684 31396
rect 17678 31356 17684 31368
rect 17736 31356 17742 31408
rect 21910 31396 21916 31408
rect 21823 31368 21916 31396
rect 5166 31328 5172 31340
rect 5127 31300 5172 31328
rect 5166 31288 5172 31300
rect 5224 31288 5230 31340
rect 5258 31288 5264 31340
rect 5316 31328 5322 31340
rect 5316 31300 5361 31328
rect 5316 31288 5322 31300
rect 8846 31288 8852 31340
rect 8904 31328 8910 31340
rect 9953 31331 10011 31337
rect 9953 31328 9965 31331
rect 8904 31300 9965 31328
rect 8904 31288 8910 31300
rect 9953 31297 9965 31300
rect 9999 31328 10011 31331
rect 10410 31328 10416 31340
rect 9999 31300 10416 31328
rect 9999 31297 10011 31300
rect 9953 31291 10011 31297
rect 10410 31288 10416 31300
rect 10468 31288 10474 31340
rect 20990 31288 20996 31340
rect 21048 31328 21054 31340
rect 21836 31337 21864 31368
rect 21910 31356 21916 31368
rect 21968 31396 21974 31408
rect 22189 31399 22247 31405
rect 22189 31396 22201 31399
rect 21968 31368 22201 31396
rect 21968 31356 21974 31368
rect 22189 31365 22201 31368
rect 22235 31365 22247 31399
rect 22189 31359 22247 31365
rect 21821 31331 21879 31337
rect 21048 31300 21772 31328
rect 21048 31288 21054 31300
rect 5074 31260 5080 31272
rect 5035 31232 5080 31260
rect 5074 31220 5080 31232
rect 5132 31220 5138 31272
rect 7745 31263 7803 31269
rect 7745 31229 7757 31263
rect 7791 31260 7803 31263
rect 8018 31260 8024 31272
rect 7791 31232 8024 31260
rect 7791 31229 7803 31232
rect 7745 31223 7803 31229
rect 8018 31220 8024 31232
rect 8076 31260 8082 31272
rect 8297 31263 8355 31269
rect 8297 31260 8309 31263
rect 8076 31232 8309 31260
rect 8076 31220 8082 31232
rect 8297 31229 8309 31232
rect 8343 31229 8355 31263
rect 8297 31223 8355 31229
rect 12437 31263 12495 31269
rect 12437 31229 12449 31263
rect 12483 31260 12495 31263
rect 13170 31260 13176 31272
rect 12483 31232 13176 31260
rect 12483 31229 12495 31232
rect 12437 31223 12495 31229
rect 13170 31220 13176 31232
rect 13228 31220 13234 31272
rect 13633 31263 13691 31269
rect 13633 31229 13645 31263
rect 13679 31260 13691 31263
rect 14274 31260 14280 31272
rect 13679 31232 14280 31260
rect 13679 31229 13691 31232
rect 13633 31223 13691 31229
rect 14274 31220 14280 31232
rect 14332 31220 14338 31272
rect 14829 31263 14887 31269
rect 14829 31229 14841 31263
rect 14875 31260 14887 31263
rect 15289 31263 15347 31269
rect 15289 31260 15301 31263
rect 14875 31232 15301 31260
rect 14875 31229 14887 31232
rect 14829 31223 14887 31229
rect 15289 31229 15301 31232
rect 15335 31260 15347 31263
rect 21542 31260 21548 31272
rect 15335 31232 16252 31260
rect 15335 31229 15347 31232
rect 15289 31223 15347 31229
rect 16224 31204 16252 31232
rect 20640 31232 21548 31260
rect 2924 31164 4292 31192
rect 9217 31195 9275 31201
rect 2924 31152 2930 31164
rect 9217 31161 9229 31195
rect 9263 31192 9275 31195
rect 9769 31195 9827 31201
rect 9769 31192 9781 31195
rect 9263 31164 9781 31192
rect 9263 31161 9275 31164
rect 9217 31155 9275 31161
rect 9769 31161 9781 31164
rect 9815 31192 9827 31195
rect 9950 31192 9956 31204
rect 9815 31164 9956 31192
rect 9815 31161 9827 31164
rect 9769 31155 9827 31161
rect 9950 31152 9956 31164
rect 10008 31152 10014 31204
rect 12621 31195 12679 31201
rect 12621 31161 12633 31195
rect 12667 31161 12679 31195
rect 12621 31155 12679 31161
rect 15197 31195 15255 31201
rect 15197 31161 15209 31195
rect 15243 31192 15255 31195
rect 15470 31192 15476 31204
rect 15243 31164 15476 31192
rect 15243 31161 15255 31164
rect 15197 31155 15255 31161
rect 1670 31124 1676 31136
rect 1631 31096 1676 31124
rect 1670 31084 1676 31096
rect 1728 31084 1734 31136
rect 4706 31124 4712 31136
rect 4667 31096 4712 31124
rect 4706 31084 4712 31096
rect 4764 31084 4770 31136
rect 5810 31124 5816 31136
rect 5771 31096 5816 31124
rect 5810 31084 5816 31096
rect 5868 31084 5874 31136
rect 6178 31084 6184 31136
rect 6236 31124 6242 31136
rect 6273 31127 6331 31133
rect 6273 31124 6285 31127
rect 6236 31096 6285 31124
rect 6236 31084 6242 31096
rect 6273 31093 6285 31096
rect 6319 31124 6331 31127
rect 6822 31124 6828 31136
rect 6319 31096 6828 31124
rect 6319 31093 6331 31096
rect 6273 31087 6331 31093
rect 6822 31084 6828 31096
rect 6880 31084 6886 31136
rect 8662 31084 8668 31136
rect 8720 31124 8726 31136
rect 9309 31127 9367 31133
rect 9309 31124 9321 31127
rect 8720 31096 9321 31124
rect 8720 31084 8726 31096
rect 9309 31093 9321 31096
rect 9355 31093 9367 31127
rect 9674 31124 9680 31136
rect 9635 31096 9680 31124
rect 9309 31087 9367 31093
rect 9674 31084 9680 31096
rect 9732 31084 9738 31136
rect 10410 31124 10416 31136
rect 10371 31096 10416 31124
rect 10410 31084 10416 31096
rect 10468 31084 10474 31136
rect 12250 31124 12256 31136
rect 12211 31096 12256 31124
rect 12250 31084 12256 31096
rect 12308 31124 12314 31136
rect 12636 31124 12664 31155
rect 15470 31152 15476 31164
rect 15528 31201 15534 31204
rect 15528 31195 15592 31201
rect 15528 31161 15546 31195
rect 15580 31161 15592 31195
rect 15528 31155 15592 31161
rect 15528 31152 15534 31155
rect 16206 31152 16212 31204
rect 16264 31152 16270 31204
rect 20640 31201 20668 31232
rect 21542 31220 21548 31232
rect 21600 31220 21606 31272
rect 21744 31260 21772 31300
rect 21821 31297 21833 31331
rect 21867 31297 21879 31331
rect 22557 31331 22615 31337
rect 22557 31328 22569 31331
rect 21821 31291 21879 31297
rect 21928 31300 22569 31328
rect 21928 31260 21956 31300
rect 22557 31297 22569 31300
rect 22603 31328 22615 31331
rect 24026 31328 24032 31340
rect 22603 31300 24032 31328
rect 22603 31297 22615 31300
rect 22557 31291 22615 31297
rect 24026 31288 24032 31300
rect 24084 31288 24090 31340
rect 24581 31331 24639 31337
rect 24581 31297 24593 31331
rect 24627 31328 24639 31331
rect 28166 31328 28172 31340
rect 24627 31300 24808 31328
rect 28127 31300 28172 31328
rect 24627 31297 24639 31300
rect 24581 31291 24639 31297
rect 21744 31232 21956 31260
rect 24044 31260 24072 31288
rect 24673 31263 24731 31269
rect 24673 31260 24685 31263
rect 24044 31232 24685 31260
rect 24673 31229 24685 31232
rect 24719 31229 24731 31263
rect 24780 31260 24808 31300
rect 28166 31288 28172 31300
rect 28224 31288 28230 31340
rect 24940 31263 24998 31269
rect 24940 31260 24952 31263
rect 24780 31232 24952 31260
rect 24673 31223 24731 31229
rect 24940 31229 24952 31232
rect 24986 31260 24998 31263
rect 27062 31260 27068 31272
rect 24986 31232 27068 31260
rect 24986 31229 24998 31232
rect 24940 31223 24998 31229
rect 27062 31220 27068 31232
rect 27120 31220 27126 31272
rect 20349 31195 20407 31201
rect 20349 31161 20361 31195
rect 20395 31192 20407 31195
rect 20625 31195 20683 31201
rect 20625 31192 20637 31195
rect 20395 31164 20637 31192
rect 20395 31161 20407 31164
rect 20349 31155 20407 31161
rect 20625 31161 20637 31164
rect 20671 31161 20683 31195
rect 21082 31192 21088 31204
rect 20995 31164 21088 31192
rect 20625 31155 20683 31161
rect 21082 31152 21088 31164
rect 21140 31192 21146 31204
rect 21637 31195 21695 31201
rect 21637 31192 21649 31195
rect 21140 31164 21649 31192
rect 21140 31152 21146 31164
rect 21637 31161 21649 31164
rect 21683 31161 21695 31195
rect 21637 31155 21695 31161
rect 27985 31195 28043 31201
rect 27985 31161 27997 31195
rect 28031 31192 28043 31195
rect 28031 31164 28764 31192
rect 28031 31161 28043 31164
rect 27985 31155 28043 31161
rect 28736 31136 28764 31164
rect 12308 31096 12664 31124
rect 12308 31084 12314 31096
rect 12710 31084 12716 31136
rect 12768 31124 12774 31136
rect 12805 31127 12863 31133
rect 12805 31124 12817 31127
rect 12768 31096 12817 31124
rect 12768 31084 12774 31096
rect 12805 31093 12817 31096
rect 12851 31093 12863 31127
rect 13814 31124 13820 31136
rect 13775 31096 13820 31124
rect 12805 31087 12863 31093
rect 13814 31084 13820 31096
rect 13872 31084 13878 31136
rect 16666 31124 16672 31136
rect 16627 31096 16672 31124
rect 16666 31084 16672 31096
rect 16724 31084 16730 31136
rect 17586 31084 17592 31136
rect 17644 31124 17650 31136
rect 18046 31124 18052 31136
rect 17644 31096 18052 31124
rect 17644 31084 17650 31096
rect 18046 31084 18052 31096
rect 18104 31124 18110 31136
rect 18233 31127 18291 31133
rect 18233 31124 18245 31127
rect 18104 31096 18245 31124
rect 18104 31084 18110 31096
rect 18233 31093 18245 31096
rect 18279 31093 18291 31127
rect 18233 31087 18291 31093
rect 25314 31084 25320 31136
rect 25372 31124 25378 31136
rect 26053 31127 26111 31133
rect 26053 31124 26065 31127
rect 25372 31096 26065 31124
rect 25372 31084 25378 31096
rect 26053 31093 26065 31096
rect 26099 31093 26111 31127
rect 26053 31087 26111 31093
rect 27525 31127 27583 31133
rect 27525 31093 27537 31127
rect 27571 31124 27583 31127
rect 28074 31124 28080 31136
rect 27571 31096 28080 31124
rect 27571 31093 27583 31096
rect 27525 31087 27583 31093
rect 28074 31084 28080 31096
rect 28132 31084 28138 31136
rect 28718 31124 28724 31136
rect 28679 31096 28724 31124
rect 28718 31084 28724 31096
rect 28776 31084 28782 31136
rect 28810 31084 28816 31136
rect 28868 31124 28874 31136
rect 28997 31127 29055 31133
rect 28997 31124 29009 31127
rect 28868 31096 29009 31124
rect 28868 31084 28874 31096
rect 28997 31093 29009 31096
rect 29043 31093 29055 31127
rect 28997 31087 29055 31093
rect 34698 31084 34704 31136
rect 34756 31124 34762 31136
rect 35434 31124 35440 31136
rect 34756 31096 35440 31124
rect 34756 31084 34762 31096
rect 35434 31084 35440 31096
rect 35492 31084 35498 31136
rect 1104 31034 38824 31056
rect 1104 30982 19606 31034
rect 19658 30982 19670 31034
rect 19722 30982 19734 31034
rect 19786 30982 19798 31034
rect 19850 30982 38824 31034
rect 1104 30960 38824 30982
rect 2866 30920 2872 30932
rect 2827 30892 2872 30920
rect 2866 30880 2872 30892
rect 2924 30880 2930 30932
rect 4341 30923 4399 30929
rect 4341 30889 4353 30923
rect 4387 30920 4399 30923
rect 4982 30920 4988 30932
rect 4387 30892 4988 30920
rect 4387 30889 4399 30892
rect 4341 30883 4399 30889
rect 4982 30880 4988 30892
rect 5040 30880 5046 30932
rect 5074 30880 5080 30932
rect 5132 30920 5138 30932
rect 5445 30923 5503 30929
rect 5445 30920 5457 30923
rect 5132 30892 5457 30920
rect 5132 30880 5138 30892
rect 5445 30889 5457 30892
rect 5491 30889 5503 30923
rect 5445 30883 5503 30889
rect 6181 30923 6239 30929
rect 6181 30889 6193 30923
rect 6227 30920 6239 30923
rect 6454 30920 6460 30932
rect 6227 30892 6460 30920
rect 6227 30889 6239 30892
rect 6181 30883 6239 30889
rect 6454 30880 6460 30892
rect 6512 30880 6518 30932
rect 9858 30920 9864 30932
rect 9819 30892 9864 30920
rect 9858 30880 9864 30892
rect 9916 30880 9922 30932
rect 14734 30920 14740 30932
rect 14695 30892 14740 30920
rect 14734 30880 14740 30892
rect 14792 30880 14798 30932
rect 15194 30880 15200 30932
rect 15252 30920 15258 30932
rect 15565 30923 15623 30929
rect 15565 30920 15577 30923
rect 15252 30892 15577 30920
rect 15252 30880 15258 30892
rect 15565 30889 15577 30892
rect 15611 30889 15623 30923
rect 15565 30883 15623 30889
rect 17678 30880 17684 30932
rect 17736 30920 17742 30932
rect 18966 30920 18972 30932
rect 17736 30892 18972 30920
rect 17736 30880 17742 30892
rect 18966 30880 18972 30892
rect 19024 30880 19030 30932
rect 21542 30880 21548 30932
rect 21600 30920 21606 30932
rect 22281 30923 22339 30929
rect 22281 30920 22293 30923
rect 21600 30892 22293 30920
rect 21600 30880 21606 30892
rect 22281 30889 22293 30892
rect 22327 30889 22339 30923
rect 22281 30883 22339 30889
rect 24026 30880 24032 30932
rect 24084 30920 24090 30932
rect 24121 30923 24179 30929
rect 24121 30920 24133 30923
rect 24084 30892 24133 30920
rect 24084 30880 24090 30892
rect 24121 30889 24133 30892
rect 24167 30889 24179 30923
rect 24121 30883 24179 30889
rect 4706 30812 4712 30864
rect 4764 30852 4770 30864
rect 13449 30855 13507 30861
rect 4764 30824 6040 30852
rect 4764 30812 4770 30824
rect 6012 30796 6040 30824
rect 13449 30821 13461 30855
rect 13495 30852 13507 30855
rect 13630 30852 13636 30864
rect 13495 30824 13636 30852
rect 13495 30821 13507 30824
rect 13449 30815 13507 30821
rect 13630 30812 13636 30824
rect 13688 30812 13694 30864
rect 21082 30812 21088 30864
rect 21140 30861 21146 30864
rect 21140 30855 21204 30861
rect 21140 30821 21158 30855
rect 21192 30821 21204 30855
rect 24136 30852 24164 30883
rect 24670 30880 24676 30932
rect 24728 30920 24734 30932
rect 25133 30923 25191 30929
rect 25133 30920 25145 30923
rect 24728 30892 25145 30920
rect 24728 30880 24734 30892
rect 25133 30889 25145 30892
rect 25179 30920 25191 30923
rect 26697 30923 26755 30929
rect 26697 30920 26709 30923
rect 25179 30892 26709 30920
rect 25179 30889 25191 30892
rect 25133 30883 25191 30889
rect 26697 30889 26709 30892
rect 26743 30889 26755 30923
rect 26697 30883 26755 30889
rect 28077 30923 28135 30929
rect 28077 30889 28089 30923
rect 28123 30920 28135 30923
rect 28166 30920 28172 30932
rect 28123 30892 28172 30920
rect 28123 30889 28135 30892
rect 28077 30883 28135 30889
rect 28166 30880 28172 30892
rect 28224 30880 28230 30932
rect 28718 30880 28724 30932
rect 28776 30920 28782 30932
rect 29733 30923 29791 30929
rect 29733 30920 29745 30923
rect 28776 30892 29745 30920
rect 28776 30880 28782 30892
rect 29733 30889 29745 30892
rect 29779 30889 29791 30923
rect 35618 30920 35624 30932
rect 35579 30892 35624 30920
rect 29733 30883 29791 30889
rect 35618 30880 35624 30892
rect 35676 30880 35682 30932
rect 25685 30855 25743 30861
rect 25685 30852 25697 30855
rect 24136 30824 25697 30852
rect 21140 30815 21204 30821
rect 25685 30821 25697 30824
rect 25731 30821 25743 30855
rect 25685 30815 25743 30821
rect 27709 30855 27767 30861
rect 27709 30821 27721 30855
rect 27755 30852 27767 30855
rect 28736 30852 28764 30880
rect 27755 30824 28764 30852
rect 27755 30821 27767 30824
rect 27709 30815 27767 30821
rect 21140 30812 21146 30815
rect 1756 30787 1814 30793
rect 1756 30753 1768 30787
rect 1802 30784 1814 30787
rect 2038 30784 2044 30796
rect 1802 30756 2044 30784
rect 1802 30753 1814 30756
rect 1756 30747 1814 30753
rect 2038 30744 2044 30756
rect 2096 30744 2102 30796
rect 4798 30784 4804 30796
rect 4759 30756 4804 30784
rect 4798 30744 4804 30756
rect 4856 30744 4862 30796
rect 5994 30784 6000 30796
rect 5907 30756 6000 30784
rect 5994 30744 6000 30756
rect 6052 30744 6058 30796
rect 8386 30784 8392 30796
rect 8347 30756 8392 30784
rect 8386 30744 8392 30756
rect 8444 30744 8450 30796
rect 9401 30787 9459 30793
rect 9401 30753 9413 30787
rect 9447 30784 9459 30787
rect 9674 30784 9680 30796
rect 9447 30756 9680 30784
rect 9447 30753 9459 30756
rect 9401 30747 9459 30753
rect 9674 30744 9680 30756
rect 9732 30784 9738 30796
rect 10594 30784 10600 30796
rect 9732 30756 10600 30784
rect 9732 30744 9738 30756
rect 10594 30744 10600 30756
rect 10652 30784 10658 30796
rect 10761 30787 10819 30793
rect 10761 30784 10773 30787
rect 10652 30756 10773 30784
rect 10652 30744 10658 30756
rect 10761 30753 10773 30756
rect 10807 30753 10819 30787
rect 10761 30747 10819 30753
rect 13357 30787 13415 30793
rect 13357 30753 13369 30787
rect 13403 30784 13415 30787
rect 13722 30784 13728 30796
rect 13403 30756 13728 30784
rect 13403 30753 13415 30756
rect 13357 30747 13415 30753
rect 13722 30744 13728 30756
rect 13780 30744 13786 30796
rect 15105 30787 15163 30793
rect 15105 30753 15117 30787
rect 15151 30784 15163 30787
rect 15930 30784 15936 30796
rect 15151 30756 15936 30784
rect 15151 30753 15163 30756
rect 15105 30747 15163 30753
rect 15930 30744 15936 30756
rect 15988 30744 15994 30796
rect 17865 30787 17923 30793
rect 17865 30784 17877 30787
rect 16040 30756 17877 30784
rect 16040 30728 16068 30756
rect 17865 30753 17877 30756
rect 17911 30753 17923 30787
rect 17865 30747 17923 30753
rect 20162 30744 20168 30796
rect 20220 30784 20226 30796
rect 20257 30787 20315 30793
rect 20257 30784 20269 30787
rect 20220 30756 20269 30784
rect 20220 30744 20226 30756
rect 20257 30753 20269 30756
rect 20303 30784 20315 30787
rect 20901 30787 20959 30793
rect 20901 30784 20913 30787
rect 20303 30756 20913 30784
rect 20303 30753 20315 30756
rect 20257 30747 20315 30753
rect 20901 30753 20913 30756
rect 20947 30784 20959 30787
rect 20990 30784 20996 30796
rect 20947 30756 20996 30784
rect 20947 30753 20959 30756
rect 20901 30747 20959 30753
rect 20990 30744 20996 30756
rect 21048 30744 21054 30796
rect 23474 30744 23480 30796
rect 23532 30784 23538 30796
rect 23569 30787 23627 30793
rect 23569 30784 23581 30787
rect 23532 30756 23581 30784
rect 23532 30744 23538 30756
rect 23569 30753 23581 30756
rect 23615 30784 23627 30787
rect 24210 30784 24216 30796
rect 23615 30756 24216 30784
rect 23615 30753 23627 30756
rect 23569 30747 23627 30753
rect 24210 30744 24216 30756
rect 24268 30744 24274 30796
rect 24578 30784 24584 30796
rect 24491 30756 24584 30784
rect 24578 30744 24584 30756
rect 24636 30784 24642 30796
rect 24762 30784 24768 30796
rect 24636 30756 24768 30784
rect 24636 30744 24642 30756
rect 24762 30744 24768 30756
rect 24820 30744 24826 30796
rect 25038 30784 25044 30796
rect 24999 30756 25044 30784
rect 25038 30744 25044 30756
rect 25096 30744 25102 30796
rect 26510 30784 26516 30796
rect 26471 30756 26516 30784
rect 26510 30744 26516 30756
rect 26568 30744 26574 30796
rect 28074 30744 28080 30796
rect 28132 30784 28138 30796
rect 28620 30787 28678 30793
rect 28620 30784 28632 30787
rect 28132 30756 28632 30784
rect 28132 30744 28138 30756
rect 28620 30753 28632 30756
rect 28666 30784 28678 30787
rect 28902 30784 28908 30796
rect 28666 30756 28908 30784
rect 28666 30753 28678 30756
rect 28620 30747 28678 30753
rect 28902 30744 28908 30756
rect 28960 30744 28966 30796
rect 35437 30787 35495 30793
rect 35437 30753 35449 30787
rect 35483 30784 35495 30787
rect 35526 30784 35532 30796
rect 35483 30756 35532 30784
rect 35483 30753 35495 30756
rect 35437 30747 35495 30753
rect 35526 30744 35532 30756
rect 35584 30744 35590 30796
rect 1394 30676 1400 30728
rect 1452 30716 1458 30728
rect 1489 30719 1547 30725
rect 1489 30716 1501 30719
rect 1452 30688 1501 30716
rect 1452 30676 1458 30688
rect 1489 30685 1501 30688
rect 1535 30685 1547 30719
rect 4890 30716 4896 30728
rect 4851 30688 4896 30716
rect 1489 30679 1547 30685
rect 4890 30676 4896 30688
rect 4948 30676 4954 30728
rect 4985 30719 5043 30725
rect 4985 30685 4997 30719
rect 5031 30716 5043 30719
rect 5258 30716 5264 30728
rect 5031 30688 5264 30716
rect 5031 30685 5043 30688
rect 4985 30679 5043 30685
rect 3970 30608 3976 30660
rect 4028 30648 4034 30660
rect 5000 30648 5028 30679
rect 5258 30676 5264 30688
rect 5316 30676 5322 30728
rect 8478 30716 8484 30728
rect 8439 30688 8484 30716
rect 8478 30676 8484 30688
rect 8536 30676 8542 30728
rect 8665 30719 8723 30725
rect 8665 30685 8677 30719
rect 8711 30716 8723 30719
rect 8846 30716 8852 30728
rect 8711 30688 8852 30716
rect 8711 30685 8723 30688
rect 8665 30679 8723 30685
rect 4028 30620 5028 30648
rect 7929 30651 7987 30657
rect 4028 30608 4034 30620
rect 7929 30617 7941 30651
rect 7975 30648 7987 30651
rect 8110 30648 8116 30660
rect 7975 30620 8116 30648
rect 7975 30617 7987 30620
rect 7929 30611 7987 30617
rect 8110 30608 8116 30620
rect 8168 30648 8174 30660
rect 8680 30648 8708 30679
rect 8846 30676 8852 30688
rect 8904 30676 8910 30728
rect 9582 30676 9588 30728
rect 9640 30716 9646 30728
rect 10502 30716 10508 30728
rect 9640 30688 10508 30716
rect 9640 30676 9646 30688
rect 10502 30676 10508 30688
rect 10560 30676 10566 30728
rect 13538 30676 13544 30728
rect 13596 30716 13602 30728
rect 16022 30716 16028 30728
rect 13596 30688 13641 30716
rect 15983 30688 16028 30716
rect 13596 30676 13602 30688
rect 16022 30676 16028 30688
rect 16080 30676 16086 30728
rect 16117 30719 16175 30725
rect 16117 30685 16129 30719
rect 16163 30716 16175 30719
rect 16666 30716 16672 30728
rect 16163 30688 16672 30716
rect 16163 30685 16175 30688
rect 16117 30679 16175 30685
rect 8168 30620 8708 30648
rect 8168 30608 8174 30620
rect 14918 30608 14924 30660
rect 14976 30648 14982 30660
rect 16132 30648 16160 30679
rect 16666 30676 16672 30688
rect 16724 30676 16730 30728
rect 16942 30676 16948 30728
rect 17000 30716 17006 30728
rect 17494 30725 17500 30728
rect 17129 30719 17187 30725
rect 17129 30716 17141 30719
rect 17000 30688 17141 30716
rect 17000 30676 17006 30688
rect 17129 30685 17141 30688
rect 17175 30685 17187 30719
rect 17129 30679 17187 30685
rect 17452 30719 17500 30725
rect 17452 30685 17464 30719
rect 17498 30685 17500 30719
rect 17452 30679 17500 30685
rect 14976 30620 16160 30648
rect 14976 30608 14982 30620
rect 4433 30583 4491 30589
rect 4433 30549 4445 30583
rect 4479 30580 4491 30583
rect 5350 30580 5356 30592
rect 4479 30552 5356 30580
rect 4479 30549 4491 30552
rect 4433 30543 4491 30549
rect 5350 30540 5356 30552
rect 5408 30540 5414 30592
rect 8018 30580 8024 30592
rect 7979 30552 8024 30580
rect 8018 30540 8024 30552
rect 8076 30540 8082 30592
rect 11885 30583 11943 30589
rect 11885 30549 11897 30583
rect 11931 30580 11943 30583
rect 12250 30580 12256 30592
rect 11931 30552 12256 30580
rect 11931 30549 11943 30552
rect 11885 30543 11943 30549
rect 12250 30540 12256 30552
rect 12308 30540 12314 30592
rect 12529 30583 12587 30589
rect 12529 30549 12541 30583
rect 12575 30580 12587 30583
rect 12618 30580 12624 30592
rect 12575 30552 12624 30580
rect 12575 30549 12587 30552
rect 12529 30543 12587 30549
rect 12618 30540 12624 30552
rect 12676 30540 12682 30592
rect 12802 30580 12808 30592
rect 12763 30552 12808 30580
rect 12802 30540 12808 30552
rect 12860 30540 12866 30592
rect 12986 30580 12992 30592
rect 12947 30552 12992 30580
rect 12986 30540 12992 30552
rect 13044 30540 13050 30592
rect 14642 30540 14648 30592
rect 14700 30580 14706 30592
rect 16114 30580 16120 30592
rect 14700 30552 16120 30580
rect 14700 30540 14706 30552
rect 16114 30540 16120 30552
rect 16172 30540 16178 30592
rect 17037 30583 17095 30589
rect 17037 30549 17049 30583
rect 17083 30580 17095 30583
rect 17144 30580 17172 30679
rect 17494 30676 17500 30679
rect 17552 30676 17558 30728
rect 17586 30676 17592 30728
rect 17644 30716 17650 30728
rect 25314 30716 25320 30728
rect 17644 30688 17689 30716
rect 25275 30688 25320 30716
rect 17644 30676 17650 30688
rect 25314 30676 25320 30688
rect 25372 30676 25378 30728
rect 28353 30719 28411 30725
rect 28353 30685 28365 30719
rect 28399 30685 28411 30719
rect 28353 30679 28411 30685
rect 17770 30580 17776 30592
rect 17083 30552 17776 30580
rect 17083 30549 17095 30552
rect 17037 30543 17095 30549
rect 17770 30540 17776 30552
rect 17828 30540 17834 30592
rect 23750 30580 23756 30592
rect 23711 30552 23756 30580
rect 23750 30540 23756 30552
rect 23808 30540 23814 30592
rect 24673 30583 24731 30589
rect 24673 30549 24685 30583
rect 24719 30580 24731 30583
rect 24762 30580 24768 30592
rect 24719 30552 24768 30580
rect 24719 30549 24731 30552
rect 24673 30543 24731 30549
rect 24762 30540 24768 30552
rect 24820 30540 24826 30592
rect 28368 30580 28396 30679
rect 28718 30580 28724 30592
rect 28368 30552 28724 30580
rect 28718 30540 28724 30552
rect 28776 30540 28782 30592
rect 1104 30490 38824 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 34966 30490
rect 35018 30438 35030 30490
rect 35082 30438 35094 30490
rect 35146 30438 35158 30490
rect 35210 30438 38824 30490
rect 1104 30416 38824 30438
rect 4617 30379 4675 30385
rect 4617 30345 4629 30379
rect 4663 30376 4675 30379
rect 4798 30376 4804 30388
rect 4663 30348 4804 30376
rect 4663 30345 4675 30348
rect 4617 30339 4675 30345
rect 3789 30311 3847 30317
rect 3789 30277 3801 30311
rect 3835 30308 3847 30311
rect 4632 30308 4660 30339
rect 4798 30336 4804 30348
rect 4856 30336 4862 30388
rect 5994 30376 6000 30388
rect 5955 30348 6000 30376
rect 5994 30336 6000 30348
rect 6052 30336 6058 30388
rect 6822 30336 6828 30388
rect 6880 30336 6886 30388
rect 8478 30376 8484 30388
rect 8312 30348 8484 30376
rect 3835 30280 4660 30308
rect 6840 30308 6868 30336
rect 7009 30311 7067 30317
rect 7009 30308 7021 30311
rect 6840 30280 7021 30308
rect 3835 30277 3847 30280
rect 3789 30271 3847 30277
rect 7009 30277 7021 30280
rect 7055 30277 7067 30311
rect 7009 30271 7067 30277
rect 8113 30311 8171 30317
rect 8113 30277 8125 30311
rect 8159 30308 8171 30311
rect 8202 30308 8208 30320
rect 8159 30280 8208 30308
rect 8159 30277 8171 30280
rect 8113 30271 8171 30277
rect 8202 30268 8208 30280
rect 8260 30308 8266 30320
rect 8312 30308 8340 30348
rect 8478 30336 8484 30348
rect 8536 30336 8542 30388
rect 9950 30376 9956 30388
rect 9911 30348 9956 30376
rect 9950 30336 9956 30348
rect 10008 30336 10014 30388
rect 14642 30336 14648 30388
rect 14700 30376 14706 30388
rect 14737 30379 14795 30385
rect 14737 30376 14749 30379
rect 14700 30348 14749 30376
rect 14700 30336 14706 30348
rect 14737 30345 14749 30348
rect 14783 30345 14795 30379
rect 14737 30339 14795 30345
rect 15197 30379 15255 30385
rect 15197 30345 15209 30379
rect 15243 30376 15255 30379
rect 15654 30376 15660 30388
rect 15243 30348 15660 30376
rect 15243 30345 15255 30348
rect 15197 30339 15255 30345
rect 15654 30336 15660 30348
rect 15712 30376 15718 30388
rect 15838 30376 15844 30388
rect 15712 30348 15844 30376
rect 15712 30336 15718 30348
rect 15838 30336 15844 30348
rect 15896 30376 15902 30388
rect 17494 30376 17500 30388
rect 15896 30348 17500 30376
rect 15896 30336 15902 30348
rect 17494 30336 17500 30348
rect 17552 30336 17558 30388
rect 21082 30336 21088 30388
rect 21140 30376 21146 30388
rect 21545 30379 21603 30385
rect 21545 30376 21557 30379
rect 21140 30348 21557 30376
rect 21140 30336 21146 30348
rect 21545 30345 21557 30348
rect 21591 30345 21603 30379
rect 23474 30376 23480 30388
rect 23435 30348 23480 30376
rect 21545 30339 21603 30345
rect 23474 30336 23480 30348
rect 23532 30336 23538 30388
rect 23750 30336 23756 30388
rect 23808 30376 23814 30388
rect 24489 30379 24547 30385
rect 24489 30376 24501 30379
rect 23808 30348 24501 30376
rect 23808 30336 23814 30348
rect 24489 30345 24501 30348
rect 24535 30376 24547 30379
rect 25038 30376 25044 30388
rect 24535 30348 25044 30376
rect 24535 30345 24547 30348
rect 24489 30339 24547 30345
rect 25038 30336 25044 30348
rect 25096 30336 25102 30388
rect 26510 30336 26516 30388
rect 26568 30376 26574 30388
rect 26605 30379 26663 30385
rect 26605 30376 26617 30379
rect 26568 30348 26617 30376
rect 26568 30336 26574 30348
rect 26605 30345 26617 30348
rect 26651 30345 26663 30379
rect 26605 30339 26663 30345
rect 28074 30336 28080 30388
rect 28132 30376 28138 30388
rect 28353 30379 28411 30385
rect 28353 30376 28365 30379
rect 28132 30348 28365 30376
rect 28132 30336 28138 30348
rect 28353 30345 28365 30348
rect 28399 30345 28411 30379
rect 28353 30339 28411 30345
rect 8260 30280 8340 30308
rect 24213 30311 24271 30317
rect 8260 30268 8266 30280
rect 24213 30277 24225 30311
rect 24259 30308 24271 30311
rect 24670 30308 24676 30320
rect 24259 30280 24676 30308
rect 24259 30277 24271 30280
rect 24213 30271 24271 30277
rect 24670 30268 24676 30280
rect 24728 30268 24734 30320
rect 34606 30268 34612 30320
rect 34664 30308 34670 30320
rect 35342 30308 35348 30320
rect 34664 30280 35348 30308
rect 34664 30268 34670 30280
rect 35342 30268 35348 30280
rect 35400 30268 35406 30320
rect 35621 30311 35679 30317
rect 35621 30277 35633 30311
rect 35667 30308 35679 30311
rect 35710 30308 35716 30320
rect 35667 30280 35716 30308
rect 35667 30277 35679 30280
rect 35621 30271 35679 30277
rect 35710 30268 35716 30280
rect 35768 30268 35774 30320
rect 4982 30200 4988 30252
rect 5040 30240 5046 30252
rect 5169 30243 5227 30249
rect 5169 30240 5181 30243
rect 5040 30212 5181 30240
rect 5040 30200 5046 30212
rect 5169 30209 5181 30212
rect 5215 30240 5227 30243
rect 5350 30240 5356 30252
rect 5215 30212 5356 30240
rect 5215 30209 5227 30212
rect 5169 30203 5227 30209
rect 5350 30200 5356 30212
rect 5408 30240 5414 30252
rect 5629 30243 5687 30249
rect 5629 30240 5641 30243
rect 5408 30212 5641 30240
rect 5408 30200 5414 30212
rect 5629 30209 5641 30212
rect 5675 30209 5687 30243
rect 8570 30240 8576 30252
rect 8531 30212 8576 30240
rect 5629 30203 5687 30209
rect 8570 30200 8576 30212
rect 8628 30200 8634 30252
rect 11882 30240 11888 30252
rect 11256 30212 11888 30240
rect 1394 30172 1400 30184
rect 1355 30144 1400 30172
rect 1394 30132 1400 30144
rect 1452 30132 1458 30184
rect 5534 30132 5540 30184
rect 5592 30172 5598 30184
rect 11256 30181 11284 30212
rect 11882 30200 11888 30212
rect 11940 30200 11946 30252
rect 12802 30200 12808 30252
rect 12860 30240 12866 30252
rect 12989 30243 13047 30249
rect 12989 30240 13001 30243
rect 12860 30212 13001 30240
rect 12860 30200 12866 30212
rect 12989 30209 13001 30212
rect 13035 30209 13047 30243
rect 12989 30203 13047 30209
rect 15746 30200 15752 30252
rect 15804 30249 15810 30252
rect 15804 30243 15826 30249
rect 15814 30209 15826 30243
rect 15804 30203 15826 30209
rect 16025 30243 16083 30249
rect 16025 30209 16037 30243
rect 16071 30240 16083 30243
rect 16114 30240 16120 30252
rect 16071 30212 16120 30240
rect 16071 30209 16083 30212
rect 16025 30203 16083 30209
rect 15804 30200 15810 30203
rect 16114 30200 16120 30212
rect 16172 30240 16178 30252
rect 17773 30243 17831 30249
rect 17773 30240 17785 30243
rect 16172 30212 17785 30240
rect 16172 30200 16178 30212
rect 17773 30209 17785 30212
rect 17819 30209 17831 30243
rect 18506 30240 18512 30252
rect 18467 30212 18512 30240
rect 17773 30203 17831 30209
rect 6825 30175 6883 30181
rect 6825 30172 6837 30175
rect 5592 30144 6837 30172
rect 5592 30132 5598 30144
rect 6825 30141 6837 30144
rect 6871 30172 6883 30175
rect 7377 30175 7435 30181
rect 7377 30172 7389 30175
rect 6871 30144 7389 30172
rect 6871 30141 6883 30144
rect 6825 30135 6883 30141
rect 7377 30141 7389 30144
rect 7423 30141 7435 30175
rect 7377 30135 7435 30141
rect 11241 30175 11299 30181
rect 11241 30141 11253 30175
rect 11287 30141 11299 30175
rect 14182 30172 14188 30184
rect 11241 30135 11299 30141
rect 13004 30144 14188 30172
rect 1670 30113 1676 30116
rect 1664 30104 1676 30113
rect 1631 30076 1676 30104
rect 1664 30067 1676 30076
rect 1670 30064 1676 30067
rect 1728 30064 1734 30116
rect 4525 30107 4583 30113
rect 4525 30073 4537 30107
rect 4571 30104 4583 30107
rect 5074 30104 5080 30116
rect 4571 30076 5080 30104
rect 4571 30073 4583 30076
rect 4525 30067 4583 30073
rect 5074 30064 5080 30076
rect 5132 30064 5138 30116
rect 7926 30064 7932 30116
rect 7984 30104 7990 30116
rect 8386 30104 8392 30116
rect 7984 30076 8392 30104
rect 7984 30064 7990 30076
rect 8386 30064 8392 30076
rect 8444 30104 8450 30116
rect 8481 30107 8539 30113
rect 8481 30104 8493 30107
rect 8444 30076 8493 30104
rect 8444 30064 8450 30076
rect 8481 30073 8493 30076
rect 8527 30104 8539 30107
rect 8840 30107 8898 30113
rect 8840 30104 8852 30107
rect 8527 30076 8852 30104
rect 8527 30073 8539 30076
rect 8481 30067 8539 30073
rect 8840 30073 8852 30076
rect 8886 30104 8898 30107
rect 9306 30104 9312 30116
rect 8886 30076 9312 30104
rect 8886 30073 8898 30076
rect 8840 30067 8898 30073
rect 9306 30064 9312 30076
rect 9364 30064 9370 30116
rect 10502 30064 10508 30116
rect 10560 30104 10566 30116
rect 10965 30107 11023 30113
rect 10965 30104 10977 30107
rect 10560 30076 10977 30104
rect 10560 30064 10566 30076
rect 10965 30073 10977 30076
rect 11011 30104 11023 30107
rect 12066 30104 12072 30116
rect 11011 30076 12072 30104
rect 11011 30073 11023 30076
rect 10965 30067 11023 30073
rect 12066 30064 12072 30076
rect 12124 30064 12130 30116
rect 12897 30107 12955 30113
rect 12897 30104 12909 30107
rect 12360 30076 12909 30104
rect 12360 30048 12388 30076
rect 12897 30073 12909 30076
rect 12943 30073 12955 30107
rect 12897 30067 12955 30073
rect 2038 29996 2044 30048
rect 2096 30036 2102 30048
rect 2777 30039 2835 30045
rect 2777 30036 2789 30039
rect 2096 30008 2789 30036
rect 2096 29996 2102 30008
rect 2777 30005 2789 30008
rect 2823 30005 2835 30039
rect 2777 29999 2835 30005
rect 2958 29996 2964 30048
rect 3016 30036 3022 30048
rect 3329 30039 3387 30045
rect 3329 30036 3341 30039
rect 3016 30008 3341 30036
rect 3016 29996 3022 30008
rect 3329 30005 3341 30008
rect 3375 30036 3387 30039
rect 3970 30036 3976 30048
rect 3375 30008 3976 30036
rect 3375 30005 3387 30008
rect 3329 29999 3387 30005
rect 3970 29996 3976 30008
rect 4028 29996 4034 30048
rect 4154 30036 4160 30048
rect 4115 30008 4160 30036
rect 4154 29996 4160 30008
rect 4212 30036 4218 30048
rect 4985 30039 5043 30045
rect 4985 30036 4997 30039
rect 4212 30008 4997 30036
rect 4212 29996 4218 30008
rect 4985 30005 4997 30008
rect 5031 30036 5043 30039
rect 5534 30036 5540 30048
rect 5031 30008 5540 30036
rect 5031 30005 5043 30008
rect 4985 29999 5043 30005
rect 5534 29996 5540 30008
rect 5592 29996 5598 30048
rect 10594 30036 10600 30048
rect 10555 30008 10600 30036
rect 10594 29996 10600 30008
rect 10652 29996 10658 30048
rect 11330 29996 11336 30048
rect 11388 30036 11394 30048
rect 11425 30039 11483 30045
rect 11425 30036 11437 30039
rect 11388 30008 11437 30036
rect 11388 29996 11394 30008
rect 11425 30005 11437 30008
rect 11471 30005 11483 30039
rect 11425 29999 11483 30005
rect 12253 30039 12311 30045
rect 12253 30005 12265 30039
rect 12299 30036 12311 30039
rect 12342 30036 12348 30048
rect 12299 30008 12348 30036
rect 12299 30005 12311 30008
rect 12253 29999 12311 30005
rect 12342 29996 12348 30008
rect 12400 29996 12406 30048
rect 12434 29996 12440 30048
rect 12492 30036 12498 30048
rect 12492 30008 12537 30036
rect 12492 29996 12498 30008
rect 12618 29996 12624 30048
rect 12676 30036 12682 30048
rect 12805 30039 12863 30045
rect 12805 30036 12817 30039
rect 12676 30008 12817 30036
rect 12676 29996 12682 30008
rect 12805 30005 12817 30008
rect 12851 30036 12863 30039
rect 13004 30036 13032 30144
rect 14182 30132 14188 30144
rect 14240 30132 14246 30184
rect 15286 30172 15292 30184
rect 15247 30144 15292 30172
rect 15286 30132 15292 30144
rect 15344 30132 15350 30184
rect 17788 30172 17816 30203
rect 18506 30200 18512 30212
rect 18564 30200 18570 30252
rect 18690 30240 18696 30252
rect 18603 30212 18696 30240
rect 18690 30200 18696 30212
rect 18748 30240 18754 30252
rect 19242 30240 19248 30252
rect 18748 30212 19248 30240
rect 18748 30200 18754 30212
rect 19242 30200 19248 30212
rect 19300 30200 19306 30252
rect 20162 30240 20168 30252
rect 20123 30212 20168 30240
rect 20162 30200 20168 30212
rect 20220 30200 20226 30252
rect 18417 30175 18475 30181
rect 18417 30172 18429 30175
rect 17788 30144 18429 30172
rect 18417 30141 18429 30144
rect 18463 30141 18475 30175
rect 18524 30172 18552 30200
rect 19061 30175 19119 30181
rect 19061 30172 19073 30175
rect 18524 30144 19073 30172
rect 18417 30135 18475 30141
rect 19061 30141 19073 30144
rect 19107 30141 19119 30175
rect 19061 30135 19119 30141
rect 24026 30132 24032 30184
rect 24084 30172 24090 30184
rect 24673 30175 24731 30181
rect 24673 30172 24685 30175
rect 24084 30144 24685 30172
rect 24084 30132 24090 30144
rect 24673 30141 24685 30144
rect 24719 30141 24731 30175
rect 24673 30135 24731 30141
rect 24940 30175 24998 30181
rect 24940 30141 24952 30175
rect 24986 30172 24998 30175
rect 25314 30172 25320 30184
rect 24986 30144 25320 30172
rect 24986 30141 24998 30144
rect 24940 30135 24998 30141
rect 25314 30132 25320 30144
rect 25372 30132 25378 30184
rect 35342 30132 35348 30184
rect 35400 30172 35406 30184
rect 35437 30175 35495 30181
rect 35437 30172 35449 30175
rect 35400 30144 35449 30172
rect 35400 30132 35406 30144
rect 35437 30141 35449 30144
rect 35483 30172 35495 30175
rect 35989 30175 36047 30181
rect 35989 30172 36001 30175
rect 35483 30144 36001 30172
rect 35483 30141 35495 30144
rect 35437 30135 35495 30141
rect 35989 30141 36001 30144
rect 36035 30141 36047 30175
rect 35989 30135 36047 30141
rect 13630 30064 13636 30116
rect 13688 30104 13694 30116
rect 13817 30107 13875 30113
rect 13817 30104 13829 30107
rect 13688 30076 13829 30104
rect 13688 30064 13694 30076
rect 13817 30073 13829 30076
rect 13863 30073 13875 30107
rect 17494 30104 17500 30116
rect 17407 30076 17500 30104
rect 13817 30067 13875 30073
rect 17494 30064 17500 30076
rect 17552 30104 17558 30116
rect 17954 30104 17960 30116
rect 17552 30076 17960 30104
rect 17552 30064 17558 30076
rect 17954 30064 17960 30076
rect 18012 30064 18018 30116
rect 20410 30107 20468 30113
rect 20410 30104 20422 30107
rect 19996 30076 20422 30104
rect 19996 30048 20024 30076
rect 20410 30073 20422 30076
rect 20456 30073 20468 30107
rect 20410 30067 20468 30073
rect 12851 30008 13032 30036
rect 13541 30039 13599 30045
rect 12851 30005 12863 30008
rect 12805 29999 12863 30005
rect 13541 30005 13553 30039
rect 13587 30036 13599 30039
rect 13722 30036 13728 30048
rect 13587 30008 13728 30036
rect 13587 30005 13599 30008
rect 13541 29999 13599 30005
rect 13722 29996 13728 30008
rect 13780 29996 13786 30048
rect 14366 30036 14372 30048
rect 14327 30008 14372 30036
rect 14366 29996 14372 30008
rect 14424 29996 14430 30048
rect 15654 29996 15660 30048
rect 15712 30036 15718 30048
rect 15755 30039 15813 30045
rect 15755 30036 15767 30039
rect 15712 30008 15767 30036
rect 15712 29996 15718 30008
rect 15755 30005 15767 30008
rect 15801 30005 15813 30039
rect 15755 29999 15813 30005
rect 16022 29996 16028 30048
rect 16080 30036 16086 30048
rect 17126 30036 17132 30048
rect 16080 30008 17132 30036
rect 16080 29996 16086 30008
rect 17126 29996 17132 30008
rect 17184 29996 17190 30048
rect 18046 30036 18052 30048
rect 18007 30008 18052 30036
rect 18046 29996 18052 30008
rect 18104 29996 18110 30048
rect 19978 30036 19984 30048
rect 19939 30008 19984 30036
rect 19978 29996 19984 30008
rect 20036 29996 20042 30048
rect 25774 29996 25780 30048
rect 25832 30036 25838 30048
rect 26053 30039 26111 30045
rect 26053 30036 26065 30039
rect 25832 30008 26065 30036
rect 25832 29996 25838 30008
rect 26053 30005 26065 30008
rect 26099 30005 26111 30039
rect 28718 30036 28724 30048
rect 28679 30008 28724 30036
rect 26053 29999 26111 30005
rect 28718 29996 28724 30008
rect 28776 29996 28782 30048
rect 35345 30039 35403 30045
rect 35345 30005 35357 30039
rect 35391 30036 35403 30039
rect 35526 30036 35532 30048
rect 35391 30008 35532 30036
rect 35391 30005 35403 30008
rect 35345 29999 35403 30005
rect 35526 29996 35532 30008
rect 35584 29996 35590 30048
rect 1104 29946 38824 29968
rect 1104 29894 19606 29946
rect 19658 29894 19670 29946
rect 19722 29894 19734 29946
rect 19786 29894 19798 29946
rect 19850 29894 38824 29946
rect 1104 29872 38824 29894
rect 1670 29792 1676 29844
rect 1728 29832 1734 29844
rect 2777 29835 2835 29841
rect 2777 29832 2789 29835
rect 1728 29804 2789 29832
rect 1728 29792 1734 29804
rect 2777 29801 2789 29804
rect 2823 29801 2835 29835
rect 2777 29795 2835 29801
rect 4525 29835 4583 29841
rect 4525 29801 4537 29835
rect 4571 29832 4583 29835
rect 4890 29832 4896 29844
rect 4571 29804 4896 29832
rect 4571 29801 4583 29804
rect 4525 29795 4583 29801
rect 4890 29792 4896 29804
rect 4948 29792 4954 29844
rect 5534 29792 5540 29844
rect 5592 29832 5598 29844
rect 6089 29835 6147 29841
rect 6089 29832 6101 29835
rect 5592 29804 6101 29832
rect 5592 29792 5598 29804
rect 6089 29801 6101 29804
rect 6135 29801 6147 29835
rect 7926 29832 7932 29844
rect 7887 29804 7932 29832
rect 6089 29795 6147 29801
rect 7926 29792 7932 29804
rect 7984 29792 7990 29844
rect 8570 29792 8576 29844
rect 8628 29832 8634 29844
rect 9033 29835 9091 29841
rect 9033 29832 9045 29835
rect 8628 29804 9045 29832
rect 8628 29792 8634 29804
rect 9033 29801 9045 29804
rect 9079 29801 9091 29835
rect 9033 29795 9091 29801
rect 10594 29792 10600 29844
rect 10652 29832 10658 29844
rect 11057 29835 11115 29841
rect 11057 29832 11069 29835
rect 10652 29804 11069 29832
rect 10652 29792 10658 29804
rect 11057 29801 11069 29804
rect 11103 29801 11115 29835
rect 13538 29832 13544 29844
rect 13499 29804 13544 29832
rect 11057 29795 11115 29801
rect 13538 29792 13544 29804
rect 13596 29792 13602 29844
rect 14182 29832 14188 29844
rect 14143 29804 14188 29832
rect 14182 29792 14188 29804
rect 14240 29792 14246 29844
rect 14737 29835 14795 29841
rect 14737 29801 14749 29835
rect 14783 29832 14795 29835
rect 14918 29832 14924 29844
rect 14783 29804 14924 29832
rect 14783 29801 14795 29804
rect 14737 29795 14795 29801
rect 14918 29792 14924 29804
rect 14976 29792 14982 29844
rect 15565 29835 15623 29841
rect 15565 29801 15577 29835
rect 15611 29832 15623 29835
rect 16022 29832 16028 29844
rect 15611 29804 16028 29832
rect 15611 29801 15623 29804
rect 15565 29795 15623 29801
rect 16022 29792 16028 29804
rect 16080 29792 16086 29844
rect 17126 29792 17132 29844
rect 17184 29832 17190 29844
rect 17957 29835 18015 29841
rect 17957 29832 17969 29835
rect 17184 29804 17969 29832
rect 17184 29792 17190 29804
rect 17957 29801 17969 29804
rect 18003 29801 18015 29835
rect 18690 29832 18696 29844
rect 18651 29804 18696 29832
rect 17957 29795 18015 29801
rect 18690 29792 18696 29804
rect 18748 29792 18754 29844
rect 21082 29832 21088 29844
rect 21043 29804 21088 29832
rect 21082 29792 21088 29804
rect 21140 29792 21146 29844
rect 23753 29835 23811 29841
rect 23753 29801 23765 29835
rect 23799 29832 23811 29835
rect 24118 29832 24124 29844
rect 23799 29804 24124 29832
rect 23799 29801 23811 29804
rect 23753 29795 23811 29801
rect 24118 29792 24124 29804
rect 24176 29792 24182 29844
rect 24213 29835 24271 29841
rect 24213 29801 24225 29835
rect 24259 29832 24271 29835
rect 24581 29835 24639 29841
rect 24581 29832 24593 29835
rect 24259 29804 24593 29832
rect 24259 29801 24271 29804
rect 24213 29795 24271 29801
rect 24581 29801 24593 29804
rect 24627 29832 24639 29835
rect 25314 29832 25320 29844
rect 24627 29804 25320 29832
rect 24627 29801 24639 29804
rect 24581 29795 24639 29801
rect 25314 29792 25320 29804
rect 25372 29792 25378 29844
rect 25774 29832 25780 29844
rect 25735 29804 25780 29832
rect 25774 29792 25780 29804
rect 25832 29792 25838 29844
rect 35618 29832 35624 29844
rect 35579 29804 35624 29832
rect 35618 29792 35624 29804
rect 35676 29792 35682 29844
rect 4976 29767 5034 29773
rect 4976 29733 4988 29767
rect 5022 29764 5034 29767
rect 5074 29764 5080 29776
rect 5022 29736 5080 29764
rect 5022 29733 5034 29736
rect 4976 29727 5034 29733
rect 5074 29724 5080 29736
rect 5132 29724 5138 29776
rect 7098 29724 7104 29776
rect 7156 29764 7162 29776
rect 8389 29767 8447 29773
rect 8389 29764 8401 29767
rect 7156 29736 8401 29764
rect 7156 29724 7162 29736
rect 8389 29733 8401 29736
rect 8435 29764 8447 29767
rect 8662 29764 8668 29776
rect 8435 29736 8668 29764
rect 8435 29733 8447 29736
rect 8389 29727 8447 29733
rect 8662 29724 8668 29736
rect 8720 29724 8726 29776
rect 9950 29773 9956 29776
rect 9944 29764 9956 29773
rect 9911 29736 9956 29764
rect 9944 29727 9956 29736
rect 9950 29724 9956 29727
rect 10008 29724 10014 29776
rect 14366 29724 14372 29776
rect 14424 29764 14430 29776
rect 17586 29764 17592 29776
rect 14424 29736 17592 29764
rect 14424 29724 14430 29736
rect 17586 29724 17592 29736
rect 17644 29724 17650 29776
rect 20990 29724 20996 29776
rect 21048 29764 21054 29776
rect 21453 29767 21511 29773
rect 21453 29764 21465 29767
rect 21048 29736 21465 29764
rect 21048 29724 21054 29736
rect 21453 29733 21465 29736
rect 21499 29733 21511 29767
rect 21453 29727 21511 29733
rect 32484 29767 32542 29773
rect 32484 29733 32496 29767
rect 32530 29764 32542 29767
rect 32674 29764 32680 29776
rect 32530 29736 32680 29764
rect 32530 29733 32542 29736
rect 32484 29727 32542 29733
rect 32674 29724 32680 29736
rect 32732 29724 32738 29776
rect 1670 29705 1676 29708
rect 1664 29696 1676 29705
rect 1631 29668 1676 29696
rect 1664 29659 1676 29668
rect 1670 29656 1676 29659
rect 1728 29656 1734 29708
rect 3421 29699 3479 29705
rect 3421 29665 3433 29699
rect 3467 29696 3479 29699
rect 3881 29699 3939 29705
rect 3881 29696 3893 29699
rect 3467 29668 3893 29696
rect 3467 29665 3479 29668
rect 3421 29659 3479 29665
rect 3881 29665 3893 29668
rect 3927 29696 3939 29699
rect 4709 29699 4767 29705
rect 4709 29696 4721 29699
rect 3927 29668 4721 29696
rect 3927 29665 3939 29668
rect 3881 29659 3939 29665
rect 4709 29665 4721 29668
rect 4755 29696 4767 29699
rect 5258 29696 5264 29708
rect 4755 29668 5264 29696
rect 4755 29665 4767 29668
rect 4709 29659 4767 29665
rect 5258 29656 5264 29668
rect 5316 29656 5322 29708
rect 7561 29699 7619 29705
rect 7561 29665 7573 29699
rect 7607 29696 7619 29699
rect 9674 29696 9680 29708
rect 7607 29668 8708 29696
rect 9587 29668 9680 29696
rect 7607 29665 7619 29668
rect 7561 29659 7619 29665
rect 8680 29640 8708 29668
rect 9674 29656 9680 29668
rect 9732 29696 9738 29708
rect 10502 29696 10508 29708
rect 9732 29668 10508 29696
rect 9732 29656 9738 29668
rect 10502 29656 10508 29668
rect 10560 29656 10566 29708
rect 12250 29656 12256 29708
rect 12308 29696 12314 29708
rect 12417 29699 12475 29705
rect 12417 29696 12429 29699
rect 12308 29668 12429 29696
rect 12308 29656 12314 29668
rect 12417 29665 12429 29668
rect 12463 29665 12475 29699
rect 12417 29659 12475 29665
rect 15105 29699 15163 29705
rect 15105 29665 15117 29699
rect 15151 29696 15163 29699
rect 15194 29696 15200 29708
rect 15151 29668 15200 29696
rect 15151 29665 15163 29668
rect 15105 29659 15163 29665
rect 15194 29656 15200 29668
rect 15252 29696 15258 29708
rect 15746 29696 15752 29708
rect 15252 29668 15752 29696
rect 15252 29656 15258 29668
rect 15746 29656 15752 29668
rect 15804 29656 15810 29708
rect 15924 29699 15982 29705
rect 15924 29665 15936 29699
rect 15970 29696 15982 29699
rect 17034 29696 17040 29708
rect 15970 29668 17040 29696
rect 15970 29665 15982 29668
rect 15924 29659 15982 29665
rect 17034 29656 17040 29668
rect 17092 29656 17098 29708
rect 19518 29696 19524 29708
rect 19479 29668 19524 29696
rect 19518 29656 19524 29668
rect 19576 29656 19582 29708
rect 23566 29696 23572 29708
rect 23527 29668 23572 29696
rect 23566 29656 23572 29668
rect 23624 29656 23630 29708
rect 25038 29696 25044 29708
rect 24999 29668 25044 29696
rect 25038 29656 25044 29668
rect 25096 29656 25102 29708
rect 27706 29696 27712 29708
rect 27667 29668 27712 29696
rect 27706 29656 27712 29668
rect 27764 29656 27770 29708
rect 34514 29656 34520 29708
rect 34572 29696 34578 29708
rect 35437 29699 35495 29705
rect 35437 29696 35449 29699
rect 34572 29668 35449 29696
rect 34572 29656 34578 29668
rect 35437 29665 35449 29668
rect 35483 29665 35495 29699
rect 35437 29659 35495 29665
rect 1394 29628 1400 29640
rect 1355 29600 1400 29628
rect 1394 29588 1400 29600
rect 1452 29588 1458 29640
rect 7466 29588 7472 29640
rect 7524 29628 7530 29640
rect 8018 29628 8024 29640
rect 7524 29600 8024 29628
rect 7524 29588 7530 29600
rect 8018 29588 8024 29600
rect 8076 29628 8082 29640
rect 8481 29631 8539 29637
rect 8481 29628 8493 29631
rect 8076 29600 8493 29628
rect 8076 29588 8082 29600
rect 8481 29597 8493 29600
rect 8527 29597 8539 29631
rect 8481 29591 8539 29597
rect 8662 29588 8668 29640
rect 8720 29628 8726 29640
rect 8720 29600 8813 29628
rect 8720 29588 8726 29600
rect 12066 29588 12072 29640
rect 12124 29628 12130 29640
rect 12161 29631 12219 29637
rect 12161 29628 12173 29631
rect 12124 29600 12173 29628
rect 12124 29588 12130 29600
rect 12161 29597 12173 29600
rect 12207 29597 12219 29631
rect 12161 29591 12219 29597
rect 15657 29631 15715 29637
rect 15657 29597 15669 29631
rect 15703 29597 15715 29631
rect 18138 29628 18144 29640
rect 18099 29600 18144 29628
rect 15657 29591 15715 29597
rect 7193 29495 7251 29501
rect 7193 29461 7205 29495
rect 7239 29492 7251 29495
rect 7834 29492 7840 29504
rect 7239 29464 7840 29492
rect 7239 29461 7251 29464
rect 7193 29455 7251 29461
rect 7834 29452 7840 29464
rect 7892 29452 7898 29504
rect 8018 29492 8024 29504
rect 7979 29464 8024 29492
rect 8018 29452 8024 29464
rect 8076 29452 8082 29504
rect 15010 29452 15016 29504
rect 15068 29492 15074 29504
rect 15672 29492 15700 29591
rect 18138 29588 18144 29600
rect 18196 29588 18202 29640
rect 19242 29588 19248 29640
rect 19300 29628 19306 29640
rect 19613 29631 19671 29637
rect 19613 29628 19625 29631
rect 19300 29600 19625 29628
rect 19300 29588 19306 29600
rect 19613 29597 19625 29600
rect 19659 29597 19671 29631
rect 19613 29591 19671 29597
rect 19705 29631 19763 29637
rect 19705 29597 19717 29631
rect 19751 29628 19763 29631
rect 19978 29628 19984 29640
rect 19751 29600 19984 29628
rect 19751 29597 19763 29600
rect 19705 29591 19763 29597
rect 18874 29520 18880 29572
rect 18932 29560 18938 29572
rect 19720 29560 19748 29591
rect 19978 29588 19984 29600
rect 20036 29588 20042 29640
rect 24854 29588 24860 29640
rect 24912 29628 24918 29640
rect 25133 29631 25191 29637
rect 25133 29628 25145 29631
rect 24912 29600 25145 29628
rect 24912 29588 24918 29600
rect 25133 29597 25145 29600
rect 25179 29597 25191 29631
rect 25314 29628 25320 29640
rect 25227 29600 25320 29628
rect 25133 29591 25191 29597
rect 25314 29588 25320 29600
rect 25372 29628 25378 29640
rect 25774 29628 25780 29640
rect 25372 29600 25780 29628
rect 25372 29588 25378 29600
rect 25774 29588 25780 29600
rect 25832 29588 25838 29640
rect 26142 29588 26148 29640
rect 26200 29628 26206 29640
rect 26513 29631 26571 29637
rect 26513 29628 26525 29631
rect 26200 29600 26525 29628
rect 26200 29588 26206 29600
rect 26513 29597 26525 29600
rect 26559 29597 26571 29631
rect 31294 29628 31300 29640
rect 31255 29600 31300 29628
rect 26513 29591 26571 29597
rect 31294 29588 31300 29600
rect 31352 29628 31358 29640
rect 32217 29631 32275 29637
rect 32217 29628 32229 29631
rect 31352 29600 32229 29628
rect 31352 29588 31358 29600
rect 32217 29597 32229 29600
rect 32263 29597 32275 29631
rect 32217 29591 32275 29597
rect 18932 29532 19748 29560
rect 18932 29520 18938 29532
rect 16022 29492 16028 29504
rect 15068 29464 16028 29492
rect 15068 29452 15074 29464
rect 16022 29452 16028 29464
rect 16080 29452 16086 29504
rect 16574 29452 16580 29504
rect 16632 29492 16638 29504
rect 17037 29495 17095 29501
rect 17037 29492 17049 29495
rect 16632 29464 17049 29492
rect 16632 29452 16638 29464
rect 17037 29461 17049 29464
rect 17083 29461 17095 29495
rect 17037 29455 17095 29461
rect 19058 29452 19064 29504
rect 19116 29492 19122 29504
rect 19153 29495 19211 29501
rect 19153 29492 19165 29495
rect 19116 29464 19165 29492
rect 19116 29452 19122 29464
rect 19153 29461 19165 29464
rect 19199 29461 19211 29495
rect 19153 29455 19211 29461
rect 19886 29452 19892 29504
rect 19944 29492 19950 29504
rect 20165 29495 20223 29501
rect 20165 29492 20177 29495
rect 19944 29464 20177 29492
rect 19944 29452 19950 29464
rect 20165 29461 20177 29464
rect 20211 29461 20223 29495
rect 20165 29455 20223 29461
rect 24486 29452 24492 29504
rect 24544 29492 24550 29504
rect 24673 29495 24731 29501
rect 24673 29492 24685 29495
rect 24544 29464 24685 29492
rect 24544 29452 24550 29464
rect 24673 29461 24685 29464
rect 24719 29461 24731 29495
rect 24673 29455 24731 29461
rect 26510 29452 26516 29504
rect 26568 29492 26574 29504
rect 27525 29495 27583 29501
rect 27525 29492 27537 29495
rect 26568 29464 27537 29492
rect 26568 29452 26574 29464
rect 27525 29461 27537 29464
rect 27571 29492 27583 29495
rect 28718 29492 28724 29504
rect 27571 29464 28724 29492
rect 27571 29461 27583 29464
rect 27525 29455 27583 29461
rect 28718 29452 28724 29464
rect 28776 29452 28782 29504
rect 33134 29452 33140 29504
rect 33192 29492 33198 29504
rect 33597 29495 33655 29501
rect 33597 29492 33609 29495
rect 33192 29464 33609 29492
rect 33192 29452 33198 29464
rect 33597 29461 33609 29464
rect 33643 29492 33655 29495
rect 34790 29492 34796 29504
rect 33643 29464 34796 29492
rect 33643 29461 33655 29464
rect 33597 29455 33655 29461
rect 34790 29452 34796 29464
rect 34848 29492 34854 29504
rect 34885 29495 34943 29501
rect 34885 29492 34897 29495
rect 34848 29464 34897 29492
rect 34848 29452 34854 29464
rect 34885 29461 34897 29464
rect 34931 29461 34943 29495
rect 34885 29455 34943 29461
rect 1104 29402 38824 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 34966 29402
rect 35018 29350 35030 29402
rect 35082 29350 35094 29402
rect 35146 29350 35158 29402
rect 35210 29350 38824 29402
rect 1104 29328 38824 29350
rect 1670 29288 1676 29300
rect 1631 29260 1676 29288
rect 1670 29248 1676 29260
rect 1728 29248 1734 29300
rect 2038 29288 2044 29300
rect 1999 29260 2044 29288
rect 2038 29248 2044 29260
rect 2096 29248 2102 29300
rect 3326 29288 3332 29300
rect 3287 29260 3332 29288
rect 3326 29248 3332 29260
rect 3384 29248 3390 29300
rect 5166 29248 5172 29300
rect 5224 29288 5230 29300
rect 5629 29291 5687 29297
rect 5629 29288 5641 29291
rect 5224 29260 5641 29288
rect 5224 29248 5230 29260
rect 5629 29257 5641 29260
rect 5675 29288 5687 29291
rect 6181 29291 6239 29297
rect 6181 29288 6193 29291
rect 5675 29260 6193 29288
rect 5675 29257 5687 29260
rect 5629 29251 5687 29257
rect 6181 29257 6193 29260
rect 6227 29257 6239 29291
rect 7098 29288 7104 29300
rect 7059 29260 7104 29288
rect 6181 29251 6239 29257
rect 7098 29248 7104 29260
rect 7156 29248 7162 29300
rect 7466 29288 7472 29300
rect 7427 29260 7472 29288
rect 7466 29248 7472 29260
rect 7524 29248 7530 29300
rect 9306 29288 9312 29300
rect 9267 29260 9312 29288
rect 9306 29248 9312 29260
rect 9364 29248 9370 29300
rect 9950 29288 9956 29300
rect 9911 29260 9956 29288
rect 9950 29248 9956 29260
rect 10008 29248 10014 29300
rect 10410 29288 10416 29300
rect 10371 29260 10416 29288
rect 10410 29248 10416 29260
rect 10468 29248 10474 29300
rect 12250 29288 12256 29300
rect 12211 29260 12256 29288
rect 12250 29248 12256 29260
rect 12308 29248 12314 29300
rect 14829 29291 14887 29297
rect 14829 29257 14841 29291
rect 14875 29288 14887 29291
rect 15470 29288 15476 29300
rect 14875 29260 15476 29288
rect 14875 29257 14887 29260
rect 14829 29251 14887 29257
rect 15470 29248 15476 29260
rect 15528 29288 15534 29300
rect 15528 29260 16528 29288
rect 15528 29248 15534 29260
rect 11517 29223 11575 29229
rect 11517 29189 11529 29223
rect 11563 29220 11575 29223
rect 12066 29220 12072 29232
rect 11563 29192 12072 29220
rect 11563 29189 11575 29192
rect 11517 29183 11575 29189
rect 12066 29180 12072 29192
rect 12124 29220 12130 29232
rect 12621 29223 12679 29229
rect 12621 29220 12633 29223
rect 12124 29192 12633 29220
rect 12124 29180 12130 29192
rect 12621 29189 12633 29192
rect 12667 29189 12679 29223
rect 15930 29220 15936 29232
rect 15891 29192 15936 29220
rect 12621 29183 12679 29189
rect 15930 29180 15936 29192
rect 15988 29180 15994 29232
rect 1394 29112 1400 29164
rect 1452 29152 1458 29164
rect 1946 29152 1952 29164
rect 1452 29124 1952 29152
rect 1452 29112 1458 29124
rect 1946 29112 1952 29124
rect 2004 29152 2010 29164
rect 2409 29155 2467 29161
rect 2409 29152 2421 29155
rect 2004 29124 2421 29152
rect 2004 29112 2010 29124
rect 2409 29121 2421 29124
rect 2455 29152 2467 29155
rect 2777 29155 2835 29161
rect 2777 29152 2789 29155
rect 2455 29124 2789 29152
rect 2455 29121 2467 29124
rect 2409 29115 2467 29121
rect 2777 29121 2789 29124
rect 2823 29152 2835 29155
rect 7837 29155 7895 29161
rect 2823 29124 4108 29152
rect 2823 29121 2835 29124
rect 2777 29115 2835 29121
rect 4080 29096 4108 29124
rect 7837 29121 7849 29155
rect 7883 29152 7895 29155
rect 10962 29152 10968 29164
rect 7883 29124 8064 29152
rect 10923 29124 10968 29152
rect 7883 29121 7895 29124
rect 7837 29115 7895 29121
rect 2682 29044 2688 29096
rect 2740 29084 2746 29096
rect 3145 29087 3203 29093
rect 3145 29084 3157 29087
rect 2740 29056 3157 29084
rect 2740 29044 2746 29056
rect 3145 29053 3157 29056
rect 3191 29084 3203 29087
rect 3697 29087 3755 29093
rect 3697 29084 3709 29087
rect 3191 29056 3709 29084
rect 3191 29053 3203 29056
rect 3145 29047 3203 29053
rect 3697 29053 3709 29056
rect 3743 29053 3755 29087
rect 3697 29047 3755 29053
rect 4062 29044 4068 29096
rect 4120 29084 4126 29096
rect 4249 29087 4307 29093
rect 4249 29084 4261 29087
rect 4120 29056 4261 29084
rect 4120 29044 4126 29056
rect 4249 29053 4261 29056
rect 4295 29084 4307 29087
rect 5258 29084 5264 29096
rect 4295 29056 5264 29084
rect 4295 29053 4307 29056
rect 4249 29047 4307 29053
rect 5258 29044 5264 29056
rect 5316 29044 5322 29096
rect 7926 29084 7932 29096
rect 7887 29056 7932 29084
rect 7926 29044 7932 29056
rect 7984 29044 7990 29096
rect 8036 29084 8064 29124
rect 10962 29112 10968 29124
rect 11020 29112 11026 29164
rect 13081 29155 13139 29161
rect 13081 29121 13093 29155
rect 13127 29152 13139 29155
rect 16390 29152 16396 29164
rect 13127 29124 13584 29152
rect 16351 29124 16396 29152
rect 13127 29121 13139 29124
rect 13081 29115 13139 29121
rect 13556 29096 13584 29124
rect 16390 29112 16396 29124
rect 16448 29112 16454 29164
rect 16500 29161 16528 29260
rect 18230 29248 18236 29300
rect 18288 29288 18294 29300
rect 19245 29291 19303 29297
rect 19245 29288 19257 29291
rect 18288 29260 19257 29288
rect 18288 29248 18294 29260
rect 19245 29257 19257 29260
rect 19291 29288 19303 29291
rect 19518 29288 19524 29300
rect 19291 29260 19524 29288
rect 19291 29257 19303 29260
rect 19245 29251 19303 29257
rect 19518 29248 19524 29260
rect 19576 29248 19582 29300
rect 19978 29248 19984 29300
rect 20036 29288 20042 29300
rect 20993 29291 21051 29297
rect 20993 29288 21005 29291
rect 20036 29260 21005 29288
rect 20036 29248 20042 29260
rect 20993 29257 21005 29260
rect 21039 29257 21051 29291
rect 20993 29251 21051 29257
rect 23477 29291 23535 29297
rect 23477 29257 23489 29291
rect 23523 29288 23535 29291
rect 23566 29288 23572 29300
rect 23523 29260 23572 29288
rect 23523 29257 23535 29260
rect 23477 29251 23535 29257
rect 23566 29248 23572 29260
rect 23624 29248 23630 29300
rect 27706 29248 27712 29300
rect 27764 29288 27770 29300
rect 27985 29291 28043 29297
rect 27985 29288 27997 29291
rect 27764 29260 27997 29288
rect 27764 29248 27770 29260
rect 27985 29257 27997 29260
rect 28031 29257 28043 29291
rect 27985 29251 28043 29257
rect 17034 29220 17040 29232
rect 16947 29192 17040 29220
rect 17034 29180 17040 29192
rect 17092 29220 17098 29232
rect 18690 29220 18696 29232
rect 17092 29192 18696 29220
rect 17092 29180 17098 29192
rect 18690 29180 18696 29192
rect 18748 29180 18754 29232
rect 18874 29220 18880 29232
rect 18835 29192 18880 29220
rect 18874 29180 18880 29192
rect 18932 29180 18938 29232
rect 25038 29180 25044 29232
rect 25096 29180 25102 29232
rect 32674 29220 32680 29232
rect 32635 29192 32680 29220
rect 32674 29180 32680 29192
rect 32732 29220 32738 29232
rect 33229 29223 33287 29229
rect 33229 29220 33241 29223
rect 32732 29192 33241 29220
rect 32732 29180 32738 29192
rect 33229 29189 33241 29192
rect 33275 29189 33287 29223
rect 33229 29183 33287 29189
rect 16485 29155 16543 29161
rect 16485 29121 16497 29155
rect 16531 29121 16543 29155
rect 16485 29115 16543 29121
rect 24765 29155 24823 29161
rect 24765 29121 24777 29155
rect 24811 29152 24823 29155
rect 25056 29152 25084 29180
rect 31294 29152 31300 29164
rect 24811 29124 25176 29152
rect 31255 29124 31300 29152
rect 24811 29121 24823 29124
rect 24765 29115 24823 29121
rect 8202 29093 8208 29096
rect 8196 29084 8208 29093
rect 8036 29056 8208 29084
rect 8196 29047 8208 29056
rect 8202 29044 8208 29047
rect 8260 29044 8266 29096
rect 13449 29087 13507 29093
rect 13449 29053 13461 29087
rect 13495 29053 13507 29087
rect 13449 29047 13507 29053
rect 4157 29019 4215 29025
rect 4157 28985 4169 29019
rect 4203 29016 4215 29019
rect 4494 29019 4552 29025
rect 4494 29016 4506 29019
rect 4203 28988 4506 29016
rect 4203 28985 4215 28988
rect 4157 28979 4215 28985
rect 4494 28985 4506 28988
rect 4540 29016 4552 29019
rect 5442 29016 5448 29028
rect 4540 28988 5448 29016
rect 4540 28985 4552 28988
rect 4494 28979 4552 28985
rect 5442 28976 5448 28988
rect 5500 28976 5506 29028
rect 10229 29019 10287 29025
rect 10229 29016 10241 29019
rect 9600 28988 10241 29016
rect 9600 28960 9628 28988
rect 10229 28985 10241 28988
rect 10275 29016 10287 29019
rect 10873 29019 10931 29025
rect 10873 29016 10885 29019
rect 10275 28988 10885 29016
rect 10275 28985 10287 28988
rect 10229 28979 10287 28985
rect 10873 28985 10885 28988
rect 10919 28985 10931 29019
rect 13464 29016 13492 29047
rect 13538 29044 13544 29096
rect 13596 29084 13602 29096
rect 13705 29087 13763 29093
rect 13705 29084 13717 29087
rect 13596 29056 13717 29084
rect 13596 29044 13602 29056
rect 13705 29053 13717 29056
rect 13751 29053 13763 29087
rect 13705 29047 13763 29053
rect 16206 29044 16212 29096
rect 16264 29084 16270 29096
rect 17126 29084 17132 29096
rect 16264 29056 17132 29084
rect 16264 29044 16270 29056
rect 17126 29044 17132 29056
rect 17184 29084 17190 29096
rect 17405 29087 17463 29093
rect 17405 29084 17417 29087
rect 17184 29056 17417 29084
rect 17184 29044 17190 29056
rect 17405 29053 17417 29056
rect 17451 29084 17463 29087
rect 19613 29087 19671 29093
rect 19613 29084 19625 29087
rect 17451 29056 19625 29084
rect 17451 29053 17463 29056
rect 17405 29047 17463 29053
rect 19613 29053 19625 29056
rect 19659 29084 19671 29087
rect 20162 29084 20168 29096
rect 19659 29056 20168 29084
rect 19659 29053 19671 29056
rect 19613 29047 19671 29053
rect 20162 29044 20168 29056
rect 20220 29044 20226 29096
rect 23937 29087 23995 29093
rect 23937 29053 23949 29087
rect 23983 29084 23995 29087
rect 24026 29084 24032 29096
rect 23983 29056 24032 29084
rect 23983 29053 23995 29056
rect 23937 29047 23995 29053
rect 24026 29044 24032 29056
rect 24084 29084 24090 29096
rect 24578 29084 24584 29096
rect 24084 29056 24584 29084
rect 24084 29044 24090 29056
rect 24578 29044 24584 29056
rect 24636 29044 24642 29096
rect 25038 29084 25044 29096
rect 24999 29056 25044 29084
rect 25038 29044 25044 29056
rect 25096 29044 25102 29096
rect 25148 29084 25176 29124
rect 31294 29112 31300 29124
rect 31352 29112 31358 29164
rect 27525 29087 27583 29093
rect 27525 29084 27537 29087
rect 25148 29056 27537 29084
rect 27525 29053 27537 29056
rect 27571 29053 27583 29087
rect 31312 29084 31340 29112
rect 31938 29084 31944 29096
rect 31312 29056 31944 29084
rect 27525 29047 27583 29053
rect 31938 29044 31944 29056
rect 31996 29044 32002 29096
rect 34885 29087 34943 29093
rect 34885 29084 34897 29087
rect 34348 29056 34897 29084
rect 15749 29019 15807 29025
rect 15749 29016 15761 29019
rect 13464 28988 13860 29016
rect 10873 28979 10931 28985
rect 9582 28908 9588 28960
rect 9640 28908 9646 28960
rect 10502 28908 10508 28960
rect 10560 28948 10566 28960
rect 10781 28951 10839 28957
rect 10781 28948 10793 28951
rect 10560 28920 10793 28948
rect 10560 28908 10566 28920
rect 10781 28917 10793 28920
rect 10827 28917 10839 28951
rect 13832 28948 13860 28988
rect 15120 28988 15761 29016
rect 15120 28960 15148 28988
rect 15749 28985 15761 28988
rect 15795 29016 15807 29019
rect 16301 29019 16359 29025
rect 16301 29016 16313 29019
rect 15795 28988 16313 29016
rect 15795 28985 15807 28988
rect 15749 28979 15807 28985
rect 16301 28985 16313 28988
rect 16347 28985 16359 29019
rect 16301 28979 16359 28985
rect 17770 28976 17776 29028
rect 17828 29016 17834 29028
rect 18509 29019 18567 29025
rect 17828 28988 17908 29016
rect 17828 28976 17834 28988
rect 14366 28948 14372 28960
rect 13832 28920 14372 28948
rect 10781 28911 10839 28917
rect 14366 28908 14372 28920
rect 14424 28908 14430 28960
rect 15102 28908 15108 28960
rect 15160 28908 15166 28960
rect 17880 28948 17908 28988
rect 18509 28985 18521 29019
rect 18555 29016 18567 29019
rect 19242 29016 19248 29028
rect 18555 28988 19248 29016
rect 18555 28985 18567 28988
rect 18509 28979 18567 28985
rect 19242 28976 19248 28988
rect 19300 28976 19306 29028
rect 19886 29025 19892 29028
rect 19880 29016 19892 29025
rect 19847 28988 19892 29016
rect 19880 28979 19892 28988
rect 19886 28976 19892 28979
rect 19944 28976 19950 29028
rect 24670 28976 24676 29028
rect 24728 29016 24734 29028
rect 25314 29025 25320 29028
rect 25308 29016 25320 29025
rect 24728 28988 25320 29016
rect 24728 28976 24734 28988
rect 25308 28979 25320 28988
rect 25314 28976 25320 28979
rect 25372 28976 25378 29028
rect 31570 29025 31576 29028
rect 31205 29019 31263 29025
rect 31205 28985 31217 29019
rect 31251 29016 31263 29019
rect 31564 29016 31576 29025
rect 31251 28988 31576 29016
rect 31251 28985 31263 28988
rect 31205 28979 31263 28985
rect 31564 28979 31576 28988
rect 31570 28976 31576 28979
rect 31628 28976 31634 29028
rect 34348 28960 34376 29056
rect 34885 29053 34897 29056
rect 34931 29053 34943 29087
rect 34885 29047 34943 29053
rect 34514 28976 34520 29028
rect 34572 29016 34578 29028
rect 34609 29019 34667 29025
rect 34609 29016 34621 29019
rect 34572 28988 34621 29016
rect 34572 28976 34578 28988
rect 34609 28985 34621 28988
rect 34655 28985 34667 29019
rect 34609 28979 34667 28985
rect 34790 28976 34796 29028
rect 34848 29016 34854 29028
rect 35130 29019 35188 29025
rect 35130 29016 35142 29019
rect 34848 28988 35142 29016
rect 34848 28976 34854 28988
rect 35130 28985 35142 28988
rect 35176 28985 35188 29019
rect 35130 28979 35188 28985
rect 18874 28948 18880 28960
rect 17880 28920 18880 28948
rect 18874 28908 18880 28920
rect 18932 28908 18938 28960
rect 24118 28948 24124 28960
rect 24079 28920 24124 28948
rect 24118 28908 24124 28920
rect 24176 28908 24182 28960
rect 24854 28908 24860 28960
rect 24912 28948 24918 28960
rect 26418 28948 26424 28960
rect 24912 28920 26424 28948
rect 24912 28908 24918 28920
rect 26418 28908 26424 28920
rect 26476 28908 26482 28960
rect 30561 28951 30619 28957
rect 30561 28917 30573 28951
rect 30607 28948 30619 28951
rect 30834 28948 30840 28960
rect 30607 28920 30840 28948
rect 30607 28917 30619 28920
rect 30561 28911 30619 28917
rect 30834 28908 30840 28920
rect 30892 28908 30898 28960
rect 33689 28951 33747 28957
rect 33689 28917 33701 28951
rect 33735 28948 33747 28951
rect 34330 28948 34336 28960
rect 33735 28920 34336 28948
rect 33735 28917 33747 28920
rect 33689 28911 33747 28917
rect 34330 28908 34336 28920
rect 34388 28908 34394 28960
rect 34882 28908 34888 28960
rect 34940 28948 34946 28960
rect 36265 28951 36323 28957
rect 36265 28948 36277 28951
rect 34940 28920 36277 28948
rect 34940 28908 34946 28920
rect 36265 28917 36277 28920
rect 36311 28917 36323 28951
rect 36265 28911 36323 28917
rect 1104 28858 38824 28880
rect 1104 28806 19606 28858
rect 19658 28806 19670 28858
rect 19722 28806 19734 28858
rect 19786 28806 19798 28858
rect 19850 28806 38824 28858
rect 1104 28784 38824 28806
rect 1946 28744 1952 28756
rect 1907 28716 1952 28744
rect 1946 28704 1952 28716
rect 2004 28704 2010 28756
rect 2409 28747 2467 28753
rect 2409 28713 2421 28747
rect 2455 28744 2467 28747
rect 2682 28744 2688 28756
rect 2455 28716 2688 28744
rect 2455 28713 2467 28716
rect 2409 28707 2467 28713
rect 2682 28704 2688 28716
rect 2740 28704 2746 28756
rect 5442 28744 5448 28756
rect 5403 28716 5448 28744
rect 5442 28704 5448 28716
rect 5500 28704 5506 28756
rect 8294 28704 8300 28756
rect 8352 28744 8358 28756
rect 8481 28747 8539 28753
rect 8481 28744 8493 28747
rect 8352 28716 8493 28744
rect 8352 28704 8358 28716
rect 8481 28713 8493 28716
rect 8527 28713 8539 28747
rect 8481 28707 8539 28713
rect 9861 28747 9919 28753
rect 9861 28713 9873 28747
rect 9907 28744 9919 28747
rect 10502 28744 10508 28756
rect 9907 28716 10508 28744
rect 9907 28713 9919 28716
rect 9861 28707 9919 28713
rect 10502 28704 10508 28716
rect 10560 28704 10566 28756
rect 10873 28747 10931 28753
rect 10873 28713 10885 28747
rect 10919 28744 10931 28747
rect 10962 28744 10968 28756
rect 10919 28716 10968 28744
rect 10919 28713 10931 28716
rect 10873 28707 10931 28713
rect 10962 28704 10968 28716
rect 11020 28704 11026 28756
rect 11057 28747 11115 28753
rect 11057 28713 11069 28747
rect 11103 28744 11115 28747
rect 12342 28744 12348 28756
rect 11103 28716 12348 28744
rect 11103 28713 11115 28716
rect 11057 28707 11115 28713
rect 12342 28704 12348 28716
rect 12400 28744 12406 28756
rect 12802 28744 12808 28756
rect 12400 28716 12664 28744
rect 12763 28716 12808 28744
rect 12400 28704 12406 28716
rect 7368 28679 7426 28685
rect 7368 28645 7380 28679
rect 7414 28676 7426 28679
rect 7558 28676 7564 28688
rect 7414 28648 7564 28676
rect 7414 28645 7426 28648
rect 7368 28639 7426 28645
rect 7558 28636 7564 28648
rect 7616 28636 7622 28688
rect 10980 28676 11008 28704
rect 12636 28676 12664 28716
rect 12802 28704 12808 28716
rect 12860 28704 12866 28756
rect 13538 28744 13544 28756
rect 13499 28716 13544 28744
rect 13538 28704 13544 28716
rect 13596 28704 13602 28756
rect 13814 28704 13820 28756
rect 13872 28744 13878 28756
rect 13909 28747 13967 28753
rect 13909 28744 13921 28747
rect 13872 28716 13921 28744
rect 13872 28704 13878 28716
rect 13909 28713 13921 28716
rect 13955 28713 13967 28747
rect 14366 28744 14372 28756
rect 14279 28716 14372 28744
rect 13909 28707 13967 28713
rect 14366 28704 14372 28716
rect 14424 28744 14430 28756
rect 15010 28744 15016 28756
rect 14424 28716 15016 28744
rect 14424 28704 14430 28716
rect 15010 28704 15016 28716
rect 15068 28704 15074 28756
rect 15194 28704 15200 28756
rect 15252 28744 15258 28756
rect 15381 28747 15439 28753
rect 15381 28744 15393 28747
rect 15252 28716 15393 28744
rect 15252 28704 15258 28716
rect 15381 28713 15393 28716
rect 15427 28713 15439 28747
rect 15838 28744 15844 28756
rect 15799 28716 15844 28744
rect 15381 28707 15439 28713
rect 15838 28704 15844 28716
rect 15896 28704 15902 28756
rect 16390 28744 16396 28756
rect 16351 28716 16396 28744
rect 16390 28704 16396 28716
rect 16448 28704 16454 28756
rect 18230 28744 18236 28756
rect 18191 28716 18236 28744
rect 18230 28704 18236 28716
rect 18288 28704 18294 28756
rect 18966 28744 18972 28756
rect 18927 28716 18972 28744
rect 18966 28704 18972 28716
rect 19024 28704 19030 28756
rect 19242 28744 19248 28756
rect 19203 28716 19248 28744
rect 19242 28704 19248 28716
rect 19300 28704 19306 28756
rect 20162 28704 20168 28756
rect 20220 28744 20226 28756
rect 20257 28747 20315 28753
rect 20257 28744 20269 28747
rect 20220 28716 20269 28744
rect 20220 28704 20226 28716
rect 20257 28713 20269 28716
rect 20303 28744 20315 28747
rect 20625 28747 20683 28753
rect 20625 28744 20637 28747
rect 20303 28716 20637 28744
rect 20303 28713 20315 28716
rect 20257 28707 20315 28713
rect 20625 28713 20637 28716
rect 20671 28713 20683 28747
rect 24026 28744 24032 28756
rect 23987 28716 24032 28744
rect 20625 28707 20683 28713
rect 15746 28676 15752 28688
rect 10980 28648 11652 28676
rect 12636 28648 13768 28676
rect 15707 28648 15752 28676
rect 2774 28568 2780 28620
rect 2832 28608 2838 28620
rect 3878 28608 3884 28620
rect 2832 28580 2877 28608
rect 3791 28580 3884 28608
rect 2832 28568 2838 28580
rect 3878 28568 3884 28580
rect 3936 28608 3942 28620
rect 4062 28608 4068 28620
rect 3936 28580 4068 28608
rect 3936 28568 3942 28580
rect 4062 28568 4068 28580
rect 4120 28568 4126 28620
rect 4332 28611 4390 28617
rect 4332 28577 4344 28611
rect 4378 28608 4390 28611
rect 4614 28608 4620 28620
rect 4378 28580 4620 28608
rect 4378 28577 4390 28580
rect 4332 28571 4390 28577
rect 4614 28568 4620 28580
rect 4672 28568 4678 28620
rect 5258 28568 5264 28620
rect 5316 28608 5322 28620
rect 6638 28608 6644 28620
rect 5316 28580 6644 28608
rect 5316 28568 5322 28580
rect 6638 28568 6644 28580
rect 6696 28608 6702 28620
rect 7101 28611 7159 28617
rect 7101 28608 7113 28611
rect 6696 28580 7113 28608
rect 6696 28568 6702 28580
rect 7101 28577 7113 28580
rect 7147 28608 7159 28611
rect 7926 28608 7932 28620
rect 7147 28580 7932 28608
rect 7147 28577 7159 28580
rect 7101 28571 7159 28577
rect 7926 28568 7932 28580
rect 7984 28568 7990 28620
rect 9674 28608 9680 28620
rect 9635 28580 9680 28608
rect 9674 28568 9680 28580
rect 9732 28568 9738 28620
rect 11422 28608 11428 28620
rect 11383 28580 11428 28608
rect 11422 28568 11428 28580
rect 11480 28568 11486 28620
rect 1854 28500 1860 28552
rect 1912 28540 1918 28552
rect 2869 28543 2927 28549
rect 2869 28540 2881 28543
rect 1912 28512 2881 28540
rect 1912 28500 1918 28512
rect 2869 28509 2881 28512
rect 2915 28509 2927 28543
rect 2869 28503 2927 28509
rect 2958 28500 2964 28552
rect 3016 28540 3022 28552
rect 11514 28540 11520 28552
rect 3016 28512 3109 28540
rect 11475 28512 11520 28540
rect 3016 28500 3022 28512
rect 11514 28500 11520 28512
rect 11572 28500 11578 28552
rect 11624 28549 11652 28648
rect 13740 28620 13768 28648
rect 15746 28636 15752 28648
rect 15804 28636 15810 28688
rect 18984 28676 19012 28704
rect 19613 28679 19671 28685
rect 19613 28676 19625 28679
rect 18984 28648 19625 28676
rect 19613 28645 19625 28648
rect 19659 28676 19671 28679
rect 19702 28676 19708 28688
rect 19659 28648 19708 28676
rect 19659 28645 19671 28648
rect 19613 28639 19671 28645
rect 19702 28636 19708 28648
rect 19760 28636 19766 28688
rect 12621 28611 12679 28617
rect 12621 28577 12633 28611
rect 12667 28608 12679 28611
rect 12710 28608 12716 28620
rect 12667 28580 12716 28608
rect 12667 28577 12679 28580
rect 12621 28571 12679 28577
rect 12710 28568 12716 28580
rect 12768 28568 12774 28620
rect 13722 28608 13728 28620
rect 13635 28580 13728 28608
rect 13722 28568 13728 28580
rect 13780 28568 13786 28620
rect 20640 28608 20668 28707
rect 24026 28704 24032 28716
rect 24084 28704 24090 28756
rect 24397 28747 24455 28753
rect 24397 28713 24409 28747
rect 24443 28744 24455 28747
rect 24762 28744 24768 28756
rect 24443 28716 24768 28744
rect 24443 28713 24455 28716
rect 24397 28707 24455 28713
rect 24762 28704 24768 28716
rect 24820 28704 24826 28756
rect 24857 28747 24915 28753
rect 24857 28713 24869 28747
rect 24903 28744 24915 28747
rect 25130 28744 25136 28756
rect 24903 28716 25136 28744
rect 24903 28713 24915 28716
rect 24857 28707 24915 28713
rect 25130 28704 25136 28716
rect 25188 28704 25194 28756
rect 25225 28747 25283 28753
rect 25225 28713 25237 28747
rect 25271 28744 25283 28747
rect 25682 28744 25688 28756
rect 25271 28716 25688 28744
rect 25271 28713 25283 28716
rect 25225 28707 25283 28713
rect 25682 28704 25688 28716
rect 25740 28744 25746 28756
rect 26142 28744 26148 28756
rect 25740 28716 26148 28744
rect 25740 28704 25746 28716
rect 26142 28704 26148 28716
rect 26200 28704 26206 28756
rect 30377 28747 30435 28753
rect 30377 28713 30389 28747
rect 30423 28744 30435 28747
rect 30837 28747 30895 28753
rect 30837 28744 30849 28747
rect 30423 28716 30849 28744
rect 30423 28713 30435 28716
rect 30377 28707 30435 28713
rect 30837 28713 30849 28716
rect 30883 28744 30895 28747
rect 31570 28744 31576 28756
rect 30883 28716 31576 28744
rect 30883 28713 30895 28716
rect 30837 28707 30895 28713
rect 31570 28704 31576 28716
rect 31628 28704 31634 28756
rect 33502 28744 33508 28756
rect 33463 28716 33508 28744
rect 33502 28704 33508 28716
rect 33560 28704 33566 28756
rect 24670 28676 24676 28688
rect 24631 28648 24676 28676
rect 24670 28636 24676 28648
rect 24728 28636 24734 28688
rect 26418 28636 26424 28688
rect 26476 28676 26482 28688
rect 34882 28685 34888 28688
rect 26758 28679 26816 28685
rect 26758 28676 26770 28679
rect 26476 28648 26770 28676
rect 26476 28636 26482 28648
rect 26758 28645 26770 28648
rect 26804 28645 26816 28679
rect 34876 28676 34888 28685
rect 34843 28648 34888 28676
rect 26758 28639 26816 28645
rect 34876 28639 34888 28648
rect 34882 28636 34888 28639
rect 34940 28636 34946 28688
rect 20714 28608 20720 28620
rect 20627 28580 20720 28608
rect 20714 28568 20720 28580
rect 20772 28608 20778 28620
rect 21174 28617 21180 28620
rect 20901 28611 20959 28617
rect 20901 28608 20913 28611
rect 20772 28580 20913 28608
rect 20772 28568 20778 28580
rect 20901 28577 20913 28580
rect 20947 28577 20959 28611
rect 21168 28608 21180 28617
rect 21135 28580 21180 28608
rect 20901 28571 20959 28577
rect 21168 28571 21180 28580
rect 21174 28568 21180 28571
rect 21232 28568 21238 28620
rect 32214 28568 32220 28620
rect 32272 28608 32278 28620
rect 32381 28611 32439 28617
rect 32381 28608 32393 28611
rect 32272 28580 32393 28608
rect 32272 28568 32278 28580
rect 32381 28577 32393 28580
rect 32427 28577 32439 28611
rect 32381 28571 32439 28577
rect 11609 28543 11667 28549
rect 11609 28509 11621 28543
rect 11655 28540 11667 28543
rect 11790 28540 11796 28552
rect 11655 28512 11796 28540
rect 11655 28509 11667 28512
rect 11609 28503 11667 28509
rect 11790 28500 11796 28512
rect 11848 28500 11854 28552
rect 16022 28540 16028 28552
rect 15935 28512 16028 28540
rect 16022 28500 16028 28512
rect 16080 28540 16086 28552
rect 16482 28540 16488 28552
rect 16080 28512 16488 28540
rect 16080 28500 16086 28512
rect 16482 28500 16488 28512
rect 16540 28500 16546 28552
rect 19705 28543 19763 28549
rect 19705 28509 19717 28543
rect 19751 28509 19763 28543
rect 19886 28540 19892 28552
rect 19847 28512 19892 28540
rect 19705 28503 19763 28509
rect 2317 28475 2375 28481
rect 2317 28441 2329 28475
rect 2363 28472 2375 28475
rect 2976 28472 3004 28500
rect 2363 28444 3004 28472
rect 19720 28472 19748 28503
rect 19886 28500 19892 28512
rect 19944 28500 19950 28552
rect 24578 28500 24584 28552
rect 24636 28540 24642 28552
rect 25317 28543 25375 28549
rect 25317 28540 25329 28543
rect 24636 28512 25329 28540
rect 24636 28500 24642 28512
rect 25317 28509 25329 28512
rect 25363 28509 25375 28543
rect 25498 28540 25504 28552
rect 25459 28512 25504 28540
rect 25317 28503 25375 28509
rect 25498 28500 25504 28512
rect 25556 28500 25562 28552
rect 26510 28540 26516 28552
rect 26252 28512 26516 28540
rect 19978 28472 19984 28484
rect 19720 28444 19984 28472
rect 2363 28441 2375 28444
rect 2317 28435 2375 28441
rect 19978 28432 19984 28444
rect 20036 28432 20042 28484
rect 22278 28472 22284 28484
rect 22239 28444 22284 28472
rect 22278 28432 22284 28444
rect 22336 28432 22342 28484
rect 25038 28364 25044 28416
rect 25096 28404 25102 28416
rect 25961 28407 26019 28413
rect 25961 28404 25973 28407
rect 25096 28376 25973 28404
rect 25096 28364 25102 28376
rect 25961 28373 25973 28376
rect 26007 28404 26019 28407
rect 26142 28404 26148 28416
rect 26007 28376 26148 28404
rect 26007 28373 26019 28376
rect 25961 28367 26019 28373
rect 26142 28364 26148 28376
rect 26200 28404 26206 28416
rect 26252 28413 26280 28512
rect 26510 28500 26516 28512
rect 26568 28500 26574 28552
rect 30926 28540 30932 28552
rect 30887 28512 30932 28540
rect 30926 28500 30932 28512
rect 30984 28500 30990 28552
rect 31021 28543 31079 28549
rect 31021 28509 31033 28543
rect 31067 28509 31079 28543
rect 31021 28503 31079 28509
rect 32125 28543 32183 28549
rect 32125 28509 32137 28543
rect 32171 28509 32183 28543
rect 34609 28543 34667 28549
rect 34609 28540 34621 28543
rect 32125 28503 32183 28509
rect 34440 28512 34621 28540
rect 30834 28432 30840 28484
rect 30892 28472 30898 28484
rect 31036 28472 31064 28503
rect 30892 28444 31064 28472
rect 30892 28432 30898 28444
rect 26237 28407 26295 28413
rect 26237 28404 26249 28407
rect 26200 28376 26249 28404
rect 26200 28364 26206 28376
rect 26237 28373 26249 28376
rect 26283 28373 26295 28407
rect 27890 28404 27896 28416
rect 27851 28376 27896 28404
rect 26237 28367 26295 28373
rect 27890 28364 27896 28376
rect 27948 28364 27954 28416
rect 30006 28404 30012 28416
rect 29967 28376 30012 28404
rect 30006 28364 30012 28376
rect 30064 28364 30070 28416
rect 30466 28404 30472 28416
rect 30427 28376 30472 28404
rect 30466 28364 30472 28376
rect 30524 28364 30530 28416
rect 31938 28404 31944 28416
rect 31851 28376 31944 28404
rect 31938 28364 31944 28376
rect 31996 28404 32002 28416
rect 32140 28404 32168 28503
rect 34330 28404 34336 28416
rect 31996 28376 34336 28404
rect 31996 28364 32002 28376
rect 34330 28364 34336 28376
rect 34388 28404 34394 28416
rect 34440 28413 34468 28512
rect 34609 28509 34621 28512
rect 34655 28509 34667 28543
rect 34609 28503 34667 28509
rect 34425 28407 34483 28413
rect 34425 28404 34437 28407
rect 34388 28376 34437 28404
rect 34388 28364 34394 28376
rect 34425 28373 34437 28376
rect 34471 28373 34483 28407
rect 35986 28404 35992 28416
rect 35947 28376 35992 28404
rect 34425 28367 34483 28373
rect 35986 28364 35992 28376
rect 36044 28364 36050 28416
rect 1104 28314 38824 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 34966 28314
rect 35018 28262 35030 28314
rect 35082 28262 35094 28314
rect 35146 28262 35158 28314
rect 35210 28262 38824 28314
rect 1104 28240 38824 28262
rect 1854 28200 1860 28212
rect 1815 28172 1860 28200
rect 1854 28160 1860 28172
rect 1912 28160 1918 28212
rect 4801 28203 4859 28209
rect 4801 28169 4813 28203
rect 4847 28200 4859 28203
rect 4890 28200 4896 28212
rect 4847 28172 4896 28200
rect 4847 28169 4859 28172
rect 4801 28163 4859 28169
rect 4890 28160 4896 28172
rect 4948 28160 4954 28212
rect 6638 28200 6644 28212
rect 6599 28172 6644 28200
rect 6638 28160 6644 28172
rect 6696 28160 6702 28212
rect 9217 28203 9275 28209
rect 9217 28169 9229 28203
rect 9263 28200 9275 28203
rect 9582 28200 9588 28212
rect 9263 28172 9588 28200
rect 9263 28169 9275 28172
rect 9217 28163 9275 28169
rect 9582 28160 9588 28172
rect 9640 28160 9646 28212
rect 9674 28160 9680 28212
rect 9732 28200 9738 28212
rect 9953 28203 10011 28209
rect 9953 28200 9965 28203
rect 9732 28172 9965 28200
rect 9732 28160 9738 28172
rect 9953 28169 9965 28172
rect 9999 28169 10011 28203
rect 11146 28200 11152 28212
rect 11059 28172 11152 28200
rect 9953 28163 10011 28169
rect 11146 28160 11152 28172
rect 11204 28200 11210 28212
rect 11514 28200 11520 28212
rect 11204 28172 11520 28200
rect 11204 28160 11210 28172
rect 11514 28160 11520 28172
rect 11572 28160 11578 28212
rect 11790 28200 11796 28212
rect 11751 28172 11796 28200
rect 11790 28160 11796 28172
rect 11848 28160 11854 28212
rect 12710 28160 12716 28212
rect 12768 28200 12774 28212
rect 13357 28203 13415 28209
rect 13357 28200 13369 28203
rect 12768 28172 13369 28200
rect 12768 28160 12774 28172
rect 13357 28169 13369 28172
rect 13403 28169 13415 28203
rect 13722 28200 13728 28212
rect 13683 28172 13728 28200
rect 13357 28163 13415 28169
rect 13722 28160 13728 28172
rect 13780 28160 13786 28212
rect 15473 28203 15531 28209
rect 15473 28169 15485 28203
rect 15519 28200 15531 28203
rect 15746 28200 15752 28212
rect 15519 28172 15752 28200
rect 15519 28169 15531 28172
rect 15473 28163 15531 28169
rect 15746 28160 15752 28172
rect 15804 28160 15810 28212
rect 15841 28203 15899 28209
rect 15841 28169 15853 28203
rect 15887 28200 15899 28203
rect 16022 28200 16028 28212
rect 15887 28172 16028 28200
rect 15887 28169 15899 28172
rect 15841 28163 15899 28169
rect 16022 28160 16028 28172
rect 16080 28160 16086 28212
rect 21634 28200 21640 28212
rect 21595 28172 21640 28200
rect 21634 28160 21640 28172
rect 21692 28160 21698 28212
rect 23477 28203 23535 28209
rect 23477 28169 23489 28203
rect 23523 28200 23535 28203
rect 24578 28200 24584 28212
rect 23523 28172 24584 28200
rect 23523 28169 23535 28172
rect 23477 28163 23535 28169
rect 24578 28160 24584 28172
rect 24636 28160 24642 28212
rect 25682 28200 25688 28212
rect 25643 28172 25688 28200
rect 25682 28160 25688 28172
rect 25740 28160 25746 28212
rect 26418 28160 26424 28212
rect 26476 28200 26482 28212
rect 28077 28203 28135 28209
rect 28077 28200 28089 28203
rect 26476 28172 28089 28200
rect 26476 28160 26482 28172
rect 28077 28169 28089 28172
rect 28123 28169 28135 28203
rect 28077 28163 28135 28169
rect 29733 28203 29791 28209
rect 29733 28169 29745 28203
rect 29779 28200 29791 28203
rect 30926 28200 30932 28212
rect 29779 28172 30932 28200
rect 29779 28169 29791 28172
rect 29733 28163 29791 28169
rect 30926 28160 30932 28172
rect 30984 28200 30990 28212
rect 31573 28203 31631 28209
rect 31573 28200 31585 28203
rect 30984 28172 31585 28200
rect 30984 28160 30990 28172
rect 31573 28169 31585 28172
rect 31619 28200 31631 28203
rect 32214 28200 32220 28212
rect 31619 28172 32220 28200
rect 31619 28169 31631 28172
rect 31573 28163 31631 28169
rect 32214 28160 32220 28172
rect 32272 28160 32278 28212
rect 33962 28160 33968 28212
rect 34020 28200 34026 28212
rect 34606 28200 34612 28212
rect 34020 28172 34612 28200
rect 34020 28160 34026 28172
rect 34606 28160 34612 28172
rect 34664 28160 34670 28212
rect 34701 28203 34759 28209
rect 34701 28169 34713 28203
rect 34747 28200 34759 28203
rect 34790 28200 34796 28212
rect 34747 28172 34796 28200
rect 34747 28169 34759 28172
rect 34701 28163 34759 28169
rect 12621 28135 12679 28141
rect 12621 28101 12633 28135
rect 12667 28132 12679 28135
rect 13630 28132 13636 28144
rect 12667 28104 13636 28132
rect 12667 28101 12679 28104
rect 12621 28095 12679 28101
rect 13630 28092 13636 28104
rect 13688 28092 13694 28144
rect 24121 28135 24179 28141
rect 24121 28101 24133 28135
rect 24167 28132 24179 28135
rect 33229 28135 33287 28141
rect 24167 28104 25544 28132
rect 24167 28101 24179 28104
rect 24121 28095 24179 28101
rect 25516 28076 25544 28104
rect 33229 28101 33241 28135
rect 33275 28132 33287 28135
rect 34514 28132 34520 28144
rect 33275 28104 34520 28132
rect 33275 28101 33287 28104
rect 33229 28095 33287 28101
rect 34514 28092 34520 28104
rect 34572 28092 34578 28144
rect 1946 28024 1952 28076
rect 2004 28064 2010 28076
rect 2317 28067 2375 28073
rect 2317 28064 2329 28067
rect 2004 28036 2329 28064
rect 2004 28024 2010 28036
rect 2317 28033 2329 28036
rect 2363 28033 2375 28067
rect 5350 28064 5356 28076
rect 5311 28036 5356 28064
rect 2317 28027 2375 28033
rect 5350 28024 5356 28036
rect 5408 28064 5414 28076
rect 6181 28067 6239 28073
rect 6181 28064 6193 28067
rect 5408 28036 6193 28064
rect 5408 28024 5414 28036
rect 6181 28033 6193 28036
rect 6227 28033 6239 28067
rect 8110 28064 8116 28076
rect 8071 28036 8116 28064
rect 6181 28027 6239 28033
rect 8110 28024 8116 28036
rect 8168 28024 8174 28076
rect 14369 28067 14427 28073
rect 14369 28033 14381 28067
rect 14415 28064 14427 28067
rect 15102 28064 15108 28076
rect 14415 28036 15108 28064
rect 14415 28033 14427 28036
rect 14369 28027 14427 28033
rect 15102 28024 15108 28036
rect 15160 28024 15166 28076
rect 15838 28024 15844 28076
rect 15896 28064 15902 28076
rect 16117 28067 16175 28073
rect 16117 28064 16129 28067
rect 15896 28036 16129 28064
rect 15896 28024 15902 28036
rect 16117 28033 16129 28036
rect 16163 28033 16175 28067
rect 16117 28027 16175 28033
rect 18509 28067 18567 28073
rect 18509 28033 18521 28067
rect 18555 28064 18567 28067
rect 19432 28067 19490 28073
rect 19432 28064 19444 28067
rect 18555 28036 19444 28064
rect 18555 28033 18567 28036
rect 18509 28027 18567 28033
rect 19076 28008 19104 28036
rect 19432 28033 19444 28036
rect 19478 28033 19490 28067
rect 19702 28064 19708 28076
rect 19663 28036 19708 28064
rect 19432 28027 19490 28033
rect 19702 28024 19708 28036
rect 19760 28024 19766 28076
rect 21174 28064 21180 28076
rect 21087 28036 21180 28064
rect 21174 28024 21180 28036
rect 21232 28064 21238 28076
rect 22281 28067 22339 28073
rect 22281 28064 22293 28067
rect 21232 28036 22293 28064
rect 21232 28024 21238 28036
rect 22281 28033 22293 28036
rect 22327 28064 22339 28067
rect 22462 28064 22468 28076
rect 22327 28036 22468 28064
rect 22327 28033 22339 28036
rect 22281 28027 22339 28033
rect 22462 28024 22468 28036
rect 22520 28064 22526 28076
rect 22649 28067 22707 28073
rect 22649 28064 22661 28067
rect 22520 28036 22661 28064
rect 22520 28024 22526 28036
rect 22649 28033 22661 28036
rect 22695 28033 22707 28067
rect 22649 28027 22707 28033
rect 24854 28024 24860 28076
rect 24912 28064 24918 28076
rect 25133 28067 25191 28073
rect 25133 28064 25145 28067
rect 24912 28036 25145 28064
rect 24912 28024 24918 28036
rect 25133 28033 25145 28036
rect 25179 28033 25191 28067
rect 25133 28027 25191 28033
rect 25498 28024 25504 28076
rect 25556 28064 25562 28076
rect 26053 28067 26111 28073
rect 26053 28064 26065 28067
rect 25556 28036 26065 28064
rect 25556 28024 25562 28036
rect 26053 28033 26065 28036
rect 26099 28064 26111 28067
rect 26099 28036 26280 28064
rect 26099 28033 26111 28036
rect 26053 28027 26111 28033
rect 5169 27999 5227 28005
rect 5169 27965 5181 27999
rect 5215 27996 5227 27999
rect 5442 27996 5448 28008
rect 5215 27968 5448 27996
rect 5215 27965 5227 27968
rect 5169 27959 5227 27965
rect 5442 27956 5448 27968
rect 5500 27996 5506 28008
rect 5813 27999 5871 28005
rect 5813 27996 5825 27999
rect 5500 27968 5825 27996
rect 5500 27956 5506 27968
rect 5813 27965 5825 27968
rect 5859 27965 5871 27999
rect 5813 27959 5871 27965
rect 8202 27956 8208 28008
rect 8260 27996 8266 28008
rect 9033 27999 9091 28005
rect 9033 27996 9045 27999
rect 8260 27968 9045 27996
rect 8260 27956 8266 27968
rect 9033 27965 9045 27968
rect 9079 27996 9091 27999
rect 9585 27999 9643 28005
rect 9585 27996 9597 27999
rect 9079 27968 9597 27996
rect 9079 27965 9091 27968
rect 9033 27959 9091 27965
rect 9585 27965 9597 27968
rect 9631 27965 9643 27999
rect 9585 27959 9643 27965
rect 12434 27956 12440 28008
rect 12492 27996 12498 28008
rect 12989 27999 13047 28005
rect 12989 27996 13001 27999
rect 12492 27968 13001 27996
rect 12492 27956 12498 27968
rect 12989 27965 13001 27968
rect 13035 27965 13047 27999
rect 12989 27959 13047 27965
rect 18874 27956 18880 28008
rect 18932 27996 18938 28008
rect 18969 27999 19027 28005
rect 18969 27996 18981 27999
rect 18932 27968 18981 27996
rect 18932 27956 18938 27968
rect 18969 27965 18981 27968
rect 19015 27965 19027 27999
rect 18969 27959 19027 27965
rect 19058 27956 19064 28008
rect 19116 27956 19122 28008
rect 19334 27956 19340 28008
rect 19392 27996 19398 28008
rect 19720 27996 19748 28024
rect 26142 27996 26148 28008
rect 19392 27968 19748 27996
rect 26103 27968 26148 27996
rect 19392 27956 19398 27968
rect 26142 27956 26148 27968
rect 26200 27956 26206 28008
rect 26252 27996 26280 28036
rect 30006 28024 30012 28076
rect 30064 28064 30070 28076
rect 30193 28067 30251 28073
rect 30193 28064 30205 28067
rect 30064 28036 30205 28064
rect 30064 28024 30070 28036
rect 30193 28033 30205 28036
rect 30239 28033 30251 28067
rect 30193 28027 30251 28033
rect 32950 28024 32956 28076
rect 33008 28064 33014 28076
rect 33781 28067 33839 28073
rect 33781 28064 33793 28067
rect 33008 28036 33793 28064
rect 33008 28024 33014 28036
rect 33781 28033 33793 28036
rect 33827 28033 33839 28067
rect 33781 28027 33839 28033
rect 26412 27999 26470 28005
rect 26412 27996 26424 27999
rect 26252 27968 26424 27996
rect 26412 27965 26424 27968
rect 26458 27996 26470 27999
rect 27890 27996 27896 28008
rect 26458 27968 27896 27996
rect 26458 27965 26470 27968
rect 26412 27959 26470 27965
rect 27890 27956 27896 27968
rect 27948 27956 27954 28008
rect 33137 27999 33195 28005
rect 33137 27965 33149 27999
rect 33183 27996 33195 27999
rect 33689 27999 33747 28005
rect 33689 27996 33701 27999
rect 33183 27968 33701 27996
rect 33183 27965 33195 27968
rect 33137 27959 33195 27965
rect 33689 27965 33701 27968
rect 33735 27996 33747 27999
rect 34716 27996 34744 28163
rect 34790 28160 34796 28172
rect 34848 28160 34854 28212
rect 34974 27996 34980 28008
rect 33735 27968 34744 27996
rect 34935 27968 34980 27996
rect 33735 27965 33747 27968
rect 33689 27959 33747 27965
rect 34974 27956 34980 27968
rect 35032 27956 35038 28008
rect 35066 27956 35072 28008
rect 35124 27996 35130 28008
rect 35244 27999 35302 28005
rect 35244 27996 35256 27999
rect 35124 27968 35256 27996
rect 35124 27956 35130 27968
rect 35244 27965 35256 27968
rect 35290 27996 35302 27999
rect 35986 27996 35992 28008
rect 35290 27968 35992 27996
rect 35290 27965 35302 27968
rect 35244 27959 35302 27965
rect 35986 27956 35992 27968
rect 36044 27956 36050 28008
rect 2225 27931 2283 27937
rect 2225 27897 2237 27931
rect 2271 27928 2283 27931
rect 2562 27931 2620 27937
rect 2562 27928 2574 27931
rect 2271 27900 2574 27928
rect 2271 27897 2283 27900
rect 2225 27891 2283 27897
rect 2562 27897 2574 27900
rect 2608 27928 2620 27931
rect 2682 27928 2688 27940
rect 2608 27900 2688 27928
rect 2608 27897 2620 27900
rect 2562 27891 2620 27897
rect 2682 27888 2688 27900
rect 2740 27888 2746 27940
rect 4341 27931 4399 27937
rect 4341 27897 4353 27931
rect 4387 27928 4399 27931
rect 4614 27928 4620 27940
rect 4387 27900 4620 27928
rect 4387 27897 4399 27900
rect 4341 27891 4399 27897
rect 4614 27888 4620 27900
rect 4672 27928 4678 27940
rect 4709 27931 4767 27937
rect 4709 27928 4721 27931
rect 4672 27900 4721 27928
rect 4672 27888 4678 27900
rect 4709 27897 4721 27900
rect 4755 27928 4767 27931
rect 7929 27931 7987 27937
rect 7929 27928 7941 27931
rect 4755 27900 5304 27928
rect 4755 27897 4767 27900
rect 4709 27891 4767 27897
rect 3697 27863 3755 27869
rect 3697 27829 3709 27863
rect 3743 27860 3755 27863
rect 4154 27860 4160 27872
rect 3743 27832 4160 27860
rect 3743 27829 3755 27832
rect 3697 27823 3755 27829
rect 4154 27820 4160 27832
rect 4212 27820 4218 27872
rect 5276 27869 5304 27900
rect 7300 27900 7941 27928
rect 7300 27872 7328 27900
rect 7929 27897 7941 27900
rect 7975 27897 7987 27931
rect 22005 27931 22063 27937
rect 22005 27928 22017 27931
rect 7929 27891 7987 27897
rect 21468 27900 22017 27928
rect 21468 27872 21496 27900
rect 22005 27897 22017 27900
rect 22051 27897 22063 27931
rect 22005 27891 22063 27897
rect 22097 27931 22155 27937
rect 22097 27897 22109 27931
rect 22143 27928 22155 27931
rect 23017 27931 23075 27937
rect 23017 27928 23029 27931
rect 22143 27900 23029 27928
rect 22143 27897 22155 27900
rect 22097 27891 22155 27897
rect 23017 27897 23029 27900
rect 23063 27897 23075 27931
rect 23017 27891 23075 27897
rect 24489 27931 24547 27937
rect 24489 27897 24501 27931
rect 24535 27928 24547 27931
rect 25041 27931 25099 27937
rect 25041 27928 25053 27931
rect 24535 27900 25053 27928
rect 24535 27897 24547 27900
rect 24489 27891 24547 27897
rect 25041 27897 25053 27900
rect 25087 27928 25099 27931
rect 26326 27928 26332 27940
rect 25087 27900 26332 27928
rect 25087 27897 25099 27900
rect 25041 27891 25099 27897
rect 5261 27863 5319 27869
rect 5261 27829 5273 27863
rect 5307 27860 5319 27863
rect 5442 27860 5448 27872
rect 5307 27832 5448 27860
rect 5307 27829 5319 27832
rect 5261 27823 5319 27829
rect 5442 27820 5448 27832
rect 5500 27820 5506 27872
rect 7282 27860 7288 27872
rect 7243 27832 7288 27860
rect 7282 27820 7288 27832
rect 7340 27820 7346 27872
rect 7466 27860 7472 27872
rect 7427 27832 7472 27860
rect 7466 27820 7472 27832
rect 7524 27820 7530 27872
rect 7558 27820 7564 27872
rect 7616 27860 7622 27872
rect 7837 27863 7895 27869
rect 7837 27860 7849 27863
rect 7616 27832 7849 27860
rect 7616 27820 7622 27832
rect 7837 27829 7849 27832
rect 7883 27829 7895 27863
rect 7837 27823 7895 27829
rect 11054 27820 11060 27872
rect 11112 27860 11118 27872
rect 11422 27860 11428 27872
rect 11112 27832 11428 27860
rect 11112 27820 11118 27832
rect 11422 27820 11428 27832
rect 11480 27820 11486 27872
rect 17954 27820 17960 27872
rect 18012 27860 18018 27872
rect 18877 27863 18935 27869
rect 18877 27860 18889 27863
rect 18012 27832 18889 27860
rect 18012 27820 18018 27832
rect 18877 27829 18889 27832
rect 18923 27860 18935 27863
rect 19435 27863 19493 27869
rect 19435 27860 19447 27863
rect 18923 27832 19447 27860
rect 18923 27829 18935 27832
rect 18877 27823 18935 27829
rect 19435 27829 19447 27832
rect 19481 27860 19493 27863
rect 20622 27860 20628 27872
rect 19481 27832 20628 27860
rect 19481 27829 19493 27832
rect 19435 27823 19493 27829
rect 20622 27820 20628 27832
rect 20680 27820 20686 27872
rect 20806 27860 20812 27872
rect 20767 27832 20812 27860
rect 20806 27820 20812 27832
rect 20864 27820 20870 27872
rect 21450 27860 21456 27872
rect 21411 27832 21456 27860
rect 21450 27820 21456 27832
rect 21508 27820 21514 27872
rect 21634 27820 21640 27872
rect 21692 27860 21698 27872
rect 22112 27860 22140 27891
rect 26326 27888 26332 27900
rect 26384 27888 26390 27940
rect 30101 27931 30159 27937
rect 30101 27897 30113 27931
rect 30147 27928 30159 27931
rect 30460 27931 30518 27937
rect 30460 27928 30472 27931
rect 30147 27900 30472 27928
rect 30147 27897 30159 27900
rect 30101 27891 30159 27897
rect 30460 27897 30472 27900
rect 30506 27928 30518 27931
rect 30926 27928 30932 27940
rect 30506 27900 30932 27928
rect 30506 27897 30518 27900
rect 30460 27891 30518 27897
rect 30926 27888 30932 27900
rect 30984 27888 30990 27940
rect 33318 27888 33324 27940
rect 33376 27928 33382 27940
rect 33597 27931 33655 27937
rect 33597 27928 33609 27931
rect 33376 27900 33609 27928
rect 33376 27888 33382 27900
rect 33597 27897 33609 27900
rect 33643 27928 33655 27931
rect 35084 27928 35112 27956
rect 33643 27900 35112 27928
rect 33643 27897 33655 27900
rect 33597 27891 33655 27897
rect 21692 27832 22140 27860
rect 21692 27820 21698 27832
rect 24578 27820 24584 27872
rect 24636 27860 24642 27872
rect 24949 27863 25007 27869
rect 24949 27860 24961 27863
rect 24636 27832 24961 27860
rect 24636 27820 24642 27832
rect 24949 27829 24961 27832
rect 24995 27829 25007 27863
rect 24949 27823 25007 27829
rect 27246 27820 27252 27872
rect 27304 27860 27310 27872
rect 27525 27863 27583 27869
rect 27525 27860 27537 27863
rect 27304 27832 27537 27860
rect 27304 27820 27310 27832
rect 27525 27829 27537 27832
rect 27571 27829 27583 27863
rect 27525 27823 27583 27829
rect 32769 27863 32827 27869
rect 32769 27829 32781 27863
rect 32815 27860 32827 27863
rect 32950 27860 32956 27872
rect 32815 27832 32956 27860
rect 32815 27829 32827 27832
rect 32769 27823 32827 27829
rect 32950 27820 32956 27832
rect 33008 27820 33014 27872
rect 34330 27860 34336 27872
rect 34243 27832 34336 27860
rect 34330 27820 34336 27832
rect 34388 27860 34394 27872
rect 34974 27860 34980 27872
rect 34388 27832 34980 27860
rect 34388 27820 34394 27832
rect 34974 27820 34980 27832
rect 35032 27820 35038 27872
rect 36354 27860 36360 27872
rect 36315 27832 36360 27860
rect 36354 27820 36360 27832
rect 36412 27820 36418 27872
rect 1104 27770 38824 27792
rect 1104 27718 19606 27770
rect 19658 27718 19670 27770
rect 19722 27718 19734 27770
rect 19786 27718 19798 27770
rect 19850 27718 38824 27770
rect 1104 27696 38824 27718
rect 1854 27616 1860 27668
rect 1912 27656 1918 27668
rect 2133 27659 2191 27665
rect 2133 27656 2145 27659
rect 1912 27628 2145 27656
rect 1912 27616 1918 27628
rect 2133 27625 2145 27628
rect 2179 27625 2191 27659
rect 2133 27619 2191 27625
rect 2774 27616 2780 27668
rect 2832 27656 2838 27668
rect 3145 27659 3203 27665
rect 3145 27656 3157 27659
rect 2832 27628 3157 27656
rect 2832 27616 2838 27628
rect 3145 27625 3157 27628
rect 3191 27656 3203 27659
rect 4062 27656 4068 27668
rect 3191 27628 4068 27656
rect 3191 27625 3203 27628
rect 3145 27619 3203 27625
rect 4062 27616 4068 27628
rect 4120 27616 4126 27668
rect 5442 27656 5448 27668
rect 5403 27628 5448 27656
rect 5442 27616 5448 27628
rect 5500 27616 5506 27668
rect 7466 27616 7472 27668
rect 7524 27656 7530 27668
rect 11146 27656 11152 27668
rect 7524 27628 8248 27656
rect 11107 27628 11152 27656
rect 7524 27616 7530 27628
rect 2222 27548 2228 27600
rect 2280 27588 2286 27600
rect 3878 27588 3884 27600
rect 2280 27560 2728 27588
rect 3839 27560 3884 27588
rect 2280 27548 2286 27560
rect 1949 27523 2007 27529
rect 1949 27489 1961 27523
rect 1995 27520 2007 27523
rect 2130 27520 2136 27532
rect 1995 27492 2136 27520
rect 1995 27489 2007 27492
rect 1949 27483 2007 27489
rect 2130 27480 2136 27492
rect 2188 27520 2194 27532
rect 2501 27523 2559 27529
rect 2501 27520 2513 27523
rect 2188 27492 2513 27520
rect 2188 27480 2194 27492
rect 2501 27489 2513 27492
rect 2547 27489 2559 27523
rect 2501 27483 2559 27489
rect 2700 27520 2728 27560
rect 3878 27548 3884 27560
rect 3936 27548 3942 27600
rect 4154 27548 4160 27600
rect 4212 27588 4218 27600
rect 4310 27591 4368 27597
rect 4310 27588 4322 27591
rect 4212 27560 4322 27588
rect 4212 27548 4218 27560
rect 4310 27557 4322 27560
rect 4356 27588 4368 27591
rect 4614 27588 4620 27600
rect 4356 27560 4620 27588
rect 4356 27557 4368 27560
rect 4310 27551 4368 27557
rect 4614 27548 4620 27560
rect 4672 27548 4678 27600
rect 7929 27591 7987 27597
rect 7929 27557 7941 27591
rect 7975 27588 7987 27591
rect 8110 27588 8116 27600
rect 7975 27560 8116 27588
rect 7975 27557 7987 27560
rect 7929 27551 7987 27557
rect 8110 27548 8116 27560
rect 8168 27548 8174 27600
rect 8220 27588 8248 27628
rect 11146 27616 11152 27628
rect 11204 27616 11210 27668
rect 14366 27656 14372 27668
rect 13832 27628 14372 27656
rect 8389 27591 8447 27597
rect 8389 27588 8401 27591
rect 8220 27560 8401 27588
rect 8389 27557 8401 27560
rect 8435 27588 8447 27591
rect 9214 27588 9220 27600
rect 8435 27560 9220 27588
rect 8435 27557 8447 27560
rect 8389 27551 8447 27557
rect 9214 27548 9220 27560
rect 9272 27548 9278 27600
rect 13446 27548 13452 27600
rect 13504 27588 13510 27600
rect 13541 27591 13599 27597
rect 13541 27588 13553 27591
rect 13504 27560 13553 27588
rect 13504 27548 13510 27560
rect 13541 27557 13553 27560
rect 13587 27588 13599 27591
rect 13832 27588 13860 27628
rect 14366 27616 14372 27628
rect 14424 27616 14430 27668
rect 19334 27656 19340 27668
rect 19295 27628 19340 27656
rect 19334 27616 19340 27628
rect 19392 27616 19398 27668
rect 21450 27656 21456 27668
rect 20640 27628 21456 27656
rect 13587 27560 13860 27588
rect 15832 27591 15890 27597
rect 13587 27557 13599 27560
rect 13541 27551 13599 27557
rect 15832 27557 15844 27591
rect 15878 27588 15890 27591
rect 16022 27588 16028 27600
rect 15878 27560 16028 27588
rect 15878 27557 15890 27560
rect 15832 27551 15890 27557
rect 16022 27548 16028 27560
rect 16080 27548 16086 27600
rect 18966 27588 18972 27600
rect 18927 27560 18972 27588
rect 18966 27548 18972 27560
rect 19024 27548 19030 27600
rect 19797 27591 19855 27597
rect 19797 27557 19809 27591
rect 19843 27588 19855 27591
rect 20640 27588 20668 27628
rect 21450 27616 21456 27628
rect 21508 27616 21514 27668
rect 22462 27656 22468 27668
rect 22423 27628 22468 27656
rect 22462 27616 22468 27628
rect 22520 27616 22526 27668
rect 26142 27616 26148 27668
rect 26200 27656 26206 27668
rect 29457 27659 29515 27665
rect 26200 27628 26372 27656
rect 26200 27616 26206 27628
rect 19843 27560 20668 27588
rect 19843 27557 19855 27560
rect 19797 27551 19855 27557
rect 20714 27548 20720 27600
rect 20772 27588 20778 27600
rect 20898 27588 20904 27600
rect 20772 27560 20904 27588
rect 20772 27548 20778 27560
rect 20898 27548 20904 27560
rect 20956 27588 20962 27600
rect 24305 27591 24363 27597
rect 20956 27560 21128 27588
rect 20956 27548 20962 27560
rect 5350 27520 5356 27532
rect 2700 27492 5356 27520
rect 1762 27412 1768 27464
rect 1820 27452 1826 27464
rect 2700 27461 2728 27492
rect 5350 27480 5356 27492
rect 5408 27480 5414 27532
rect 8481 27523 8539 27529
rect 8481 27489 8493 27523
rect 8527 27520 8539 27523
rect 8846 27520 8852 27532
rect 8527 27492 8852 27520
rect 8527 27489 8539 27492
rect 8481 27483 8539 27489
rect 8846 27480 8852 27492
rect 8904 27480 8910 27532
rect 10965 27523 11023 27529
rect 10965 27489 10977 27523
rect 11011 27520 11023 27523
rect 11054 27520 11060 27532
rect 11011 27492 11060 27520
rect 11011 27489 11023 27492
rect 10965 27483 11023 27489
rect 11054 27480 11060 27492
rect 11112 27480 11118 27532
rect 21100 27529 21128 27560
rect 24305 27557 24317 27591
rect 24351 27588 24363 27591
rect 24762 27588 24768 27600
rect 24351 27560 24768 27588
rect 24351 27557 24363 27560
rect 24305 27551 24363 27557
rect 24762 27548 24768 27560
rect 24820 27548 24826 27600
rect 21085 27523 21143 27529
rect 21085 27489 21097 27523
rect 21131 27489 21143 27523
rect 21085 27483 21143 27489
rect 21352 27523 21410 27529
rect 21352 27489 21364 27523
rect 21398 27520 21410 27523
rect 21726 27520 21732 27532
rect 21398 27492 21732 27520
rect 21398 27489 21410 27492
rect 21352 27483 21410 27489
rect 21726 27480 21732 27492
rect 21784 27480 21790 27532
rect 25130 27480 25136 27532
rect 25188 27520 25194 27532
rect 25225 27523 25283 27529
rect 25225 27520 25237 27523
rect 25188 27492 25237 27520
rect 25188 27480 25194 27492
rect 25225 27489 25237 27492
rect 25271 27489 25283 27523
rect 25225 27483 25283 27489
rect 25317 27523 25375 27529
rect 25317 27489 25329 27523
rect 25363 27520 25375 27523
rect 25406 27520 25412 27532
rect 25363 27492 25412 27520
rect 25363 27489 25375 27492
rect 25317 27483 25375 27489
rect 25406 27480 25412 27492
rect 25464 27520 25470 27532
rect 26142 27520 26148 27532
rect 25464 27492 26148 27520
rect 25464 27480 25470 27492
rect 26142 27480 26148 27492
rect 26200 27480 26206 27532
rect 2593 27455 2651 27461
rect 2593 27452 2605 27455
rect 1820 27424 2605 27452
rect 1820 27412 1826 27424
rect 2593 27421 2605 27424
rect 2639 27421 2651 27455
rect 2593 27415 2651 27421
rect 2685 27455 2743 27461
rect 2685 27421 2697 27455
rect 2731 27421 2743 27455
rect 2685 27415 2743 27421
rect 4065 27455 4123 27461
rect 4065 27421 4077 27455
rect 4111 27421 4123 27455
rect 8662 27452 8668 27464
rect 8623 27424 8668 27452
rect 4065 27415 4123 27421
rect 1946 27344 1952 27396
rect 2004 27384 2010 27396
rect 3970 27384 3976 27396
rect 2004 27356 3976 27384
rect 2004 27344 2010 27356
rect 3970 27344 3976 27356
rect 4028 27384 4034 27396
rect 4080 27384 4108 27415
rect 8662 27412 8668 27424
rect 8720 27412 8726 27464
rect 15562 27452 15568 27464
rect 15523 27424 15568 27452
rect 15562 27412 15568 27424
rect 15620 27412 15626 27464
rect 25498 27452 25504 27464
rect 25459 27424 25504 27452
rect 25498 27412 25504 27424
rect 25556 27412 25562 27464
rect 26344 27461 26372 27628
rect 29457 27625 29469 27659
rect 29503 27656 29515 27659
rect 29822 27656 29828 27668
rect 29503 27628 29828 27656
rect 29503 27625 29515 27628
rect 29457 27619 29515 27625
rect 29822 27616 29828 27628
rect 29880 27656 29886 27668
rect 30006 27656 30012 27668
rect 29880 27628 30012 27656
rect 29880 27616 29886 27628
rect 30006 27616 30012 27628
rect 30064 27616 30070 27668
rect 30466 27616 30472 27668
rect 30524 27656 30530 27668
rect 33318 27656 33324 27668
rect 30524 27628 31708 27656
rect 33279 27628 33324 27656
rect 30524 27616 30530 27628
rect 31680 27588 31708 27628
rect 33318 27616 33324 27628
rect 33376 27616 33382 27668
rect 35066 27656 35072 27668
rect 35027 27628 35072 27656
rect 35066 27616 35072 27628
rect 35124 27616 35130 27668
rect 32582 27588 32588 27600
rect 31680 27560 32588 27588
rect 32582 27548 32588 27560
rect 32640 27548 32646 27600
rect 26780 27523 26838 27529
rect 26780 27489 26792 27523
rect 26826 27520 26838 27523
rect 27246 27520 27252 27532
rect 26826 27492 27252 27520
rect 26826 27489 26838 27492
rect 26780 27483 26838 27489
rect 27246 27480 27252 27492
rect 27304 27480 27310 27532
rect 29086 27480 29092 27532
rect 29144 27520 29150 27532
rect 29805 27523 29863 27529
rect 29805 27520 29817 27523
rect 29144 27492 29817 27520
rect 29144 27480 29150 27492
rect 29805 27489 29817 27492
rect 29851 27520 29863 27523
rect 30742 27520 30748 27532
rect 29851 27492 30748 27520
rect 29851 27489 29863 27492
rect 29805 27483 29863 27489
rect 30742 27480 30748 27492
rect 30800 27480 30806 27532
rect 32490 27520 32496 27532
rect 32451 27492 32496 27520
rect 32490 27480 32496 27492
rect 32548 27480 32554 27532
rect 34057 27523 34115 27529
rect 34057 27489 34069 27523
rect 34103 27520 34115 27523
rect 34146 27520 34152 27532
rect 34103 27492 34152 27520
rect 34103 27489 34115 27492
rect 34057 27483 34115 27489
rect 34146 27480 34152 27492
rect 34204 27520 34210 27532
rect 34606 27520 34612 27532
rect 34204 27492 34612 27520
rect 34204 27480 34210 27492
rect 34606 27480 34612 27492
rect 34664 27480 34670 27532
rect 35428 27523 35486 27529
rect 35428 27489 35440 27523
rect 35474 27520 35486 27523
rect 36354 27520 36360 27532
rect 35474 27492 36360 27520
rect 35474 27489 35486 27492
rect 35428 27483 35486 27489
rect 36354 27480 36360 27492
rect 36412 27480 36418 27532
rect 26329 27455 26387 27461
rect 26329 27421 26341 27455
rect 26375 27452 26387 27455
rect 26510 27452 26516 27464
rect 26375 27424 26516 27452
rect 26375 27421 26387 27424
rect 26329 27415 26387 27421
rect 26510 27412 26516 27424
rect 26568 27412 26574 27464
rect 29546 27452 29552 27464
rect 29507 27424 29552 27452
rect 29546 27412 29552 27424
rect 29604 27412 29610 27464
rect 32677 27455 32735 27461
rect 32677 27452 32689 27455
rect 31864 27424 32689 27452
rect 4028 27356 4108 27384
rect 8021 27387 8079 27393
rect 4028 27344 4034 27356
rect 8021 27353 8033 27387
rect 8067 27384 8079 27387
rect 8202 27384 8208 27396
rect 8067 27356 8208 27384
rect 8067 27353 8079 27356
rect 8021 27347 8079 27353
rect 8202 27344 8208 27356
rect 8260 27344 8266 27396
rect 18601 27387 18659 27393
rect 18601 27353 18613 27387
rect 18647 27384 18659 27387
rect 18874 27384 18880 27396
rect 18647 27356 18880 27384
rect 18647 27353 18659 27356
rect 18601 27347 18659 27353
rect 18874 27344 18880 27356
rect 18932 27384 18938 27396
rect 20346 27384 20352 27396
rect 18932 27356 20352 27384
rect 18932 27344 18938 27356
rect 20346 27344 20352 27356
rect 20404 27344 20410 27396
rect 24857 27387 24915 27393
rect 24857 27353 24869 27387
rect 24903 27384 24915 27387
rect 24946 27384 24952 27396
rect 24903 27356 24952 27384
rect 24903 27353 24915 27356
rect 24857 27347 24915 27353
rect 24946 27344 24952 27356
rect 25004 27344 25010 27396
rect 27890 27384 27896 27396
rect 27851 27356 27896 27384
rect 27890 27344 27896 27356
rect 27948 27344 27954 27396
rect 7193 27319 7251 27325
rect 7193 27285 7205 27319
rect 7239 27316 7251 27319
rect 7558 27316 7564 27328
rect 7239 27288 7564 27316
rect 7239 27285 7251 27288
rect 7193 27279 7251 27285
rect 7558 27276 7564 27288
rect 7616 27276 7622 27328
rect 16942 27316 16948 27328
rect 16903 27288 16948 27316
rect 16942 27276 16948 27288
rect 17000 27276 17006 27328
rect 19705 27319 19763 27325
rect 19705 27285 19717 27319
rect 19751 27316 19763 27319
rect 19978 27316 19984 27328
rect 19751 27288 19984 27316
rect 19751 27285 19763 27288
rect 19705 27279 19763 27285
rect 19978 27276 19984 27288
rect 20036 27276 20042 27328
rect 24578 27316 24584 27328
rect 24539 27288 24584 27316
rect 24578 27276 24584 27288
rect 24636 27276 24642 27328
rect 25222 27276 25228 27328
rect 25280 27316 25286 27328
rect 25869 27319 25927 27325
rect 25869 27316 25881 27319
rect 25280 27288 25881 27316
rect 25280 27276 25286 27288
rect 25869 27285 25881 27288
rect 25915 27285 25927 27319
rect 30926 27316 30932 27328
rect 30887 27288 30932 27316
rect 25869 27279 25927 27285
rect 30926 27276 30932 27288
rect 30984 27276 30990 27328
rect 31570 27276 31576 27328
rect 31628 27316 31634 27328
rect 31864 27325 31892 27424
rect 32677 27421 32689 27424
rect 32723 27452 32735 27455
rect 34698 27452 34704 27464
rect 32723 27424 34704 27452
rect 32723 27421 32735 27424
rect 32677 27415 32735 27421
rect 34698 27412 34704 27424
rect 34756 27412 34762 27464
rect 34974 27412 34980 27464
rect 35032 27452 35038 27464
rect 35161 27455 35219 27461
rect 35161 27452 35173 27455
rect 35032 27424 35173 27452
rect 35032 27412 35038 27424
rect 35161 27421 35173 27424
rect 35207 27421 35219 27455
rect 35161 27415 35219 27421
rect 31849 27319 31907 27325
rect 31849 27316 31861 27319
rect 31628 27288 31861 27316
rect 31628 27276 31634 27288
rect 31849 27285 31861 27288
rect 31895 27285 31907 27319
rect 32122 27316 32128 27328
rect 32083 27288 32128 27316
rect 31849 27279 31907 27285
rect 32122 27276 32128 27288
rect 32180 27276 32186 27328
rect 34238 27316 34244 27328
rect 34199 27288 34244 27316
rect 34238 27276 34244 27288
rect 34296 27276 34302 27328
rect 35176 27316 35204 27415
rect 35526 27316 35532 27328
rect 35176 27288 35532 27316
rect 35526 27276 35532 27288
rect 35584 27276 35590 27328
rect 36541 27319 36599 27325
rect 36541 27285 36553 27319
rect 36587 27316 36599 27319
rect 36814 27316 36820 27328
rect 36587 27288 36820 27316
rect 36587 27285 36599 27288
rect 36541 27279 36599 27285
rect 36814 27276 36820 27288
rect 36872 27276 36878 27328
rect 1104 27226 38824 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 34966 27226
rect 35018 27174 35030 27226
rect 35082 27174 35094 27226
rect 35146 27174 35158 27226
rect 35210 27174 38824 27226
rect 1104 27152 38824 27174
rect 1762 27112 1768 27124
rect 1723 27084 1768 27112
rect 1762 27072 1768 27084
rect 1820 27072 1826 27124
rect 2774 27072 2780 27124
rect 2832 27112 2838 27124
rect 3237 27115 3295 27121
rect 3237 27112 3249 27115
rect 2832 27084 3249 27112
rect 2832 27072 2838 27084
rect 3237 27081 3249 27084
rect 3283 27112 3295 27115
rect 4157 27115 4215 27121
rect 4157 27112 4169 27115
rect 3283 27084 4169 27112
rect 3283 27081 3295 27084
rect 3237 27075 3295 27081
rect 4157 27081 4169 27084
rect 4203 27112 4215 27115
rect 5350 27112 5356 27124
rect 4203 27084 4844 27112
rect 5311 27084 5356 27112
rect 4203 27081 4215 27084
rect 4157 27075 4215 27081
rect 4062 27004 4068 27056
rect 4120 27044 4126 27056
rect 4341 27047 4399 27053
rect 4341 27044 4353 27047
rect 4120 27016 4353 27044
rect 4120 27004 4126 27016
rect 4341 27013 4353 27016
rect 4387 27013 4399 27047
rect 4341 27007 4399 27013
rect 4816 26985 4844 27084
rect 5350 27072 5356 27084
rect 5408 27072 5414 27124
rect 5718 27112 5724 27124
rect 5679 27084 5724 27112
rect 5718 27072 5724 27084
rect 5776 27112 5782 27124
rect 6181 27115 6239 27121
rect 6181 27112 6193 27115
rect 5776 27084 6193 27112
rect 5776 27072 5782 27084
rect 6181 27081 6193 27084
rect 6227 27081 6239 27115
rect 6181 27075 6239 27081
rect 4801 26979 4859 26985
rect 4801 26945 4813 26979
rect 4847 26945 4859 26979
rect 4801 26939 4859 26945
rect 4985 26979 5043 26985
rect 4985 26945 4997 26979
rect 5031 26976 5043 26979
rect 5368 26976 5396 27072
rect 5031 26948 5396 26976
rect 6196 26976 6224 27075
rect 7558 27072 7564 27124
rect 7616 27112 7622 27124
rect 8297 27115 8355 27121
rect 8297 27112 8309 27115
rect 7616 27084 8309 27112
rect 7616 27072 7622 27084
rect 8297 27081 8309 27084
rect 8343 27081 8355 27115
rect 9214 27112 9220 27124
rect 9175 27084 9220 27112
rect 8297 27075 8355 27081
rect 9214 27072 9220 27084
rect 9272 27072 9278 27124
rect 10229 27115 10287 27121
rect 10229 27081 10241 27115
rect 10275 27112 10287 27115
rect 10962 27112 10968 27124
rect 10275 27084 10968 27112
rect 10275 27081 10287 27084
rect 10229 27075 10287 27081
rect 10962 27072 10968 27084
rect 11020 27072 11026 27124
rect 15657 27115 15715 27121
rect 15657 27081 15669 27115
rect 15703 27112 15715 27115
rect 16022 27112 16028 27124
rect 15703 27084 16028 27112
rect 15703 27081 15715 27084
rect 15657 27075 15715 27081
rect 16022 27072 16028 27084
rect 16080 27072 16086 27124
rect 18690 27112 18696 27124
rect 18651 27084 18696 27112
rect 18690 27072 18696 27084
rect 18748 27072 18754 27124
rect 21177 27115 21235 27121
rect 21177 27081 21189 27115
rect 21223 27112 21235 27115
rect 21634 27112 21640 27124
rect 21223 27084 21640 27112
rect 21223 27081 21235 27084
rect 21177 27075 21235 27081
rect 21634 27072 21640 27084
rect 21692 27072 21698 27124
rect 24213 27115 24271 27121
rect 24213 27081 24225 27115
rect 24259 27112 24271 27115
rect 25406 27112 25412 27124
rect 24259 27084 25412 27112
rect 24259 27081 24271 27084
rect 24213 27075 24271 27081
rect 25406 27072 25412 27084
rect 25464 27072 25470 27124
rect 29086 27112 29092 27124
rect 29047 27084 29092 27112
rect 29086 27072 29092 27084
rect 29144 27072 29150 27124
rect 32582 27072 32588 27124
rect 32640 27112 32646 27124
rect 33321 27115 33379 27121
rect 33321 27112 33333 27115
rect 32640 27084 33333 27112
rect 32640 27072 32646 27084
rect 33321 27081 33333 27084
rect 33367 27081 33379 27115
rect 34146 27112 34152 27124
rect 34107 27084 34152 27112
rect 33321 27075 33379 27081
rect 34146 27072 34152 27084
rect 34204 27072 34210 27124
rect 34514 27072 34520 27124
rect 34572 27112 34578 27124
rect 34609 27115 34667 27121
rect 34609 27112 34621 27115
rect 34572 27084 34621 27112
rect 34572 27072 34578 27084
rect 34609 27081 34621 27084
rect 34655 27081 34667 27115
rect 34609 27075 34667 27081
rect 35989 27115 36047 27121
rect 35989 27081 36001 27115
rect 36035 27112 36047 27115
rect 36354 27112 36360 27124
rect 36035 27084 36360 27112
rect 36035 27081 36047 27084
rect 35989 27075 36047 27081
rect 8662 27004 8668 27056
rect 8720 27044 8726 27056
rect 9585 27047 9643 27053
rect 9585 27044 9597 27047
rect 8720 27016 9597 27044
rect 8720 27004 8726 27016
rect 9585 27013 9597 27016
rect 9631 27044 9643 27047
rect 9858 27044 9864 27056
rect 9631 27016 9864 27044
rect 9631 27013 9643 27016
rect 9585 27007 9643 27013
rect 9858 27004 9864 27016
rect 9916 27044 9922 27056
rect 11330 27044 11336 27056
rect 9916 27016 11336 27044
rect 9916 27004 9922 27016
rect 11330 27004 11336 27016
rect 11388 27004 11394 27056
rect 26510 27004 26516 27056
rect 26568 27044 26574 27056
rect 27617 27047 27675 27053
rect 27617 27044 27629 27047
rect 26568 27016 27629 27044
rect 26568 27004 26574 27016
rect 27617 27013 27629 27016
rect 27663 27044 27675 27047
rect 29546 27044 29552 27056
rect 27663 27016 29552 27044
rect 27663 27013 27675 27016
rect 27617 27007 27675 27013
rect 29546 27004 29552 27016
rect 29604 27004 29610 27056
rect 32309 27047 32367 27053
rect 32309 27013 32321 27047
rect 32355 27044 32367 27047
rect 32490 27044 32496 27056
rect 32355 27016 32496 27044
rect 32355 27013 32367 27016
rect 32309 27007 32367 27013
rect 32490 27004 32496 27016
rect 32548 27044 32554 27056
rect 33689 27047 33747 27053
rect 33689 27044 33701 27047
rect 32548 27016 33701 27044
rect 32548 27004 32554 27016
rect 33689 27013 33701 27016
rect 33735 27013 33747 27047
rect 33689 27007 33747 27013
rect 6914 26976 6920 26988
rect 6196 26948 6920 26976
rect 5031 26945 5043 26948
rect 4985 26939 5043 26945
rect 6914 26936 6920 26948
rect 6972 26936 6978 26988
rect 13357 26979 13415 26985
rect 13357 26945 13369 26979
rect 13403 26976 13415 26979
rect 13403 26948 13584 26976
rect 13403 26945 13415 26948
rect 13357 26939 13415 26945
rect 1486 26868 1492 26920
rect 1544 26908 1550 26920
rect 1857 26911 1915 26917
rect 1857 26908 1869 26911
rect 1544 26880 1869 26908
rect 1544 26868 1550 26880
rect 1857 26877 1869 26880
rect 1903 26908 1915 26911
rect 1946 26908 1952 26920
rect 1903 26880 1952 26908
rect 1903 26877 1915 26880
rect 1857 26871 1915 26877
rect 1946 26868 1952 26880
rect 2004 26868 2010 26920
rect 2130 26917 2136 26920
rect 2124 26908 2136 26917
rect 2091 26880 2136 26908
rect 2124 26871 2136 26880
rect 2188 26908 2194 26920
rect 3789 26911 3847 26917
rect 3789 26908 3801 26911
rect 2188 26880 3801 26908
rect 2130 26868 2136 26871
rect 2188 26868 2194 26880
rect 3789 26877 3801 26880
rect 3835 26877 3847 26911
rect 3789 26871 3847 26877
rect 4614 26868 4620 26920
rect 4672 26908 4678 26920
rect 4709 26911 4767 26917
rect 4709 26908 4721 26911
rect 4672 26880 4721 26908
rect 4672 26868 4678 26880
rect 4709 26877 4721 26880
rect 4755 26877 4767 26911
rect 4709 26871 4767 26877
rect 9674 26868 9680 26920
rect 9732 26908 9738 26920
rect 10045 26911 10103 26917
rect 10045 26908 10057 26911
rect 9732 26880 10057 26908
rect 9732 26868 9738 26880
rect 10045 26877 10057 26880
rect 10091 26908 10103 26911
rect 10597 26911 10655 26917
rect 10597 26908 10609 26911
rect 10091 26880 10609 26908
rect 10091 26877 10103 26880
rect 10045 26871 10103 26877
rect 10597 26877 10609 26880
rect 10643 26877 10655 26911
rect 13446 26908 13452 26920
rect 13407 26880 13452 26908
rect 10597 26871 10655 26877
rect 13446 26868 13452 26880
rect 13504 26868 13510 26920
rect 13556 26908 13584 26948
rect 15562 26936 15568 26988
rect 15620 26976 15626 26988
rect 16025 26979 16083 26985
rect 16025 26976 16037 26979
rect 15620 26948 16037 26976
rect 15620 26936 15626 26948
rect 16025 26945 16037 26948
rect 16071 26976 16083 26979
rect 17126 26976 17132 26988
rect 16071 26948 17132 26976
rect 16071 26945 16083 26948
rect 16025 26939 16083 26945
rect 17126 26936 17132 26948
rect 17184 26936 17190 26988
rect 21726 26976 21732 26988
rect 21687 26948 21732 26976
rect 21726 26936 21732 26948
rect 21784 26976 21790 26988
rect 22278 26976 22284 26988
rect 21784 26948 22284 26976
rect 21784 26936 21790 26948
rect 22278 26936 22284 26948
rect 22336 26936 22342 26988
rect 24949 26979 25007 26985
rect 24949 26945 24961 26979
rect 24995 26976 25007 26979
rect 25130 26976 25136 26988
rect 24995 26948 25136 26976
rect 24995 26945 25007 26948
rect 24949 26939 25007 26945
rect 25130 26936 25136 26948
rect 25188 26976 25194 26988
rect 29822 26976 29828 26988
rect 25188 26948 25360 26976
rect 29783 26948 29828 26976
rect 25188 26936 25194 26948
rect 13722 26917 13728 26920
rect 13716 26908 13728 26917
rect 13556 26880 13728 26908
rect 13716 26871 13728 26880
rect 13722 26868 13728 26871
rect 13780 26868 13786 26920
rect 18049 26911 18107 26917
rect 18049 26877 18061 26911
rect 18095 26908 18107 26911
rect 18690 26908 18696 26920
rect 18095 26880 18696 26908
rect 18095 26877 18107 26880
rect 18049 26871 18107 26877
rect 18690 26868 18696 26880
rect 18748 26868 18754 26920
rect 25222 26908 25228 26920
rect 25183 26880 25228 26908
rect 25222 26868 25228 26880
rect 25280 26868 25286 26920
rect 25332 26908 25360 26948
rect 29822 26936 29828 26948
rect 29880 26936 29886 26988
rect 32217 26979 32275 26985
rect 32217 26945 32229 26979
rect 32263 26976 32275 26979
rect 32674 26976 32680 26988
rect 32263 26948 32680 26976
rect 32263 26945 32275 26948
rect 32217 26939 32275 26945
rect 32674 26936 32680 26948
rect 32732 26976 32738 26988
rect 32769 26979 32827 26985
rect 32769 26976 32781 26979
rect 32732 26948 32781 26976
rect 32732 26936 32738 26948
rect 32769 26945 32781 26948
rect 32815 26945 32827 26979
rect 32950 26976 32956 26988
rect 32911 26948 32956 26976
rect 32769 26939 32827 26945
rect 32950 26936 32956 26948
rect 33008 26936 33014 26988
rect 27709 26911 27767 26917
rect 27709 26908 27721 26911
rect 25332 26880 27721 26908
rect 27709 26877 27721 26880
rect 27755 26877 27767 26911
rect 34624 26908 34652 27075
rect 36354 27072 36360 27084
rect 36412 27072 36418 27124
rect 34698 26936 34704 26988
rect 34756 26976 34762 26988
rect 35437 26979 35495 26985
rect 35437 26976 35449 26979
rect 34756 26948 35449 26976
rect 34756 26936 34762 26948
rect 35437 26945 35449 26948
rect 35483 26945 35495 26979
rect 36998 26976 37004 26988
rect 36959 26948 37004 26976
rect 35437 26939 35495 26945
rect 36998 26936 37004 26948
rect 37056 26936 37062 26988
rect 35345 26911 35403 26917
rect 35345 26908 35357 26911
rect 34624 26880 35357 26908
rect 27709 26871 27767 26877
rect 35345 26877 35357 26880
rect 35391 26877 35403 26911
rect 35345 26871 35403 26877
rect 36354 26868 36360 26920
rect 36412 26908 36418 26920
rect 36909 26911 36967 26917
rect 36909 26908 36921 26911
rect 36412 26880 36921 26908
rect 36412 26868 36418 26880
rect 36909 26877 36921 26880
rect 36955 26877 36967 26911
rect 36909 26871 36967 26877
rect 6641 26843 6699 26849
rect 6641 26809 6653 26843
rect 6687 26840 6699 26843
rect 7184 26843 7242 26849
rect 7184 26840 7196 26843
rect 6687 26812 7196 26840
rect 6687 26809 6699 26812
rect 6641 26803 6699 26809
rect 7184 26809 7196 26812
rect 7230 26840 7242 26843
rect 7282 26840 7288 26852
rect 7230 26812 7288 26840
rect 7230 26809 7242 26812
rect 7184 26803 7242 26809
rect 7282 26800 7288 26812
rect 7340 26840 7346 26852
rect 8202 26840 8208 26852
rect 7340 26812 8208 26840
rect 7340 26800 7346 26812
rect 8202 26800 8208 26812
rect 8260 26800 8266 26852
rect 21085 26843 21143 26849
rect 21085 26809 21097 26843
rect 21131 26840 21143 26843
rect 21637 26843 21695 26849
rect 21637 26840 21649 26843
rect 21131 26812 21649 26840
rect 21131 26809 21143 26812
rect 21085 26803 21143 26809
rect 21637 26809 21649 26812
rect 21683 26840 21695 26843
rect 21910 26840 21916 26852
rect 21683 26812 21916 26840
rect 21683 26809 21695 26812
rect 21637 26803 21695 26809
rect 21910 26800 21916 26812
rect 21968 26800 21974 26852
rect 25498 26849 25504 26852
rect 24581 26843 24639 26849
rect 24581 26809 24593 26843
rect 24627 26840 24639 26843
rect 25492 26840 25504 26849
rect 24627 26812 25504 26840
rect 24627 26809 24639 26812
rect 24581 26803 24639 26809
rect 25492 26803 25504 26812
rect 25498 26800 25504 26803
rect 25556 26800 25562 26852
rect 29730 26840 29736 26852
rect 29643 26812 29736 26840
rect 29730 26800 29736 26812
rect 29788 26840 29794 26852
rect 30070 26843 30128 26849
rect 30070 26840 30082 26843
rect 29788 26812 30082 26840
rect 29788 26800 29794 26812
rect 30070 26809 30082 26812
rect 30116 26809 30128 26843
rect 30070 26803 30128 26809
rect 31849 26843 31907 26849
rect 31849 26809 31861 26843
rect 31895 26840 31907 26843
rect 32677 26843 32735 26849
rect 32677 26840 32689 26843
rect 31895 26812 32689 26840
rect 31895 26809 31907 26812
rect 31849 26803 31907 26809
rect 32677 26809 32689 26812
rect 32723 26840 32735 26843
rect 33042 26840 33048 26852
rect 32723 26812 33048 26840
rect 32723 26809 32735 26812
rect 32677 26803 32735 26809
rect 33042 26800 33048 26812
rect 33100 26800 33106 26852
rect 34974 26800 34980 26852
rect 35032 26840 35038 26852
rect 35253 26843 35311 26849
rect 35253 26840 35265 26843
rect 35032 26812 35265 26840
rect 35032 26800 35038 26812
rect 35253 26809 35265 26812
rect 35299 26840 35311 26843
rect 35299 26812 36492 26840
rect 35299 26809 35311 26812
rect 35253 26803 35311 26809
rect 8846 26772 8852 26784
rect 8807 26744 8852 26772
rect 8846 26732 8852 26744
rect 8904 26732 8910 26784
rect 11054 26772 11060 26784
rect 11015 26744 11060 26772
rect 11054 26732 11060 26744
rect 11112 26732 11118 26784
rect 14826 26772 14832 26784
rect 14787 26744 14832 26772
rect 14826 26732 14832 26744
rect 14884 26732 14890 26784
rect 17954 26732 17960 26784
rect 18012 26772 18018 26784
rect 18233 26775 18291 26781
rect 18233 26772 18245 26775
rect 18012 26744 18245 26772
rect 18012 26732 18018 26744
rect 18233 26741 18245 26744
rect 18279 26741 18291 26775
rect 19334 26772 19340 26784
rect 19295 26744 19340 26772
rect 18233 26735 18291 26741
rect 19334 26732 19340 26744
rect 19392 26732 19398 26784
rect 20162 26772 20168 26784
rect 20123 26744 20168 26772
rect 20162 26732 20168 26744
rect 20220 26732 20226 26784
rect 20717 26775 20775 26781
rect 20717 26741 20729 26775
rect 20763 26772 20775 26775
rect 21266 26772 21272 26784
rect 20763 26744 21272 26772
rect 20763 26741 20775 26744
rect 20717 26735 20775 26741
rect 21266 26732 21272 26744
rect 21324 26772 21330 26784
rect 21545 26775 21603 26781
rect 21545 26772 21557 26775
rect 21324 26744 21557 26772
rect 21324 26732 21330 26744
rect 21545 26741 21557 26744
rect 21591 26741 21603 26775
rect 22278 26772 22284 26784
rect 22191 26744 22284 26772
rect 21545 26735 21603 26741
rect 22278 26732 22284 26744
rect 22336 26772 22342 26784
rect 22557 26775 22615 26781
rect 22557 26772 22569 26775
rect 22336 26744 22569 26772
rect 22336 26732 22342 26744
rect 22557 26741 22569 26744
rect 22603 26741 22615 26775
rect 22557 26735 22615 26741
rect 25314 26732 25320 26784
rect 25372 26772 25378 26784
rect 26605 26775 26663 26781
rect 26605 26772 26617 26775
rect 25372 26744 26617 26772
rect 25372 26732 25378 26744
rect 26605 26741 26617 26744
rect 26651 26741 26663 26775
rect 27246 26772 27252 26784
rect 27207 26744 27252 26772
rect 26605 26735 26663 26741
rect 27246 26732 27252 26744
rect 27304 26732 27310 26784
rect 30742 26732 30748 26784
rect 30800 26772 30806 26784
rect 31205 26775 31263 26781
rect 31205 26772 31217 26775
rect 30800 26744 31217 26772
rect 30800 26732 30806 26744
rect 31205 26741 31217 26744
rect 31251 26772 31263 26775
rect 31662 26772 31668 26784
rect 31251 26744 31668 26772
rect 31251 26741 31263 26744
rect 31205 26735 31263 26741
rect 31662 26732 31668 26744
rect 31720 26732 31726 26784
rect 34422 26732 34428 26784
rect 34480 26772 34486 26784
rect 36464 26781 36492 26812
rect 34885 26775 34943 26781
rect 34885 26772 34897 26775
rect 34480 26744 34897 26772
rect 34480 26732 34486 26744
rect 34885 26741 34897 26744
rect 34931 26741 34943 26775
rect 34885 26735 34943 26741
rect 36449 26775 36507 26781
rect 36449 26741 36461 26775
rect 36495 26741 36507 26775
rect 36814 26772 36820 26784
rect 36775 26744 36820 26772
rect 36449 26735 36507 26741
rect 36814 26732 36820 26744
rect 36872 26772 36878 26784
rect 37461 26775 37519 26781
rect 37461 26772 37473 26775
rect 36872 26744 37473 26772
rect 36872 26732 36878 26744
rect 37461 26741 37473 26744
rect 37507 26741 37519 26775
rect 37826 26772 37832 26784
rect 37787 26744 37832 26772
rect 37461 26735 37519 26741
rect 37826 26732 37832 26744
rect 37884 26732 37890 26784
rect 1104 26682 38824 26704
rect 1104 26630 19606 26682
rect 19658 26630 19670 26682
rect 19722 26630 19734 26682
rect 19786 26630 19798 26682
rect 19850 26630 38824 26682
rect 1104 26608 38824 26630
rect 2130 26528 2136 26580
rect 2188 26568 2194 26580
rect 2869 26571 2927 26577
rect 2869 26568 2881 26571
rect 2188 26540 2881 26568
rect 2188 26528 2194 26540
rect 2869 26537 2881 26540
rect 2915 26537 2927 26571
rect 2869 26531 2927 26537
rect 4341 26571 4399 26577
rect 4341 26537 4353 26571
rect 4387 26568 4399 26571
rect 4614 26568 4620 26580
rect 4387 26540 4620 26568
rect 4387 26537 4399 26540
rect 4341 26531 4399 26537
rect 4614 26528 4620 26540
rect 4672 26528 4678 26580
rect 6454 26568 6460 26580
rect 6415 26540 6460 26568
rect 6454 26528 6460 26540
rect 6512 26528 6518 26580
rect 6638 26528 6644 26580
rect 6696 26568 6702 26580
rect 6914 26568 6920 26580
rect 6696 26540 6920 26568
rect 6696 26528 6702 26540
rect 6914 26528 6920 26540
rect 6972 26568 6978 26580
rect 7469 26571 7527 26577
rect 7469 26568 7481 26571
rect 6972 26540 7481 26568
rect 6972 26528 6978 26540
rect 7469 26537 7481 26540
rect 7515 26537 7527 26571
rect 7469 26531 7527 26537
rect 11054 26528 11060 26580
rect 11112 26568 11118 26580
rect 11241 26571 11299 26577
rect 11241 26568 11253 26571
rect 11112 26540 11253 26568
rect 11112 26528 11118 26540
rect 11241 26537 11253 26540
rect 11287 26537 11299 26571
rect 11241 26531 11299 26537
rect 11330 26528 11336 26580
rect 11388 26568 11394 26580
rect 11701 26571 11759 26577
rect 11701 26568 11713 26571
rect 11388 26540 11713 26568
rect 11388 26528 11394 26540
rect 11701 26537 11713 26540
rect 11747 26568 11759 26571
rect 12805 26571 12863 26577
rect 12805 26568 12817 26571
rect 11747 26540 12817 26568
rect 11747 26537 11759 26540
rect 11701 26531 11759 26537
rect 12805 26537 12817 26540
rect 12851 26537 12863 26571
rect 12805 26531 12863 26537
rect 13265 26571 13323 26577
rect 13265 26537 13277 26571
rect 13311 26568 13323 26571
rect 13538 26568 13544 26580
rect 13311 26540 13544 26568
rect 13311 26537 13323 26540
rect 13265 26531 13323 26537
rect 13538 26528 13544 26540
rect 13596 26568 13602 26580
rect 14826 26568 14832 26580
rect 13596 26540 14832 26568
rect 13596 26528 13602 26540
rect 14826 26528 14832 26540
rect 14884 26528 14890 26580
rect 19150 26528 19156 26580
rect 19208 26568 19214 26580
rect 19245 26571 19303 26577
rect 19245 26568 19257 26571
rect 19208 26540 19257 26568
rect 19208 26528 19214 26540
rect 19245 26537 19257 26540
rect 19291 26537 19303 26571
rect 19245 26531 19303 26537
rect 19334 26528 19340 26580
rect 19392 26568 19398 26580
rect 19705 26571 19763 26577
rect 19705 26568 19717 26571
rect 19392 26540 19717 26568
rect 19392 26528 19398 26540
rect 19705 26537 19717 26540
rect 19751 26537 19763 26571
rect 22278 26568 22284 26580
rect 22239 26540 22284 26568
rect 19705 26531 19763 26537
rect 22278 26528 22284 26540
rect 22336 26528 22342 26580
rect 25498 26528 25504 26580
rect 25556 26568 25562 26580
rect 25685 26571 25743 26577
rect 25685 26568 25697 26571
rect 25556 26540 25697 26568
rect 25556 26528 25562 26540
rect 25685 26537 25697 26540
rect 25731 26537 25743 26571
rect 29362 26568 29368 26580
rect 29323 26540 29368 26568
rect 25685 26531 25743 26537
rect 29362 26528 29368 26540
rect 29420 26528 29426 26580
rect 29546 26528 29552 26580
rect 29604 26568 29610 26580
rect 29733 26571 29791 26577
rect 29733 26568 29745 26571
rect 29604 26540 29745 26568
rect 29604 26528 29610 26540
rect 29733 26537 29745 26540
rect 29779 26537 29791 26571
rect 30742 26568 30748 26580
rect 30703 26540 30748 26568
rect 29733 26531 29791 26537
rect 30742 26528 30748 26540
rect 30800 26528 30806 26580
rect 30834 26528 30840 26580
rect 30892 26568 30898 26580
rect 32674 26568 32680 26580
rect 30892 26540 32680 26568
rect 30892 26528 30898 26540
rect 32674 26528 32680 26540
rect 32732 26568 32738 26580
rect 32950 26568 32956 26580
rect 32732 26540 32956 26568
rect 32732 26528 32738 26540
rect 32950 26528 32956 26540
rect 33008 26568 33014 26580
rect 33229 26571 33287 26577
rect 33229 26568 33241 26571
rect 33008 26540 33241 26568
rect 33008 26528 33014 26540
rect 33229 26537 33241 26540
rect 33275 26568 33287 26571
rect 34238 26568 34244 26580
rect 33275 26540 34244 26568
rect 33275 26537 33287 26540
rect 33229 26531 33287 26537
rect 34238 26528 34244 26540
rect 34296 26528 34302 26580
rect 34974 26568 34980 26580
rect 34935 26540 34980 26568
rect 34974 26528 34980 26540
rect 35032 26528 35038 26580
rect 36998 26528 37004 26580
rect 37056 26568 37062 26580
rect 37093 26571 37151 26577
rect 37093 26568 37105 26571
rect 37056 26540 37105 26568
rect 37056 26528 37062 26540
rect 37093 26537 37105 26540
rect 37139 26537 37151 26571
rect 37093 26531 37151 26537
rect 1762 26509 1768 26512
rect 1756 26500 1768 26509
rect 1723 26472 1768 26500
rect 1756 26463 1768 26472
rect 1762 26460 1768 26463
rect 1820 26460 1826 26512
rect 15832 26503 15890 26509
rect 15832 26469 15844 26503
rect 15878 26500 15890 26503
rect 16114 26500 16120 26512
rect 15878 26472 16120 26500
rect 15878 26469 15890 26472
rect 15832 26463 15890 26469
rect 16114 26460 16120 26472
rect 16172 26500 16178 26512
rect 16942 26500 16948 26512
rect 16172 26472 16948 26500
rect 16172 26460 16178 26472
rect 16942 26460 16948 26472
rect 17000 26460 17006 26512
rect 19426 26460 19432 26512
rect 19484 26500 19490 26512
rect 19613 26503 19671 26509
rect 19613 26500 19625 26503
rect 19484 26472 19625 26500
rect 19484 26460 19490 26472
rect 19613 26469 19625 26472
rect 19659 26500 19671 26503
rect 20162 26500 20168 26512
rect 19659 26472 20168 26500
rect 19659 26469 19671 26472
rect 19613 26463 19671 26469
rect 20162 26460 20168 26472
rect 20220 26460 20226 26512
rect 24121 26503 24179 26509
rect 24121 26469 24133 26503
rect 24167 26500 24179 26503
rect 25314 26500 25320 26512
rect 24167 26472 25320 26500
rect 24167 26469 24179 26472
rect 24121 26463 24179 26469
rect 25314 26460 25320 26472
rect 25372 26460 25378 26512
rect 31938 26500 31944 26512
rect 31851 26472 31944 26500
rect 31938 26460 31944 26472
rect 31996 26500 32002 26512
rect 32585 26503 32643 26509
rect 32585 26500 32597 26503
rect 31996 26472 32597 26500
rect 31996 26460 32002 26472
rect 32585 26469 32597 26472
rect 32631 26469 32643 26503
rect 35526 26500 35532 26512
rect 32585 26463 32643 26469
rect 35176 26472 35532 26500
rect 1486 26432 1492 26444
rect 1447 26404 1492 26432
rect 1486 26392 1492 26404
rect 1544 26392 1550 26444
rect 6730 26392 6736 26444
rect 6788 26432 6794 26444
rect 6825 26435 6883 26441
rect 6825 26432 6837 26435
rect 6788 26404 6837 26432
rect 6788 26392 6794 26404
rect 6825 26401 6837 26404
rect 6871 26401 6883 26435
rect 6825 26395 6883 26401
rect 8389 26435 8447 26441
rect 8389 26401 8401 26435
rect 8435 26432 8447 26435
rect 9030 26432 9036 26444
rect 8435 26404 9036 26432
rect 8435 26401 8447 26404
rect 8389 26395 8447 26401
rect 9030 26392 9036 26404
rect 9088 26392 9094 26444
rect 11606 26432 11612 26444
rect 11567 26404 11612 26432
rect 11606 26392 11612 26404
rect 11664 26392 11670 26444
rect 13170 26432 13176 26444
rect 13131 26404 13176 26432
rect 13170 26392 13176 26404
rect 13228 26392 13234 26444
rect 15562 26432 15568 26444
rect 15523 26404 15568 26432
rect 15562 26392 15568 26404
rect 15620 26392 15626 26444
rect 18049 26435 18107 26441
rect 18049 26401 18061 26435
rect 18095 26432 18107 26435
rect 18322 26432 18328 26444
rect 18095 26404 18328 26432
rect 18095 26401 18107 26404
rect 18049 26395 18107 26401
rect 18322 26392 18328 26404
rect 18380 26432 18386 26444
rect 19242 26432 19248 26444
rect 18380 26404 19248 26432
rect 18380 26392 18386 26404
rect 19242 26392 19248 26404
rect 19300 26392 19306 26444
rect 20070 26432 20076 26444
rect 19904 26404 20076 26432
rect 6917 26367 6975 26373
rect 6917 26364 6929 26367
rect 6840 26336 6929 26364
rect 6840 26308 6868 26336
rect 6917 26333 6929 26336
rect 6963 26333 6975 26367
rect 6917 26327 6975 26333
rect 7101 26367 7159 26373
rect 7101 26333 7113 26367
rect 7147 26364 7159 26367
rect 8110 26364 8116 26376
rect 7147 26336 8116 26364
rect 7147 26333 7159 26336
rect 7101 26327 7159 26333
rect 6822 26256 6828 26308
rect 6880 26256 6886 26308
rect 7116 26296 7144 26327
rect 8110 26324 8116 26336
rect 8168 26324 8174 26376
rect 8478 26364 8484 26376
rect 8439 26336 8484 26364
rect 8478 26324 8484 26336
rect 8536 26324 8542 26376
rect 8570 26324 8576 26376
rect 8628 26364 8634 26376
rect 8628 26336 8673 26364
rect 8628 26324 8634 26336
rect 11422 26324 11428 26376
rect 11480 26364 11486 26376
rect 19904 26373 19932 26404
rect 20070 26392 20076 26404
rect 20128 26432 20134 26444
rect 20717 26435 20775 26441
rect 20717 26432 20729 26435
rect 20128 26404 20729 26432
rect 20128 26392 20134 26404
rect 20717 26401 20729 26404
rect 20763 26432 20775 26435
rect 21168 26435 21226 26441
rect 21168 26432 21180 26435
rect 20763 26404 21180 26432
rect 20763 26401 20775 26404
rect 20717 26395 20775 26401
rect 21168 26401 21180 26404
rect 21214 26432 21226 26435
rect 22002 26432 22008 26444
rect 21214 26404 22008 26432
rect 21214 26401 21226 26404
rect 21168 26395 21226 26401
rect 22002 26392 22008 26404
rect 22060 26392 22066 26444
rect 24946 26392 24952 26444
rect 25004 26432 25010 26444
rect 25041 26435 25099 26441
rect 25041 26432 25053 26435
rect 25004 26404 25053 26432
rect 25004 26392 25010 26404
rect 25041 26401 25053 26404
rect 25087 26401 25099 26435
rect 25041 26395 25099 26401
rect 26418 26392 26424 26444
rect 26476 26432 26482 26444
rect 27249 26435 27307 26441
rect 27249 26432 27261 26435
rect 26476 26404 27261 26432
rect 26476 26392 26482 26404
rect 27249 26401 27261 26404
rect 27295 26401 27307 26435
rect 27249 26395 27307 26401
rect 28902 26392 28908 26444
rect 28960 26432 28966 26444
rect 29178 26432 29184 26444
rect 28960 26404 29184 26432
rect 28960 26392 28966 26404
rect 29178 26392 29184 26404
rect 29236 26392 29242 26444
rect 30653 26435 30711 26441
rect 30653 26401 30665 26435
rect 30699 26432 30711 26435
rect 30926 26432 30932 26444
rect 30699 26404 30932 26432
rect 30699 26401 30711 26404
rect 30653 26395 30711 26401
rect 30926 26392 30932 26404
rect 30984 26432 30990 26444
rect 31478 26432 31484 26444
rect 30984 26404 31484 26432
rect 30984 26392 30990 26404
rect 31478 26392 31484 26404
rect 31536 26392 31542 26444
rect 32493 26435 32551 26441
rect 32493 26401 32505 26435
rect 32539 26401 32551 26435
rect 34054 26432 34060 26444
rect 34015 26404 34060 26432
rect 32493 26395 32551 26401
rect 11793 26367 11851 26373
rect 11793 26364 11805 26367
rect 11480 26336 11805 26364
rect 11480 26324 11486 26336
rect 11793 26333 11805 26336
rect 11839 26333 11851 26367
rect 11793 26327 11851 26333
rect 13357 26367 13415 26373
rect 13357 26333 13369 26367
rect 13403 26333 13415 26367
rect 13357 26327 13415 26333
rect 19889 26367 19947 26373
rect 19889 26333 19901 26367
rect 19935 26333 19947 26367
rect 20898 26364 20904 26376
rect 20859 26336 20904 26364
rect 19889 26327 19947 26333
rect 6932 26268 7144 26296
rect 8021 26299 8079 26305
rect 5810 26188 5816 26240
rect 5868 26228 5874 26240
rect 6932 26228 6960 26268
rect 8021 26265 8033 26299
rect 8067 26296 8079 26299
rect 9309 26299 9367 26305
rect 9309 26296 9321 26299
rect 8067 26268 9321 26296
rect 8067 26265 8079 26268
rect 8021 26259 8079 26265
rect 9309 26265 9321 26268
rect 9355 26296 9367 26299
rect 9674 26296 9680 26308
rect 9355 26268 9680 26296
rect 9355 26265 9367 26268
rect 9309 26259 9367 26265
rect 9674 26256 9680 26268
rect 9732 26256 9738 26308
rect 12713 26299 12771 26305
rect 12713 26296 12725 26299
rect 12268 26268 12725 26296
rect 5868 26200 6960 26228
rect 5868 26188 5874 26200
rect 8570 26188 8576 26240
rect 8628 26228 8634 26240
rect 10594 26228 10600 26240
rect 8628 26200 10600 26228
rect 8628 26188 8634 26200
rect 10594 26188 10600 26200
rect 10652 26228 10658 26240
rect 12268 26228 12296 26268
rect 12713 26265 12725 26268
rect 12759 26296 12771 26299
rect 13372 26296 13400 26327
rect 20898 26324 20904 26336
rect 20956 26324 20962 26376
rect 24118 26324 24124 26376
rect 24176 26364 24182 26376
rect 24578 26364 24584 26376
rect 24176 26336 24584 26364
rect 24176 26324 24182 26336
rect 24578 26324 24584 26336
rect 24636 26364 24642 26376
rect 25133 26367 25191 26373
rect 25133 26364 25145 26367
rect 24636 26336 25145 26364
rect 24636 26324 24642 26336
rect 25133 26333 25145 26336
rect 25179 26333 25191 26367
rect 25314 26364 25320 26376
rect 25275 26336 25320 26364
rect 25133 26327 25191 26333
rect 25314 26324 25320 26336
rect 25372 26324 25378 26376
rect 26513 26367 26571 26373
rect 26513 26333 26525 26367
rect 26559 26333 26571 26367
rect 26513 26327 26571 26333
rect 16945 26299 17003 26305
rect 16945 26296 16957 26299
rect 12759 26268 13400 26296
rect 16500 26268 16957 26296
rect 12759 26265 12771 26268
rect 12713 26259 12771 26265
rect 16500 26240 16528 26268
rect 16945 26265 16957 26268
rect 16991 26265 17003 26299
rect 16945 26259 17003 26265
rect 19153 26299 19211 26305
rect 19153 26265 19165 26299
rect 19199 26296 19211 26299
rect 20346 26296 20352 26308
rect 19199 26268 19288 26296
rect 20259 26268 20352 26296
rect 19199 26265 19211 26268
rect 19153 26259 19211 26265
rect 10652 26200 12296 26228
rect 12345 26231 12403 26237
rect 10652 26188 10658 26200
rect 12345 26197 12357 26231
rect 12391 26228 12403 26231
rect 12434 26228 12440 26240
rect 12391 26200 12440 26228
rect 12391 26197 12403 26200
rect 12345 26191 12403 26197
rect 12434 26188 12440 26200
rect 12492 26188 12498 26240
rect 16482 26188 16488 26240
rect 16540 26188 16546 26240
rect 17954 26188 17960 26240
rect 18012 26228 18018 26240
rect 18233 26231 18291 26237
rect 18233 26228 18245 26231
rect 18012 26200 18245 26228
rect 18012 26188 18018 26200
rect 18233 26197 18245 26200
rect 18279 26197 18291 26231
rect 19260 26228 19288 26268
rect 20346 26256 20352 26268
rect 20404 26296 20410 26308
rect 20530 26296 20536 26308
rect 20404 26268 20536 26296
rect 20404 26256 20410 26268
rect 20530 26256 20536 26268
rect 20588 26256 20594 26308
rect 19794 26228 19800 26240
rect 19260 26200 19800 26228
rect 18233 26191 18291 26197
rect 19794 26188 19800 26200
rect 19852 26188 19858 26240
rect 20916 26228 20944 26324
rect 24673 26299 24731 26305
rect 24673 26265 24685 26299
rect 24719 26296 24731 26299
rect 26234 26296 26240 26308
rect 24719 26268 24900 26296
rect 26195 26268 26240 26296
rect 24719 26265 24731 26268
rect 24673 26259 24731 26265
rect 22922 26228 22928 26240
rect 20916 26200 22928 26228
rect 22922 26188 22928 26200
rect 22980 26188 22986 26240
rect 24489 26231 24547 26237
rect 24489 26197 24501 26231
rect 24535 26228 24547 26231
rect 24578 26228 24584 26240
rect 24535 26200 24584 26228
rect 24535 26197 24547 26200
rect 24489 26191 24547 26197
rect 24578 26188 24584 26200
rect 24636 26188 24642 26240
rect 24872 26228 24900 26268
rect 26234 26256 26240 26268
rect 26292 26296 26298 26308
rect 26528 26296 26556 26327
rect 26694 26324 26700 26376
rect 26752 26364 26758 26376
rect 26836 26367 26894 26373
rect 26836 26364 26848 26367
rect 26752 26336 26848 26364
rect 26752 26324 26758 26336
rect 26836 26333 26848 26336
rect 26882 26333 26894 26367
rect 26836 26327 26894 26333
rect 26970 26324 26976 26376
rect 27028 26364 27034 26376
rect 30193 26367 30251 26373
rect 27028 26336 27073 26364
rect 27028 26324 27034 26336
rect 30193 26333 30205 26367
rect 30239 26364 30251 26367
rect 30834 26364 30840 26376
rect 30239 26336 30840 26364
rect 30239 26333 30251 26336
rect 30193 26327 30251 26333
rect 30834 26324 30840 26336
rect 30892 26324 30898 26376
rect 31662 26364 31668 26376
rect 31575 26336 31668 26364
rect 26292 26268 26556 26296
rect 26292 26256 26298 26268
rect 28258 26256 28264 26308
rect 28316 26296 28322 26308
rect 28353 26299 28411 26305
rect 28353 26296 28365 26299
rect 28316 26268 28365 26296
rect 28316 26256 28322 26268
rect 28353 26265 28365 26268
rect 28399 26265 28411 26299
rect 31588 26296 31616 26336
rect 31662 26324 31668 26336
rect 31720 26364 31726 26376
rect 32508 26364 32536 26395
rect 34054 26392 34060 26404
rect 34112 26392 34118 26444
rect 34606 26392 34612 26444
rect 34664 26432 34670 26444
rect 35176 26441 35204 26472
rect 35526 26460 35532 26472
rect 35584 26460 35590 26512
rect 35161 26435 35219 26441
rect 35161 26432 35173 26435
rect 34664 26404 35173 26432
rect 34664 26392 34670 26404
rect 35161 26401 35173 26404
rect 35207 26401 35219 26435
rect 35161 26395 35219 26401
rect 35250 26392 35256 26444
rect 35308 26432 35314 26444
rect 35417 26435 35475 26441
rect 35417 26432 35429 26435
rect 35308 26404 35429 26432
rect 35308 26392 35314 26404
rect 35417 26401 35429 26404
rect 35463 26432 35475 26435
rect 36814 26432 36820 26444
rect 35463 26404 36820 26432
rect 35463 26401 35475 26404
rect 35417 26395 35475 26401
rect 36814 26392 36820 26404
rect 36872 26392 36878 26444
rect 32677 26367 32735 26373
rect 32677 26364 32689 26367
rect 31720 26336 32536 26364
rect 32600 26336 32689 26364
rect 31720 26324 31726 26336
rect 28353 26259 28411 26265
rect 31496 26268 31616 26296
rect 32125 26299 32183 26305
rect 25038 26228 25044 26240
rect 24872 26200 25044 26228
rect 25038 26188 25044 26200
rect 25096 26188 25102 26240
rect 30285 26231 30343 26237
rect 30285 26197 30297 26231
rect 30331 26228 30343 26231
rect 31496 26228 31524 26268
rect 32125 26265 32137 26299
rect 32171 26296 32183 26299
rect 32306 26296 32312 26308
rect 32171 26268 32312 26296
rect 32171 26265 32183 26268
rect 32125 26259 32183 26265
rect 32306 26256 32312 26268
rect 32364 26256 32370 26308
rect 30331 26200 31524 26228
rect 30331 26197 30343 26200
rect 30285 26191 30343 26197
rect 31570 26188 31576 26240
rect 31628 26228 31634 26240
rect 32600 26228 32628 26336
rect 32677 26333 32689 26336
rect 32723 26333 32735 26367
rect 32677 26327 32735 26333
rect 33042 26324 33048 26376
rect 33100 26364 33106 26376
rect 33505 26367 33563 26373
rect 33505 26364 33517 26367
rect 33100 26336 33517 26364
rect 33100 26324 33106 26336
rect 33505 26333 33517 26336
rect 33551 26333 33563 26367
rect 33505 26327 33563 26333
rect 36541 26299 36599 26305
rect 36541 26296 36553 26299
rect 36096 26268 36553 26296
rect 34241 26231 34299 26237
rect 34241 26228 34253 26231
rect 31628 26200 34253 26228
rect 31628 26188 31634 26200
rect 34241 26197 34253 26200
rect 34287 26197 34299 26231
rect 34241 26191 34299 26197
rect 35526 26188 35532 26240
rect 35584 26228 35590 26240
rect 36096 26228 36124 26268
rect 36541 26265 36553 26268
rect 36587 26265 36599 26299
rect 36541 26259 36599 26265
rect 35584 26200 36124 26228
rect 35584 26188 35590 26200
rect 1104 26138 38824 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 34966 26138
rect 35018 26086 35030 26138
rect 35082 26086 35094 26138
rect 35146 26086 35158 26138
rect 35210 26086 38824 26138
rect 1104 26064 38824 26086
rect 2222 26024 2228 26036
rect 2183 25996 2228 26024
rect 2222 25984 2228 25996
rect 2280 25984 2286 26036
rect 5810 26024 5816 26036
rect 5771 25996 5816 26024
rect 5810 25984 5816 25996
rect 5868 25984 5874 26036
rect 8202 26024 8208 26036
rect 8163 25996 8208 26024
rect 8202 25984 8208 25996
rect 8260 25984 8266 26036
rect 8478 25984 8484 26036
rect 8536 26024 8542 26036
rect 8757 26027 8815 26033
rect 8757 26024 8769 26027
rect 8536 25996 8769 26024
rect 8536 25984 8542 25996
rect 8757 25993 8769 25996
rect 8803 25993 8815 26027
rect 8757 25987 8815 25993
rect 9309 26027 9367 26033
rect 9309 25993 9321 26027
rect 9355 26024 9367 26027
rect 9582 26024 9588 26036
rect 9355 25996 9588 26024
rect 9355 25993 9367 25996
rect 9309 25987 9367 25993
rect 9582 25984 9588 25996
rect 9640 25984 9646 26036
rect 11330 26024 11336 26036
rect 11291 25996 11336 26024
rect 11330 25984 11336 25996
rect 11388 25984 11394 26036
rect 16761 26027 16819 26033
rect 16761 25993 16773 26027
rect 16807 26024 16819 26027
rect 17862 26024 17868 26036
rect 16807 25996 17868 26024
rect 16807 25993 16819 25996
rect 16761 25987 16819 25993
rect 6638 25848 6644 25900
rect 6696 25888 6702 25900
rect 6825 25891 6883 25897
rect 6825 25888 6837 25891
rect 6696 25860 6837 25888
rect 6696 25848 6702 25860
rect 6825 25857 6837 25860
rect 6871 25857 6883 25891
rect 9858 25888 9864 25900
rect 9819 25860 9864 25888
rect 6825 25851 6883 25857
rect 9858 25848 9864 25860
rect 9916 25888 9922 25900
rect 10321 25891 10379 25897
rect 10321 25888 10333 25891
rect 9916 25860 10333 25888
rect 9916 25848 9922 25860
rect 10321 25857 10333 25860
rect 10367 25888 10379 25891
rect 10873 25891 10931 25897
rect 10873 25888 10885 25891
rect 10367 25860 10885 25888
rect 10367 25857 10379 25860
rect 10321 25851 10379 25857
rect 10873 25857 10885 25860
rect 10919 25857 10931 25891
rect 10873 25851 10931 25857
rect 15197 25891 15255 25897
rect 15197 25857 15209 25891
rect 15243 25888 15255 25891
rect 15565 25891 15623 25897
rect 15565 25888 15577 25891
rect 15243 25860 15577 25888
rect 15243 25857 15255 25860
rect 15197 25851 15255 25857
rect 15565 25857 15577 25860
rect 15611 25888 15623 25891
rect 16114 25888 16120 25900
rect 15611 25860 16120 25888
rect 15611 25857 15623 25860
rect 15565 25851 15623 25857
rect 16114 25848 16120 25860
rect 16172 25848 16178 25900
rect 16298 25888 16304 25900
rect 16211 25860 16304 25888
rect 16298 25848 16304 25860
rect 16356 25888 16362 25900
rect 16776 25888 16804 25987
rect 17862 25984 17868 25996
rect 17920 25984 17926 26036
rect 18322 26024 18328 26036
rect 18283 25996 18328 26024
rect 18322 25984 18328 25996
rect 18380 25984 18386 26036
rect 19150 25984 19156 26036
rect 19208 26024 19214 26036
rect 19245 26027 19303 26033
rect 19245 26024 19257 26027
rect 19208 25996 19257 26024
rect 19208 25984 19214 25996
rect 19245 25993 19257 25996
rect 19291 25993 19303 26027
rect 19245 25987 19303 25993
rect 21910 25984 21916 26036
rect 21968 26024 21974 26036
rect 22649 26027 22707 26033
rect 22649 26024 22661 26027
rect 21968 25996 22661 26024
rect 21968 25984 21974 25996
rect 22649 25993 22661 25996
rect 22695 25993 22707 26027
rect 22922 26024 22928 26036
rect 22883 25996 22928 26024
rect 22649 25987 22707 25993
rect 17126 25956 17132 25968
rect 17087 25928 17132 25956
rect 17126 25916 17132 25928
rect 17184 25916 17190 25968
rect 22664 25956 22692 25987
rect 22922 25984 22928 25996
rect 22980 25984 22986 26036
rect 26326 25984 26332 26036
rect 26384 26024 26390 26036
rect 27065 26027 27123 26033
rect 27065 26024 27077 26027
rect 26384 25996 27077 26024
rect 26384 25984 26390 25996
rect 27065 25993 27077 25996
rect 27111 25993 27123 26027
rect 27065 25987 27123 25993
rect 28813 26027 28871 26033
rect 28813 25993 28825 26027
rect 28859 26024 28871 26027
rect 28902 26024 28908 26036
rect 28859 25996 28908 26024
rect 28859 25993 28871 25996
rect 28813 25987 28871 25993
rect 28902 25984 28908 25996
rect 28960 25984 28966 26036
rect 31754 25984 31760 26036
rect 31812 26024 31818 26036
rect 32217 26027 32275 26033
rect 31812 25996 31857 26024
rect 31812 25984 31818 25996
rect 32217 25993 32229 26027
rect 32263 26024 32275 26027
rect 34054 26024 34060 26036
rect 32263 25996 33963 26024
rect 34015 25996 34060 26024
rect 32263 25993 32275 25996
rect 32217 25987 32275 25993
rect 23845 25959 23903 25965
rect 23845 25956 23857 25959
rect 22664 25928 23857 25956
rect 23845 25925 23857 25928
rect 23891 25956 23903 25959
rect 24302 25956 24308 25968
rect 23891 25928 24308 25956
rect 23891 25925 23903 25928
rect 23845 25919 23903 25925
rect 24302 25916 24308 25928
rect 24360 25916 24366 25968
rect 26237 25959 26295 25965
rect 26237 25925 26249 25959
rect 26283 25956 26295 25959
rect 26418 25956 26424 25968
rect 26283 25928 26424 25956
rect 26283 25925 26295 25928
rect 26237 25919 26295 25925
rect 26418 25916 26424 25928
rect 26476 25956 26482 25968
rect 28077 25959 28135 25965
rect 28077 25956 28089 25959
rect 26476 25928 28089 25956
rect 26476 25916 26482 25928
rect 28077 25925 28089 25928
rect 28123 25925 28135 25959
rect 28077 25919 28135 25925
rect 33045 25959 33103 25965
rect 33045 25925 33057 25959
rect 33091 25956 33103 25959
rect 33318 25956 33324 25968
rect 33091 25928 33324 25956
rect 33091 25925 33103 25928
rect 33045 25919 33103 25925
rect 33318 25916 33324 25928
rect 33376 25916 33382 25968
rect 33935 25956 33963 25996
rect 34054 25984 34060 25996
rect 34112 25984 34118 26036
rect 34606 26024 34612 26036
rect 34567 25996 34612 26024
rect 34606 25984 34612 25996
rect 34664 25984 34670 26036
rect 35710 25984 35716 26036
rect 35768 26024 35774 26036
rect 36081 26027 36139 26033
rect 36081 26024 36093 26027
rect 35768 25996 36093 26024
rect 35768 25984 35774 25996
rect 36081 25993 36093 25996
rect 36127 25993 36139 26027
rect 36081 25987 36139 25993
rect 34624 25956 34652 25984
rect 33935 25928 34652 25956
rect 16356 25860 16804 25888
rect 19153 25891 19211 25897
rect 16356 25848 16362 25860
rect 19153 25857 19165 25891
rect 19199 25888 19211 25891
rect 19242 25888 19248 25900
rect 19199 25860 19248 25888
rect 19199 25857 19211 25860
rect 19153 25851 19211 25857
rect 19242 25848 19248 25860
rect 19300 25848 19306 25900
rect 19794 25888 19800 25900
rect 19755 25860 19800 25888
rect 19794 25848 19800 25860
rect 19852 25848 19858 25900
rect 20530 25848 20536 25900
rect 20588 25888 20594 25900
rect 20809 25891 20867 25897
rect 20809 25888 20821 25891
rect 20588 25860 20821 25888
rect 20588 25848 20594 25860
rect 20809 25857 20821 25860
rect 20855 25888 20867 25891
rect 20990 25888 20996 25900
rect 20855 25860 20996 25888
rect 20855 25857 20867 25860
rect 20809 25851 20867 25857
rect 20990 25848 20996 25860
rect 21048 25848 21054 25900
rect 21266 25848 21272 25900
rect 21324 25888 21330 25900
rect 24320 25888 24348 25916
rect 21324 25860 21369 25888
rect 24320 25860 24532 25888
rect 21324 25848 21330 25860
rect 9674 25820 9680 25832
rect 9635 25792 9680 25820
rect 9674 25780 9680 25792
rect 9732 25780 9738 25832
rect 12434 25780 12440 25832
rect 12492 25820 12498 25832
rect 12704 25823 12762 25829
rect 12704 25820 12716 25823
rect 12492 25792 12537 25820
rect 12636 25792 12716 25820
rect 12492 25780 12498 25792
rect 1673 25755 1731 25761
rect 1673 25721 1685 25755
rect 1719 25752 1731 25755
rect 1762 25752 1768 25764
rect 1719 25724 1768 25752
rect 1719 25721 1731 25724
rect 1673 25715 1731 25721
rect 1762 25712 1768 25724
rect 1820 25752 1826 25764
rect 2682 25752 2688 25764
rect 1820 25724 2688 25752
rect 1820 25712 1826 25724
rect 2682 25712 2688 25724
rect 2740 25712 2746 25764
rect 6181 25755 6239 25761
rect 6181 25721 6193 25755
rect 6227 25752 6239 25755
rect 6730 25752 6736 25764
rect 6227 25724 6736 25752
rect 6227 25721 6239 25724
rect 6181 25715 6239 25721
rect 6730 25712 6736 25724
rect 6788 25752 6794 25764
rect 7098 25761 7104 25764
rect 7092 25752 7104 25761
rect 6788 25724 7104 25752
rect 6788 25712 6794 25724
rect 7092 25715 7104 25724
rect 7098 25712 7104 25715
rect 7156 25712 7162 25764
rect 12253 25755 12311 25761
rect 12253 25721 12265 25755
rect 12299 25752 12311 25755
rect 12636 25752 12664 25792
rect 12704 25789 12716 25792
rect 12750 25820 12762 25823
rect 13538 25820 13544 25832
rect 12750 25792 13544 25820
rect 12750 25789 12762 25792
rect 12704 25783 12762 25789
rect 13538 25780 13544 25792
rect 13596 25780 13602 25832
rect 14829 25823 14887 25829
rect 14829 25789 14841 25823
rect 14875 25820 14887 25823
rect 15102 25820 15108 25832
rect 14875 25792 15108 25820
rect 14875 25789 14887 25792
rect 14829 25783 14887 25789
rect 15102 25780 15108 25792
rect 15160 25820 15166 25832
rect 16022 25820 16028 25832
rect 15160 25792 16028 25820
rect 15160 25780 15166 25792
rect 16022 25780 16028 25792
rect 16080 25820 16086 25832
rect 16482 25820 16488 25832
rect 16080 25792 16488 25820
rect 16080 25780 16086 25792
rect 16482 25780 16488 25792
rect 16540 25780 16546 25832
rect 18785 25823 18843 25829
rect 18785 25789 18797 25823
rect 18831 25820 18843 25823
rect 19613 25823 19671 25829
rect 19613 25820 19625 25823
rect 18831 25792 19625 25820
rect 18831 25789 18843 25792
rect 18785 25783 18843 25789
rect 19613 25789 19625 25792
rect 19659 25820 19671 25823
rect 19978 25820 19984 25832
rect 19659 25792 19984 25820
rect 19659 25789 19671 25792
rect 19613 25783 19671 25789
rect 19978 25780 19984 25792
rect 20036 25820 20042 25832
rect 20622 25820 20628 25832
rect 20036 25792 20628 25820
rect 20036 25780 20042 25792
rect 20622 25780 20628 25792
rect 20680 25780 20686 25832
rect 20898 25780 20904 25832
rect 20956 25820 20962 25832
rect 21545 25823 21603 25829
rect 21545 25820 21557 25823
rect 20956 25792 21557 25820
rect 20956 25780 20962 25792
rect 21545 25789 21557 25792
rect 21591 25789 21603 25823
rect 23474 25820 23480 25832
rect 23435 25792 23480 25820
rect 21545 25783 21603 25789
rect 23474 25780 23480 25792
rect 23532 25820 23538 25832
rect 24394 25820 24400 25832
rect 23532 25792 24400 25820
rect 23532 25780 23538 25792
rect 24394 25780 24400 25792
rect 24452 25780 24458 25832
rect 24504 25820 24532 25860
rect 24578 25848 24584 25900
rect 24636 25888 24642 25900
rect 24860 25891 24918 25897
rect 24860 25888 24872 25891
rect 24636 25860 24872 25888
rect 24636 25848 24642 25860
rect 24860 25857 24872 25860
rect 24906 25857 24918 25891
rect 24860 25851 24918 25857
rect 27246 25848 27252 25900
rect 27304 25888 27310 25900
rect 27706 25888 27712 25900
rect 27304 25860 27712 25888
rect 27304 25848 27310 25860
rect 27706 25848 27712 25860
rect 27764 25848 27770 25900
rect 31478 25848 31484 25900
rect 31536 25888 31542 25900
rect 32033 25891 32091 25897
rect 32033 25888 32045 25891
rect 31536 25860 32045 25888
rect 31536 25848 31542 25860
rect 32033 25857 32045 25860
rect 32079 25857 32091 25891
rect 33686 25888 33692 25900
rect 33647 25860 33692 25888
rect 32033 25851 32091 25857
rect 33686 25848 33692 25860
rect 33744 25848 33750 25900
rect 24946 25820 24952 25832
rect 24504 25792 24952 25820
rect 24946 25780 24952 25792
rect 25004 25820 25010 25832
rect 25133 25823 25191 25829
rect 25133 25820 25145 25823
rect 25004 25792 25145 25820
rect 25004 25780 25010 25792
rect 25133 25789 25145 25792
rect 25179 25789 25191 25823
rect 25133 25783 25191 25789
rect 27062 25780 27068 25832
rect 27120 25820 27126 25832
rect 27433 25823 27491 25829
rect 27433 25820 27445 25823
rect 27120 25792 27445 25820
rect 27120 25780 27126 25792
rect 27433 25789 27445 25792
rect 27479 25789 27491 25823
rect 27433 25783 27491 25789
rect 29089 25823 29147 25829
rect 29089 25789 29101 25823
rect 29135 25820 29147 25823
rect 29178 25820 29184 25832
rect 29135 25792 29184 25820
rect 29135 25789 29147 25792
rect 29089 25783 29147 25789
rect 29178 25780 29184 25792
rect 29236 25780 29242 25832
rect 29733 25823 29791 25829
rect 29733 25789 29745 25823
rect 29779 25820 29791 25823
rect 29822 25820 29828 25832
rect 29779 25792 29828 25820
rect 29779 25789 29791 25792
rect 29733 25783 29791 25789
rect 29822 25780 29828 25792
rect 29880 25780 29886 25832
rect 31754 25780 31760 25832
rect 31812 25820 31818 25832
rect 32401 25823 32459 25829
rect 32401 25820 32413 25823
rect 31812 25792 32413 25820
rect 31812 25780 31818 25792
rect 32401 25789 32413 25792
rect 32447 25820 32459 25823
rect 33042 25820 33048 25832
rect 32447 25792 33048 25820
rect 32447 25789 32459 25792
rect 32401 25783 32459 25789
rect 33042 25780 33048 25792
rect 33100 25780 33106 25832
rect 35345 25823 35403 25829
rect 35345 25789 35357 25823
rect 35391 25820 35403 25823
rect 35526 25820 35532 25832
rect 35391 25792 35532 25820
rect 35391 25789 35403 25792
rect 35345 25783 35403 25789
rect 35526 25780 35532 25792
rect 35584 25820 35590 25832
rect 35621 25823 35679 25829
rect 35621 25820 35633 25823
rect 35584 25792 35633 25820
rect 35584 25780 35590 25792
rect 35621 25789 35633 25792
rect 35667 25789 35679 25823
rect 35621 25783 35679 25789
rect 35805 25823 35863 25829
rect 35805 25789 35817 25823
rect 35851 25820 35863 25823
rect 36633 25823 36691 25829
rect 36633 25820 36645 25823
rect 35851 25792 36645 25820
rect 35851 25789 35863 25792
rect 35805 25783 35863 25789
rect 36633 25789 36645 25792
rect 36679 25820 36691 25823
rect 37185 25823 37243 25829
rect 37185 25820 37197 25823
rect 36679 25792 37197 25820
rect 36679 25789 36691 25792
rect 36633 25783 36691 25789
rect 37185 25789 37197 25792
rect 37231 25789 37243 25823
rect 37185 25783 37243 25789
rect 12299 25724 12664 25752
rect 12299 25721 12311 25724
rect 12253 25715 12311 25721
rect 19334 25712 19340 25764
rect 19392 25752 19398 25764
rect 19705 25755 19763 25761
rect 19705 25752 19717 25755
rect 19392 25724 19717 25752
rect 19392 25712 19398 25724
rect 19705 25721 19717 25724
rect 19751 25752 19763 25755
rect 20916 25752 20944 25780
rect 19751 25724 20944 25752
rect 26973 25755 27031 25761
rect 19751 25721 19763 25724
rect 19705 25715 19763 25721
rect 26973 25721 26985 25755
rect 27019 25752 27031 25755
rect 27525 25755 27583 25761
rect 27525 25752 27537 25755
rect 27019 25724 27537 25752
rect 27019 25721 27031 25724
rect 26973 25715 27031 25721
rect 27525 25721 27537 25724
rect 27571 25752 27583 25755
rect 28258 25752 28264 25764
rect 27571 25724 28264 25752
rect 27571 25721 27583 25724
rect 27525 25715 27583 25721
rect 28258 25712 28264 25724
rect 28316 25712 28322 25764
rect 30006 25761 30012 25764
rect 29641 25755 29699 25761
rect 29641 25721 29653 25755
rect 29687 25752 29699 25755
rect 30000 25752 30012 25761
rect 29687 25724 30012 25752
rect 29687 25721 29699 25724
rect 29641 25715 29699 25721
rect 30000 25715 30012 25724
rect 30006 25712 30012 25715
rect 30064 25712 30070 25764
rect 33505 25755 33563 25761
rect 33505 25752 33517 25755
rect 32876 25724 33517 25752
rect 32876 25696 32904 25724
rect 33505 25721 33517 25724
rect 33551 25721 33563 25755
rect 33505 25715 33563 25721
rect 35437 25755 35495 25761
rect 35437 25721 35449 25755
rect 35483 25752 35495 25755
rect 35710 25752 35716 25764
rect 35483 25724 35716 25752
rect 35483 25721 35495 25724
rect 35437 25715 35495 25721
rect 35710 25712 35716 25724
rect 35768 25712 35774 25764
rect 1946 25644 1952 25696
rect 2004 25684 2010 25696
rect 2501 25687 2559 25693
rect 2501 25684 2513 25687
rect 2004 25656 2513 25684
rect 2004 25644 2010 25656
rect 2501 25653 2513 25656
rect 2547 25653 2559 25687
rect 2501 25647 2559 25653
rect 6549 25687 6607 25693
rect 6549 25653 6561 25687
rect 6595 25684 6607 25687
rect 6822 25684 6828 25696
rect 6595 25656 6828 25684
rect 6595 25653 6607 25656
rect 6549 25647 6607 25653
rect 6822 25644 6828 25656
rect 6880 25644 6886 25696
rect 9030 25644 9036 25696
rect 9088 25684 9094 25696
rect 9125 25687 9183 25693
rect 9125 25684 9137 25687
rect 9088 25656 9137 25684
rect 9088 25644 9094 25656
rect 9125 25653 9137 25656
rect 9171 25653 9183 25687
rect 9125 25647 9183 25653
rect 9674 25644 9680 25696
rect 9732 25684 9738 25696
rect 9769 25687 9827 25693
rect 9769 25684 9781 25687
rect 9732 25656 9781 25684
rect 9732 25644 9738 25656
rect 9769 25653 9781 25656
rect 9815 25653 9827 25687
rect 11606 25684 11612 25696
rect 11567 25656 11612 25684
rect 9769 25647 9827 25653
rect 11606 25644 11612 25656
rect 11664 25644 11670 25696
rect 13814 25684 13820 25696
rect 13775 25656 13820 25684
rect 13814 25644 13820 25656
rect 13872 25684 13878 25696
rect 14369 25687 14427 25693
rect 14369 25684 14381 25687
rect 13872 25656 14381 25684
rect 13872 25644 13878 25656
rect 14369 25653 14381 25656
rect 14415 25653 14427 25687
rect 15654 25684 15660 25696
rect 15615 25656 15660 25684
rect 14369 25647 14427 25653
rect 15654 25644 15660 25656
rect 15712 25644 15718 25696
rect 20254 25684 20260 25696
rect 20215 25656 20260 25684
rect 20254 25644 20260 25656
rect 20312 25644 20318 25696
rect 20714 25684 20720 25696
rect 20627 25656 20720 25684
rect 20714 25644 20720 25656
rect 20772 25684 20778 25696
rect 21275 25687 21333 25693
rect 21275 25684 21287 25687
rect 20772 25656 21287 25684
rect 20772 25644 20778 25656
rect 21275 25653 21287 25656
rect 21321 25684 21333 25687
rect 24305 25687 24363 25693
rect 24305 25684 24317 25687
rect 21321 25656 24317 25684
rect 21321 25653 21333 25656
rect 21275 25647 21333 25653
rect 24305 25653 24317 25656
rect 24351 25684 24363 25687
rect 24863 25687 24921 25693
rect 24863 25684 24875 25687
rect 24351 25656 24875 25684
rect 24351 25653 24363 25656
rect 24305 25647 24363 25653
rect 24863 25653 24875 25656
rect 24909 25684 24921 25687
rect 26602 25684 26608 25696
rect 24909 25656 26608 25684
rect 24909 25653 24921 25656
rect 24863 25647 24921 25653
rect 26602 25644 26608 25656
rect 26660 25644 26666 25696
rect 28902 25684 28908 25696
rect 28863 25656 28908 25684
rect 28902 25644 28908 25656
rect 28960 25644 28966 25696
rect 31110 25684 31116 25696
rect 31071 25656 31116 25684
rect 31110 25644 31116 25656
rect 31168 25644 31174 25696
rect 32858 25684 32864 25696
rect 32819 25656 32864 25684
rect 32858 25644 32864 25656
rect 32916 25644 32922 25696
rect 33134 25644 33140 25696
rect 33192 25684 33198 25696
rect 33413 25687 33471 25693
rect 33413 25684 33425 25687
rect 33192 25656 33425 25684
rect 33192 25644 33198 25656
rect 33413 25653 33425 25656
rect 33459 25653 33471 25687
rect 36814 25684 36820 25696
rect 36775 25656 36820 25684
rect 33413 25647 33471 25653
rect 36814 25644 36820 25656
rect 36872 25644 36878 25696
rect 1104 25594 38824 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 38824 25594
rect 1104 25520 38824 25542
rect 6549 25483 6607 25489
rect 6549 25449 6561 25483
rect 6595 25480 6607 25483
rect 7098 25480 7104 25492
rect 6595 25452 7104 25480
rect 6595 25449 6607 25452
rect 6549 25443 6607 25449
rect 7098 25440 7104 25452
rect 7156 25480 7162 25492
rect 8113 25483 8171 25489
rect 8113 25480 8125 25483
rect 7156 25452 8125 25480
rect 7156 25440 7162 25452
rect 8113 25449 8125 25452
rect 8159 25449 8171 25483
rect 8113 25443 8171 25449
rect 8570 25440 8576 25492
rect 8628 25480 8634 25492
rect 8665 25483 8723 25489
rect 8665 25480 8677 25483
rect 8628 25452 8677 25480
rect 8628 25440 8634 25452
rect 8665 25449 8677 25452
rect 8711 25449 8723 25483
rect 8665 25443 8723 25449
rect 10045 25483 10103 25489
rect 10045 25449 10057 25483
rect 10091 25480 10103 25483
rect 11606 25480 11612 25492
rect 10091 25452 11612 25480
rect 10091 25449 10103 25452
rect 10045 25443 10103 25449
rect 11606 25440 11612 25452
rect 11664 25440 11670 25492
rect 13538 25480 13544 25492
rect 13499 25452 13544 25480
rect 13538 25440 13544 25452
rect 13596 25440 13602 25492
rect 14550 25480 14556 25492
rect 14511 25452 14556 25480
rect 14550 25440 14556 25452
rect 14608 25440 14614 25492
rect 18414 25480 18420 25492
rect 18375 25452 18420 25480
rect 18414 25440 18420 25452
rect 18472 25440 18478 25492
rect 19334 25480 19340 25492
rect 19295 25452 19340 25480
rect 19334 25440 19340 25452
rect 19392 25440 19398 25492
rect 20070 25480 20076 25492
rect 20031 25452 20076 25480
rect 20070 25440 20076 25452
rect 20128 25440 20134 25492
rect 20717 25483 20775 25489
rect 20717 25449 20729 25483
rect 20763 25480 20775 25483
rect 20806 25480 20812 25492
rect 20763 25452 20812 25480
rect 20763 25449 20775 25452
rect 20717 25443 20775 25449
rect 20806 25440 20812 25452
rect 20864 25440 20870 25492
rect 22094 25440 22100 25492
rect 22152 25480 22158 25492
rect 22281 25483 22339 25489
rect 22281 25480 22293 25483
rect 22152 25452 22293 25480
rect 22152 25440 22158 25452
rect 22281 25449 22293 25452
rect 22327 25449 22339 25483
rect 24118 25480 24124 25492
rect 24079 25452 24124 25480
rect 22281 25443 22339 25449
rect 24118 25440 24124 25452
rect 24176 25440 24182 25492
rect 24302 25440 24308 25492
rect 24360 25480 24366 25492
rect 24397 25483 24455 25489
rect 24397 25480 24409 25483
rect 24360 25452 24409 25480
rect 24360 25440 24366 25452
rect 24397 25449 24409 25452
rect 24443 25449 24455 25483
rect 24578 25480 24584 25492
rect 24539 25452 24584 25480
rect 24397 25443 24455 25449
rect 24578 25440 24584 25452
rect 24636 25440 24642 25492
rect 25222 25440 25228 25492
rect 25280 25480 25286 25492
rect 26145 25483 26203 25489
rect 26145 25480 26157 25483
rect 25280 25452 26157 25480
rect 25280 25440 25286 25452
rect 26145 25449 26157 25452
rect 26191 25449 26203 25483
rect 26145 25443 26203 25449
rect 26789 25483 26847 25489
rect 26789 25449 26801 25483
rect 26835 25480 26847 25483
rect 26970 25480 26976 25492
rect 26835 25452 26976 25480
rect 26835 25449 26847 25452
rect 26789 25443 26847 25449
rect 26970 25440 26976 25452
rect 27028 25480 27034 25492
rect 27065 25483 27123 25489
rect 27065 25480 27077 25483
rect 27028 25452 27077 25480
rect 27028 25440 27034 25452
rect 27065 25449 27077 25452
rect 27111 25449 27123 25483
rect 27065 25443 27123 25449
rect 27249 25483 27307 25489
rect 27249 25449 27261 25483
rect 27295 25480 27307 25483
rect 27522 25480 27528 25492
rect 27295 25452 27528 25480
rect 27295 25449 27307 25452
rect 27249 25443 27307 25449
rect 12434 25412 12440 25424
rect 11624 25384 12440 25412
rect 6638 25304 6644 25356
rect 6696 25344 6702 25356
rect 6733 25347 6791 25353
rect 6733 25344 6745 25347
rect 6696 25316 6745 25344
rect 6696 25304 6702 25316
rect 6733 25313 6745 25316
rect 6779 25313 6791 25347
rect 6733 25307 6791 25313
rect 6822 25304 6828 25356
rect 6880 25344 6886 25356
rect 6989 25347 7047 25353
rect 6989 25344 7001 25347
rect 6880 25316 7001 25344
rect 6880 25304 6886 25316
rect 6989 25313 7001 25316
rect 7035 25313 7047 25347
rect 6989 25307 7047 25313
rect 10134 25304 10140 25356
rect 10192 25344 10198 25356
rect 11624 25353 11652 25384
rect 12434 25372 12440 25384
rect 12492 25372 12498 25424
rect 15740 25415 15798 25421
rect 15740 25381 15752 25415
rect 15786 25412 15798 25415
rect 16022 25412 16028 25424
rect 15786 25384 16028 25412
rect 15786 25381 15798 25384
rect 15740 25375 15798 25381
rect 16022 25372 16028 25384
rect 16080 25372 16086 25424
rect 19886 25372 19892 25424
rect 19944 25412 19950 25424
rect 21146 25415 21204 25421
rect 21146 25412 21158 25415
rect 19944 25384 21158 25412
rect 19944 25372 19950 25384
rect 21146 25381 21158 25384
rect 21192 25412 21204 25415
rect 21450 25412 21456 25424
rect 21192 25384 21456 25412
rect 21192 25381 21204 25384
rect 21146 25375 21204 25381
rect 21450 25372 21456 25384
rect 21508 25372 21514 25424
rect 11882 25353 11888 25356
rect 10413 25347 10471 25353
rect 10413 25344 10425 25347
rect 10192 25316 10425 25344
rect 10192 25304 10198 25316
rect 10413 25313 10425 25316
rect 10459 25313 10471 25347
rect 10413 25307 10471 25313
rect 11609 25347 11667 25353
rect 11609 25313 11621 25347
rect 11655 25313 11667 25347
rect 11876 25344 11888 25353
rect 11843 25316 11888 25344
rect 11609 25307 11667 25313
rect 11876 25307 11888 25316
rect 11882 25304 11888 25307
rect 11940 25304 11946 25356
rect 14458 25304 14464 25356
rect 14516 25344 14522 25356
rect 14737 25347 14795 25353
rect 14737 25344 14749 25347
rect 14516 25316 14749 25344
rect 14516 25304 14522 25316
rect 14737 25313 14749 25316
rect 14783 25313 14795 25347
rect 14737 25307 14795 25313
rect 18325 25347 18383 25353
rect 18325 25313 18337 25347
rect 18371 25344 18383 25347
rect 18598 25344 18604 25356
rect 18371 25316 18604 25344
rect 18371 25313 18383 25316
rect 18325 25307 18383 25313
rect 18598 25304 18604 25316
rect 18656 25304 18662 25356
rect 24762 25304 24768 25356
rect 24820 25344 24826 25356
rect 24949 25347 25007 25353
rect 24949 25344 24961 25347
rect 24820 25316 24961 25344
rect 24820 25304 24826 25316
rect 24949 25313 24961 25316
rect 24995 25313 25007 25347
rect 24949 25307 25007 25313
rect 26234 25304 26240 25356
rect 26292 25344 26298 25356
rect 26329 25347 26387 25353
rect 26329 25344 26341 25347
rect 26292 25316 26341 25344
rect 26292 25304 26298 25316
rect 26329 25313 26341 25316
rect 26375 25344 26387 25347
rect 27264 25344 27292 25443
rect 27522 25440 27528 25452
rect 27580 25440 27586 25492
rect 27706 25480 27712 25492
rect 27667 25452 27712 25480
rect 27706 25440 27712 25452
rect 27764 25440 27770 25492
rect 29730 25480 29736 25492
rect 29691 25452 29736 25480
rect 29730 25440 29736 25452
rect 29788 25440 29794 25492
rect 30190 25480 30196 25492
rect 30151 25452 30196 25480
rect 30190 25440 30196 25452
rect 30248 25440 30254 25492
rect 31662 25480 31668 25492
rect 31623 25452 31668 25480
rect 31662 25440 31668 25452
rect 31720 25440 31726 25492
rect 31754 25440 31760 25492
rect 31812 25480 31818 25492
rect 33781 25483 33839 25489
rect 31812 25452 31857 25480
rect 31812 25440 31818 25452
rect 33781 25449 33793 25483
rect 33827 25449 33839 25483
rect 34238 25480 34244 25492
rect 34199 25452 34244 25480
rect 33781 25443 33839 25449
rect 29748 25412 29776 25440
rect 30561 25415 30619 25421
rect 30561 25412 30573 25415
rect 29748 25384 30573 25412
rect 30561 25381 30573 25384
rect 30607 25412 30619 25415
rect 31110 25412 31116 25424
rect 30607 25384 31116 25412
rect 30607 25381 30619 25384
rect 30561 25375 30619 25381
rect 31110 25372 31116 25384
rect 31168 25372 31174 25424
rect 31297 25415 31355 25421
rect 31297 25381 31309 25415
rect 31343 25412 31355 25415
rect 31570 25412 31576 25424
rect 31343 25384 31576 25412
rect 31343 25381 31355 25384
rect 31297 25375 31355 25381
rect 31570 25372 31576 25384
rect 31628 25372 31634 25424
rect 33796 25412 33824 25443
rect 34238 25440 34244 25452
rect 34296 25440 34302 25492
rect 34606 25440 34612 25492
rect 34664 25480 34670 25492
rect 34793 25483 34851 25489
rect 34793 25480 34805 25483
rect 34664 25452 34805 25480
rect 34664 25440 34670 25452
rect 34793 25449 34805 25452
rect 34839 25449 34851 25483
rect 35250 25480 35256 25492
rect 35211 25452 35256 25480
rect 34793 25443 34851 25449
rect 35250 25440 35256 25452
rect 35308 25440 35314 25492
rect 33870 25412 33876 25424
rect 33783 25384 33876 25412
rect 33870 25372 33876 25384
rect 33928 25412 33934 25424
rect 33928 25384 35756 25412
rect 33928 25372 33934 25384
rect 26375 25316 27292 25344
rect 26375 25313 26387 25316
rect 26329 25307 26387 25313
rect 27338 25304 27344 25356
rect 27396 25344 27402 25356
rect 27433 25347 27491 25353
rect 27433 25344 27445 25347
rect 27396 25316 27445 25344
rect 27396 25304 27402 25316
rect 27433 25313 27445 25316
rect 27479 25344 27491 25347
rect 28902 25344 28908 25356
rect 27479 25316 28908 25344
rect 27479 25313 27491 25316
rect 27433 25307 27491 25313
rect 28902 25304 28908 25316
rect 28960 25304 28966 25356
rect 29365 25347 29423 25353
rect 29365 25313 29377 25347
rect 29411 25344 29423 25347
rect 29822 25344 29828 25356
rect 29411 25316 29828 25344
rect 29411 25313 29423 25316
rect 29365 25307 29423 25313
rect 29822 25304 29828 25316
rect 29880 25304 29886 25356
rect 30006 25304 30012 25356
rect 30064 25344 30070 25356
rect 30101 25347 30159 25353
rect 30101 25344 30113 25347
rect 30064 25316 30113 25344
rect 30064 25304 30070 25316
rect 30101 25313 30113 25316
rect 30147 25344 30159 25347
rect 30650 25344 30656 25356
rect 30147 25316 30656 25344
rect 30147 25313 30159 25316
rect 30101 25307 30159 25313
rect 30650 25304 30656 25316
rect 30708 25304 30714 25356
rect 31938 25353 31944 25356
rect 31933 25344 31944 25353
rect 31899 25316 31944 25344
rect 31933 25307 31944 25316
rect 31938 25304 31944 25307
rect 31996 25304 32002 25356
rect 32490 25344 32496 25356
rect 32451 25316 32496 25344
rect 32490 25304 32496 25316
rect 32548 25304 32554 25356
rect 34054 25304 34060 25356
rect 34112 25344 34118 25356
rect 35728 25353 35756 25384
rect 34149 25347 34207 25353
rect 34149 25344 34161 25347
rect 34112 25316 34161 25344
rect 34112 25304 34118 25316
rect 34149 25313 34161 25316
rect 34195 25313 34207 25347
rect 34149 25307 34207 25313
rect 35713 25347 35771 25353
rect 35713 25313 35725 25347
rect 35759 25344 35771 25347
rect 35894 25344 35900 25356
rect 35759 25316 35900 25344
rect 35759 25313 35771 25316
rect 35713 25307 35771 25313
rect 35894 25304 35900 25316
rect 35952 25304 35958 25356
rect 10502 25276 10508 25288
rect 10463 25248 10508 25276
rect 10502 25236 10508 25248
rect 10560 25236 10566 25288
rect 10594 25236 10600 25288
rect 10652 25276 10658 25288
rect 10652 25248 10697 25276
rect 10652 25236 10658 25248
rect 15378 25236 15384 25288
rect 15436 25276 15442 25288
rect 15473 25279 15531 25285
rect 15473 25276 15485 25279
rect 15436 25248 15485 25276
rect 15436 25236 15442 25248
rect 15473 25245 15485 25248
rect 15519 25245 15531 25279
rect 15473 25239 15531 25245
rect 17954 25236 17960 25288
rect 18012 25276 18018 25288
rect 18509 25279 18567 25285
rect 18509 25276 18521 25279
rect 18012 25248 18521 25276
rect 18012 25236 18018 25248
rect 18509 25245 18521 25248
rect 18555 25245 18567 25279
rect 18509 25239 18567 25245
rect 19613 25279 19671 25285
rect 19613 25245 19625 25279
rect 19659 25276 19671 25279
rect 20714 25276 20720 25288
rect 19659 25248 20720 25276
rect 19659 25245 19671 25248
rect 19613 25239 19671 25245
rect 20714 25236 20720 25248
rect 20772 25236 20778 25288
rect 20898 25276 20904 25288
rect 20859 25248 20904 25276
rect 20898 25236 20904 25248
rect 20956 25236 20962 25288
rect 25038 25276 25044 25288
rect 24999 25248 25044 25276
rect 25038 25236 25044 25248
rect 25096 25236 25102 25288
rect 25225 25279 25283 25285
rect 25225 25245 25237 25279
rect 25271 25276 25283 25279
rect 26142 25276 26148 25288
rect 25271 25248 26148 25276
rect 25271 25245 25283 25248
rect 25225 25239 25283 25245
rect 24854 25168 24860 25220
rect 24912 25208 24918 25220
rect 25240 25208 25268 25239
rect 26142 25236 26148 25248
rect 26200 25236 26206 25288
rect 30834 25276 30840 25288
rect 30795 25248 30840 25276
rect 30834 25236 30840 25248
rect 30892 25236 30898 25288
rect 32122 25236 32128 25288
rect 32180 25276 32186 25288
rect 32585 25279 32643 25285
rect 32585 25276 32597 25279
rect 32180 25248 32597 25276
rect 32180 25236 32186 25248
rect 32585 25245 32597 25248
rect 32631 25245 32643 25279
rect 32585 25239 32643 25245
rect 32677 25279 32735 25285
rect 32677 25245 32689 25279
rect 32723 25245 32735 25279
rect 32677 25239 32735 25245
rect 24912 25180 25268 25208
rect 24912 25168 24918 25180
rect 31570 25168 31576 25220
rect 31628 25208 31634 25220
rect 32692 25208 32720 25239
rect 34330 25236 34336 25288
rect 34388 25276 34394 25288
rect 35805 25279 35863 25285
rect 34388 25248 34433 25276
rect 34388 25236 34394 25248
rect 35805 25245 35817 25279
rect 35851 25245 35863 25279
rect 35805 25239 35863 25245
rect 35989 25279 36047 25285
rect 35989 25245 36001 25279
rect 36035 25276 36047 25279
rect 36814 25276 36820 25288
rect 36035 25248 36820 25276
rect 36035 25245 36047 25248
rect 35989 25239 36047 25245
rect 31628 25180 32720 25208
rect 33597 25211 33655 25217
rect 31628 25168 31634 25180
rect 33597 25177 33609 25211
rect 33643 25208 33655 25211
rect 33686 25208 33692 25220
rect 33643 25180 33692 25208
rect 33643 25177 33655 25180
rect 33597 25171 33655 25177
rect 33686 25168 33692 25180
rect 33744 25208 33750 25220
rect 34348 25208 34376 25236
rect 33744 25180 34376 25208
rect 33744 25168 33750 25180
rect 34514 25168 34520 25220
rect 34572 25208 34578 25220
rect 35345 25211 35403 25217
rect 35345 25208 35357 25211
rect 34572 25180 35357 25208
rect 34572 25168 34578 25180
rect 35345 25177 35357 25180
rect 35391 25177 35403 25211
rect 35345 25171 35403 25177
rect 35710 25168 35716 25220
rect 35768 25208 35774 25220
rect 35820 25208 35848 25239
rect 36814 25236 36820 25248
rect 36872 25236 36878 25288
rect 35768 25180 35848 25208
rect 35768 25168 35774 25180
rect 1673 25143 1731 25149
rect 1673 25109 1685 25143
rect 1719 25140 1731 25143
rect 1946 25140 1952 25152
rect 1719 25112 1952 25140
rect 1719 25109 1731 25112
rect 1673 25103 1731 25109
rect 1946 25100 1952 25112
rect 2004 25100 2010 25152
rect 9401 25143 9459 25149
rect 9401 25109 9413 25143
rect 9447 25140 9459 25143
rect 9674 25140 9680 25152
rect 9447 25112 9680 25140
rect 9447 25109 9459 25112
rect 9401 25103 9459 25109
rect 9674 25100 9680 25112
rect 9732 25100 9738 25152
rect 9953 25143 10011 25149
rect 9953 25109 9965 25143
rect 9999 25140 10011 25143
rect 10134 25140 10140 25152
rect 9999 25112 10140 25140
rect 9999 25109 10011 25112
rect 9953 25103 10011 25109
rect 10134 25100 10140 25112
rect 10192 25100 10198 25152
rect 12986 25140 12992 25152
rect 12947 25112 12992 25140
rect 12986 25100 12992 25112
rect 13044 25100 13050 25152
rect 16574 25100 16580 25152
rect 16632 25140 16638 25152
rect 16853 25143 16911 25149
rect 16853 25140 16865 25143
rect 16632 25112 16865 25140
rect 16632 25100 16638 25112
rect 16853 25109 16865 25112
rect 16899 25109 16911 25143
rect 16853 25103 16911 25109
rect 17862 25100 17868 25152
rect 17920 25140 17926 25152
rect 17957 25143 18015 25149
rect 17957 25140 17969 25143
rect 17920 25112 17969 25140
rect 17920 25100 17926 25112
rect 17957 25109 17969 25112
rect 18003 25109 18015 25143
rect 17957 25103 18015 25109
rect 28997 25143 29055 25149
rect 28997 25109 29009 25143
rect 29043 25140 29055 25143
rect 29178 25140 29184 25152
rect 29043 25112 29184 25140
rect 29043 25109 29055 25112
rect 28997 25103 29055 25109
rect 29178 25100 29184 25112
rect 29236 25100 29242 25152
rect 32125 25143 32183 25149
rect 32125 25109 32137 25143
rect 32171 25140 32183 25143
rect 32214 25140 32220 25152
rect 32171 25112 32220 25140
rect 32171 25109 32183 25112
rect 32125 25103 32183 25109
rect 32214 25100 32220 25112
rect 32272 25100 32278 25152
rect 33134 25140 33140 25152
rect 33095 25112 33140 25140
rect 33134 25100 33140 25112
rect 33192 25100 33198 25152
rect 1104 25050 38824 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 34966 25050
rect 35018 24998 35030 25050
rect 35082 24998 35094 25050
rect 35146 24998 35158 25050
rect 35210 24998 38824 25050
rect 1104 24976 38824 24998
rect 5905 24939 5963 24945
rect 5905 24905 5917 24939
rect 5951 24936 5963 24939
rect 6181 24939 6239 24945
rect 6181 24936 6193 24939
rect 5951 24908 6193 24936
rect 5951 24905 5963 24908
rect 5905 24899 5963 24905
rect 6181 24905 6193 24908
rect 6227 24936 6239 24939
rect 6638 24936 6644 24948
rect 6227 24908 6644 24936
rect 6227 24905 6239 24908
rect 6181 24899 6239 24905
rect 6564 24732 6592 24908
rect 6638 24896 6644 24908
rect 6696 24896 6702 24948
rect 6822 24896 6828 24948
rect 6880 24936 6886 24948
rect 8297 24939 8355 24945
rect 8297 24936 8309 24939
rect 6880 24908 8309 24936
rect 6880 24896 6886 24908
rect 8297 24905 8309 24908
rect 8343 24905 8355 24939
rect 8297 24899 8355 24905
rect 8570 24896 8576 24948
rect 8628 24936 8634 24948
rect 8941 24939 8999 24945
rect 8941 24936 8953 24939
rect 8628 24908 8953 24936
rect 8628 24896 8634 24908
rect 8941 24905 8953 24908
rect 8987 24905 8999 24939
rect 8941 24899 8999 24905
rect 9769 24939 9827 24945
rect 9769 24905 9781 24939
rect 9815 24936 9827 24939
rect 10502 24936 10508 24948
rect 9815 24908 10508 24936
rect 9815 24905 9827 24908
rect 9769 24899 9827 24905
rect 10502 24896 10508 24908
rect 10560 24896 10566 24948
rect 11882 24936 11888 24948
rect 11843 24908 11888 24936
rect 11882 24896 11888 24908
rect 11940 24896 11946 24948
rect 12710 24936 12716 24948
rect 12268 24908 12716 24936
rect 6641 24803 6699 24809
rect 6641 24769 6653 24803
rect 6687 24800 6699 24803
rect 9401 24803 9459 24809
rect 6687 24772 7052 24800
rect 6687 24769 6699 24772
rect 6641 24763 6699 24769
rect 6914 24732 6920 24744
rect 6564 24704 6920 24732
rect 6914 24692 6920 24704
rect 6972 24692 6978 24744
rect 7024 24732 7052 24772
rect 9401 24769 9413 24803
rect 9447 24800 9459 24803
rect 9447 24772 9996 24800
rect 9447 24769 9459 24772
rect 9401 24763 9459 24769
rect 7184 24735 7242 24741
rect 7184 24732 7196 24735
rect 7024 24704 7196 24732
rect 7184 24701 7196 24704
rect 7230 24732 7242 24735
rect 9030 24732 9036 24744
rect 7230 24704 9036 24732
rect 7230 24701 7242 24704
rect 7184 24695 7242 24701
rect 9030 24692 9036 24704
rect 9088 24692 9094 24744
rect 9858 24732 9864 24744
rect 9819 24704 9864 24732
rect 9858 24692 9864 24704
rect 9916 24692 9922 24744
rect 9968 24732 9996 24772
rect 10134 24741 10140 24744
rect 10128 24732 10140 24741
rect 9968 24704 10140 24732
rect 10128 24695 10140 24704
rect 10134 24692 10140 24695
rect 10192 24692 10198 24744
rect 10502 24692 10508 24744
rect 10560 24732 10566 24744
rect 12161 24735 12219 24741
rect 12161 24732 12173 24735
rect 10560 24704 12173 24732
rect 10560 24692 10566 24704
rect 12161 24701 12173 24704
rect 12207 24732 12219 24735
rect 12268 24732 12296 24908
rect 12710 24896 12716 24908
rect 12768 24896 12774 24948
rect 15102 24936 15108 24948
rect 15063 24908 15108 24936
rect 15102 24896 15108 24908
rect 15160 24896 15166 24948
rect 18325 24939 18383 24945
rect 18325 24905 18337 24939
rect 18371 24936 18383 24939
rect 18414 24936 18420 24948
rect 18371 24908 18420 24936
rect 18371 24905 18383 24908
rect 18325 24899 18383 24905
rect 18414 24896 18420 24908
rect 18472 24896 18478 24948
rect 19153 24939 19211 24945
rect 19153 24905 19165 24939
rect 19199 24936 19211 24939
rect 20254 24936 20260 24948
rect 19199 24908 20260 24936
rect 19199 24905 19211 24908
rect 19153 24899 19211 24905
rect 20254 24896 20260 24908
rect 20312 24936 20318 24948
rect 21266 24936 21272 24948
rect 20312 24908 21272 24936
rect 20312 24896 20318 24908
rect 21266 24896 21272 24908
rect 21324 24896 21330 24948
rect 21450 24936 21456 24948
rect 21411 24908 21456 24936
rect 21450 24896 21456 24908
rect 21508 24936 21514 24948
rect 22005 24939 22063 24945
rect 22005 24936 22017 24939
rect 21508 24908 22017 24936
rect 21508 24896 21514 24908
rect 22005 24905 22017 24908
rect 22051 24905 22063 24939
rect 27338 24936 27344 24948
rect 27299 24908 27344 24936
rect 22005 24899 22063 24905
rect 27338 24896 27344 24908
rect 27396 24896 27402 24948
rect 30650 24896 30656 24948
rect 30708 24936 30714 24948
rect 31021 24939 31079 24945
rect 31021 24936 31033 24939
rect 30708 24908 31033 24936
rect 30708 24896 30714 24908
rect 31021 24905 31033 24908
rect 31067 24905 31079 24939
rect 31021 24899 31079 24905
rect 31938 24896 31944 24948
rect 31996 24936 32002 24948
rect 32125 24939 32183 24945
rect 32125 24936 32137 24939
rect 31996 24908 32137 24936
rect 31996 24896 32002 24908
rect 32125 24905 32137 24908
rect 32171 24936 32183 24939
rect 32490 24936 32496 24948
rect 32171 24908 32496 24936
rect 32171 24905 32183 24908
rect 32125 24899 32183 24905
rect 32490 24896 32496 24908
rect 32548 24896 32554 24948
rect 33597 24939 33655 24945
rect 33597 24905 33609 24939
rect 33643 24936 33655 24939
rect 33873 24939 33931 24945
rect 33873 24936 33885 24939
rect 33643 24908 33885 24936
rect 33643 24905 33655 24908
rect 33597 24899 33655 24905
rect 33873 24905 33885 24908
rect 33919 24936 33931 24939
rect 34054 24936 34060 24948
rect 33919 24908 34060 24936
rect 33919 24905 33931 24908
rect 33873 24899 33931 24905
rect 34054 24896 34060 24908
rect 34112 24896 34118 24948
rect 34238 24936 34244 24948
rect 34199 24908 34244 24936
rect 34238 24896 34244 24908
rect 34296 24896 34302 24948
rect 36814 24896 36820 24948
rect 36872 24936 36878 24948
rect 37001 24939 37059 24945
rect 37001 24936 37013 24939
rect 36872 24908 37013 24936
rect 36872 24896 36878 24908
rect 37001 24905 37013 24908
rect 37047 24905 37059 24939
rect 37001 24899 37059 24905
rect 25038 24868 25044 24880
rect 24596 24840 25044 24868
rect 23937 24803 23995 24809
rect 23937 24769 23949 24803
rect 23983 24800 23995 24803
rect 24596 24800 24624 24840
rect 25038 24828 25044 24840
rect 25096 24828 25102 24880
rect 23983 24772 24624 24800
rect 24673 24803 24731 24809
rect 23983 24769 23995 24772
rect 23937 24763 23995 24769
rect 24673 24769 24685 24803
rect 24719 24800 24731 24803
rect 24762 24800 24768 24812
rect 24719 24772 24768 24800
rect 24719 24769 24731 24772
rect 24673 24763 24731 24769
rect 24762 24760 24768 24772
rect 24820 24760 24826 24812
rect 32674 24800 32680 24812
rect 32635 24772 32680 24800
rect 32674 24760 32680 24772
rect 32732 24760 32738 24812
rect 34606 24760 34612 24812
rect 34664 24800 34670 24812
rect 35069 24803 35127 24809
rect 35069 24800 35081 24803
rect 34664 24772 35081 24800
rect 34664 24760 34670 24772
rect 35069 24769 35081 24772
rect 35115 24769 35127 24803
rect 35069 24763 35127 24769
rect 12710 24741 12716 24744
rect 12437 24735 12495 24741
rect 12437 24732 12449 24735
rect 12207 24704 12296 24732
rect 12360 24704 12449 24732
rect 12207 24701 12219 24704
rect 12161 24695 12219 24701
rect 12360 24664 12388 24704
rect 12437 24701 12449 24704
rect 12483 24701 12495 24735
rect 12704 24732 12716 24741
rect 12623 24704 12716 24732
rect 12437 24695 12495 24701
rect 12704 24695 12716 24704
rect 12768 24732 12774 24744
rect 12986 24732 12992 24744
rect 12768 24704 12992 24732
rect 12710 24692 12716 24695
rect 12768 24692 12774 24704
rect 12986 24692 12992 24704
rect 13044 24692 13050 24744
rect 15289 24735 15347 24741
rect 15289 24701 15301 24735
rect 15335 24732 15347 24735
rect 15378 24732 15384 24744
rect 15335 24704 15384 24732
rect 15335 24701 15347 24704
rect 15289 24695 15347 24701
rect 15378 24692 15384 24704
rect 15436 24732 15442 24744
rect 18966 24732 18972 24744
rect 15436 24704 17356 24732
rect 18927 24704 18972 24732
rect 15436 24692 15442 24704
rect 14829 24667 14887 24673
rect 12360 24636 12572 24664
rect 11238 24596 11244 24608
rect 11199 24568 11244 24596
rect 11238 24556 11244 24568
rect 11296 24556 11302 24608
rect 12434 24556 12440 24608
rect 12492 24596 12498 24608
rect 12544 24596 12572 24636
rect 14829 24633 14841 24667
rect 14875 24664 14887 24667
rect 15556 24667 15614 24673
rect 15556 24664 15568 24667
rect 14875 24636 15568 24664
rect 14875 24633 14887 24636
rect 14829 24627 14887 24633
rect 15556 24633 15568 24636
rect 15602 24664 15614 24667
rect 15930 24664 15936 24676
rect 15602 24636 15936 24664
rect 15602 24633 15614 24636
rect 15556 24627 15614 24633
rect 15930 24624 15936 24636
rect 15988 24624 15994 24676
rect 17328 24673 17356 24704
rect 18966 24692 18972 24704
rect 19024 24732 19030 24744
rect 19521 24735 19579 24741
rect 19521 24732 19533 24735
rect 19024 24704 19533 24732
rect 19024 24692 19030 24704
rect 19521 24701 19533 24704
rect 19567 24701 19579 24735
rect 19521 24695 19579 24701
rect 19886 24692 19892 24744
rect 19944 24732 19950 24744
rect 20073 24735 20131 24741
rect 20073 24732 20085 24735
rect 19944 24704 20085 24732
rect 19944 24692 19950 24704
rect 20073 24701 20085 24704
rect 20119 24732 20131 24735
rect 20898 24732 20904 24744
rect 20119 24704 20904 24732
rect 20119 24701 20131 24704
rect 20073 24695 20131 24701
rect 20898 24692 20904 24704
rect 20956 24692 20962 24744
rect 24305 24735 24363 24741
rect 24305 24701 24317 24735
rect 24351 24732 24363 24735
rect 24854 24732 24860 24744
rect 24351 24704 24860 24732
rect 24351 24701 24363 24704
rect 24305 24695 24363 24701
rect 24854 24692 24860 24704
rect 24912 24692 24918 24744
rect 25041 24735 25099 24741
rect 25041 24701 25053 24735
rect 25087 24732 25099 24735
rect 25130 24732 25136 24744
rect 25087 24704 25136 24732
rect 25087 24701 25099 24704
rect 25041 24695 25099 24701
rect 25130 24692 25136 24704
rect 25188 24692 25194 24744
rect 25314 24741 25320 24744
rect 25308 24732 25320 24741
rect 25275 24704 25320 24732
rect 25308 24695 25320 24704
rect 25314 24692 25320 24695
rect 25372 24692 25378 24744
rect 29641 24735 29699 24741
rect 29641 24701 29653 24735
rect 29687 24732 29699 24735
rect 29730 24732 29736 24744
rect 29687 24704 29736 24732
rect 29687 24701 29699 24704
rect 29641 24695 29699 24701
rect 29730 24692 29736 24704
rect 29788 24692 29794 24744
rect 32493 24735 32551 24741
rect 32493 24732 32505 24735
rect 31588 24704 32505 24732
rect 17313 24667 17371 24673
rect 17313 24633 17325 24667
rect 17359 24664 17371 24667
rect 19904 24664 19932 24692
rect 17359 24636 19932 24664
rect 19981 24667 20039 24673
rect 17359 24633 17371 24636
rect 17313 24627 17371 24633
rect 19981 24633 19993 24667
rect 20027 24664 20039 24667
rect 20254 24664 20260 24676
rect 20027 24636 20260 24664
rect 20027 24633 20039 24636
rect 19981 24627 20039 24633
rect 20254 24624 20260 24636
rect 20312 24673 20318 24676
rect 20312 24667 20376 24673
rect 20312 24633 20330 24667
rect 20364 24633 20376 24667
rect 20312 24627 20376 24633
rect 29549 24667 29607 24673
rect 29549 24633 29561 24667
rect 29595 24664 29607 24667
rect 29886 24667 29944 24673
rect 29886 24664 29898 24667
rect 29595 24636 29898 24664
rect 29595 24633 29607 24636
rect 29549 24627 29607 24633
rect 29886 24633 29898 24636
rect 29932 24664 29944 24667
rect 30926 24664 30932 24676
rect 29932 24636 30932 24664
rect 29932 24633 29944 24636
rect 29886 24627 29944 24633
rect 20312 24624 20318 24627
rect 30926 24624 30932 24636
rect 30984 24664 30990 24676
rect 31588 24673 31616 24704
rect 32493 24701 32505 24704
rect 32539 24701 32551 24735
rect 32493 24695 32551 24701
rect 33689 24735 33747 24741
rect 33689 24701 33701 24735
rect 33735 24732 33747 24735
rect 33778 24732 33784 24744
rect 33735 24704 33784 24732
rect 33735 24701 33747 24704
rect 33689 24695 33747 24701
rect 33778 24692 33784 24704
rect 33836 24732 33842 24744
rect 34422 24732 34428 24744
rect 33836 24704 34428 24732
rect 33836 24692 33842 24704
rect 34422 24692 34428 24704
rect 34480 24692 34486 24744
rect 31573 24667 31631 24673
rect 31573 24664 31585 24667
rect 30984 24636 31585 24664
rect 30984 24624 30990 24636
rect 31573 24633 31585 24636
rect 31619 24633 31631 24667
rect 31573 24627 31631 24633
rect 32033 24667 32091 24673
rect 32033 24633 32045 24667
rect 32079 24664 32091 24667
rect 32585 24667 32643 24673
rect 32585 24664 32597 24667
rect 32079 24636 32597 24664
rect 32079 24633 32091 24636
rect 32033 24627 32091 24633
rect 32585 24633 32597 24636
rect 32631 24633 32643 24667
rect 32585 24627 32643 24633
rect 34701 24667 34759 24673
rect 34701 24633 34713 24667
rect 34747 24664 34759 24667
rect 35336 24667 35394 24673
rect 35336 24664 35348 24667
rect 34747 24636 35348 24664
rect 34747 24633 34759 24636
rect 34701 24627 34759 24633
rect 35336 24633 35348 24636
rect 35382 24664 35394 24667
rect 35526 24664 35532 24676
rect 35382 24636 35532 24664
rect 35382 24633 35394 24636
rect 35336 24627 35394 24633
rect 13814 24596 13820 24608
rect 12492 24568 12572 24596
rect 13775 24568 13820 24596
rect 12492 24556 12498 24568
rect 13814 24556 13820 24568
rect 13872 24556 13878 24608
rect 14458 24596 14464 24608
rect 14419 24568 14464 24596
rect 14458 24556 14464 24568
rect 14516 24556 14522 24608
rect 16666 24596 16672 24608
rect 16627 24568 16672 24596
rect 16666 24556 16672 24568
rect 16724 24556 16730 24608
rect 17770 24596 17776 24608
rect 17731 24568 17776 24596
rect 17770 24556 17776 24568
rect 17828 24556 17834 24608
rect 18598 24596 18604 24608
rect 18559 24568 18604 24596
rect 18598 24556 18604 24568
rect 18656 24556 18662 24608
rect 22370 24596 22376 24608
rect 22331 24568 22376 24596
rect 22370 24556 22376 24568
rect 22428 24556 22434 24608
rect 26142 24556 26148 24608
rect 26200 24596 26206 24608
rect 26418 24596 26424 24608
rect 26200 24568 26424 24596
rect 26200 24556 26206 24568
rect 26418 24556 26424 24568
rect 26476 24556 26482 24608
rect 29089 24599 29147 24605
rect 29089 24565 29101 24599
rect 29135 24596 29147 24599
rect 30834 24596 30840 24608
rect 29135 24568 30840 24596
rect 29135 24565 29147 24568
rect 29089 24559 29147 24565
rect 30834 24556 30840 24568
rect 30892 24556 30898 24608
rect 31110 24556 31116 24608
rect 31168 24596 31174 24608
rect 32048 24596 32076 24627
rect 35526 24624 35532 24636
rect 35584 24624 35590 24676
rect 31168 24568 32076 24596
rect 31168 24556 31174 24568
rect 32122 24556 32128 24608
rect 32180 24596 32186 24608
rect 33137 24599 33195 24605
rect 33137 24596 33149 24599
rect 32180 24568 33149 24596
rect 32180 24556 32186 24568
rect 33137 24565 33149 24568
rect 33183 24565 33195 24599
rect 33137 24559 33195 24565
rect 35158 24556 35164 24608
rect 35216 24596 35222 24608
rect 36449 24599 36507 24605
rect 36449 24596 36461 24599
rect 35216 24568 36461 24596
rect 35216 24556 35222 24568
rect 36449 24565 36461 24568
rect 36495 24565 36507 24599
rect 36449 24559 36507 24565
rect 1104 24506 38824 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 38824 24506
rect 1104 24432 38824 24454
rect 6822 24392 6828 24404
rect 6783 24364 6828 24392
rect 6822 24352 6828 24364
rect 6880 24352 6886 24404
rect 8478 24392 8484 24404
rect 8439 24364 8484 24392
rect 8478 24352 8484 24364
rect 8536 24352 8542 24404
rect 11793 24395 11851 24401
rect 11793 24361 11805 24395
rect 11839 24392 11851 24395
rect 15470 24392 15476 24404
rect 11839 24364 12480 24392
rect 15431 24364 15476 24392
rect 11839 24361 11851 24364
rect 11793 24355 11851 24361
rect 12452 24336 12480 24364
rect 15470 24352 15476 24364
rect 15528 24352 15534 24404
rect 15930 24392 15936 24404
rect 15843 24364 15936 24392
rect 15930 24352 15936 24364
rect 15988 24392 15994 24404
rect 16482 24392 16488 24404
rect 15988 24364 16488 24392
rect 15988 24352 15994 24364
rect 16482 24352 16488 24364
rect 16540 24352 16546 24404
rect 20806 24352 20812 24404
rect 20864 24392 20870 24404
rect 20901 24395 20959 24401
rect 20901 24392 20913 24395
rect 20864 24364 20913 24392
rect 20864 24352 20870 24364
rect 20901 24361 20913 24364
rect 20947 24361 20959 24395
rect 20901 24355 20959 24361
rect 24673 24395 24731 24401
rect 24673 24361 24685 24395
rect 24719 24392 24731 24395
rect 24762 24392 24768 24404
rect 24719 24364 24768 24392
rect 24719 24361 24731 24364
rect 24673 24355 24731 24361
rect 24762 24352 24768 24364
rect 24820 24352 24826 24404
rect 25130 24352 25136 24404
rect 25188 24392 25194 24404
rect 25501 24395 25559 24401
rect 25501 24392 25513 24395
rect 25188 24364 25513 24392
rect 25188 24352 25194 24364
rect 25501 24361 25513 24364
rect 25547 24361 25559 24395
rect 26234 24392 26240 24404
rect 26195 24364 26240 24392
rect 25501 24355 25559 24361
rect 26234 24352 26240 24364
rect 26292 24352 26298 24404
rect 30926 24392 30932 24404
rect 30887 24364 30932 24392
rect 30926 24352 30932 24364
rect 30984 24352 30990 24404
rect 31938 24392 31944 24404
rect 31899 24364 31944 24392
rect 31938 24352 31944 24364
rect 31996 24352 32002 24404
rect 32122 24392 32128 24404
rect 32083 24364 32128 24392
rect 32122 24352 32128 24364
rect 32180 24352 32186 24404
rect 33778 24392 33784 24404
rect 33739 24364 33784 24392
rect 33778 24352 33784 24364
rect 33836 24352 33842 24404
rect 34149 24395 34207 24401
rect 34149 24361 34161 24395
rect 34195 24392 34207 24395
rect 34330 24392 34336 24404
rect 34195 24364 34336 24392
rect 34195 24361 34207 24364
rect 34149 24355 34207 24361
rect 34330 24352 34336 24364
rect 34388 24392 34394 24404
rect 36265 24395 36323 24401
rect 36265 24392 36277 24395
rect 34388 24364 36277 24392
rect 34388 24352 34394 24364
rect 36265 24361 36277 24364
rect 36311 24361 36323 24395
rect 36265 24355 36323 24361
rect 10036 24327 10094 24333
rect 7116 24296 7788 24324
rect 7116 24265 7144 24296
rect 7760 24268 7788 24296
rect 10036 24293 10048 24327
rect 10082 24324 10094 24327
rect 10594 24324 10600 24336
rect 10082 24296 10600 24324
rect 10082 24293 10094 24296
rect 10036 24287 10094 24293
rect 10594 24284 10600 24296
rect 10652 24324 10658 24336
rect 11238 24324 11244 24336
rect 10652 24296 11244 24324
rect 10652 24284 10658 24296
rect 11238 24284 11244 24296
rect 11296 24284 11302 24336
rect 12434 24284 12440 24336
rect 12492 24324 12498 24336
rect 12492 24296 12585 24324
rect 12492 24284 12498 24296
rect 14550 24284 14556 24336
rect 14608 24324 14614 24336
rect 14645 24327 14703 24333
rect 14645 24324 14657 24327
rect 14608 24296 14657 24324
rect 14608 24284 14614 24296
rect 14645 24293 14657 24296
rect 14691 24324 14703 24327
rect 15105 24327 15163 24333
rect 15105 24324 15117 24327
rect 14691 24296 15117 24324
rect 14691 24293 14703 24296
rect 14645 24287 14703 24293
rect 15105 24293 15117 24296
rect 15151 24324 15163 24327
rect 15378 24324 15384 24336
rect 15151 24296 15384 24324
rect 15151 24293 15163 24296
rect 15105 24287 15163 24293
rect 15378 24284 15384 24296
rect 15436 24284 15442 24336
rect 20714 24284 20720 24336
rect 20772 24324 20778 24336
rect 21269 24327 21327 24333
rect 21269 24324 21281 24327
rect 20772 24296 21281 24324
rect 20772 24284 20778 24296
rect 21269 24293 21281 24296
rect 21315 24293 21327 24327
rect 21269 24287 21327 24293
rect 25225 24327 25283 24333
rect 25225 24293 25237 24327
rect 25271 24324 25283 24327
rect 25314 24324 25320 24336
rect 25271 24296 25320 24324
rect 25271 24293 25283 24296
rect 25225 24287 25283 24293
rect 25314 24284 25320 24296
rect 25372 24284 25378 24336
rect 32030 24284 32036 24336
rect 32088 24324 32094 24336
rect 33137 24327 33195 24333
rect 33137 24324 33149 24327
rect 32088 24296 33149 24324
rect 32088 24284 32094 24296
rect 33137 24293 33149 24296
rect 33183 24293 33195 24327
rect 35894 24324 35900 24336
rect 35855 24296 35900 24324
rect 33137 24287 33195 24293
rect 35894 24284 35900 24296
rect 35952 24284 35958 24336
rect 7101 24259 7159 24265
rect 7101 24225 7113 24259
rect 7147 24225 7159 24259
rect 7101 24219 7159 24225
rect 7190 24216 7196 24268
rect 7248 24256 7254 24268
rect 7357 24259 7415 24265
rect 7357 24256 7369 24259
rect 7248 24228 7369 24256
rect 7248 24216 7254 24228
rect 7357 24225 7369 24228
rect 7403 24225 7415 24259
rect 7357 24219 7415 24225
rect 7742 24216 7748 24268
rect 7800 24256 7806 24268
rect 9493 24259 9551 24265
rect 9493 24256 9505 24259
rect 7800 24228 9505 24256
rect 7800 24216 7806 24228
rect 9493 24225 9505 24228
rect 9539 24256 9551 24259
rect 9769 24259 9827 24265
rect 9769 24256 9781 24259
rect 9539 24228 9781 24256
rect 9539 24225 9551 24228
rect 9493 24219 9551 24225
rect 9769 24225 9781 24228
rect 9815 24256 9827 24259
rect 9858 24256 9864 24268
rect 9815 24228 9864 24256
rect 9815 24225 9827 24228
rect 9769 24219 9827 24225
rect 9858 24216 9864 24228
rect 9916 24256 9922 24268
rect 10410 24256 10416 24268
rect 9916 24228 10416 24256
rect 9916 24216 9922 24228
rect 10410 24216 10416 24228
rect 10468 24216 10474 24268
rect 12452 24120 12480 24284
rect 15841 24259 15899 24265
rect 15841 24225 15853 24259
rect 15887 24256 15899 24259
rect 16666 24256 16672 24268
rect 15887 24228 16672 24256
rect 15887 24225 15899 24228
rect 15841 24219 15899 24225
rect 16666 24216 16672 24228
rect 16724 24216 16730 24268
rect 17037 24259 17095 24265
rect 17037 24225 17049 24259
rect 17083 24256 17095 24259
rect 17126 24256 17132 24268
rect 17083 24228 17132 24256
rect 17083 24225 17095 24228
rect 17037 24219 17095 24225
rect 17126 24216 17132 24228
rect 17184 24256 17190 24268
rect 17862 24256 17868 24268
rect 17184 24228 17868 24256
rect 17184 24216 17190 24228
rect 17862 24216 17868 24228
rect 17920 24216 17926 24268
rect 18506 24216 18512 24268
rect 18564 24256 18570 24268
rect 18966 24256 18972 24268
rect 18564 24228 18972 24256
rect 18564 24216 18570 24228
rect 18966 24216 18972 24228
rect 19024 24216 19030 24268
rect 20898 24216 20904 24268
rect 20956 24256 20962 24268
rect 22005 24259 22063 24265
rect 22005 24256 22017 24259
rect 20956 24228 22017 24256
rect 20956 24216 20962 24228
rect 22005 24225 22017 24228
rect 22051 24256 22063 24259
rect 22370 24256 22376 24268
rect 22051 24228 22376 24256
rect 22051 24225 22063 24228
rect 22005 24219 22063 24225
rect 22370 24216 22376 24228
rect 22428 24216 22434 24268
rect 29086 24216 29092 24268
rect 29144 24256 29150 24268
rect 29816 24259 29874 24265
rect 29816 24256 29828 24259
rect 29144 24228 29828 24256
rect 29144 24216 29150 24228
rect 29816 24225 29828 24228
rect 29862 24256 29874 24259
rect 31110 24256 31116 24268
rect 29862 24228 31116 24256
rect 29862 24225 29874 24228
rect 29816 24219 29874 24225
rect 31110 24216 31116 24228
rect 31168 24216 31174 24268
rect 32122 24216 32128 24268
rect 32180 24256 32186 24268
rect 32493 24259 32551 24265
rect 32493 24256 32505 24259
rect 32180 24228 32505 24256
rect 32180 24216 32186 24228
rect 32493 24225 32505 24228
rect 32539 24225 32551 24259
rect 32493 24219 32551 24225
rect 34606 24216 34612 24268
rect 34664 24256 34670 24268
rect 34885 24259 34943 24265
rect 34885 24256 34897 24259
rect 34664 24228 34897 24256
rect 34664 24216 34670 24228
rect 34885 24225 34897 24228
rect 34931 24225 34943 24259
rect 34885 24219 34943 24225
rect 36081 24259 36139 24265
rect 36081 24225 36093 24259
rect 36127 24256 36139 24259
rect 36906 24256 36912 24268
rect 36127 24228 36912 24256
rect 36127 24225 36139 24228
rect 36081 24219 36139 24225
rect 36906 24216 36912 24228
rect 36964 24216 36970 24268
rect 16117 24191 16175 24197
rect 16117 24157 16129 24191
rect 16163 24188 16175 24191
rect 16298 24188 16304 24200
rect 16163 24160 16304 24188
rect 16163 24157 16175 24160
rect 16117 24151 16175 24157
rect 16298 24148 16304 24160
rect 16356 24148 16362 24200
rect 18782 24148 18788 24200
rect 18840 24188 18846 24200
rect 19061 24191 19119 24197
rect 19061 24188 19073 24191
rect 18840 24160 19073 24188
rect 18840 24148 18846 24160
rect 19061 24157 19073 24160
rect 19107 24157 19119 24191
rect 19061 24151 19119 24157
rect 19153 24191 19211 24197
rect 19153 24157 19165 24191
rect 19199 24157 19211 24191
rect 19153 24151 19211 24157
rect 12529 24123 12587 24129
rect 12529 24120 12541 24123
rect 12452 24092 12541 24120
rect 12529 24089 12541 24092
rect 12575 24120 12587 24123
rect 12986 24120 12992 24132
rect 12575 24092 12992 24120
rect 12575 24089 12587 24092
rect 12529 24083 12587 24089
rect 12986 24080 12992 24092
rect 13044 24080 13050 24132
rect 18049 24123 18107 24129
rect 18049 24089 18061 24123
rect 18095 24120 18107 24123
rect 18230 24120 18236 24132
rect 18095 24092 18236 24120
rect 18095 24089 18107 24092
rect 18049 24083 18107 24089
rect 18230 24080 18236 24092
rect 18288 24120 18294 24132
rect 19168 24120 19196 24151
rect 21082 24148 21088 24200
rect 21140 24188 21146 24200
rect 21361 24191 21419 24197
rect 21361 24188 21373 24191
rect 21140 24160 21373 24188
rect 21140 24148 21146 24160
rect 21361 24157 21373 24160
rect 21407 24157 21419 24191
rect 21361 24151 21419 24157
rect 21453 24191 21511 24197
rect 21453 24157 21465 24191
rect 21499 24157 21511 24191
rect 21453 24151 21511 24157
rect 29549 24191 29607 24197
rect 29549 24157 29561 24191
rect 29595 24157 29607 24191
rect 32582 24188 32588 24200
rect 32543 24160 32588 24188
rect 29549 24151 29607 24157
rect 18288 24092 19196 24120
rect 18288 24080 18294 24092
rect 19334 24080 19340 24132
rect 19392 24120 19398 24132
rect 19981 24123 20039 24129
rect 19981 24120 19993 24123
rect 19392 24092 19993 24120
rect 19392 24080 19398 24092
rect 19981 24089 19993 24092
rect 20027 24089 20039 24123
rect 19981 24083 20039 24089
rect 20254 24080 20260 24132
rect 20312 24120 20318 24132
rect 21468 24120 21496 24151
rect 20312 24092 21496 24120
rect 20312 24080 20318 24092
rect 11146 24052 11152 24064
rect 11107 24024 11152 24052
rect 11146 24012 11152 24024
rect 11204 24012 11210 24064
rect 17218 24052 17224 24064
rect 17179 24024 17224 24052
rect 17218 24012 17224 24024
rect 17276 24012 17282 24064
rect 18414 24052 18420 24064
rect 18375 24024 18420 24052
rect 18414 24012 18420 24024
rect 18472 24012 18478 24064
rect 18598 24052 18604 24064
rect 18559 24024 18604 24052
rect 18598 24012 18604 24024
rect 18656 24012 18662 24064
rect 19518 24012 19524 24064
rect 19576 24052 19582 24064
rect 19613 24055 19671 24061
rect 19613 24052 19625 24055
rect 19576 24024 19625 24052
rect 19576 24012 19582 24024
rect 19613 24021 19625 24024
rect 19659 24021 19671 24055
rect 19613 24015 19671 24021
rect 19794 24012 19800 24064
rect 19852 24052 19858 24064
rect 20349 24055 20407 24061
rect 20349 24052 20361 24055
rect 19852 24024 20361 24052
rect 19852 24012 19858 24024
rect 20349 24021 20361 24024
rect 20395 24021 20407 24055
rect 20349 24015 20407 24021
rect 29457 24055 29515 24061
rect 29457 24021 29469 24055
rect 29503 24052 29515 24055
rect 29564 24052 29592 24151
rect 32582 24148 32588 24160
rect 32640 24148 32646 24200
rect 32674 24148 32680 24200
rect 32732 24188 32738 24200
rect 32732 24160 32777 24188
rect 32732 24148 32738 24160
rect 34422 24148 34428 24200
rect 34480 24188 34486 24200
rect 34977 24191 35035 24197
rect 34977 24188 34989 24191
rect 34480 24160 34989 24188
rect 34480 24148 34486 24160
rect 34977 24157 34989 24160
rect 35023 24157 35035 24191
rect 35158 24188 35164 24200
rect 35119 24160 35164 24188
rect 34977 24151 35035 24157
rect 35158 24148 35164 24160
rect 35216 24148 35222 24200
rect 31573 24123 31631 24129
rect 31573 24089 31585 24123
rect 31619 24120 31631 24123
rect 32692 24120 32720 24148
rect 31619 24092 32720 24120
rect 31619 24089 31631 24092
rect 31573 24083 31631 24089
rect 33318 24080 33324 24132
rect 33376 24120 33382 24132
rect 35529 24123 35587 24129
rect 35529 24120 35541 24123
rect 33376 24092 35541 24120
rect 33376 24080 33382 24092
rect 35529 24089 35541 24092
rect 35575 24120 35587 24123
rect 35710 24120 35716 24132
rect 35575 24092 35716 24120
rect 35575 24089 35587 24092
rect 35529 24083 35587 24089
rect 35710 24080 35716 24092
rect 35768 24080 35774 24132
rect 29730 24052 29736 24064
rect 29503 24024 29736 24052
rect 29503 24021 29515 24024
rect 29457 24015 29515 24021
rect 29730 24012 29736 24024
rect 29788 24012 29794 24064
rect 34514 24052 34520 24064
rect 34475 24024 34520 24052
rect 34514 24012 34520 24024
rect 34572 24012 34578 24064
rect 1104 23962 38824 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 34966 23962
rect 35018 23910 35030 23962
rect 35082 23910 35094 23962
rect 35146 23910 35158 23962
rect 35210 23910 38824 23962
rect 1104 23888 38824 23910
rect 7190 23848 7196 23860
rect 7151 23820 7196 23848
rect 7190 23808 7196 23820
rect 7248 23808 7254 23860
rect 9030 23848 9036 23860
rect 8991 23820 9036 23848
rect 9030 23808 9036 23820
rect 9088 23808 9094 23860
rect 9674 23808 9680 23860
rect 9732 23848 9738 23860
rect 10137 23851 10195 23857
rect 10137 23848 10149 23851
rect 9732 23820 10149 23848
rect 9732 23808 9738 23820
rect 10137 23817 10149 23820
rect 10183 23817 10195 23851
rect 10137 23811 10195 23817
rect 14461 23851 14519 23857
rect 14461 23817 14473 23851
rect 14507 23848 14519 23851
rect 16577 23851 16635 23857
rect 16577 23848 16589 23851
rect 14507 23820 16589 23848
rect 14507 23817 14519 23820
rect 14461 23811 14519 23817
rect 7561 23715 7619 23721
rect 7561 23681 7573 23715
rect 7607 23712 7619 23715
rect 9861 23715 9919 23721
rect 7607 23684 7788 23712
rect 7607 23681 7619 23684
rect 7561 23675 7619 23681
rect 7653 23647 7711 23653
rect 7653 23613 7665 23647
rect 7699 23613 7711 23647
rect 7760 23644 7788 23684
rect 9861 23681 9873 23715
rect 9907 23712 9919 23715
rect 10226 23712 10232 23724
rect 9907 23684 10232 23712
rect 9907 23681 9919 23684
rect 9861 23675 9919 23681
rect 10226 23672 10232 23684
rect 10284 23712 10290 23724
rect 10594 23712 10600 23724
rect 10284 23684 10600 23712
rect 10284 23672 10290 23684
rect 10594 23672 10600 23684
rect 10652 23672 10658 23724
rect 10686 23672 10692 23724
rect 10744 23712 10750 23724
rect 14568 23712 14596 23820
rect 16577 23817 16589 23820
rect 16623 23848 16635 23851
rect 16666 23848 16672 23860
rect 16623 23820 16672 23848
rect 16623 23817 16635 23820
rect 16577 23811 16635 23817
rect 16666 23808 16672 23820
rect 16724 23808 16730 23860
rect 17126 23848 17132 23860
rect 17087 23820 17132 23848
rect 17126 23808 17132 23820
rect 17184 23808 17190 23860
rect 19058 23848 19064 23860
rect 19019 23820 19064 23848
rect 19058 23808 19064 23820
rect 19116 23808 19122 23860
rect 20254 23848 20260 23860
rect 20215 23820 20260 23848
rect 20254 23808 20260 23820
rect 20312 23808 20318 23860
rect 20714 23848 20720 23860
rect 20675 23820 20720 23848
rect 20714 23808 20720 23820
rect 20772 23808 20778 23860
rect 22002 23808 22008 23860
rect 22060 23848 22066 23860
rect 22097 23851 22155 23857
rect 22097 23848 22109 23851
rect 22060 23820 22109 23848
rect 22060 23808 22066 23820
rect 22097 23817 22109 23820
rect 22143 23817 22155 23851
rect 29086 23848 29092 23860
rect 29047 23820 29092 23848
rect 22097 23811 22155 23817
rect 29086 23808 29092 23820
rect 29144 23808 29150 23860
rect 31110 23848 31116 23860
rect 31071 23820 31116 23848
rect 31110 23808 31116 23820
rect 31168 23808 31174 23860
rect 32122 23848 32128 23860
rect 32083 23820 32128 23848
rect 32122 23808 32128 23820
rect 32180 23808 32186 23860
rect 32401 23851 32459 23857
rect 32401 23817 32413 23851
rect 32447 23848 32459 23851
rect 33042 23848 33048 23860
rect 32447 23820 33048 23848
rect 32447 23817 32459 23820
rect 32401 23811 32459 23817
rect 33042 23808 33048 23820
rect 33100 23808 33106 23860
rect 34238 23808 34244 23860
rect 34296 23848 34302 23860
rect 34606 23848 34612 23860
rect 34296 23820 34612 23848
rect 34296 23808 34302 23820
rect 34606 23808 34612 23820
rect 34664 23808 34670 23860
rect 36906 23848 36912 23860
rect 36867 23820 36912 23848
rect 36906 23808 36912 23820
rect 36964 23808 36970 23860
rect 19076 23712 19104 23808
rect 32674 23740 32680 23792
rect 32732 23780 32738 23792
rect 33137 23783 33195 23789
rect 33137 23780 33149 23783
rect 32732 23752 33149 23780
rect 32732 23740 32738 23752
rect 33137 23749 33149 23752
rect 33183 23749 33195 23783
rect 33137 23743 33195 23749
rect 33597 23783 33655 23789
rect 33597 23749 33609 23783
rect 33643 23780 33655 23783
rect 34330 23780 34336 23792
rect 33643 23752 34336 23780
rect 33643 23749 33655 23752
rect 33597 23743 33655 23749
rect 10744 23684 10789 23712
rect 14568 23684 14688 23712
rect 10744 23672 10750 23684
rect 7920 23647 7978 23653
rect 7920 23644 7932 23647
rect 7760 23616 7932 23644
rect 7653 23607 7711 23613
rect 7920 23613 7932 23616
rect 7966 23644 7978 23647
rect 8478 23644 8484 23656
rect 7966 23616 8484 23644
rect 7966 23613 7978 23616
rect 7920 23607 7978 23613
rect 7668 23576 7696 23607
rect 8478 23604 8484 23616
rect 8536 23604 8542 23656
rect 10502 23644 10508 23656
rect 10463 23616 10508 23644
rect 10502 23604 10508 23616
rect 10560 23644 10566 23656
rect 11146 23644 11152 23656
rect 10560 23616 11152 23644
rect 10560 23604 10566 23616
rect 11146 23604 11152 23616
rect 11204 23604 11210 23656
rect 12986 23604 12992 23656
rect 13044 23644 13050 23656
rect 14550 23644 14556 23656
rect 13044 23616 14556 23644
rect 13044 23604 13050 23616
rect 14550 23604 14556 23616
rect 14608 23604 14614 23656
rect 14660 23644 14688 23684
rect 18340 23684 19104 23712
rect 18340 23653 18368 23684
rect 19426 23672 19432 23724
rect 19484 23712 19490 23724
rect 19794 23712 19800 23724
rect 19484 23684 19800 23712
rect 19484 23672 19490 23684
rect 19794 23672 19800 23684
rect 19852 23672 19858 23724
rect 14809 23647 14867 23653
rect 14809 23644 14821 23647
rect 14660 23616 14821 23644
rect 14809 23613 14821 23616
rect 14855 23613 14867 23647
rect 14809 23607 14867 23613
rect 18325 23647 18383 23653
rect 18325 23613 18337 23647
rect 18371 23613 18383 23647
rect 18325 23607 18383 23613
rect 18414 23604 18420 23656
rect 18472 23644 18478 23656
rect 18509 23647 18567 23653
rect 18509 23644 18521 23647
rect 18472 23616 18521 23644
rect 18472 23604 18478 23616
rect 18509 23613 18521 23616
rect 18555 23613 18567 23647
rect 18509 23607 18567 23613
rect 19058 23604 19064 23656
rect 19116 23644 19122 23656
rect 19518 23644 19524 23656
rect 19116 23616 19524 23644
rect 19116 23604 19122 23616
rect 19518 23604 19524 23616
rect 19576 23604 19582 23656
rect 29730 23644 29736 23656
rect 29691 23616 29736 23644
rect 29730 23604 29736 23616
rect 29788 23604 29794 23656
rect 31757 23647 31815 23653
rect 31757 23613 31769 23647
rect 31803 23644 31815 23647
rect 32217 23647 32275 23653
rect 32217 23644 32229 23647
rect 31803 23616 32229 23644
rect 31803 23613 31815 23616
rect 31757 23607 31815 23613
rect 32217 23613 32229 23616
rect 32263 23644 32275 23647
rect 32306 23644 32312 23656
rect 32263 23616 32312 23644
rect 32263 23613 32275 23616
rect 32217 23607 32275 23613
rect 32306 23604 32312 23616
rect 32364 23604 32370 23656
rect 33704 23653 33732 23752
rect 34330 23740 34336 23752
rect 34388 23740 34394 23792
rect 33689 23647 33747 23653
rect 33689 23613 33701 23647
rect 33735 23613 33747 23647
rect 33689 23607 33747 23613
rect 34885 23647 34943 23653
rect 34885 23613 34897 23647
rect 34931 23644 34943 23647
rect 36538 23644 36544 23656
rect 34931 23616 36544 23644
rect 34931 23613 34943 23616
rect 34885 23607 34943 23613
rect 36538 23604 36544 23616
rect 36596 23604 36602 23656
rect 7742 23576 7748 23588
rect 7668 23548 7748 23576
rect 7742 23536 7748 23548
rect 7800 23536 7806 23588
rect 20809 23579 20867 23585
rect 20809 23545 20821 23579
rect 20855 23576 20867 23579
rect 21542 23576 21548 23588
rect 20855 23548 21548 23576
rect 20855 23545 20867 23548
rect 20809 23539 20867 23545
rect 21542 23536 21548 23548
rect 21600 23536 21606 23588
rect 29641 23579 29699 23585
rect 29641 23545 29653 23579
rect 29687 23576 29699 23579
rect 30000 23579 30058 23585
rect 30000 23576 30012 23579
rect 29687 23548 30012 23576
rect 29687 23545 29699 23548
rect 29641 23539 29699 23545
rect 30000 23545 30012 23548
rect 30046 23576 30058 23579
rect 30926 23576 30932 23588
rect 30046 23548 30932 23576
rect 30046 23545 30058 23548
rect 30000 23539 30058 23545
rect 30926 23536 30932 23548
rect 30984 23536 30990 23588
rect 32582 23576 32588 23588
rect 31772 23548 32588 23576
rect 31772 23520 31800 23548
rect 32582 23536 32588 23548
rect 32640 23576 32646 23588
rect 32769 23579 32827 23585
rect 32769 23576 32781 23579
rect 32640 23548 32781 23576
rect 32640 23536 32646 23548
rect 32769 23545 32781 23548
rect 32815 23545 32827 23579
rect 32769 23539 32827 23545
rect 34330 23536 34336 23588
rect 34388 23576 34394 23588
rect 35152 23579 35210 23585
rect 35152 23576 35164 23579
rect 34388 23548 35164 23576
rect 34388 23536 34394 23548
rect 35152 23545 35164 23548
rect 35198 23576 35210 23579
rect 35250 23576 35256 23588
rect 35198 23548 35256 23576
rect 35198 23545 35210 23548
rect 35152 23539 35210 23545
rect 35250 23536 35256 23548
rect 35308 23576 35314 23588
rect 35894 23576 35900 23588
rect 35308 23548 35900 23576
rect 35308 23536 35314 23548
rect 35894 23536 35900 23548
rect 35952 23536 35958 23588
rect 10410 23468 10416 23520
rect 10468 23508 10474 23520
rect 11609 23511 11667 23517
rect 11609 23508 11621 23511
rect 10468 23480 11621 23508
rect 10468 23468 10474 23480
rect 11609 23477 11621 23480
rect 11655 23508 11667 23511
rect 12342 23508 12348 23520
rect 11655 23480 12348 23508
rect 11655 23477 11667 23480
rect 11609 23471 11667 23477
rect 12342 23468 12348 23480
rect 12400 23468 12406 23520
rect 15194 23468 15200 23520
rect 15252 23508 15258 23520
rect 15933 23511 15991 23517
rect 15933 23508 15945 23511
rect 15252 23480 15945 23508
rect 15252 23468 15258 23480
rect 15933 23477 15945 23480
rect 15979 23477 15991 23511
rect 15933 23471 15991 23477
rect 16574 23468 16580 23520
rect 16632 23508 16638 23520
rect 17773 23511 17831 23517
rect 17773 23508 17785 23511
rect 16632 23480 17785 23508
rect 16632 23468 16638 23480
rect 17773 23477 17785 23480
rect 17819 23508 17831 23511
rect 18506 23508 18512 23520
rect 17819 23480 18512 23508
rect 17819 23477 17831 23480
rect 17773 23471 17831 23477
rect 18506 23468 18512 23480
rect 18564 23468 18570 23520
rect 18690 23508 18696 23520
rect 18651 23480 18696 23508
rect 18690 23468 18696 23480
rect 18748 23468 18754 23520
rect 19150 23508 19156 23520
rect 19111 23480 19156 23508
rect 19150 23468 19156 23480
rect 19208 23468 19214 23520
rect 19334 23468 19340 23520
rect 19392 23508 19398 23520
rect 19613 23511 19671 23517
rect 19613 23508 19625 23511
rect 19392 23480 19625 23508
rect 19392 23468 19398 23480
rect 19613 23477 19625 23480
rect 19659 23477 19671 23511
rect 28718 23508 28724 23520
rect 28679 23480 28724 23508
rect 19613 23471 19671 23477
rect 28718 23468 28724 23480
rect 28776 23468 28782 23520
rect 31754 23468 31760 23520
rect 31812 23468 31818 23520
rect 33873 23511 33931 23517
rect 33873 23477 33885 23511
rect 33919 23508 33931 23511
rect 34422 23508 34428 23520
rect 33919 23480 34428 23508
rect 33919 23477 33931 23480
rect 33873 23471 33931 23477
rect 34422 23468 34428 23480
rect 34480 23468 34486 23520
rect 36262 23508 36268 23520
rect 36223 23480 36268 23508
rect 36262 23468 36268 23480
rect 36320 23468 36326 23520
rect 1104 23418 38824 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 38824 23418
rect 1104 23344 38824 23366
rect 7193 23307 7251 23313
rect 7193 23273 7205 23307
rect 7239 23304 7251 23307
rect 7742 23304 7748 23316
rect 7239 23276 7748 23304
rect 7239 23273 7251 23276
rect 7193 23267 7251 23273
rect 7742 23264 7748 23276
rect 7800 23264 7806 23316
rect 10226 23304 10232 23316
rect 10187 23276 10232 23304
rect 10226 23264 10232 23276
rect 10284 23264 10290 23316
rect 10410 23304 10416 23316
rect 10371 23276 10416 23304
rect 10410 23264 10416 23276
rect 10468 23264 10474 23316
rect 10686 23264 10692 23316
rect 10744 23304 10750 23316
rect 10873 23307 10931 23313
rect 10873 23304 10885 23307
rect 10744 23276 10885 23304
rect 10744 23264 10750 23276
rect 10873 23273 10885 23276
rect 10919 23273 10931 23307
rect 14090 23304 14096 23316
rect 14003 23276 14096 23304
rect 10873 23267 10931 23273
rect 14090 23264 14096 23276
rect 14148 23304 14154 23316
rect 15102 23304 15108 23316
rect 14148 23276 15108 23304
rect 14148 23264 14154 23276
rect 15102 23264 15108 23276
rect 15160 23264 15166 23316
rect 15473 23307 15531 23313
rect 15473 23273 15485 23307
rect 15519 23304 15531 23307
rect 16390 23304 16396 23316
rect 15519 23276 16396 23304
rect 15519 23273 15531 23276
rect 15473 23267 15531 23273
rect 16390 23264 16396 23276
rect 16448 23304 16454 23316
rect 16761 23307 16819 23313
rect 16761 23304 16773 23307
rect 16448 23276 16773 23304
rect 16448 23264 16454 23276
rect 16761 23273 16773 23276
rect 16807 23273 16819 23307
rect 16761 23267 16819 23273
rect 16853 23307 16911 23313
rect 16853 23273 16865 23307
rect 16899 23304 16911 23307
rect 17218 23304 17224 23316
rect 16899 23276 17224 23304
rect 16899 23273 16911 23276
rect 16853 23267 16911 23273
rect 17218 23264 17224 23276
rect 17276 23264 17282 23316
rect 18230 23304 18236 23316
rect 18191 23276 18236 23304
rect 18230 23264 18236 23276
rect 18288 23264 18294 23316
rect 18693 23307 18751 23313
rect 18693 23273 18705 23307
rect 18739 23304 18751 23307
rect 18782 23304 18788 23316
rect 18739 23276 18788 23304
rect 18739 23273 18751 23276
rect 18693 23267 18751 23273
rect 18782 23264 18788 23276
rect 18840 23264 18846 23316
rect 20254 23264 20260 23316
rect 20312 23304 20318 23316
rect 20441 23307 20499 23313
rect 20441 23304 20453 23307
rect 20312 23276 20453 23304
rect 20312 23264 20318 23276
rect 20441 23273 20453 23276
rect 20487 23273 20499 23307
rect 21082 23304 21088 23316
rect 21043 23276 21088 23304
rect 20441 23267 20499 23273
rect 21082 23264 21088 23276
rect 21140 23264 21146 23316
rect 25130 23304 25136 23316
rect 25091 23276 25136 23304
rect 25130 23264 25136 23276
rect 25188 23264 25194 23316
rect 30926 23304 30932 23316
rect 30839 23276 30932 23304
rect 30926 23264 30932 23276
rect 30984 23304 30990 23316
rect 32122 23304 32128 23316
rect 30984 23276 32128 23304
rect 30984 23264 30990 23276
rect 32122 23264 32128 23276
rect 32180 23264 32186 23316
rect 32309 23307 32367 23313
rect 32309 23273 32321 23307
rect 32355 23304 32367 23307
rect 32858 23304 32864 23316
rect 32355 23276 32864 23304
rect 32355 23273 32367 23276
rect 32309 23267 32367 23273
rect 32858 23264 32864 23276
rect 32916 23264 32922 23316
rect 33597 23307 33655 23313
rect 33597 23273 33609 23307
rect 33643 23304 33655 23307
rect 34238 23304 34244 23316
rect 33643 23276 34244 23304
rect 33643 23273 33655 23276
rect 33597 23267 33655 23273
rect 34238 23264 34244 23276
rect 34296 23264 34302 23316
rect 34422 23304 34428 23316
rect 34383 23276 34428 23304
rect 34422 23264 34428 23276
rect 34480 23264 34486 23316
rect 34514 23264 34520 23316
rect 34572 23304 34578 23316
rect 34977 23307 35035 23313
rect 34977 23304 34989 23307
rect 34572 23276 34989 23304
rect 34572 23264 34578 23276
rect 34977 23273 34989 23276
rect 35023 23273 35035 23307
rect 35894 23304 35900 23316
rect 35855 23276 35900 23304
rect 34977 23267 35035 23273
rect 35894 23264 35900 23276
rect 35952 23264 35958 23316
rect 15930 23236 15936 23248
rect 15891 23208 15936 23236
rect 15930 23196 15936 23208
rect 15988 23196 15994 23248
rect 16298 23236 16304 23248
rect 16259 23208 16304 23236
rect 16298 23196 16304 23208
rect 16356 23196 16362 23248
rect 19328 23239 19386 23245
rect 19328 23205 19340 23239
rect 19374 23236 19386 23239
rect 19426 23236 19432 23248
rect 19374 23208 19432 23236
rect 19374 23205 19386 23208
rect 19328 23199 19386 23205
rect 19426 23196 19432 23208
rect 19484 23196 19490 23248
rect 26513 23239 26571 23245
rect 26513 23205 26525 23239
rect 26559 23236 26571 23239
rect 27154 23236 27160 23248
rect 26559 23208 27160 23236
rect 26559 23205 26571 23208
rect 26513 23199 26571 23205
rect 27154 23196 27160 23208
rect 27212 23196 27218 23248
rect 29730 23236 29736 23248
rect 29564 23208 29736 23236
rect 10594 23168 10600 23180
rect 10555 23140 10600 23168
rect 10594 23128 10600 23140
rect 10652 23128 10658 23180
rect 13998 23168 14004 23180
rect 13959 23140 14004 23168
rect 13998 23128 14004 23140
rect 14056 23128 14062 23180
rect 15286 23168 15292 23180
rect 15247 23140 15292 23168
rect 15286 23128 15292 23140
rect 15344 23128 15350 23180
rect 13538 23100 13544 23112
rect 13451 23072 13544 23100
rect 13538 23060 13544 23072
rect 13596 23100 13602 23112
rect 14277 23103 14335 23109
rect 14277 23100 14289 23103
rect 13596 23072 14289 23100
rect 13596 23060 13602 23072
rect 14277 23069 14289 23072
rect 14323 23100 14335 23103
rect 16316 23100 16344 23196
rect 18049 23171 18107 23177
rect 18049 23137 18061 23171
rect 18095 23168 18107 23171
rect 18138 23168 18144 23180
rect 18095 23140 18144 23168
rect 18095 23137 18107 23140
rect 18049 23131 18107 23137
rect 18138 23128 18144 23140
rect 18196 23168 18202 23180
rect 18690 23168 18696 23180
rect 18196 23140 18696 23168
rect 18196 23128 18202 23140
rect 18690 23128 18696 23140
rect 18748 23128 18754 23180
rect 19061 23171 19119 23177
rect 19061 23137 19073 23171
rect 19107 23168 19119 23171
rect 19150 23168 19156 23180
rect 19107 23140 19156 23168
rect 19107 23137 19119 23140
rect 19061 23131 19119 23137
rect 19150 23128 19156 23140
rect 19208 23168 19214 23180
rect 19886 23168 19892 23180
rect 19208 23140 19892 23168
rect 19208 23128 19214 23140
rect 19886 23128 19892 23140
rect 19944 23128 19950 23180
rect 26697 23171 26755 23177
rect 26697 23137 26709 23171
rect 26743 23168 26755 23171
rect 26786 23168 26792 23180
rect 26743 23140 26792 23168
rect 26743 23137 26755 23140
rect 26697 23131 26755 23137
rect 26786 23128 26792 23140
rect 26844 23128 26850 23180
rect 29564 23177 29592 23208
rect 29730 23196 29736 23208
rect 29788 23196 29794 23248
rect 34057 23239 34115 23245
rect 34057 23205 34069 23239
rect 34103 23236 34115 23239
rect 34330 23236 34336 23248
rect 34103 23208 34336 23236
rect 34103 23205 34115 23208
rect 34057 23199 34115 23205
rect 34330 23196 34336 23208
rect 34388 23196 34394 23248
rect 29457 23171 29515 23177
rect 29457 23137 29469 23171
rect 29503 23168 29515 23171
rect 29549 23171 29607 23177
rect 29549 23168 29561 23171
rect 29503 23140 29561 23168
rect 29503 23137 29515 23140
rect 29457 23131 29515 23137
rect 29549 23137 29561 23140
rect 29595 23137 29607 23171
rect 29549 23131 29607 23137
rect 29638 23128 29644 23180
rect 29696 23168 29702 23180
rect 29816 23171 29874 23177
rect 29816 23168 29828 23171
rect 29696 23140 29828 23168
rect 29696 23128 29702 23140
rect 29816 23137 29828 23140
rect 29862 23168 29874 23171
rect 31018 23168 31024 23180
rect 29862 23140 31024 23168
rect 29862 23137 29874 23140
rect 29816 23131 29874 23137
rect 31018 23128 31024 23140
rect 31076 23128 31082 23180
rect 32125 23171 32183 23177
rect 32125 23137 32137 23171
rect 32171 23168 32183 23171
rect 32214 23168 32220 23180
rect 32171 23140 32220 23168
rect 32171 23137 32183 23140
rect 32125 23131 32183 23137
rect 32214 23128 32220 23140
rect 32272 23128 32278 23180
rect 33318 23128 33324 23180
rect 33376 23168 33382 23180
rect 33413 23171 33471 23177
rect 33413 23168 33425 23171
rect 33376 23140 33425 23168
rect 33376 23128 33382 23140
rect 33413 23137 33425 23140
rect 33459 23137 33471 23171
rect 33413 23131 33471 23137
rect 34698 23128 34704 23180
rect 34756 23168 34762 23180
rect 34885 23171 34943 23177
rect 34885 23168 34897 23171
rect 34756 23140 34897 23168
rect 34756 23128 34762 23140
rect 34885 23137 34897 23140
rect 34931 23168 34943 23171
rect 36081 23171 36139 23177
rect 36081 23168 36093 23171
rect 34931 23140 36093 23168
rect 34931 23137 34943 23140
rect 34885 23131 34943 23137
rect 36081 23137 36093 23140
rect 36127 23137 36139 23171
rect 36081 23131 36139 23137
rect 17034 23100 17040 23112
rect 14323 23072 16344 23100
rect 16947 23072 17040 23100
rect 14323 23069 14335 23072
rect 14277 23063 14335 23069
rect 17034 23060 17040 23072
rect 17092 23100 17098 23112
rect 17402 23100 17408 23112
rect 17092 23072 17408 23100
rect 17092 23060 17098 23072
rect 17402 23060 17408 23072
rect 17460 23060 17466 23112
rect 35161 23103 35219 23109
rect 35161 23069 35173 23103
rect 35207 23100 35219 23103
rect 35250 23100 35256 23112
rect 35207 23072 35256 23100
rect 35207 23069 35219 23072
rect 35161 23063 35219 23069
rect 35250 23060 35256 23072
rect 35308 23100 35314 23112
rect 36262 23100 36268 23112
rect 35308 23072 36268 23100
rect 35308 23060 35314 23072
rect 36262 23060 36268 23072
rect 36320 23060 36326 23112
rect 16393 23035 16451 23041
rect 16393 23001 16405 23035
rect 16439 23032 16451 23035
rect 18782 23032 18788 23044
rect 16439 23004 18788 23032
rect 16439 23001 16451 23004
rect 16393 22995 16451 23001
rect 18782 22992 18788 23004
rect 18840 22992 18846 23044
rect 13630 22964 13636 22976
rect 13591 22936 13636 22964
rect 13630 22924 13636 22936
rect 13688 22924 13694 22976
rect 21542 22964 21548 22976
rect 21503 22936 21548 22964
rect 21542 22924 21548 22936
rect 21600 22924 21606 22976
rect 26142 22924 26148 22976
rect 26200 22964 26206 22976
rect 26881 22967 26939 22973
rect 26881 22964 26893 22967
rect 26200 22936 26893 22964
rect 26200 22924 26206 22936
rect 26881 22933 26893 22936
rect 26927 22933 26939 22967
rect 34514 22964 34520 22976
rect 34475 22936 34520 22964
rect 26881 22927 26939 22933
rect 34514 22924 34520 22936
rect 34572 22924 34578 22976
rect 35526 22964 35532 22976
rect 35487 22936 35532 22964
rect 35526 22924 35532 22936
rect 35584 22924 35590 22976
rect 36538 22964 36544 22976
rect 36499 22936 36544 22964
rect 36538 22924 36544 22936
rect 36596 22924 36602 22976
rect 1104 22874 38824 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 34966 22874
rect 35018 22822 35030 22874
rect 35082 22822 35094 22874
rect 35146 22822 35158 22874
rect 35210 22822 38824 22874
rect 1104 22800 38824 22822
rect 6914 22720 6920 22772
rect 6972 22760 6978 22772
rect 7561 22763 7619 22769
rect 7561 22760 7573 22763
rect 6972 22732 7573 22760
rect 6972 22720 6978 22732
rect 7561 22729 7573 22732
rect 7607 22729 7619 22763
rect 7561 22723 7619 22729
rect 8113 22763 8171 22769
rect 8113 22729 8125 22763
rect 8159 22760 8171 22763
rect 8570 22760 8576 22772
rect 8159 22732 8576 22760
rect 8159 22729 8171 22732
rect 8113 22723 8171 22729
rect 7745 22559 7803 22565
rect 7745 22525 7757 22559
rect 7791 22556 7803 22559
rect 8128 22556 8156 22723
rect 8570 22720 8576 22732
rect 8628 22760 8634 22772
rect 10505 22763 10563 22769
rect 10505 22760 10517 22763
rect 8628 22732 10517 22760
rect 8628 22720 8634 22732
rect 10505 22729 10517 22732
rect 10551 22760 10563 22763
rect 10594 22760 10600 22772
rect 10551 22732 10600 22760
rect 10551 22729 10563 22732
rect 10505 22723 10563 22729
rect 10594 22720 10600 22732
rect 10652 22720 10658 22772
rect 12989 22763 13047 22769
rect 12989 22729 13001 22763
rect 13035 22760 13047 22763
rect 13170 22760 13176 22772
rect 13035 22732 13176 22760
rect 13035 22729 13047 22732
rect 12989 22723 13047 22729
rect 13170 22720 13176 22732
rect 13228 22760 13234 22772
rect 13998 22760 14004 22772
rect 13228 22732 14004 22760
rect 13228 22720 13234 22732
rect 13998 22720 14004 22732
rect 14056 22760 14062 22772
rect 15197 22763 15255 22769
rect 15197 22760 15209 22763
rect 14056 22732 15209 22760
rect 14056 22720 14062 22732
rect 15197 22729 15209 22732
rect 15243 22729 15255 22763
rect 15197 22723 15255 22729
rect 16301 22763 16359 22769
rect 16301 22729 16313 22763
rect 16347 22760 16359 22763
rect 17218 22760 17224 22772
rect 16347 22732 17224 22760
rect 16347 22729 16359 22732
rect 16301 22723 16359 22729
rect 17218 22720 17224 22732
rect 17276 22720 17282 22772
rect 18233 22763 18291 22769
rect 18233 22729 18245 22763
rect 18279 22760 18291 22763
rect 19058 22760 19064 22772
rect 18279 22732 19064 22760
rect 18279 22729 18291 22732
rect 18233 22723 18291 22729
rect 19058 22720 19064 22732
rect 19116 22720 19122 22772
rect 19426 22720 19432 22772
rect 19484 22760 19490 22772
rect 20533 22763 20591 22769
rect 20533 22760 20545 22763
rect 19484 22732 20545 22760
rect 19484 22720 19490 22732
rect 20533 22729 20545 22732
rect 20579 22729 20591 22763
rect 27154 22760 27160 22772
rect 27115 22732 27160 22760
rect 20533 22723 20591 22729
rect 27154 22720 27160 22732
rect 27212 22720 27218 22772
rect 31018 22760 31024 22772
rect 30931 22732 31024 22760
rect 31018 22720 31024 22732
rect 31076 22760 31082 22772
rect 31662 22760 31668 22772
rect 31076 22732 31668 22760
rect 31076 22720 31082 22732
rect 31662 22720 31668 22732
rect 31720 22720 31726 22772
rect 32214 22720 32220 22772
rect 32272 22760 32278 22772
rect 32585 22763 32643 22769
rect 32585 22760 32597 22763
rect 32272 22732 32597 22760
rect 32272 22720 32278 22732
rect 32585 22729 32597 22732
rect 32631 22729 32643 22763
rect 32950 22760 32956 22772
rect 32911 22732 32956 22760
rect 32585 22723 32643 22729
rect 32950 22720 32956 22732
rect 33008 22720 33014 22772
rect 33318 22720 33324 22772
rect 33376 22760 33382 22772
rect 33413 22763 33471 22769
rect 33413 22760 33425 22763
rect 33376 22732 33425 22760
rect 33376 22720 33382 22732
rect 33413 22729 33425 22732
rect 33459 22729 33471 22763
rect 33413 22723 33471 22729
rect 34609 22763 34667 22769
rect 34609 22729 34621 22763
rect 34655 22760 34667 22763
rect 34698 22760 34704 22772
rect 34655 22732 34704 22760
rect 34655 22729 34667 22732
rect 34609 22723 34667 22729
rect 34698 22720 34704 22732
rect 34756 22720 34762 22772
rect 35069 22763 35127 22769
rect 35069 22729 35081 22763
rect 35115 22760 35127 22763
rect 35434 22760 35440 22772
rect 35115 22732 35440 22760
rect 35115 22729 35127 22732
rect 35069 22723 35127 22729
rect 35434 22720 35440 22732
rect 35492 22720 35498 22772
rect 36173 22763 36231 22769
rect 36173 22729 36185 22763
rect 36219 22760 36231 22763
rect 36262 22760 36268 22772
rect 36219 22732 36268 22760
rect 36219 22729 36231 22732
rect 36173 22723 36231 22729
rect 36262 22720 36268 22732
rect 36320 22720 36326 22772
rect 16393 22695 16451 22701
rect 16393 22661 16405 22695
rect 16439 22692 16451 22695
rect 16482 22692 16488 22704
rect 16439 22664 16488 22692
rect 16439 22661 16451 22664
rect 16393 22655 16451 22661
rect 16482 22652 16488 22664
rect 16540 22652 16546 22704
rect 18414 22652 18420 22704
rect 18472 22692 18478 22704
rect 18969 22695 19027 22701
rect 18969 22692 18981 22695
rect 18472 22664 18981 22692
rect 18472 22652 18478 22664
rect 18969 22661 18981 22664
rect 19015 22661 19027 22695
rect 18969 22655 19027 22661
rect 26513 22695 26571 22701
rect 26513 22661 26525 22695
rect 26559 22692 26571 22695
rect 26786 22692 26792 22704
rect 26559 22664 26792 22692
rect 26559 22661 26571 22664
rect 26513 22655 26571 22661
rect 17034 22624 17040 22636
rect 16995 22596 17040 22624
rect 17034 22584 17040 22596
rect 17092 22624 17098 22636
rect 17402 22624 17408 22636
rect 17092 22596 17408 22624
rect 17092 22584 17098 22596
rect 17402 22584 17408 22596
rect 17460 22624 17466 22636
rect 17773 22627 17831 22633
rect 17773 22624 17785 22627
rect 17460 22596 17785 22624
rect 17460 22584 17466 22596
rect 17773 22593 17785 22596
rect 17819 22593 17831 22627
rect 17773 22587 17831 22593
rect 18693 22627 18751 22633
rect 18693 22593 18705 22627
rect 18739 22624 18751 22627
rect 18782 22624 18788 22636
rect 18739 22596 18788 22624
rect 18739 22593 18751 22596
rect 18693 22587 18751 22593
rect 7791 22528 8156 22556
rect 13817 22559 13875 22565
rect 7791 22525 7803 22528
rect 7745 22519 7803 22525
rect 13817 22525 13829 22559
rect 13863 22556 13875 22559
rect 13906 22556 13912 22568
rect 13863 22528 13912 22556
rect 13863 22525 13875 22528
rect 13817 22519 13875 22525
rect 13906 22516 13912 22528
rect 13964 22556 13970 22568
rect 14642 22556 14648 22568
rect 13964 22528 14648 22556
rect 13964 22516 13970 22528
rect 14642 22516 14648 22528
rect 14700 22516 14706 22568
rect 18074 22559 18132 22565
rect 18074 22525 18086 22559
rect 18120 22556 18132 22559
rect 18708 22556 18736 22587
rect 18782 22584 18788 22596
rect 18840 22584 18846 22636
rect 18984 22624 19012 22655
rect 26786 22652 26792 22664
rect 26844 22692 26850 22704
rect 27433 22695 27491 22701
rect 27433 22692 27445 22695
rect 26844 22664 27445 22692
rect 26844 22652 26850 22664
rect 27433 22661 27445 22664
rect 27479 22661 27491 22695
rect 27433 22655 27491 22661
rect 25130 22624 25136 22636
rect 18984 22596 19288 22624
rect 25091 22596 25136 22624
rect 19150 22556 19156 22568
rect 18120 22528 18736 22556
rect 19111 22528 19156 22556
rect 18120 22525 18132 22528
rect 18074 22519 18132 22525
rect 19150 22516 19156 22528
rect 19208 22516 19214 22568
rect 19260 22556 19288 22596
rect 25130 22584 25136 22596
rect 25188 22584 25194 22636
rect 35713 22627 35771 22633
rect 35713 22593 35725 22627
rect 35759 22624 35771 22627
rect 36078 22624 36084 22636
rect 35759 22596 36084 22624
rect 35759 22593 35771 22596
rect 35713 22587 35771 22593
rect 36078 22584 36084 22596
rect 36136 22624 36142 22636
rect 36449 22627 36507 22633
rect 36449 22624 36461 22627
rect 36136 22596 36461 22624
rect 36136 22584 36142 22596
rect 36449 22593 36461 22596
rect 36495 22593 36507 22627
rect 36449 22587 36507 22593
rect 19409 22559 19467 22565
rect 19409 22556 19421 22559
rect 19260 22528 19421 22556
rect 19409 22525 19421 22528
rect 19455 22556 19467 22559
rect 19978 22556 19984 22568
rect 19455 22528 19984 22556
rect 19455 22525 19467 22528
rect 19409 22519 19467 22525
rect 19978 22516 19984 22528
rect 20036 22516 20042 22568
rect 28718 22556 28724 22568
rect 28631 22528 28724 22556
rect 28718 22516 28724 22528
rect 28776 22556 28782 22568
rect 29089 22559 29147 22565
rect 29089 22556 29101 22559
rect 28776 22528 29101 22556
rect 28776 22516 28782 22528
rect 29089 22525 29101 22528
rect 29135 22556 29147 22559
rect 29641 22559 29699 22565
rect 29641 22556 29653 22559
rect 29135 22528 29653 22556
rect 29135 22525 29147 22528
rect 29089 22519 29147 22525
rect 29641 22525 29653 22528
rect 29687 22556 29699 22559
rect 29730 22556 29736 22568
rect 29687 22528 29736 22556
rect 29687 22525 29699 22528
rect 29641 22519 29699 22525
rect 29730 22516 29736 22528
rect 29788 22516 29794 22568
rect 32309 22559 32367 22565
rect 32309 22525 32321 22559
rect 32355 22556 32367 22559
rect 32950 22556 32956 22568
rect 32355 22528 32956 22556
rect 32355 22525 32367 22528
rect 32309 22519 32367 22525
rect 32950 22516 32956 22528
rect 33008 22516 33014 22568
rect 33689 22559 33747 22565
rect 33689 22525 33701 22559
rect 33735 22556 33747 22559
rect 33870 22556 33876 22568
rect 33735 22528 33876 22556
rect 33735 22525 33747 22528
rect 33689 22519 33747 22525
rect 33870 22516 33876 22528
rect 33928 22516 33934 22568
rect 35437 22559 35495 22565
rect 35437 22525 35449 22559
rect 35483 22556 35495 22559
rect 35526 22556 35532 22568
rect 35483 22528 35532 22556
rect 35483 22525 35495 22528
rect 35437 22519 35495 22525
rect 35526 22516 35532 22528
rect 35584 22556 35590 22568
rect 35894 22556 35900 22568
rect 35584 22528 35900 22556
rect 35584 22516 35590 22528
rect 35894 22516 35900 22528
rect 35952 22516 35958 22568
rect 14090 22497 14096 22500
rect 13357 22491 13415 22497
rect 13357 22457 13369 22491
rect 13403 22488 13415 22491
rect 13725 22491 13783 22497
rect 13725 22488 13737 22491
rect 13403 22460 13737 22488
rect 13403 22457 13415 22460
rect 13357 22451 13415 22457
rect 13725 22457 13737 22460
rect 13771 22488 13783 22491
rect 14084 22488 14096 22497
rect 13771 22460 14096 22488
rect 13771 22457 13783 22460
rect 13725 22451 13783 22457
rect 14084 22451 14096 22460
rect 14090 22448 14096 22451
rect 14148 22448 14154 22500
rect 15933 22491 15991 22497
rect 15933 22457 15945 22491
rect 15979 22488 15991 22491
rect 16761 22491 16819 22497
rect 15979 22460 16712 22488
rect 15979 22457 15991 22460
rect 15933 22451 15991 22457
rect 16684 22420 16712 22460
rect 16761 22457 16773 22491
rect 16807 22488 16819 22491
rect 17034 22488 17040 22500
rect 16807 22460 17040 22488
rect 16807 22457 16819 22460
rect 16761 22451 16819 22457
rect 17034 22448 17040 22460
rect 17092 22488 17098 22500
rect 17405 22491 17463 22497
rect 17405 22488 17417 22491
rect 17092 22460 17417 22488
rect 17092 22448 17098 22460
rect 17405 22457 17417 22460
rect 17451 22457 17463 22491
rect 17405 22451 17463 22457
rect 25041 22491 25099 22497
rect 25041 22457 25053 22491
rect 25087 22488 25099 22491
rect 25314 22488 25320 22500
rect 25087 22460 25320 22488
rect 25087 22457 25099 22460
rect 25041 22451 25099 22457
rect 25314 22448 25320 22460
rect 25372 22497 25378 22500
rect 25372 22491 25436 22497
rect 25372 22457 25390 22491
rect 25424 22457 25436 22491
rect 29546 22488 29552 22500
rect 29459 22460 29552 22488
rect 25372 22451 25436 22457
rect 25372 22448 25378 22451
rect 29546 22448 29552 22460
rect 29604 22488 29610 22500
rect 29886 22491 29944 22497
rect 29886 22488 29898 22491
rect 29604 22460 29898 22488
rect 29604 22448 29610 22460
rect 29886 22457 29898 22460
rect 29932 22457 29944 22491
rect 29886 22451 29944 22457
rect 16850 22420 16856 22432
rect 16684 22392 16856 22420
rect 16850 22380 16856 22392
rect 16908 22380 16914 22432
rect 22370 22420 22376 22432
rect 22331 22392 22376 22420
rect 22370 22380 22376 22392
rect 22428 22380 22434 22432
rect 32122 22420 32128 22432
rect 32083 22392 32128 22420
rect 32122 22380 32128 22392
rect 32180 22380 32186 22432
rect 33873 22423 33931 22429
rect 33873 22389 33885 22423
rect 33919 22420 33931 22423
rect 34422 22420 34428 22432
rect 33919 22392 34428 22420
rect 33919 22389 33931 22392
rect 33873 22383 33931 22389
rect 34422 22380 34428 22392
rect 34480 22380 34486 22432
rect 35158 22380 35164 22432
rect 35216 22420 35222 22432
rect 35529 22423 35587 22429
rect 35529 22420 35541 22423
rect 35216 22392 35541 22420
rect 35216 22380 35222 22392
rect 35529 22389 35541 22392
rect 35575 22420 35587 22423
rect 36817 22423 36875 22429
rect 36817 22420 36829 22423
rect 35575 22392 36829 22420
rect 35575 22389 35587 22392
rect 35529 22383 35587 22389
rect 36817 22389 36829 22392
rect 36863 22389 36875 22423
rect 36817 22383 36875 22389
rect 1104 22330 38824 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 38824 22330
rect 1104 22256 38824 22278
rect 13538 22216 13544 22228
rect 13499 22188 13544 22216
rect 13538 22176 13544 22188
rect 13596 22176 13602 22228
rect 14001 22219 14059 22225
rect 14001 22185 14013 22219
rect 14047 22216 14059 22219
rect 14090 22216 14096 22228
rect 14047 22188 14096 22216
rect 14047 22185 14059 22188
rect 14001 22179 14059 22185
rect 14090 22176 14096 22188
rect 14148 22176 14154 22228
rect 14642 22216 14648 22228
rect 14603 22188 14648 22216
rect 14642 22176 14648 22188
rect 14700 22176 14706 22228
rect 15105 22219 15163 22225
rect 15105 22185 15117 22219
rect 15151 22216 15163 22219
rect 15286 22216 15292 22228
rect 15151 22188 15292 22216
rect 15151 22185 15163 22188
rect 15105 22179 15163 22185
rect 15286 22176 15292 22188
rect 15344 22176 15350 22228
rect 16390 22216 16396 22228
rect 16351 22188 16396 22216
rect 16390 22176 16396 22188
rect 16448 22176 16454 22228
rect 17034 22216 17040 22228
rect 16995 22188 17040 22216
rect 17034 22176 17040 22188
rect 17092 22176 17098 22228
rect 17402 22216 17408 22228
rect 17363 22188 17408 22216
rect 17402 22176 17408 22188
rect 17460 22176 17466 22228
rect 18138 22216 18144 22228
rect 18099 22188 18144 22216
rect 18138 22176 18144 22188
rect 18196 22176 18202 22228
rect 29638 22216 29644 22228
rect 29599 22188 29644 22216
rect 29638 22176 29644 22188
rect 29696 22176 29702 22228
rect 33781 22219 33839 22225
rect 33781 22185 33793 22219
rect 33827 22216 33839 22219
rect 33870 22216 33876 22228
rect 33827 22188 33876 22216
rect 33827 22185 33839 22188
rect 33781 22179 33839 22185
rect 33870 22176 33876 22188
rect 33928 22176 33934 22228
rect 34517 22219 34575 22225
rect 34517 22185 34529 22219
rect 34563 22216 34575 22219
rect 34606 22216 34612 22228
rect 34563 22188 34612 22216
rect 34563 22185 34575 22188
rect 34517 22179 34575 22185
rect 34606 22176 34612 22188
rect 34664 22176 34670 22228
rect 35158 22216 35164 22228
rect 34716 22188 35164 22216
rect 19426 22148 19432 22160
rect 19260 22120 19432 22148
rect 12250 22040 12256 22092
rect 12308 22080 12314 22092
rect 13173 22083 13231 22089
rect 13173 22080 13185 22083
rect 12308 22052 13185 22080
rect 12308 22040 12314 22052
rect 13173 22049 13185 22052
rect 13219 22049 13231 22083
rect 13173 22043 13231 22049
rect 14093 22083 14151 22089
rect 14093 22049 14105 22083
rect 14139 22080 14151 22083
rect 14642 22080 14648 22092
rect 14139 22052 14648 22080
rect 14139 22049 14151 22052
rect 14093 22043 14151 22049
rect 14642 22040 14648 22052
rect 14700 22040 14706 22092
rect 15657 22083 15715 22089
rect 15657 22049 15669 22083
rect 15703 22049 15715 22083
rect 16850 22080 16856 22092
rect 16811 22052 16856 22080
rect 15657 22043 15715 22049
rect 12434 21972 12440 22024
rect 12492 22012 12498 22024
rect 12805 22015 12863 22021
rect 12805 22012 12817 22015
rect 12492 21984 12817 22012
rect 12492 21972 12498 21984
rect 12805 21981 12817 21984
rect 12851 21981 12863 22015
rect 12805 21975 12863 21981
rect 13538 21972 13544 22024
rect 13596 22012 13602 22024
rect 14185 22015 14243 22021
rect 14185 22012 14197 22015
rect 13596 21984 14197 22012
rect 13596 21972 13602 21984
rect 14185 21981 14197 21984
rect 14231 22012 14243 22015
rect 15010 22012 15016 22024
rect 14231 21984 15016 22012
rect 14231 21981 14243 21984
rect 14185 21975 14243 21981
rect 15010 21972 15016 21984
rect 15068 21972 15074 22024
rect 12986 21944 12992 21956
rect 12947 21916 12992 21944
rect 12986 21904 12992 21916
rect 13044 21904 13050 21956
rect 13633 21947 13691 21953
rect 13633 21913 13645 21947
rect 13679 21944 13691 21947
rect 15672 21944 15700 22043
rect 16850 22040 16856 22052
rect 16908 22040 16914 22092
rect 18598 22080 18604 22092
rect 18559 22052 18604 22080
rect 18598 22040 18604 22052
rect 18656 22040 18662 22092
rect 19153 22083 19211 22089
rect 19153 22049 19165 22083
rect 19199 22080 19211 22083
rect 19260 22080 19288 22120
rect 19426 22108 19432 22120
rect 19484 22108 19490 22160
rect 26786 22157 26792 22160
rect 26780 22148 26792 22157
rect 26747 22120 26792 22148
rect 26780 22111 26792 22120
rect 26786 22108 26792 22111
rect 26844 22108 26850 22160
rect 34330 22108 34336 22160
rect 34388 22148 34394 22160
rect 34716 22148 34744 22188
rect 35158 22176 35164 22188
rect 35216 22176 35222 22228
rect 34388 22120 34744 22148
rect 34876 22151 34934 22157
rect 34388 22108 34394 22120
rect 34876 22117 34888 22151
rect 34922 22148 34934 22151
rect 35250 22148 35256 22160
rect 34922 22120 35256 22148
rect 34922 22117 34934 22120
rect 34876 22111 34934 22117
rect 35250 22108 35256 22120
rect 35308 22108 35314 22160
rect 35618 22108 35624 22160
rect 35676 22108 35682 22160
rect 35802 22108 35808 22160
rect 35860 22148 35866 22160
rect 36170 22148 36176 22160
rect 35860 22120 36176 22148
rect 35860 22108 35866 22120
rect 36170 22108 36176 22120
rect 36228 22108 36234 22160
rect 19199 22052 19288 22080
rect 19199 22049 19211 22052
rect 19153 22043 19211 22049
rect 22278 22040 22284 22092
rect 22336 22080 22342 22092
rect 22741 22083 22799 22089
rect 22741 22080 22753 22083
rect 22336 22052 22753 22080
rect 22336 22040 22342 22052
rect 22741 22049 22753 22052
rect 22787 22049 22799 22083
rect 22741 22043 22799 22049
rect 22833 22083 22891 22089
rect 22833 22049 22845 22083
rect 22879 22080 22891 22083
rect 23106 22080 23112 22092
rect 22879 22052 23112 22080
rect 22879 22049 22891 22052
rect 22833 22043 22891 22049
rect 23106 22040 23112 22052
rect 23164 22040 23170 22092
rect 24026 22040 24032 22092
rect 24084 22080 24090 22092
rect 24193 22083 24251 22089
rect 24193 22080 24205 22083
rect 24084 22052 24205 22080
rect 24084 22040 24090 22052
rect 24193 22049 24205 22052
rect 24239 22049 24251 22083
rect 35636 22080 35664 22108
rect 35710 22080 35716 22092
rect 35636 22052 35716 22080
rect 24193 22043 24251 22049
rect 35710 22040 35716 22052
rect 35768 22040 35774 22092
rect 15746 21972 15752 22024
rect 15804 22012 15810 22024
rect 15933 22015 15991 22021
rect 15804 21984 15849 22012
rect 15804 21972 15810 21984
rect 15933 21981 15945 22015
rect 15979 22012 15991 22015
rect 16022 22012 16028 22024
rect 15979 21984 16028 22012
rect 15979 21981 15991 21984
rect 15933 21975 15991 21981
rect 16022 21972 16028 21984
rect 16080 21972 16086 22024
rect 22370 21972 22376 22024
rect 22428 22012 22434 22024
rect 23014 22012 23020 22024
rect 22428 21984 23020 22012
rect 22428 21972 22434 21984
rect 23014 21972 23020 21984
rect 23072 21972 23078 22024
rect 23937 22015 23995 22021
rect 23937 21981 23949 22015
rect 23983 21981 23995 22015
rect 26510 22012 26516 22024
rect 26471 21984 26516 22012
rect 23937 21975 23995 21981
rect 15838 21944 15844 21956
rect 13679 21916 15844 21944
rect 13679 21913 13691 21916
rect 13633 21907 13691 21913
rect 15838 21904 15844 21916
rect 15896 21904 15902 21956
rect 18785 21947 18843 21953
rect 18785 21913 18797 21947
rect 18831 21944 18843 21947
rect 19242 21944 19248 21956
rect 18831 21916 19248 21944
rect 18831 21913 18843 21916
rect 18785 21907 18843 21913
rect 19242 21904 19248 21916
rect 19300 21904 19306 21956
rect 19150 21836 19156 21888
rect 19208 21876 19214 21888
rect 19613 21879 19671 21885
rect 19613 21876 19625 21879
rect 19208 21848 19625 21876
rect 19208 21836 19214 21848
rect 19613 21845 19625 21848
rect 19659 21876 19671 21879
rect 19981 21879 20039 21885
rect 19981 21876 19993 21879
rect 19659 21848 19993 21876
rect 19659 21845 19671 21848
rect 19613 21839 19671 21845
rect 19981 21845 19993 21848
rect 20027 21876 20039 21879
rect 21082 21876 21088 21888
rect 20027 21848 21088 21876
rect 20027 21845 20039 21848
rect 19981 21839 20039 21845
rect 21082 21836 21088 21848
rect 21140 21836 21146 21888
rect 22278 21876 22284 21888
rect 22239 21848 22284 21876
rect 22278 21836 22284 21848
rect 22336 21836 22342 21888
rect 22373 21879 22431 21885
rect 22373 21845 22385 21879
rect 22419 21876 22431 21879
rect 23474 21876 23480 21888
rect 22419 21848 23480 21876
rect 22419 21845 22431 21848
rect 22373 21839 22431 21845
rect 23474 21836 23480 21848
rect 23532 21836 23538 21888
rect 23658 21836 23664 21888
rect 23716 21876 23722 21888
rect 23753 21879 23811 21885
rect 23753 21876 23765 21879
rect 23716 21848 23765 21876
rect 23716 21836 23722 21848
rect 23753 21845 23765 21848
rect 23799 21876 23811 21879
rect 23952 21876 23980 21975
rect 26510 21972 26516 21984
rect 26568 21972 26574 22024
rect 32122 21972 32128 22024
rect 32180 22012 32186 22024
rect 34149 22015 34207 22021
rect 34149 22012 34161 22015
rect 32180 21984 34161 22012
rect 32180 21972 32186 21984
rect 34149 21981 34161 21984
rect 34195 22012 34207 22015
rect 34606 22012 34612 22024
rect 34195 21984 34612 22012
rect 34195 21981 34207 21984
rect 34149 21975 34207 21981
rect 34606 21972 34612 21984
rect 34664 21972 34670 22024
rect 36170 21944 36176 21956
rect 35820 21916 36176 21944
rect 25130 21876 25136 21888
rect 23799 21848 25136 21876
rect 23799 21845 23811 21848
rect 23753 21839 23811 21845
rect 25130 21836 25136 21848
rect 25188 21836 25194 21888
rect 25314 21876 25320 21888
rect 25275 21848 25320 21876
rect 25314 21836 25320 21848
rect 25372 21836 25378 21888
rect 27154 21836 27160 21888
rect 27212 21876 27218 21888
rect 27893 21879 27951 21885
rect 27893 21876 27905 21879
rect 27212 21848 27905 21876
rect 27212 21836 27218 21848
rect 27893 21845 27905 21848
rect 27939 21845 27951 21879
rect 27893 21839 27951 21845
rect 29730 21836 29736 21888
rect 29788 21876 29794 21888
rect 30009 21879 30067 21885
rect 30009 21876 30021 21879
rect 29788 21848 30021 21876
rect 29788 21836 29794 21848
rect 30009 21845 30021 21848
rect 30055 21876 30067 21879
rect 30558 21876 30564 21888
rect 30055 21848 30564 21876
rect 30055 21845 30067 21848
rect 30009 21839 30067 21845
rect 30558 21836 30564 21848
rect 30616 21836 30622 21888
rect 35342 21836 35348 21888
rect 35400 21876 35406 21888
rect 35820 21876 35848 21916
rect 36170 21904 36176 21916
rect 36228 21904 36234 21956
rect 35986 21876 35992 21888
rect 35400 21848 35848 21876
rect 35947 21848 35992 21876
rect 35400 21836 35406 21848
rect 35986 21836 35992 21848
rect 36044 21836 36050 21888
rect 1104 21786 38824 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 34966 21786
rect 35018 21734 35030 21786
rect 35082 21734 35094 21786
rect 35146 21734 35158 21786
rect 35210 21734 38824 21786
rect 1104 21712 38824 21734
rect 8570 21672 8576 21684
rect 8531 21644 8576 21672
rect 8570 21632 8576 21644
rect 8628 21632 8634 21684
rect 13170 21672 13176 21684
rect 13131 21644 13176 21672
rect 13170 21632 13176 21644
rect 13228 21632 13234 21684
rect 14642 21672 14648 21684
rect 14603 21644 14648 21672
rect 14642 21632 14648 21644
rect 14700 21632 14706 21684
rect 15657 21675 15715 21681
rect 15657 21641 15669 21675
rect 15703 21672 15715 21675
rect 15746 21672 15752 21684
rect 15703 21644 15752 21672
rect 15703 21641 15715 21644
rect 15657 21635 15715 21641
rect 15746 21632 15752 21644
rect 15804 21632 15810 21684
rect 15838 21632 15844 21684
rect 15896 21672 15902 21684
rect 15933 21675 15991 21681
rect 15933 21672 15945 21675
rect 15896 21644 15945 21672
rect 15896 21632 15902 21644
rect 15933 21641 15945 21644
rect 15979 21641 15991 21675
rect 15933 21635 15991 21641
rect 16393 21675 16451 21681
rect 16393 21641 16405 21675
rect 16439 21672 16451 21675
rect 16850 21672 16856 21684
rect 16439 21644 16856 21672
rect 16439 21641 16451 21644
rect 16393 21635 16451 21641
rect 16850 21632 16856 21644
rect 16908 21672 16914 21684
rect 17405 21675 17463 21681
rect 17405 21672 17417 21675
rect 16908 21644 17417 21672
rect 16908 21632 16914 21644
rect 17405 21641 17417 21644
rect 17451 21641 17463 21675
rect 19978 21672 19984 21684
rect 19939 21644 19984 21672
rect 17405 21635 17463 21641
rect 19978 21632 19984 21644
rect 20036 21632 20042 21684
rect 22278 21632 22284 21684
rect 22336 21672 22342 21684
rect 22465 21675 22523 21681
rect 22465 21672 22477 21675
rect 22336 21644 22477 21672
rect 22336 21632 22342 21644
rect 22465 21641 22477 21644
rect 22511 21672 22523 21675
rect 23385 21675 23443 21681
rect 23385 21672 23397 21675
rect 22511 21644 23397 21672
rect 22511 21641 22523 21644
rect 22465 21635 22523 21641
rect 23385 21641 23397 21644
rect 23431 21641 23443 21675
rect 23385 21635 23443 21641
rect 26053 21675 26111 21681
rect 26053 21641 26065 21675
rect 26099 21672 26111 21675
rect 26142 21672 26148 21684
rect 26099 21644 26148 21672
rect 26099 21641 26111 21644
rect 26053 21635 26111 21641
rect 13188 21536 13216 21632
rect 17037 21539 17095 21545
rect 13188 21508 13400 21536
rect 8757 21471 8815 21477
rect 8757 21437 8769 21471
rect 8803 21468 8815 21471
rect 8803 21440 9168 21468
rect 8803 21437 8815 21440
rect 8757 21431 8815 21437
rect 9140 21344 9168 21440
rect 12434 21428 12440 21480
rect 12492 21468 12498 21480
rect 13265 21471 13323 21477
rect 13265 21468 13277 21471
rect 12492 21440 13277 21468
rect 12492 21428 12498 21440
rect 13265 21437 13277 21440
rect 13311 21437 13323 21471
rect 13372 21468 13400 21508
rect 17037 21505 17049 21539
rect 17083 21536 17095 21539
rect 17126 21536 17132 21548
rect 17083 21508 17132 21536
rect 17083 21505 17095 21508
rect 17037 21499 17095 21505
rect 17126 21496 17132 21508
rect 17184 21536 17190 21548
rect 17770 21536 17776 21548
rect 17184 21508 17776 21536
rect 17184 21496 17190 21508
rect 17770 21496 17776 21508
rect 17828 21496 17834 21548
rect 23400 21536 23428 21635
rect 26142 21632 26148 21644
rect 26200 21632 26206 21684
rect 26786 21672 26792 21684
rect 26747 21644 26792 21672
rect 26786 21632 26792 21644
rect 26844 21632 26850 21684
rect 27890 21672 27896 21684
rect 27851 21644 27896 21672
rect 27890 21632 27896 21644
rect 27948 21632 27954 21684
rect 29546 21632 29552 21684
rect 29604 21672 29610 21684
rect 31113 21675 31171 21681
rect 31113 21672 31125 21675
rect 29604 21644 31125 21672
rect 29604 21632 29610 21644
rect 31113 21641 31125 21644
rect 31159 21641 31171 21675
rect 31113 21635 31171 21641
rect 34701 21675 34759 21681
rect 34701 21641 34713 21675
rect 34747 21672 34759 21675
rect 35250 21672 35256 21684
rect 34747 21644 35256 21672
rect 34747 21641 34759 21644
rect 34701 21635 34759 21641
rect 35250 21632 35256 21644
rect 35308 21632 35314 21684
rect 35802 21632 35808 21684
rect 35860 21672 35866 21684
rect 36078 21672 36084 21684
rect 35860 21644 36084 21672
rect 35860 21632 35866 21644
rect 36078 21632 36084 21644
rect 36136 21672 36142 21684
rect 36265 21675 36323 21681
rect 36265 21672 36277 21675
rect 36136 21644 36277 21672
rect 36136 21632 36142 21644
rect 36265 21641 36277 21644
rect 36311 21641 36323 21675
rect 36265 21635 36323 21641
rect 26326 21564 26332 21616
rect 26384 21604 26390 21616
rect 27433 21607 27491 21613
rect 27433 21604 27445 21607
rect 26384 21576 27445 21604
rect 26384 21564 26390 21576
rect 27433 21573 27445 21576
rect 27479 21573 27491 21607
rect 27433 21567 27491 21573
rect 23400 21508 23796 21536
rect 13521 21471 13579 21477
rect 13521 21468 13533 21471
rect 13372 21440 13533 21468
rect 13265 21431 13323 21437
rect 13521 21437 13533 21440
rect 13567 21437 13579 21471
rect 13521 21431 13579 21437
rect 17865 21471 17923 21477
rect 17865 21437 17877 21471
rect 17911 21468 17923 21471
rect 18601 21471 18659 21477
rect 18601 21468 18613 21471
rect 17911 21440 18613 21468
rect 17911 21437 17923 21440
rect 17865 21431 17923 21437
rect 18601 21437 18613 21440
rect 18647 21468 18659 21471
rect 19150 21468 19156 21480
rect 18647 21440 19156 21468
rect 18647 21437 18659 21440
rect 18601 21431 18659 21437
rect 19150 21428 19156 21440
rect 19208 21428 19214 21480
rect 21082 21468 21088 21480
rect 21043 21440 21088 21468
rect 21082 21428 21088 21440
rect 21140 21428 21146 21480
rect 23658 21468 23664 21480
rect 23619 21440 23664 21468
rect 23658 21428 23664 21440
rect 23716 21428 23722 21480
rect 23768 21468 23796 21508
rect 23917 21471 23975 21477
rect 23917 21468 23929 21471
rect 23768 21440 23929 21468
rect 23917 21437 23929 21440
rect 23963 21437 23975 21471
rect 26142 21468 26148 21480
rect 26103 21440 26148 21468
rect 23917 21431 23975 21437
rect 26142 21428 26148 21440
rect 26200 21428 26206 21480
rect 27249 21471 27307 21477
rect 27249 21437 27261 21471
rect 27295 21468 27307 21471
rect 27890 21468 27896 21480
rect 27295 21440 27896 21468
rect 27295 21437 27307 21440
rect 27249 21431 27307 21437
rect 27890 21428 27896 21440
rect 27948 21428 27954 21480
rect 29733 21471 29791 21477
rect 29733 21437 29745 21471
rect 29779 21468 29791 21471
rect 30558 21468 30564 21480
rect 29779 21440 30564 21468
rect 29779 21437 29791 21440
rect 29733 21431 29791 21437
rect 30558 21428 30564 21440
rect 30616 21428 30622 21480
rect 33965 21471 34023 21477
rect 33965 21437 33977 21471
rect 34011 21468 34023 21471
rect 34606 21468 34612 21480
rect 34011 21440 34612 21468
rect 34011 21437 34023 21440
rect 33965 21431 34023 21437
rect 34606 21428 34612 21440
rect 34664 21468 34670 21480
rect 34882 21468 34888 21480
rect 34664 21440 34888 21468
rect 34664 21428 34670 21440
rect 34882 21428 34888 21440
rect 34940 21428 34946 21480
rect 35152 21471 35210 21477
rect 35152 21468 35164 21471
rect 34992 21440 35164 21468
rect 12805 21403 12863 21409
rect 12805 21369 12817 21403
rect 12851 21400 12863 21403
rect 12986 21400 12992 21412
rect 12851 21372 12992 21400
rect 12851 21369 12863 21372
rect 12805 21363 12863 21369
rect 12986 21360 12992 21372
rect 13044 21400 13050 21412
rect 14642 21400 14648 21412
rect 13044 21372 14648 21400
rect 13044 21360 13050 21372
rect 14642 21360 14648 21372
rect 14700 21360 14706 21412
rect 18846 21403 18904 21409
rect 18846 21400 18858 21403
rect 18432 21372 18858 21400
rect 9122 21332 9128 21344
rect 9083 21304 9128 21332
rect 9122 21292 9128 21304
rect 9180 21292 9186 21344
rect 12250 21332 12256 21344
rect 12211 21304 12256 21332
rect 12250 21292 12256 21304
rect 12308 21292 12314 21344
rect 14090 21292 14096 21344
rect 14148 21332 14154 21344
rect 15197 21335 15255 21341
rect 15197 21332 15209 21335
rect 14148 21304 15209 21332
rect 14148 21292 14154 21304
rect 15197 21301 15209 21304
rect 15243 21301 15255 21335
rect 16758 21332 16764 21344
rect 16719 21304 16764 21332
rect 15197 21295 15255 21301
rect 16758 21292 16764 21304
rect 16816 21292 16822 21344
rect 16850 21292 16856 21344
rect 16908 21332 16914 21344
rect 16908 21304 16953 21332
rect 16908 21292 16914 21304
rect 17954 21292 17960 21344
rect 18012 21332 18018 21344
rect 18432 21341 18460 21372
rect 18846 21369 18858 21372
rect 18892 21400 18904 21403
rect 19242 21400 19248 21412
rect 18892 21372 19248 21400
rect 18892 21369 18904 21372
rect 18846 21363 18904 21369
rect 19242 21360 19248 21372
rect 19300 21360 19306 21412
rect 20993 21403 21051 21409
rect 20993 21369 21005 21403
rect 21039 21400 21051 21403
rect 21330 21403 21388 21409
rect 21330 21400 21342 21403
rect 21039 21372 21342 21400
rect 21039 21369 21051 21372
rect 20993 21363 21051 21369
rect 21330 21369 21342 21372
rect 21376 21400 21388 21403
rect 21376 21372 23152 21400
rect 21376 21369 21388 21372
rect 21330 21363 21388 21369
rect 23124 21344 23152 21372
rect 25130 21360 25136 21412
rect 25188 21400 25194 21412
rect 25685 21403 25743 21409
rect 25685 21400 25697 21403
rect 25188 21372 25697 21400
rect 25188 21360 25194 21372
rect 25685 21369 25697 21372
rect 25731 21400 25743 21403
rect 26510 21400 26516 21412
rect 25731 21372 26516 21400
rect 25731 21369 25743 21372
rect 25685 21363 25743 21369
rect 26510 21360 26516 21372
rect 26568 21400 26574 21412
rect 27157 21403 27215 21409
rect 27157 21400 27169 21403
rect 26568 21372 27169 21400
rect 26568 21360 26574 21372
rect 27157 21369 27169 21372
rect 27203 21400 27215 21403
rect 27614 21400 27620 21412
rect 27203 21372 27620 21400
rect 27203 21369 27215 21372
rect 27157 21363 27215 21369
rect 27614 21360 27620 21372
rect 27672 21360 27678 21412
rect 29641 21403 29699 21409
rect 29641 21369 29653 21403
rect 29687 21400 29699 21403
rect 29978 21403 30036 21409
rect 29978 21400 29990 21403
rect 29687 21372 29990 21400
rect 29687 21369 29699 21372
rect 29641 21363 29699 21369
rect 29978 21369 29990 21372
rect 30024 21400 30036 21403
rect 30190 21400 30196 21412
rect 30024 21372 30196 21400
rect 30024 21369 30036 21372
rect 29978 21363 30036 21369
rect 30190 21360 30196 21372
rect 30248 21360 30254 21412
rect 33318 21360 33324 21412
rect 33376 21400 33382 21412
rect 34333 21403 34391 21409
rect 34333 21400 34345 21403
rect 33376 21372 34345 21400
rect 33376 21360 33382 21372
rect 34333 21369 34345 21372
rect 34379 21400 34391 21403
rect 34992 21400 35020 21440
rect 35152 21437 35164 21440
rect 35198 21468 35210 21471
rect 35986 21468 35992 21480
rect 35198 21440 35992 21468
rect 35198 21437 35210 21440
rect 35152 21431 35210 21437
rect 35986 21428 35992 21440
rect 36044 21428 36050 21480
rect 34379 21372 35020 21400
rect 34379 21369 34391 21372
rect 34333 21363 34391 21369
rect 18417 21335 18475 21341
rect 18417 21332 18429 21335
rect 18012 21304 18429 21332
rect 18012 21292 18018 21304
rect 18417 21301 18429 21304
rect 18463 21301 18475 21335
rect 23106 21332 23112 21344
rect 23067 21304 23112 21332
rect 18417 21295 18475 21301
rect 23106 21292 23112 21304
rect 23164 21292 23170 21344
rect 24026 21292 24032 21344
rect 24084 21332 24090 21344
rect 24946 21332 24952 21344
rect 24084 21304 24952 21332
rect 24084 21292 24090 21304
rect 24946 21292 24952 21304
rect 25004 21332 25010 21344
rect 25041 21335 25099 21341
rect 25041 21332 25053 21335
rect 25004 21304 25053 21332
rect 25004 21292 25010 21304
rect 25041 21301 25053 21304
rect 25087 21301 25099 21335
rect 25041 21295 25099 21301
rect 26234 21292 26240 21344
rect 26292 21332 26298 21344
rect 26329 21335 26387 21341
rect 26329 21332 26341 21335
rect 26292 21304 26341 21332
rect 26292 21292 26298 21304
rect 26329 21301 26341 21304
rect 26375 21301 26387 21335
rect 26329 21295 26387 21301
rect 1104 21242 38824 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 38824 21242
rect 1104 21168 38824 21190
rect 13722 21088 13728 21140
rect 13780 21128 13786 21140
rect 14090 21128 14096 21140
rect 13780 21100 14096 21128
rect 13780 21088 13786 21100
rect 14090 21088 14096 21100
rect 14148 21088 14154 21140
rect 15286 21128 15292 21140
rect 15247 21100 15292 21128
rect 15286 21088 15292 21100
rect 15344 21088 15350 21140
rect 16758 21128 16764 21140
rect 16719 21100 16764 21128
rect 16758 21088 16764 21100
rect 16816 21128 16822 21140
rect 17681 21131 17739 21137
rect 17681 21128 17693 21131
rect 16816 21100 17693 21128
rect 16816 21088 16822 21100
rect 17681 21097 17693 21100
rect 17727 21097 17739 21131
rect 17681 21091 17739 21097
rect 18598 21088 18604 21140
rect 18656 21128 18662 21140
rect 18693 21131 18751 21137
rect 18693 21128 18705 21131
rect 18656 21100 18705 21128
rect 18656 21088 18662 21100
rect 18693 21097 18705 21100
rect 18739 21097 18751 21131
rect 18693 21091 18751 21097
rect 19334 21088 19340 21140
rect 19392 21128 19398 21140
rect 19429 21131 19487 21137
rect 19429 21128 19441 21131
rect 19392 21100 19441 21128
rect 19392 21088 19398 21100
rect 19429 21097 19441 21100
rect 19475 21097 19487 21131
rect 21082 21128 21088 21140
rect 21043 21100 21088 21128
rect 19429 21091 19487 21097
rect 21082 21088 21088 21100
rect 21140 21088 21146 21140
rect 23106 21128 23112 21140
rect 23067 21100 23112 21128
rect 23106 21088 23112 21100
rect 23164 21088 23170 21140
rect 24026 21128 24032 21140
rect 23987 21100 24032 21128
rect 24026 21088 24032 21100
rect 24084 21088 24090 21140
rect 25498 21128 25504 21140
rect 25459 21100 25504 21128
rect 25498 21088 25504 21100
rect 25556 21088 25562 21140
rect 26602 21088 26608 21140
rect 26660 21128 26666 21140
rect 26881 21131 26939 21137
rect 26881 21128 26893 21131
rect 26660 21100 26893 21128
rect 26660 21088 26666 21100
rect 26881 21097 26893 21100
rect 26927 21128 26939 21131
rect 28261 21131 28319 21137
rect 28261 21128 28273 21131
rect 26927 21100 28273 21128
rect 26927 21097 26939 21100
rect 26881 21091 26939 21097
rect 28261 21097 28273 21100
rect 28307 21097 28319 21131
rect 28261 21091 28319 21097
rect 30558 21088 30564 21140
rect 30616 21128 30622 21140
rect 30653 21131 30711 21137
rect 30653 21128 30665 21131
rect 30616 21100 30665 21128
rect 30616 21088 30622 21100
rect 30653 21097 30665 21100
rect 30699 21128 30711 21131
rect 32122 21128 32128 21140
rect 30699 21100 32128 21128
rect 30699 21097 30711 21100
rect 30653 21091 30711 21097
rect 32122 21088 32128 21100
rect 32180 21088 32186 21140
rect 33318 21128 33324 21140
rect 33279 21100 33324 21128
rect 33318 21088 33324 21100
rect 33376 21088 33382 21140
rect 35894 21088 35900 21140
rect 35952 21128 35958 21140
rect 36633 21131 36691 21137
rect 36633 21128 36645 21131
rect 35952 21100 36645 21128
rect 35952 21088 35958 21100
rect 36633 21097 36645 21100
rect 36679 21097 36691 21131
rect 36633 21091 36691 21097
rect 12986 21069 12992 21072
rect 12980 21060 12992 21069
rect 12947 21032 12992 21060
rect 12980 21023 12992 21032
rect 12986 21020 12992 21023
rect 13044 21020 13050 21072
rect 17126 21060 17132 21072
rect 17087 21032 17132 21060
rect 17126 21020 17132 21032
rect 17184 21020 17190 21072
rect 12434 20952 12440 21004
rect 12492 20992 12498 21004
rect 12713 20995 12771 21001
rect 12713 20992 12725 20995
rect 12492 20964 12725 20992
rect 12492 20952 12498 20964
rect 12713 20961 12725 20964
rect 12759 20961 12771 20995
rect 12713 20955 12771 20961
rect 15657 20995 15715 21001
rect 15657 20961 15669 20995
rect 15703 20992 15715 20995
rect 16482 20992 16488 21004
rect 15703 20964 16488 20992
rect 15703 20961 15715 20964
rect 15657 20955 15715 20961
rect 16482 20952 16488 20964
rect 16540 20952 16546 21004
rect 15746 20924 15752 20936
rect 15707 20896 15752 20924
rect 15746 20884 15752 20896
rect 15804 20884 15810 20936
rect 15933 20927 15991 20933
rect 15933 20893 15945 20927
rect 15979 20924 15991 20927
rect 16022 20924 16028 20936
rect 15979 20896 16028 20924
rect 15979 20893 15991 20896
rect 15933 20887 15991 20893
rect 14737 20859 14795 20865
rect 14737 20825 14749 20859
rect 14783 20856 14795 20859
rect 15105 20859 15163 20865
rect 15105 20856 15117 20859
rect 14783 20828 15117 20856
rect 14783 20825 14795 20828
rect 14737 20819 14795 20825
rect 15105 20825 15117 20828
rect 15151 20856 15163 20859
rect 15948 20856 15976 20887
rect 16022 20884 16028 20896
rect 16080 20924 16086 20936
rect 17144 20924 17172 21020
rect 17954 20952 17960 21004
rect 18012 20992 18018 21004
rect 18049 20995 18107 21001
rect 18049 20992 18061 20995
rect 18012 20964 18061 20992
rect 18012 20952 18018 20964
rect 18049 20961 18061 20964
rect 18095 20961 18107 20995
rect 18049 20955 18107 20961
rect 18141 20995 18199 21001
rect 18141 20961 18153 20995
rect 18187 20992 18199 20995
rect 18322 20992 18328 21004
rect 18187 20964 18328 20992
rect 18187 20961 18199 20964
rect 18141 20955 18199 20961
rect 18322 20952 18328 20964
rect 18380 20952 18386 21004
rect 19150 20952 19156 21004
rect 19208 20992 19214 21004
rect 19245 20995 19303 21001
rect 19245 20992 19257 20995
rect 19208 20964 19257 20992
rect 19208 20952 19214 20964
rect 19245 20961 19257 20964
rect 19291 20992 19303 20995
rect 19518 20992 19524 21004
rect 19291 20964 19524 20992
rect 19291 20961 19303 20964
rect 19245 20955 19303 20961
rect 19518 20952 19524 20964
rect 19576 20952 19582 21004
rect 21726 20992 21732 21004
rect 21687 20964 21732 20992
rect 21726 20952 21732 20964
rect 21784 20952 21790 21004
rect 22002 21001 22008 21004
rect 21996 20992 22008 21001
rect 21963 20964 22008 20992
rect 21996 20955 22008 20964
rect 22002 20952 22008 20955
rect 22060 20952 22066 21004
rect 24210 20992 24216 21004
rect 24171 20964 24216 20992
rect 24210 20952 24216 20964
rect 24268 20952 24274 21004
rect 28074 20992 28080 21004
rect 28035 20964 28080 20992
rect 28074 20952 28080 20964
rect 28132 20952 28138 21004
rect 29822 20992 29828 21004
rect 29783 20964 29828 20992
rect 29822 20952 29828 20964
rect 29880 20952 29886 21004
rect 29917 20995 29975 21001
rect 29917 20961 29929 20995
rect 29963 20992 29975 20995
rect 30282 20992 30288 21004
rect 29963 20964 30288 20992
rect 29963 20961 29975 20964
rect 29917 20955 29975 20961
rect 18230 20924 18236 20936
rect 16080 20896 17172 20924
rect 18191 20896 18236 20924
rect 16080 20884 16086 20896
rect 18230 20884 18236 20896
rect 18288 20884 18294 20936
rect 26970 20924 26976 20936
rect 26931 20896 26976 20924
rect 26970 20884 26976 20896
rect 27028 20884 27034 20936
rect 27154 20924 27160 20936
rect 27115 20896 27160 20924
rect 27154 20884 27160 20896
rect 27212 20884 27218 20936
rect 29365 20927 29423 20933
rect 29365 20893 29377 20927
rect 29411 20924 29423 20927
rect 29932 20924 29960 20955
rect 30282 20952 30288 20964
rect 30340 20952 30346 21004
rect 29411 20896 29960 20924
rect 30009 20927 30067 20933
rect 29411 20893 29423 20896
rect 29365 20887 29423 20893
rect 30009 20893 30021 20927
rect 30055 20893 30067 20927
rect 30009 20887 30067 20893
rect 15151 20828 15976 20856
rect 16485 20859 16543 20865
rect 15151 20825 15163 20828
rect 15105 20819 15163 20825
rect 16485 20825 16497 20859
rect 16531 20856 16543 20859
rect 16850 20856 16856 20868
rect 16531 20828 16856 20856
rect 16531 20825 16543 20828
rect 16485 20819 16543 20825
rect 16850 20816 16856 20828
rect 16908 20856 16914 20868
rect 17862 20856 17868 20868
rect 16908 20828 17868 20856
rect 16908 20816 16914 20828
rect 17862 20816 17868 20828
rect 17920 20816 17926 20868
rect 26329 20859 26387 20865
rect 26329 20825 26341 20859
rect 26375 20856 26387 20859
rect 27172 20856 27200 20884
rect 26375 20828 27200 20856
rect 26375 20825 26387 20828
rect 26329 20819 26387 20825
rect 29086 20816 29092 20868
rect 29144 20856 29150 20868
rect 29546 20856 29552 20868
rect 29144 20828 29552 20856
rect 29144 20816 29150 20828
rect 29546 20816 29552 20828
rect 29604 20856 29610 20868
rect 30024 20856 30052 20887
rect 33686 20884 33692 20936
rect 33744 20924 33750 20936
rect 33873 20927 33931 20933
rect 33873 20924 33885 20927
rect 33744 20896 33885 20924
rect 33744 20884 33750 20896
rect 33873 20893 33885 20896
rect 33919 20924 33931 20927
rect 33965 20927 34023 20933
rect 33965 20924 33977 20927
rect 33919 20896 33977 20924
rect 33919 20893 33931 20896
rect 33873 20887 33931 20893
rect 33965 20893 33977 20896
rect 34011 20893 34023 20927
rect 33965 20887 34023 20893
rect 34146 20884 34152 20936
rect 34204 20924 34210 20936
rect 34288 20927 34346 20933
rect 34288 20924 34300 20927
rect 34204 20896 34300 20924
rect 34204 20884 34210 20896
rect 34288 20893 34300 20896
rect 34334 20893 34346 20927
rect 34288 20887 34346 20893
rect 34422 20884 34428 20936
rect 34480 20924 34486 20936
rect 34480 20896 34525 20924
rect 34480 20884 34486 20896
rect 34606 20884 34612 20936
rect 34664 20924 34670 20936
rect 34701 20927 34759 20933
rect 34701 20924 34713 20927
rect 34664 20896 34713 20924
rect 34664 20884 34670 20896
rect 34701 20893 34713 20896
rect 34747 20893 34759 20927
rect 34701 20887 34759 20893
rect 34882 20884 34888 20936
rect 34940 20924 34946 20936
rect 34940 20896 35940 20924
rect 34940 20884 34946 20896
rect 29604 20828 30052 20856
rect 29604 20816 29610 20828
rect 35912 20800 35940 20896
rect 16666 20748 16672 20800
rect 16724 20788 16730 20800
rect 17497 20791 17555 20797
rect 17497 20788 17509 20791
rect 16724 20760 17509 20788
rect 16724 20748 16730 20760
rect 17497 20757 17509 20760
rect 17543 20757 17555 20791
rect 17497 20751 17555 20757
rect 20530 20748 20536 20800
rect 20588 20788 20594 20800
rect 21637 20791 21695 20797
rect 21637 20788 21649 20791
rect 20588 20760 21649 20788
rect 20588 20748 20594 20760
rect 21637 20757 21649 20760
rect 21683 20788 21695 20791
rect 23014 20788 23020 20800
rect 21683 20760 23020 20788
rect 21683 20757 21695 20760
rect 21637 20751 21695 20757
rect 23014 20748 23020 20760
rect 23072 20748 23078 20800
rect 26510 20788 26516 20800
rect 26471 20760 26516 20788
rect 26510 20748 26516 20760
rect 26568 20748 26574 20800
rect 27614 20788 27620 20800
rect 27575 20760 27620 20788
rect 27614 20748 27620 20760
rect 27672 20748 27678 20800
rect 29454 20788 29460 20800
rect 29415 20760 29460 20788
rect 29454 20748 29460 20760
rect 29512 20748 29518 20800
rect 35342 20748 35348 20800
rect 35400 20788 35406 20800
rect 35805 20791 35863 20797
rect 35805 20788 35817 20791
rect 35400 20760 35817 20788
rect 35400 20748 35406 20760
rect 35805 20757 35817 20760
rect 35851 20757 35863 20791
rect 35805 20751 35863 20757
rect 35894 20748 35900 20800
rect 35952 20788 35958 20800
rect 36081 20791 36139 20797
rect 36081 20788 36093 20791
rect 35952 20760 36093 20788
rect 35952 20748 35958 20760
rect 36081 20757 36093 20760
rect 36127 20788 36139 20791
rect 36538 20788 36544 20800
rect 36127 20760 36544 20788
rect 36127 20757 36139 20760
rect 36081 20751 36139 20757
rect 36538 20748 36544 20760
rect 36596 20748 36602 20800
rect 1104 20698 38824 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 34966 20698
rect 35018 20646 35030 20698
rect 35082 20646 35094 20698
rect 35146 20646 35158 20698
rect 35210 20646 38824 20698
rect 1104 20624 38824 20646
rect 10042 20584 10048 20596
rect 10003 20556 10048 20584
rect 10042 20544 10048 20556
rect 10100 20544 10106 20596
rect 12805 20587 12863 20593
rect 12805 20553 12817 20587
rect 12851 20584 12863 20587
rect 12986 20584 12992 20596
rect 12851 20556 12992 20584
rect 12851 20553 12863 20556
rect 12805 20547 12863 20553
rect 12986 20544 12992 20556
rect 13044 20544 13050 20596
rect 15197 20587 15255 20593
rect 15197 20553 15209 20587
rect 15243 20584 15255 20587
rect 15657 20587 15715 20593
rect 15657 20584 15669 20587
rect 15243 20556 15669 20584
rect 15243 20553 15255 20556
rect 15197 20547 15255 20553
rect 15657 20553 15669 20556
rect 15703 20584 15715 20587
rect 15746 20584 15752 20596
rect 15703 20556 15752 20584
rect 15703 20553 15715 20556
rect 15657 20547 15715 20553
rect 15746 20544 15752 20556
rect 15804 20544 15810 20596
rect 16574 20544 16580 20596
rect 16632 20584 16638 20596
rect 16669 20587 16727 20593
rect 16669 20584 16681 20587
rect 16632 20556 16681 20584
rect 16632 20544 16638 20556
rect 16669 20553 16681 20556
rect 16715 20553 16727 20587
rect 16669 20547 16727 20553
rect 17129 20587 17187 20593
rect 17129 20553 17141 20587
rect 17175 20584 17187 20587
rect 17954 20584 17960 20596
rect 17175 20556 17960 20584
rect 17175 20553 17187 20556
rect 17129 20547 17187 20553
rect 17954 20544 17960 20556
rect 18012 20544 18018 20596
rect 19334 20544 19340 20596
rect 19392 20584 19398 20596
rect 19429 20587 19487 20593
rect 19429 20584 19441 20587
rect 19392 20556 19441 20584
rect 19392 20544 19398 20556
rect 19429 20553 19441 20556
rect 19475 20553 19487 20587
rect 19429 20547 19487 20553
rect 19518 20544 19524 20596
rect 19576 20584 19582 20596
rect 19981 20587 20039 20593
rect 19981 20584 19993 20587
rect 19576 20556 19993 20584
rect 19576 20544 19582 20556
rect 19981 20553 19993 20556
rect 20027 20553 20039 20587
rect 26602 20584 26608 20596
rect 26563 20556 26608 20584
rect 19981 20547 20039 20553
rect 26602 20544 26608 20556
rect 26660 20544 26666 20596
rect 28074 20544 28080 20596
rect 28132 20584 28138 20596
rect 28629 20587 28687 20593
rect 28629 20584 28641 20587
rect 28132 20556 28641 20584
rect 28132 20544 28138 20556
rect 28629 20553 28641 20556
rect 28675 20553 28687 20587
rect 29086 20584 29092 20596
rect 29047 20556 29092 20584
rect 28629 20547 28687 20553
rect 29086 20544 29092 20556
rect 29144 20544 29150 20596
rect 29822 20544 29828 20596
rect 29880 20584 29886 20596
rect 30009 20587 30067 20593
rect 30009 20584 30021 20587
rect 29880 20556 30021 20584
rect 29880 20544 29886 20556
rect 30009 20553 30021 20556
rect 30055 20553 30067 20587
rect 30009 20547 30067 20553
rect 33229 20587 33287 20593
rect 33229 20553 33241 20587
rect 33275 20584 33287 20587
rect 34330 20584 34336 20596
rect 33275 20556 34336 20584
rect 33275 20553 33287 20556
rect 33229 20547 33287 20553
rect 34330 20544 34336 20556
rect 34388 20544 34394 20596
rect 34422 20544 34428 20596
rect 34480 20584 34486 20596
rect 34609 20587 34667 20593
rect 34609 20584 34621 20587
rect 34480 20556 34621 20584
rect 34480 20544 34486 20556
rect 34609 20553 34621 20556
rect 34655 20553 34667 20587
rect 34609 20547 34667 20553
rect 9122 20476 9128 20528
rect 9180 20516 9186 20528
rect 9493 20519 9551 20525
rect 9493 20516 9505 20519
rect 9180 20488 9505 20516
rect 9180 20476 9186 20488
rect 9493 20485 9505 20488
rect 9539 20516 9551 20519
rect 9539 20488 11652 20516
rect 9539 20485 9551 20488
rect 9493 20479 9551 20485
rect 9677 20383 9735 20389
rect 9677 20349 9689 20383
rect 9723 20380 9735 20383
rect 10042 20380 10048 20392
rect 9723 20352 10048 20380
rect 9723 20349 9735 20352
rect 9677 20343 9735 20349
rect 10042 20340 10048 20352
rect 10100 20340 10106 20392
rect 11624 20389 11652 20488
rect 23382 20476 23388 20528
rect 23440 20516 23446 20528
rect 24486 20516 24492 20528
rect 23440 20488 24492 20516
rect 23440 20476 23446 20488
rect 15010 20408 15016 20460
rect 15068 20448 15074 20460
rect 16209 20451 16267 20457
rect 16209 20448 16221 20451
rect 15068 20420 16221 20448
rect 15068 20408 15074 20420
rect 16209 20417 16221 20420
rect 16255 20448 16267 20451
rect 16390 20448 16396 20460
rect 16255 20420 16396 20448
rect 16255 20417 16267 20420
rect 16209 20411 16267 20417
rect 16390 20408 16396 20420
rect 16448 20408 16454 20460
rect 22373 20451 22431 20457
rect 22373 20417 22385 20451
rect 22419 20448 22431 20451
rect 23014 20448 23020 20460
rect 22419 20420 23020 20448
rect 22419 20417 22431 20420
rect 22373 20411 22431 20417
rect 23014 20408 23020 20420
rect 23072 20408 23078 20460
rect 23474 20408 23480 20460
rect 23532 20448 23538 20460
rect 24320 20457 24348 20488
rect 24486 20476 24492 20488
rect 24544 20516 24550 20528
rect 25685 20519 25743 20525
rect 25685 20516 25697 20519
rect 24544 20488 25697 20516
rect 24544 20476 24550 20488
rect 25685 20485 25697 20488
rect 25731 20485 25743 20519
rect 25685 20479 25743 20485
rect 24121 20451 24179 20457
rect 24121 20448 24133 20451
rect 23532 20420 24133 20448
rect 23532 20408 23538 20420
rect 24121 20417 24133 20420
rect 24167 20417 24179 20451
rect 24121 20411 24179 20417
rect 24305 20451 24363 20457
rect 24305 20417 24317 20451
rect 24351 20417 24363 20451
rect 24946 20448 24952 20460
rect 24907 20420 24952 20448
rect 24305 20411 24363 20417
rect 24946 20408 24952 20420
rect 25004 20408 25010 20460
rect 25130 20448 25136 20460
rect 25043 20420 25136 20448
rect 25130 20408 25136 20420
rect 25188 20448 25194 20460
rect 26142 20448 26148 20460
rect 25188 20420 25452 20448
rect 25188 20408 25194 20420
rect 11609 20383 11667 20389
rect 11609 20349 11621 20383
rect 11655 20380 11667 20383
rect 11885 20383 11943 20389
rect 11885 20380 11897 20383
rect 11655 20352 11897 20380
rect 11655 20349 11667 20352
rect 11609 20343 11667 20349
rect 11885 20349 11897 20352
rect 11931 20349 11943 20383
rect 11885 20343 11943 20349
rect 13173 20383 13231 20389
rect 13173 20349 13185 20383
rect 13219 20349 13231 20383
rect 13173 20343 13231 20349
rect 13188 20312 13216 20343
rect 13262 20340 13268 20392
rect 13320 20380 13326 20392
rect 13440 20383 13498 20389
rect 13440 20380 13452 20383
rect 13320 20352 13452 20380
rect 13320 20340 13326 20352
rect 13440 20349 13452 20352
rect 13486 20380 13498 20383
rect 13722 20380 13728 20392
rect 13486 20352 13728 20380
rect 13486 20349 13498 20352
rect 13440 20343 13498 20349
rect 13722 20340 13728 20352
rect 13780 20340 13786 20392
rect 18046 20380 18052 20392
rect 18007 20352 18052 20380
rect 18046 20340 18052 20352
rect 18104 20340 18110 20392
rect 20901 20383 20959 20389
rect 20901 20349 20913 20383
rect 20947 20380 20959 20383
rect 21269 20383 21327 20389
rect 21269 20380 21281 20383
rect 20947 20352 21281 20380
rect 20947 20349 20959 20352
rect 20901 20343 20959 20349
rect 21269 20349 21281 20352
rect 21315 20380 21327 20383
rect 22094 20380 22100 20392
rect 21315 20352 22100 20380
rect 21315 20349 21327 20352
rect 21269 20343 21327 20349
rect 22094 20340 22100 20352
rect 22152 20340 22158 20392
rect 23385 20383 23443 20389
rect 23385 20349 23397 20383
rect 23431 20380 23443 20383
rect 24857 20383 24915 20389
rect 24857 20380 24869 20383
rect 23431 20352 24869 20380
rect 23431 20349 23443 20352
rect 23385 20343 23443 20349
rect 24857 20349 24869 20352
rect 24903 20380 24915 20383
rect 25314 20380 25320 20392
rect 24903 20352 25320 20380
rect 24903 20349 24915 20352
rect 24857 20343 24915 20349
rect 25314 20340 25320 20352
rect 25372 20340 25378 20392
rect 13998 20312 14004 20324
rect 13188 20284 14004 20312
rect 13998 20272 14004 20284
rect 14056 20272 14062 20324
rect 18322 20321 18328 20324
rect 15565 20315 15623 20321
rect 15565 20312 15577 20315
rect 14568 20284 15577 20312
rect 11425 20247 11483 20253
rect 11425 20213 11437 20247
rect 11471 20244 11483 20247
rect 12250 20244 12256 20256
rect 11471 20216 12256 20244
rect 11471 20213 11483 20216
rect 11425 20207 11483 20213
rect 12250 20204 12256 20216
rect 12308 20244 12314 20256
rect 12618 20244 12624 20256
rect 12308 20216 12624 20244
rect 12308 20204 12314 20216
rect 12618 20204 12624 20216
rect 12676 20204 12682 20256
rect 13722 20204 13728 20256
rect 13780 20244 13786 20256
rect 14568 20253 14596 20284
rect 15565 20281 15577 20284
rect 15611 20312 15623 20315
rect 16117 20315 16175 20321
rect 16117 20312 16129 20315
rect 15611 20284 16129 20312
rect 15611 20281 15623 20284
rect 15565 20275 15623 20281
rect 16117 20281 16129 20284
rect 16163 20281 16175 20315
rect 16117 20275 16175 20281
rect 17497 20315 17555 20321
rect 17497 20281 17509 20315
rect 17543 20312 17555 20315
rect 17865 20315 17923 20321
rect 17865 20312 17877 20315
rect 17543 20284 17877 20312
rect 17543 20281 17555 20284
rect 17497 20275 17555 20281
rect 17865 20281 17877 20284
rect 17911 20312 17923 20315
rect 18316 20312 18328 20321
rect 17911 20284 18328 20312
rect 17911 20281 17923 20284
rect 17865 20275 17923 20281
rect 18316 20275 18328 20284
rect 18322 20272 18328 20275
rect 18380 20272 18386 20324
rect 22189 20315 22247 20321
rect 22189 20312 22201 20315
rect 21560 20284 22201 20312
rect 14553 20247 14611 20253
rect 14553 20244 14565 20247
rect 13780 20216 14565 20244
rect 13780 20204 13786 20216
rect 14553 20213 14565 20216
rect 14599 20213 14611 20247
rect 14553 20207 14611 20213
rect 15746 20204 15752 20256
rect 15804 20244 15810 20256
rect 16025 20247 16083 20253
rect 16025 20244 16037 20247
rect 15804 20216 16037 20244
rect 15804 20204 15810 20216
rect 16025 20213 16037 20216
rect 16071 20213 16083 20247
rect 16025 20207 16083 20213
rect 21450 20204 21456 20256
rect 21508 20244 21514 20256
rect 21560 20253 21588 20284
rect 22189 20281 22201 20284
rect 22235 20281 22247 20315
rect 22189 20275 22247 20281
rect 23109 20315 23167 20321
rect 23109 20281 23121 20315
rect 23155 20312 23167 20315
rect 24029 20315 24087 20321
rect 24029 20312 24041 20315
rect 23155 20284 24041 20312
rect 23155 20281 23167 20284
rect 23109 20275 23167 20281
rect 24029 20281 24041 20284
rect 24075 20312 24087 20315
rect 25424 20312 25452 20420
rect 25516 20420 26148 20448
rect 25516 20389 25544 20420
rect 26142 20408 26148 20420
rect 26200 20408 26206 20460
rect 29549 20451 29607 20457
rect 29549 20417 29561 20451
rect 29595 20448 29607 20451
rect 29840 20448 29868 20544
rect 33870 20476 33876 20528
rect 33928 20516 33934 20528
rect 34146 20516 34152 20528
rect 33928 20488 34152 20516
rect 33928 20476 33934 20488
rect 34146 20476 34152 20488
rect 34204 20516 34210 20528
rect 34241 20519 34299 20525
rect 34241 20516 34253 20519
rect 34204 20488 34253 20516
rect 34204 20476 34210 20488
rect 34241 20485 34253 20488
rect 34287 20485 34299 20519
rect 34241 20479 34299 20485
rect 30558 20448 30564 20460
rect 29595 20420 29868 20448
rect 30519 20420 30564 20448
rect 29595 20417 29607 20420
rect 29549 20411 29607 20417
rect 30558 20408 30564 20420
rect 30616 20408 30622 20460
rect 33318 20408 33324 20460
rect 33376 20448 33382 20460
rect 33781 20451 33839 20457
rect 33781 20448 33793 20451
rect 33376 20420 33793 20448
rect 33376 20408 33382 20420
rect 33781 20417 33793 20420
rect 33827 20417 33839 20451
rect 33781 20411 33839 20417
rect 25501 20383 25559 20389
rect 25501 20349 25513 20383
rect 25547 20349 25559 20383
rect 25501 20343 25559 20349
rect 26697 20383 26755 20389
rect 26697 20349 26709 20383
rect 26743 20380 26755 20383
rect 26743 20352 27660 20380
rect 26743 20349 26755 20352
rect 26697 20343 26755 20349
rect 27632 20324 27660 20352
rect 33410 20340 33416 20392
rect 33468 20380 33474 20392
rect 33597 20383 33655 20389
rect 33597 20380 33609 20383
rect 33468 20352 33609 20380
rect 33468 20340 33474 20352
rect 33597 20349 33609 20352
rect 33643 20380 33655 20383
rect 34238 20380 34244 20392
rect 33643 20352 34244 20380
rect 33643 20349 33655 20352
rect 33597 20343 33655 20349
rect 34238 20340 34244 20352
rect 34296 20340 34302 20392
rect 34977 20383 35035 20389
rect 34977 20349 34989 20383
rect 35023 20349 35035 20383
rect 34977 20343 35035 20349
rect 25866 20312 25872 20324
rect 24075 20284 24532 20312
rect 25424 20284 25872 20312
rect 24075 20281 24087 20284
rect 24029 20275 24087 20281
rect 21545 20247 21603 20253
rect 21545 20244 21557 20247
rect 21508 20216 21557 20244
rect 21508 20204 21514 20216
rect 21545 20213 21557 20216
rect 21591 20213 21603 20247
rect 21545 20207 21603 20213
rect 21729 20247 21787 20253
rect 21729 20213 21741 20247
rect 21775 20244 21787 20247
rect 21910 20244 21916 20256
rect 21775 20216 21916 20244
rect 21775 20213 21787 20216
rect 21729 20207 21787 20213
rect 21910 20204 21916 20216
rect 21968 20204 21974 20256
rect 22094 20204 22100 20256
rect 22152 20244 22158 20256
rect 23658 20244 23664 20256
rect 22152 20216 22197 20244
rect 23619 20216 23664 20244
rect 22152 20204 22158 20216
rect 23658 20204 23664 20216
rect 23716 20204 23722 20256
rect 24504 20253 24532 20284
rect 25866 20272 25872 20284
rect 25924 20312 25930 20324
rect 26326 20312 26332 20324
rect 25924 20284 26332 20312
rect 25924 20272 25930 20284
rect 26326 20272 26332 20284
rect 26384 20272 26390 20324
rect 26964 20315 27022 20321
rect 26964 20281 26976 20315
rect 27010 20312 27022 20315
rect 27154 20312 27160 20324
rect 27010 20284 27160 20312
rect 27010 20281 27022 20284
rect 26964 20275 27022 20281
rect 27154 20272 27160 20284
rect 27212 20272 27218 20324
rect 27614 20272 27620 20324
rect 27672 20272 27678 20324
rect 30469 20315 30527 20321
rect 30469 20281 30481 20315
rect 30515 20312 30527 20315
rect 30806 20315 30864 20321
rect 30806 20312 30818 20315
rect 30515 20284 30818 20312
rect 30515 20281 30527 20284
rect 30469 20275 30527 20281
rect 30806 20281 30818 20284
rect 30852 20312 30864 20315
rect 30926 20312 30932 20324
rect 30852 20284 30932 20312
rect 30852 20281 30864 20284
rect 30806 20275 30864 20281
rect 30926 20272 30932 20284
rect 30984 20272 30990 20324
rect 33137 20315 33195 20321
rect 33137 20281 33149 20315
rect 33183 20312 33195 20315
rect 33689 20315 33747 20321
rect 33689 20312 33701 20315
rect 33183 20284 33701 20312
rect 33183 20281 33195 20284
rect 33137 20275 33195 20281
rect 33689 20281 33701 20284
rect 33735 20312 33747 20315
rect 34606 20312 34612 20324
rect 33735 20284 34612 20312
rect 33735 20281 33747 20284
rect 33689 20275 33747 20281
rect 34606 20272 34612 20284
rect 34664 20272 34670 20324
rect 24489 20247 24547 20253
rect 24489 20213 24501 20247
rect 24535 20213 24547 20247
rect 28074 20244 28080 20256
rect 28035 20216 28080 20244
rect 24489 20207 24547 20213
rect 28074 20204 28080 20216
rect 28132 20204 28138 20256
rect 31938 20244 31944 20256
rect 31899 20216 31944 20244
rect 31938 20204 31944 20216
rect 31996 20204 32002 20256
rect 34992 20244 35020 20343
rect 35066 20340 35072 20392
rect 35124 20380 35130 20392
rect 35244 20383 35302 20389
rect 35244 20380 35256 20383
rect 35124 20352 35256 20380
rect 35124 20340 35130 20352
rect 35244 20349 35256 20352
rect 35290 20380 35302 20383
rect 35802 20380 35808 20392
rect 35290 20352 35808 20380
rect 35290 20349 35302 20352
rect 35244 20343 35302 20349
rect 35802 20340 35808 20352
rect 35860 20340 35866 20392
rect 35802 20244 35808 20256
rect 34992 20216 35808 20244
rect 35802 20204 35808 20216
rect 35860 20204 35866 20256
rect 36170 20204 36176 20256
rect 36228 20244 36234 20256
rect 36357 20247 36415 20253
rect 36357 20244 36369 20247
rect 36228 20216 36369 20244
rect 36228 20204 36234 20216
rect 36357 20213 36369 20216
rect 36403 20213 36415 20247
rect 36357 20207 36415 20213
rect 1104 20154 38824 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 38824 20154
rect 1104 20080 38824 20102
rect 2774 20040 2780 20052
rect 2735 20012 2780 20040
rect 2774 20000 2780 20012
rect 2832 20000 2838 20052
rect 12434 20000 12440 20052
rect 12492 20040 12498 20052
rect 12713 20043 12771 20049
rect 12713 20040 12725 20043
rect 12492 20012 12725 20040
rect 12492 20000 12498 20012
rect 12713 20009 12725 20012
rect 12759 20009 12771 20043
rect 13262 20040 13268 20052
rect 13223 20012 13268 20040
rect 12713 20003 12771 20009
rect 13262 20000 13268 20012
rect 13320 20000 13326 20052
rect 13446 20000 13452 20052
rect 13504 20040 13510 20052
rect 13541 20043 13599 20049
rect 13541 20040 13553 20043
rect 13504 20012 13553 20040
rect 13504 20000 13510 20012
rect 13541 20009 13553 20012
rect 13587 20040 13599 20043
rect 13998 20040 14004 20052
rect 13587 20012 14004 20040
rect 13587 20009 13599 20012
rect 13541 20003 13599 20009
rect 13998 20000 14004 20012
rect 14056 20000 14062 20052
rect 15010 20040 15016 20052
rect 14971 20012 15016 20040
rect 15010 20000 15016 20012
rect 15068 20000 15074 20052
rect 15746 20040 15752 20052
rect 15707 20012 15752 20040
rect 15746 20000 15752 20012
rect 15804 20000 15810 20052
rect 17954 20000 17960 20052
rect 18012 20040 18018 20052
rect 18417 20043 18475 20049
rect 18417 20040 18429 20043
rect 18012 20012 18429 20040
rect 18012 20000 18018 20012
rect 18417 20009 18429 20012
rect 18463 20009 18475 20043
rect 18417 20003 18475 20009
rect 21269 20043 21327 20049
rect 21269 20009 21281 20043
rect 21315 20040 21327 20043
rect 21726 20040 21732 20052
rect 21315 20012 21732 20040
rect 21315 20009 21327 20012
rect 21269 20003 21327 20009
rect 1578 19932 1584 19984
rect 1636 19981 1642 19984
rect 1636 19975 1700 19981
rect 1636 19941 1654 19975
rect 1688 19941 1700 19975
rect 1636 19935 1700 19941
rect 1636 19932 1642 19935
rect 1397 19907 1455 19913
rect 1397 19873 1409 19907
rect 1443 19904 1455 19907
rect 1946 19904 1952 19916
rect 1443 19876 1952 19904
rect 1443 19873 1455 19876
rect 1397 19867 1455 19873
rect 1946 19864 1952 19876
rect 2004 19864 2010 19916
rect 12618 19864 12624 19916
rect 12676 19904 12682 19916
rect 13538 19904 13544 19916
rect 12676 19876 13544 19904
rect 12676 19864 12682 19876
rect 13538 19864 13544 19876
rect 13596 19904 13602 19916
rect 13725 19907 13783 19913
rect 13725 19904 13737 19907
rect 13596 19876 13737 19904
rect 13596 19864 13602 19876
rect 13725 19873 13737 19876
rect 13771 19873 13783 19907
rect 14016 19904 14044 20000
rect 16666 19972 16672 19984
rect 15948 19944 16672 19972
rect 15948 19913 15976 19944
rect 16666 19932 16672 19944
rect 16724 19932 16730 19984
rect 16206 19913 16212 19916
rect 15933 19907 15991 19913
rect 15933 19904 15945 19907
rect 14016 19876 15945 19904
rect 13725 19867 13783 19873
rect 15933 19873 15945 19876
rect 15979 19873 15991 19907
rect 16200 19904 16212 19913
rect 16167 19876 16212 19904
rect 15933 19867 15991 19873
rect 16200 19867 16212 19876
rect 16206 19864 16212 19867
rect 16264 19864 16270 19916
rect 18782 19904 18788 19916
rect 18743 19876 18788 19904
rect 18782 19864 18788 19876
rect 18840 19864 18846 19916
rect 21376 19913 21404 20012
rect 21726 20000 21732 20012
rect 21784 20000 21790 20052
rect 22094 20000 22100 20052
rect 22152 20040 22158 20052
rect 22741 20043 22799 20049
rect 22741 20040 22753 20043
rect 22152 20012 22753 20040
rect 22152 20000 22158 20012
rect 22741 20009 22753 20012
rect 22787 20009 22799 20043
rect 23382 20040 23388 20052
rect 23343 20012 23388 20040
rect 22741 20003 22799 20009
rect 23382 20000 23388 20012
rect 23440 20000 23446 20052
rect 23474 20000 23480 20052
rect 23532 20040 23538 20052
rect 23661 20043 23719 20049
rect 23661 20040 23673 20043
rect 23532 20012 23673 20040
rect 23532 20000 23538 20012
rect 23661 20009 23673 20012
rect 23707 20009 23719 20043
rect 23661 20003 23719 20009
rect 24765 20043 24823 20049
rect 24765 20009 24777 20043
rect 24811 20040 24823 20043
rect 24946 20040 24952 20052
rect 24811 20012 24952 20040
rect 24811 20009 24823 20012
rect 24765 20003 24823 20009
rect 24946 20000 24952 20012
rect 25004 20000 25010 20052
rect 25317 20043 25375 20049
rect 25317 20009 25329 20043
rect 25363 20040 25375 20043
rect 25406 20040 25412 20052
rect 25363 20012 25412 20040
rect 25363 20009 25375 20012
rect 25317 20003 25375 20009
rect 25406 20000 25412 20012
rect 25464 20000 25470 20052
rect 26329 20043 26387 20049
rect 26329 20009 26341 20043
rect 26375 20040 26387 20043
rect 26970 20040 26976 20052
rect 26375 20012 26976 20040
rect 26375 20009 26387 20012
rect 26329 20003 26387 20009
rect 26970 20000 26976 20012
rect 27028 20000 27034 20052
rect 27246 20000 27252 20052
rect 27304 20040 27310 20052
rect 27433 20043 27491 20049
rect 27433 20040 27445 20043
rect 27304 20012 27445 20040
rect 27304 20000 27310 20012
rect 27433 20009 27445 20012
rect 27479 20009 27491 20043
rect 27433 20003 27491 20009
rect 29454 20000 29460 20052
rect 29512 20040 29518 20052
rect 29825 20043 29883 20049
rect 29825 20040 29837 20043
rect 29512 20012 29837 20040
rect 29512 20000 29518 20012
rect 29825 20009 29837 20012
rect 29871 20009 29883 20043
rect 30374 20040 30380 20052
rect 30335 20012 30380 20040
rect 29825 20003 29883 20009
rect 30374 20000 30380 20012
rect 30432 20000 30438 20052
rect 33321 20043 33379 20049
rect 33321 20009 33333 20043
rect 33367 20040 33379 20043
rect 33410 20040 33416 20052
rect 33367 20012 33416 20040
rect 33367 20009 33379 20012
rect 33321 20003 33379 20009
rect 33410 20000 33416 20012
rect 33468 20000 33474 20052
rect 33597 20043 33655 20049
rect 33597 20009 33609 20043
rect 33643 20040 33655 20043
rect 35621 20043 35679 20049
rect 35621 20040 35633 20043
rect 33643 20012 35633 20040
rect 33643 20009 33655 20012
rect 33597 20003 33655 20009
rect 35621 20009 35633 20012
rect 35667 20040 35679 20043
rect 36173 20043 36231 20049
rect 36173 20040 36185 20043
rect 35667 20012 36185 20040
rect 35667 20009 35679 20012
rect 35621 20003 35679 20009
rect 36173 20009 36185 20012
rect 36219 20009 36231 20043
rect 36173 20003 36231 20009
rect 27157 19975 27215 19981
rect 27157 19941 27169 19975
rect 27203 19972 27215 19975
rect 28074 19972 28080 19984
rect 27203 19944 28080 19972
rect 27203 19941 27215 19944
rect 27157 19935 27215 19941
rect 28074 19932 28080 19944
rect 28132 19981 28138 19984
rect 28132 19975 28196 19981
rect 28132 19941 28150 19975
rect 28184 19941 28196 19975
rect 28132 19935 28196 19941
rect 28132 19932 28138 19935
rect 30190 19932 30196 19984
rect 30248 19972 30254 19984
rect 31389 19975 31447 19981
rect 31389 19972 31401 19975
rect 30248 19944 31401 19972
rect 30248 19932 30254 19944
rect 21361 19907 21419 19913
rect 21361 19873 21373 19907
rect 21407 19873 21419 19907
rect 21361 19867 21419 19873
rect 21450 19864 21456 19916
rect 21508 19904 21514 19916
rect 21617 19907 21675 19913
rect 21617 19904 21629 19907
rect 21508 19876 21629 19904
rect 21508 19864 21514 19876
rect 21617 19873 21629 19876
rect 21663 19873 21675 19907
rect 21617 19867 21675 19873
rect 25225 19907 25283 19913
rect 25225 19873 25237 19907
rect 25271 19904 25283 19907
rect 25314 19904 25320 19916
rect 25271 19876 25320 19904
rect 25271 19873 25283 19876
rect 25225 19867 25283 19873
rect 25314 19864 25320 19876
rect 25372 19864 25378 19916
rect 26513 19907 26571 19913
rect 26513 19873 26525 19907
rect 26559 19904 26571 19907
rect 26602 19904 26608 19916
rect 26559 19876 26608 19904
rect 26559 19873 26571 19876
rect 26513 19867 26571 19873
rect 26602 19864 26608 19876
rect 26660 19864 26666 19916
rect 27614 19864 27620 19916
rect 27672 19904 27678 19916
rect 27893 19907 27951 19913
rect 27893 19904 27905 19907
rect 27672 19876 27905 19904
rect 27672 19864 27678 19876
rect 27893 19873 27905 19876
rect 27939 19904 27951 19907
rect 28718 19904 28724 19916
rect 27939 19876 28724 19904
rect 27939 19873 27951 19876
rect 27893 19867 27951 19873
rect 28718 19864 28724 19876
rect 28776 19864 28782 19916
rect 30742 19904 30748 19916
rect 30703 19876 30748 19904
rect 30742 19864 30748 19876
rect 30800 19864 30806 19916
rect 17862 19836 17868 19848
rect 17328 19808 17868 19836
rect 17328 19777 17356 19808
rect 17862 19796 17868 19808
rect 17920 19836 17926 19848
rect 18877 19839 18935 19845
rect 18877 19836 18889 19839
rect 17920 19808 18889 19836
rect 17920 19796 17926 19808
rect 18877 19805 18889 19808
rect 18923 19805 18935 19839
rect 18877 19799 18935 19805
rect 18969 19839 19027 19845
rect 18969 19805 18981 19839
rect 19015 19805 19027 19839
rect 23842 19836 23848 19848
rect 23803 19808 23848 19836
rect 18969 19799 19027 19805
rect 17313 19771 17371 19777
rect 17313 19737 17325 19771
rect 17359 19737 17371 19771
rect 18984 19768 19012 19799
rect 23842 19796 23848 19808
rect 23900 19796 23906 19848
rect 25501 19839 25559 19845
rect 25501 19805 25513 19839
rect 25547 19836 25559 19839
rect 26142 19836 26148 19848
rect 25547 19808 26148 19836
rect 25547 19805 25559 19808
rect 25501 19799 25559 19805
rect 17313 19731 17371 19737
rect 18248 19740 19012 19768
rect 18248 19712 18276 19740
rect 24762 19728 24768 19780
rect 24820 19768 24826 19780
rect 25516 19768 25544 19799
rect 26142 19796 26148 19808
rect 26200 19796 26206 19848
rect 29086 19796 29092 19848
rect 29144 19836 29150 19848
rect 31036 19845 31064 19944
rect 31389 19941 31401 19944
rect 31435 19941 31447 19975
rect 31389 19935 31447 19941
rect 33965 19975 34023 19981
rect 33965 19941 33977 19975
rect 34011 19972 34023 19975
rect 34054 19972 34060 19984
rect 34011 19944 34060 19972
rect 34011 19941 34023 19944
rect 33965 19935 34023 19941
rect 34054 19932 34060 19944
rect 34112 19972 34118 19984
rect 34422 19972 34428 19984
rect 34112 19944 34428 19972
rect 34112 19932 34118 19944
rect 34422 19932 34428 19944
rect 34480 19932 34486 19984
rect 35066 19972 35072 19984
rect 35027 19944 35072 19972
rect 35066 19932 35072 19944
rect 35124 19932 35130 19984
rect 35526 19904 35532 19916
rect 35487 19876 35532 19904
rect 35526 19864 35532 19876
rect 35584 19864 35590 19916
rect 30285 19839 30343 19845
rect 30285 19836 30297 19839
rect 29144 19808 30297 19836
rect 29144 19796 29150 19808
rect 30285 19805 30297 19808
rect 30331 19836 30343 19839
rect 30837 19839 30895 19845
rect 30837 19836 30849 19839
rect 30331 19808 30849 19836
rect 30331 19805 30343 19808
rect 30285 19799 30343 19805
rect 30837 19805 30849 19808
rect 30883 19805 30895 19839
rect 30837 19799 30895 19805
rect 31021 19839 31079 19845
rect 31021 19805 31033 19839
rect 31067 19836 31079 19839
rect 31938 19836 31944 19848
rect 31067 19808 31944 19836
rect 31067 19805 31079 19808
rect 31021 19799 31079 19805
rect 31938 19796 31944 19808
rect 31996 19796 32002 19848
rect 33778 19796 33784 19848
rect 33836 19836 33842 19848
rect 34057 19839 34115 19845
rect 34057 19836 34069 19839
rect 33836 19808 34069 19836
rect 33836 19796 33842 19808
rect 34057 19805 34069 19808
rect 34103 19805 34115 19839
rect 34238 19836 34244 19848
rect 34199 19808 34244 19836
rect 34057 19799 34115 19805
rect 34238 19796 34244 19808
rect 34296 19796 34302 19848
rect 35710 19836 35716 19848
rect 35671 19808 35716 19836
rect 35710 19796 35716 19808
rect 35768 19796 35774 19848
rect 24820 19740 25544 19768
rect 24820 19728 24826 19740
rect 34606 19728 34612 19780
rect 34664 19768 34670 19780
rect 34701 19771 34759 19777
rect 34701 19768 34713 19771
rect 34664 19740 34713 19768
rect 34664 19728 34670 19740
rect 34701 19737 34713 19740
rect 34747 19768 34759 19771
rect 35250 19768 35256 19780
rect 34747 19740 35256 19768
rect 34747 19737 34759 19740
rect 34701 19731 34759 19737
rect 35250 19728 35256 19740
rect 35308 19728 35314 19780
rect 17954 19700 17960 19712
rect 17915 19672 17960 19700
rect 17954 19660 17960 19672
rect 18012 19700 18018 19712
rect 18230 19700 18236 19712
rect 18012 19672 18236 19700
rect 18012 19660 18018 19672
rect 18230 19660 18236 19672
rect 18288 19660 18294 19712
rect 24210 19660 24216 19712
rect 24268 19700 24274 19712
rect 24305 19703 24363 19709
rect 24305 19700 24317 19703
rect 24268 19672 24317 19700
rect 24268 19660 24274 19672
rect 24305 19669 24317 19672
rect 24351 19669 24363 19703
rect 24305 19663 24363 19669
rect 24857 19703 24915 19709
rect 24857 19669 24869 19703
rect 24903 19700 24915 19703
rect 25774 19700 25780 19712
rect 24903 19672 25780 19700
rect 24903 19669 24915 19672
rect 24857 19663 24915 19669
rect 25774 19660 25780 19672
rect 25832 19660 25838 19712
rect 25866 19660 25872 19712
rect 25924 19700 25930 19712
rect 25924 19672 25969 19700
rect 25924 19660 25930 19672
rect 26050 19660 26056 19712
rect 26108 19700 26114 19712
rect 26697 19703 26755 19709
rect 26697 19700 26709 19703
rect 26108 19672 26709 19700
rect 26108 19660 26114 19672
rect 26697 19669 26709 19672
rect 26743 19669 26755 19703
rect 26697 19663 26755 19669
rect 28994 19660 29000 19712
rect 29052 19700 29058 19712
rect 29273 19703 29331 19709
rect 29273 19700 29285 19703
rect 29052 19672 29285 19700
rect 29052 19660 29058 19672
rect 29273 19669 29285 19672
rect 29319 19669 29331 19703
rect 29273 19663 29331 19669
rect 30926 19660 30932 19712
rect 30984 19700 30990 19712
rect 32398 19700 32404 19712
rect 30984 19672 32404 19700
rect 30984 19660 30990 19672
rect 32398 19660 32404 19672
rect 32456 19660 32462 19712
rect 35161 19703 35219 19709
rect 35161 19669 35173 19703
rect 35207 19700 35219 19703
rect 35342 19700 35348 19712
rect 35207 19672 35348 19700
rect 35207 19669 35219 19672
rect 35161 19663 35219 19669
rect 35342 19660 35348 19672
rect 35400 19660 35406 19712
rect 1104 19610 38824 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 34966 19610
rect 35018 19558 35030 19610
rect 35082 19558 35094 19610
rect 35146 19558 35158 19610
rect 35210 19558 38824 19610
rect 1104 19536 38824 19558
rect 1578 19496 1584 19508
rect 1539 19468 1584 19496
rect 1578 19456 1584 19468
rect 1636 19456 1642 19508
rect 1946 19496 1952 19508
rect 1907 19468 1952 19496
rect 1946 19456 1952 19468
rect 2004 19456 2010 19508
rect 14826 19496 14832 19508
rect 14739 19468 14832 19496
rect 14826 19456 14832 19468
rect 14884 19496 14890 19508
rect 15746 19496 15752 19508
rect 14884 19468 15752 19496
rect 14884 19456 14890 19468
rect 15746 19456 15752 19468
rect 15804 19456 15810 19508
rect 17862 19496 17868 19508
rect 17823 19468 17868 19496
rect 17862 19456 17868 19468
rect 17920 19456 17926 19508
rect 18322 19456 18328 19508
rect 18380 19496 18386 19508
rect 19429 19499 19487 19505
rect 19429 19496 19441 19499
rect 18380 19468 19441 19496
rect 18380 19456 18386 19468
rect 19429 19465 19441 19468
rect 19475 19465 19487 19499
rect 19429 19459 19487 19465
rect 24854 19456 24860 19508
rect 24912 19496 24918 19508
rect 25406 19496 25412 19508
rect 24912 19468 25412 19496
rect 24912 19456 24918 19468
rect 25406 19456 25412 19468
rect 25464 19496 25470 19508
rect 25593 19499 25651 19505
rect 25593 19496 25605 19499
rect 25464 19468 25605 19496
rect 25464 19456 25470 19468
rect 25593 19465 25605 19468
rect 25639 19465 25651 19499
rect 26050 19496 26056 19508
rect 26011 19468 26056 19496
rect 25593 19459 25651 19465
rect 26050 19456 26056 19468
rect 26108 19456 26114 19508
rect 26602 19496 26608 19508
rect 26563 19468 26608 19496
rect 26602 19456 26608 19468
rect 26660 19456 26666 19508
rect 28074 19496 28080 19508
rect 28035 19468 28080 19496
rect 28074 19456 28080 19468
rect 28132 19456 28138 19508
rect 34054 19496 34060 19508
rect 34015 19468 34060 19496
rect 34054 19456 34060 19468
rect 34112 19456 34118 19508
rect 35802 19496 35808 19508
rect 35084 19468 35808 19496
rect 12989 19363 13047 19369
rect 12989 19329 13001 19363
rect 13035 19360 13047 19363
rect 13446 19360 13452 19372
rect 13035 19332 13452 19360
rect 13035 19329 13047 19332
rect 12989 19323 13047 19329
rect 13446 19320 13452 19332
rect 13504 19320 13510 19372
rect 16390 19320 16396 19372
rect 16448 19360 16454 19372
rect 16485 19363 16543 19369
rect 16485 19360 16497 19363
rect 16448 19332 16497 19360
rect 16448 19320 16454 19332
rect 16485 19329 16497 19332
rect 16531 19360 16543 19363
rect 17954 19360 17960 19372
rect 16531 19332 17080 19360
rect 16531 19329 16543 19332
rect 16485 19323 16543 19329
rect 13722 19301 13728 19304
rect 13716 19292 13728 19301
rect 13648 19264 13728 19292
rect 13357 19227 13415 19233
rect 13357 19193 13369 19227
rect 13403 19224 13415 19227
rect 13648 19224 13676 19264
rect 13716 19255 13728 19264
rect 13722 19252 13728 19255
rect 13780 19252 13786 19304
rect 15473 19295 15531 19301
rect 15473 19261 15485 19295
rect 15519 19292 15531 19295
rect 16206 19292 16212 19304
rect 15519 19264 16212 19292
rect 15519 19261 15531 19264
rect 15473 19255 15531 19261
rect 16206 19252 16212 19264
rect 16264 19292 16270 19304
rect 16301 19295 16359 19301
rect 16301 19292 16313 19295
rect 16264 19264 16313 19292
rect 16264 19252 16270 19264
rect 16301 19261 16313 19264
rect 16347 19292 16359 19295
rect 16945 19295 17003 19301
rect 16945 19292 16957 19295
rect 16347 19264 16957 19292
rect 16347 19261 16359 19264
rect 16301 19255 16359 19261
rect 16945 19261 16957 19264
rect 16991 19261 17003 19295
rect 17052 19292 17080 19332
rect 17880 19332 17960 19360
rect 17313 19295 17371 19301
rect 17313 19292 17325 19295
rect 17052 19264 17325 19292
rect 16945 19255 17003 19261
rect 17313 19261 17325 19264
rect 17359 19292 17371 19295
rect 17880 19292 17908 19332
rect 17954 19320 17960 19332
rect 18012 19320 18018 19372
rect 25225 19363 25283 19369
rect 25225 19329 25237 19363
rect 25271 19360 25283 19363
rect 25406 19360 25412 19372
rect 25271 19332 25412 19360
rect 25271 19329 25283 19332
rect 25225 19323 25283 19329
rect 25406 19320 25412 19332
rect 25464 19360 25470 19372
rect 26068 19360 26096 19456
rect 25464 19332 26096 19360
rect 27709 19363 27767 19369
rect 25464 19320 25470 19332
rect 27709 19329 27721 19363
rect 27755 19360 27767 19363
rect 28092 19360 28120 19456
rect 27755 19332 28120 19360
rect 27755 19329 27767 19332
rect 27709 19323 27767 19329
rect 29454 19320 29460 19372
rect 29512 19360 29518 19372
rect 30104 19363 30162 19369
rect 30104 19360 30116 19363
rect 29512 19332 30116 19360
rect 29512 19320 29518 19332
rect 30104 19329 30116 19332
rect 30150 19329 30162 19363
rect 30104 19323 30162 19329
rect 30190 19320 30196 19372
rect 30248 19360 30254 19372
rect 30558 19360 30564 19372
rect 30248 19332 30564 19360
rect 30248 19320 30254 19332
rect 30558 19320 30564 19332
rect 30616 19320 30622 19372
rect 32398 19320 32404 19372
rect 32456 19360 32462 19372
rect 35084 19369 35112 19468
rect 35802 19456 35808 19468
rect 35860 19456 35866 19508
rect 32861 19363 32919 19369
rect 32861 19360 32873 19363
rect 32456 19332 32873 19360
rect 32456 19320 32462 19332
rect 32861 19329 32873 19332
rect 32907 19329 32919 19363
rect 32861 19323 32919 19329
rect 35069 19363 35127 19369
rect 35069 19329 35081 19363
rect 35115 19329 35127 19363
rect 35069 19323 35127 19329
rect 18046 19292 18052 19304
rect 17359 19264 17908 19292
rect 18007 19264 18052 19292
rect 17359 19261 17371 19264
rect 17313 19255 17371 19261
rect 18046 19252 18052 19264
rect 18104 19252 18110 19304
rect 20533 19295 20591 19301
rect 20533 19261 20545 19295
rect 20579 19292 20591 19295
rect 20622 19292 20628 19304
rect 20579 19264 20628 19292
rect 20579 19261 20591 19264
rect 20533 19255 20591 19261
rect 20622 19252 20628 19264
rect 20680 19292 20686 19304
rect 20993 19295 21051 19301
rect 20993 19292 21005 19295
rect 20680 19264 21005 19292
rect 20680 19252 20686 19264
rect 20993 19261 21005 19264
rect 21039 19292 21051 19295
rect 21726 19292 21732 19304
rect 21039 19264 21732 19292
rect 21039 19261 21051 19264
rect 20993 19255 21051 19261
rect 21726 19252 21732 19264
rect 21784 19292 21790 19304
rect 22925 19295 22983 19301
rect 22925 19292 22937 19295
rect 21784 19264 22937 19292
rect 21784 19252 21790 19264
rect 22925 19261 22937 19264
rect 22971 19261 22983 19295
rect 22925 19255 22983 19261
rect 23477 19295 23535 19301
rect 23477 19261 23489 19295
rect 23523 19292 23535 19295
rect 24762 19292 24768 19304
rect 23523 19264 24768 19292
rect 23523 19261 23535 19264
rect 23477 19255 23535 19261
rect 24762 19252 24768 19264
rect 24820 19252 24826 19304
rect 26510 19252 26516 19304
rect 26568 19292 26574 19304
rect 27525 19295 27583 19301
rect 27525 19292 27537 19295
rect 26568 19264 27537 19292
rect 26568 19252 26574 19264
rect 27525 19261 27537 19264
rect 27571 19292 27583 19295
rect 27798 19292 27804 19304
rect 27571 19264 27804 19292
rect 27571 19261 27583 19264
rect 27525 19255 27583 19261
rect 27798 19252 27804 19264
rect 27856 19252 27862 19304
rect 29641 19295 29699 19301
rect 29641 19292 29653 19295
rect 28644 19264 29653 19292
rect 15838 19224 15844 19236
rect 13403 19196 13676 19224
rect 15751 19196 15844 19224
rect 13403 19193 13415 19196
rect 13357 19187 13415 19193
rect 15838 19184 15844 19196
rect 15896 19224 15902 19236
rect 16393 19227 16451 19233
rect 16393 19224 16405 19227
rect 15896 19196 16405 19224
rect 15896 19184 15902 19196
rect 16393 19193 16405 19196
rect 16439 19193 16451 19227
rect 16393 19187 16451 19193
rect 18138 19184 18144 19236
rect 18196 19224 18202 19236
rect 18316 19227 18374 19233
rect 18316 19224 18328 19227
rect 18196 19196 18328 19224
rect 18196 19184 18202 19196
rect 18316 19193 18328 19196
rect 18362 19224 18374 19227
rect 18782 19224 18788 19236
rect 18362 19196 18788 19224
rect 18362 19193 18374 19196
rect 18316 19187 18374 19193
rect 18782 19184 18788 19196
rect 18840 19224 18846 19236
rect 18840 19196 20024 19224
rect 18840 19184 18846 19196
rect 19996 19168 20024 19196
rect 20162 19184 20168 19236
rect 20220 19224 20226 19236
rect 20809 19227 20867 19233
rect 20809 19224 20821 19227
rect 20220 19196 20821 19224
rect 20220 19184 20226 19196
rect 20809 19193 20821 19196
rect 20855 19224 20867 19227
rect 21238 19227 21296 19233
rect 21238 19224 21250 19227
rect 20855 19196 21250 19224
rect 20855 19193 20867 19196
rect 20809 19187 20867 19193
rect 21238 19193 21250 19196
rect 21284 19193 21296 19227
rect 25041 19227 25099 19233
rect 25041 19224 25053 19227
rect 21238 19187 21296 19193
rect 24412 19196 25053 19224
rect 15933 19159 15991 19165
rect 15933 19125 15945 19159
rect 15979 19156 15991 19159
rect 16482 19156 16488 19168
rect 15979 19128 16488 19156
rect 15979 19125 15991 19128
rect 15933 19119 15991 19125
rect 16482 19116 16488 19128
rect 16540 19116 16546 19168
rect 19978 19156 19984 19168
rect 19939 19128 19984 19156
rect 19978 19116 19984 19128
rect 20036 19116 20042 19168
rect 21450 19116 21456 19168
rect 21508 19156 21514 19168
rect 22373 19159 22431 19165
rect 22373 19156 22385 19159
rect 21508 19128 22385 19156
rect 21508 19116 21514 19128
rect 22373 19125 22385 19128
rect 22419 19125 22431 19159
rect 24118 19156 24124 19168
rect 24079 19128 24124 19156
rect 22373 19119 22431 19125
rect 24118 19116 24124 19128
rect 24176 19116 24182 19168
rect 24302 19116 24308 19168
rect 24360 19156 24366 19168
rect 24412 19165 24440 19196
rect 25041 19193 25053 19196
rect 25087 19193 25099 19227
rect 26878 19224 26884 19236
rect 26839 19196 26884 19224
rect 25041 19187 25099 19193
rect 26878 19184 26884 19196
rect 26936 19224 26942 19236
rect 27433 19227 27491 19233
rect 27433 19224 27445 19227
rect 26936 19196 27445 19224
rect 26936 19184 26942 19196
rect 27433 19193 27445 19196
rect 27479 19193 27491 19227
rect 27433 19187 27491 19193
rect 28644 19168 28672 19264
rect 29641 19261 29653 19264
rect 29687 19261 29699 19295
rect 30377 19295 30435 19301
rect 30377 19292 30389 19295
rect 29641 19255 29699 19261
rect 29748 19264 30389 19292
rect 29089 19227 29147 19233
rect 29089 19193 29101 19227
rect 29135 19224 29147 19227
rect 29748 19224 29776 19264
rect 30377 19261 30389 19264
rect 30423 19292 30435 19295
rect 30742 19292 30748 19304
rect 30423 19264 30748 19292
rect 30423 19261 30435 19264
rect 30377 19255 30435 19261
rect 30742 19252 30748 19264
rect 30800 19292 30806 19304
rect 31757 19295 31815 19301
rect 31757 19292 31769 19295
rect 30800 19264 31769 19292
rect 30800 19252 30806 19264
rect 31757 19261 31769 19264
rect 31803 19292 31815 19295
rect 33042 19292 33048 19304
rect 31803 19264 33048 19292
rect 31803 19261 31815 19264
rect 31757 19255 31815 19261
rect 33042 19252 33048 19264
rect 33100 19252 33106 19304
rect 35336 19295 35394 19301
rect 35336 19292 35348 19295
rect 35176 19264 35348 19292
rect 29135 19196 29776 19224
rect 29135 19193 29147 19196
rect 29089 19187 29147 19193
rect 32122 19184 32128 19236
rect 32180 19224 32186 19236
rect 32217 19227 32275 19233
rect 32217 19224 32229 19227
rect 32180 19196 32229 19224
rect 32180 19184 32186 19196
rect 32217 19193 32229 19196
rect 32263 19224 32275 19227
rect 32677 19227 32735 19233
rect 32677 19224 32689 19227
rect 32263 19196 32689 19224
rect 32263 19193 32275 19196
rect 32217 19187 32275 19193
rect 32677 19193 32689 19196
rect 32723 19193 32735 19227
rect 32677 19187 32735 19193
rect 34238 19184 34244 19236
rect 34296 19224 34302 19236
rect 35176 19224 35204 19264
rect 35336 19261 35348 19264
rect 35382 19292 35394 19295
rect 36170 19292 36176 19304
rect 35382 19264 36176 19292
rect 35382 19261 35394 19264
rect 35336 19255 35394 19261
rect 36170 19252 36176 19264
rect 36228 19252 36234 19304
rect 34296 19196 35204 19224
rect 34296 19184 34302 19196
rect 35802 19184 35808 19236
rect 35860 19224 35866 19236
rect 37001 19227 37059 19233
rect 37001 19224 37013 19227
rect 35860 19196 37013 19224
rect 35860 19184 35866 19196
rect 37001 19193 37013 19196
rect 37047 19193 37059 19227
rect 37001 19187 37059 19193
rect 24397 19159 24455 19165
rect 24397 19156 24409 19159
rect 24360 19128 24409 19156
rect 24360 19116 24366 19128
rect 24397 19125 24409 19128
rect 24443 19125 24455 19159
rect 24578 19156 24584 19168
rect 24539 19128 24584 19156
rect 24397 19119 24455 19125
rect 24578 19116 24584 19128
rect 24636 19116 24642 19168
rect 24670 19116 24676 19168
rect 24728 19156 24734 19168
rect 24949 19159 25007 19165
rect 24949 19156 24961 19159
rect 24728 19128 24961 19156
rect 24728 19116 24734 19128
rect 24949 19125 24961 19128
rect 24995 19125 25007 19159
rect 24949 19119 25007 19125
rect 27065 19159 27123 19165
rect 27065 19125 27077 19159
rect 27111 19156 27123 19159
rect 28350 19156 28356 19168
rect 27111 19128 28356 19156
rect 27111 19125 27123 19128
rect 27065 19119 27123 19125
rect 28350 19116 28356 19128
rect 28408 19116 28414 19168
rect 28626 19156 28632 19168
rect 28587 19128 28632 19156
rect 28626 19116 28632 19128
rect 28684 19116 28690 19168
rect 29362 19116 29368 19168
rect 29420 19156 29426 19168
rect 29457 19159 29515 19165
rect 29457 19156 29469 19159
rect 29420 19128 29469 19156
rect 29420 19116 29426 19128
rect 29457 19125 29469 19128
rect 29503 19156 29515 19159
rect 30107 19159 30165 19165
rect 30107 19156 30119 19159
rect 29503 19128 30119 19156
rect 29503 19125 29515 19128
rect 29457 19119 29515 19125
rect 30107 19125 30119 19128
rect 30153 19156 30165 19159
rect 30374 19156 30380 19168
rect 30153 19128 30380 19156
rect 30153 19125 30165 19128
rect 30107 19119 30165 19125
rect 30374 19116 30380 19128
rect 30432 19116 30438 19168
rect 31294 19116 31300 19168
rect 31352 19156 31358 19168
rect 31481 19159 31539 19165
rect 31481 19156 31493 19159
rect 31352 19128 31493 19156
rect 31352 19116 31358 19128
rect 31481 19125 31493 19128
rect 31527 19125 31539 19159
rect 32306 19156 32312 19168
rect 32267 19128 32312 19156
rect 31481 19119 31539 19125
rect 32306 19116 32312 19128
rect 32364 19116 32370 19168
rect 32766 19156 32772 19168
rect 32727 19128 32772 19156
rect 32766 19116 32772 19128
rect 32824 19116 32830 19168
rect 33689 19159 33747 19165
rect 33689 19125 33701 19159
rect 33735 19156 33747 19159
rect 33778 19156 33784 19168
rect 33735 19128 33784 19156
rect 33735 19125 33747 19128
rect 33689 19119 33747 19125
rect 33778 19116 33784 19128
rect 33836 19156 33842 19168
rect 33962 19156 33968 19168
rect 33836 19128 33968 19156
rect 33836 19116 33842 19128
rect 33962 19116 33968 19128
rect 34020 19116 34026 19168
rect 34701 19159 34759 19165
rect 34701 19125 34713 19159
rect 34747 19156 34759 19159
rect 35526 19156 35532 19168
rect 34747 19128 35532 19156
rect 34747 19125 34759 19128
rect 34701 19119 34759 19125
rect 35526 19116 35532 19128
rect 35584 19116 35590 19168
rect 35710 19116 35716 19168
rect 35768 19156 35774 19168
rect 36449 19159 36507 19165
rect 36449 19156 36461 19159
rect 35768 19128 36461 19156
rect 35768 19116 35774 19128
rect 36449 19125 36461 19128
rect 36495 19125 36507 19159
rect 36449 19119 36507 19125
rect 1104 19066 38824 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 38824 19066
rect 1104 18992 38824 19014
rect 13538 18952 13544 18964
rect 13499 18924 13544 18952
rect 13538 18912 13544 18924
rect 13596 18912 13602 18964
rect 16206 18912 16212 18964
rect 16264 18952 16270 18964
rect 16669 18955 16727 18961
rect 16669 18952 16681 18955
rect 16264 18924 16681 18952
rect 16264 18912 16270 18924
rect 16669 18921 16681 18924
rect 16715 18921 16727 18955
rect 18138 18952 18144 18964
rect 18099 18924 18144 18952
rect 16669 18915 16727 18921
rect 18138 18912 18144 18924
rect 18196 18912 18202 18964
rect 20530 18952 20536 18964
rect 20491 18924 20536 18952
rect 20530 18912 20536 18924
rect 20588 18912 20594 18964
rect 21450 18952 21456 18964
rect 21411 18924 21456 18952
rect 21450 18912 21456 18924
rect 21508 18912 21514 18964
rect 23937 18955 23995 18961
rect 23937 18921 23949 18955
rect 23983 18952 23995 18955
rect 24670 18952 24676 18964
rect 23983 18924 24676 18952
rect 23983 18921 23995 18924
rect 23937 18915 23995 18921
rect 24670 18912 24676 18924
rect 24728 18912 24734 18964
rect 24854 18952 24860 18964
rect 24815 18924 24860 18952
rect 24854 18912 24860 18924
rect 24912 18912 24918 18964
rect 25317 18955 25375 18961
rect 25317 18921 25329 18955
rect 25363 18952 25375 18955
rect 25498 18952 25504 18964
rect 25363 18924 25504 18952
rect 25363 18921 25375 18924
rect 25317 18915 25375 18921
rect 25498 18912 25504 18924
rect 25556 18952 25562 18964
rect 27065 18955 27123 18961
rect 27065 18952 27077 18955
rect 25556 18924 27077 18952
rect 25556 18912 25562 18924
rect 27065 18921 27077 18924
rect 27111 18921 27123 18955
rect 27798 18952 27804 18964
rect 27759 18924 27804 18952
rect 27065 18915 27123 18921
rect 27798 18912 27804 18924
rect 27856 18912 27862 18964
rect 28350 18952 28356 18964
rect 28263 18924 28356 18952
rect 28350 18912 28356 18924
rect 28408 18952 28414 18964
rect 28718 18952 28724 18964
rect 28408 18924 28724 18952
rect 28408 18912 28414 18924
rect 28718 18912 28724 18924
rect 28776 18952 28782 18964
rect 29086 18952 29092 18964
rect 28776 18924 29092 18952
rect 28776 18912 28782 18924
rect 29086 18912 29092 18924
rect 29144 18912 29150 18964
rect 30926 18952 30932 18964
rect 30887 18924 30932 18952
rect 30926 18912 30932 18924
rect 30984 18912 30990 18964
rect 32122 18952 32128 18964
rect 32083 18924 32128 18952
rect 32122 18912 32128 18924
rect 32180 18912 32186 18964
rect 33505 18955 33563 18961
rect 33505 18921 33517 18955
rect 33551 18952 33563 18955
rect 34238 18952 34244 18964
rect 33551 18924 34244 18952
rect 33551 18921 33563 18924
rect 33505 18915 33563 18921
rect 34238 18912 34244 18924
rect 34296 18912 34302 18964
rect 35250 18912 35256 18964
rect 35308 18952 35314 18964
rect 35437 18955 35495 18961
rect 35437 18952 35449 18955
rect 35308 18924 35449 18952
rect 35308 18912 35314 18924
rect 35437 18921 35449 18924
rect 35483 18921 35495 18955
rect 35437 18915 35495 18921
rect 35526 18912 35532 18964
rect 35584 18952 35590 18964
rect 36265 18955 36323 18961
rect 36265 18952 36277 18955
rect 35584 18924 36277 18952
rect 35584 18912 35590 18924
rect 36265 18921 36277 18924
rect 36311 18921 36323 18955
rect 36265 18915 36323 18921
rect 15556 18887 15614 18893
rect 15556 18853 15568 18887
rect 15602 18884 15614 18887
rect 15838 18884 15844 18896
rect 15602 18856 15844 18884
rect 15602 18853 15614 18856
rect 15556 18847 15614 18853
rect 15838 18844 15844 18856
rect 15896 18844 15902 18896
rect 22094 18844 22100 18896
rect 22152 18884 22158 18896
rect 22152 18856 22324 18884
rect 22152 18844 22158 18856
rect 18414 18816 18420 18828
rect 18375 18788 18420 18816
rect 18414 18776 18420 18788
rect 18472 18776 18478 18828
rect 22296 18825 22324 18856
rect 25590 18844 25596 18896
rect 25648 18884 25654 18896
rect 25958 18884 25964 18896
rect 25648 18856 25964 18884
rect 25648 18844 25654 18856
rect 25958 18844 25964 18856
rect 26016 18844 26022 18896
rect 28810 18844 28816 18896
rect 28868 18884 28874 18896
rect 28997 18887 29055 18893
rect 28997 18884 29009 18887
rect 28868 18856 29009 18884
rect 28868 18844 28874 18856
rect 28997 18853 29009 18856
rect 29043 18853 29055 18887
rect 28997 18847 29055 18853
rect 29457 18887 29515 18893
rect 29457 18853 29469 18887
rect 29503 18884 29515 18887
rect 29794 18887 29852 18893
rect 29794 18884 29806 18887
rect 29503 18856 29806 18884
rect 29503 18853 29515 18856
rect 29457 18847 29515 18853
rect 29794 18853 29806 18856
rect 29840 18884 29852 18887
rect 30282 18884 30288 18896
rect 29840 18856 30288 18884
rect 29840 18853 29852 18856
rect 29794 18847 29852 18853
rect 30282 18844 30288 18856
rect 30340 18844 30346 18896
rect 36170 18884 36176 18896
rect 36131 18856 36176 18884
rect 36170 18844 36176 18856
rect 36228 18844 36234 18896
rect 21821 18819 21879 18825
rect 21821 18785 21833 18819
rect 21867 18816 21879 18819
rect 22281 18819 22339 18825
rect 21867 18788 22232 18816
rect 21867 18785 21879 18788
rect 21821 18779 21879 18785
rect 13998 18708 14004 18760
rect 14056 18748 14062 18760
rect 15289 18751 15347 18757
rect 15289 18748 15301 18751
rect 14056 18720 15301 18748
rect 14056 18708 14062 18720
rect 15289 18717 15301 18720
rect 15335 18717 15347 18751
rect 15289 18711 15347 18717
rect 20070 18708 20076 18760
rect 20128 18748 20134 18760
rect 20165 18751 20223 18757
rect 20165 18748 20177 18751
rect 20128 18720 20177 18748
rect 20128 18708 20134 18720
rect 20165 18717 20177 18720
rect 20211 18748 20223 18751
rect 20254 18748 20260 18760
rect 20211 18720 20260 18748
rect 20211 18717 20223 18720
rect 20165 18711 20223 18717
rect 20254 18708 20260 18720
rect 20312 18708 20318 18760
rect 22204 18680 22232 18788
rect 22281 18785 22293 18819
rect 22327 18816 22339 18819
rect 22922 18816 22928 18828
rect 22327 18788 22928 18816
rect 22327 18785 22339 18788
rect 22281 18779 22339 18785
rect 22922 18776 22928 18788
rect 22980 18776 22986 18828
rect 23658 18776 23664 18828
rect 23716 18816 23722 18828
rect 23753 18819 23811 18825
rect 23753 18816 23765 18819
rect 23716 18788 23765 18816
rect 23716 18776 23722 18788
rect 23753 18785 23765 18788
rect 23799 18785 23811 18819
rect 25222 18816 25228 18828
rect 25183 18788 25228 18816
rect 23753 18779 23811 18785
rect 25222 18776 25228 18788
rect 25280 18776 25286 18828
rect 25774 18776 25780 18828
rect 25832 18816 25838 18828
rect 26513 18819 26571 18825
rect 26513 18816 26525 18819
rect 25832 18788 26525 18816
rect 25832 18776 25838 18788
rect 26513 18785 26525 18788
rect 26559 18785 26571 18819
rect 26878 18816 26884 18828
rect 26839 18788 26884 18816
rect 26513 18779 26571 18785
rect 26878 18776 26884 18788
rect 26936 18816 26942 18828
rect 27433 18819 27491 18825
rect 27433 18816 27445 18819
rect 26936 18788 27445 18816
rect 26936 18776 26942 18788
rect 27433 18785 27445 18788
rect 27479 18785 27491 18819
rect 30190 18816 30196 18828
rect 27433 18779 27491 18785
rect 29564 18788 30196 18816
rect 22370 18748 22376 18760
rect 22331 18720 22376 18748
rect 22370 18708 22376 18720
rect 22428 18708 22434 18760
rect 22557 18751 22615 18757
rect 22557 18748 22569 18751
rect 22480 18720 22569 18748
rect 22480 18680 22508 18720
rect 22557 18717 22569 18720
rect 22603 18748 22615 18751
rect 24486 18748 24492 18760
rect 22603 18720 24492 18748
rect 22603 18717 22615 18720
rect 22557 18711 22615 18717
rect 24486 18708 24492 18720
rect 24544 18708 24550 18760
rect 25406 18748 25412 18760
rect 25367 18720 25412 18748
rect 25406 18708 25412 18720
rect 25464 18708 25470 18760
rect 28442 18748 28448 18760
rect 28403 18720 28448 18748
rect 28442 18708 28448 18720
rect 28500 18708 28506 18760
rect 28629 18751 28687 18757
rect 28629 18717 28641 18751
rect 28675 18748 28687 18751
rect 28902 18748 28908 18760
rect 28675 18720 28908 18748
rect 28675 18717 28687 18720
rect 28629 18711 28687 18717
rect 28902 18708 28908 18720
rect 28960 18708 28966 18760
rect 29086 18708 29092 18760
rect 29144 18748 29150 18760
rect 29564 18757 29592 18788
rect 30190 18776 30196 18788
rect 30248 18776 30254 18828
rect 33597 18819 33655 18825
rect 33597 18785 33609 18819
rect 33643 18816 33655 18819
rect 33686 18816 33692 18828
rect 33643 18788 33692 18816
rect 33643 18785 33655 18788
rect 33597 18779 33655 18785
rect 29549 18751 29607 18757
rect 29549 18748 29561 18751
rect 29144 18720 29561 18748
rect 29144 18708 29150 18720
rect 29549 18717 29561 18720
rect 29595 18717 29607 18751
rect 33612 18748 33640 18779
rect 33686 18776 33692 18788
rect 33744 18776 33750 18828
rect 33870 18776 33876 18828
rect 33928 18825 33934 18828
rect 33928 18819 33978 18825
rect 33928 18785 33932 18819
rect 33966 18785 33978 18819
rect 33928 18779 33978 18785
rect 33928 18776 33934 18779
rect 34054 18748 34060 18760
rect 29549 18711 29607 18717
rect 31496 18720 33640 18748
rect 34018 18720 34060 18748
rect 22204 18652 22508 18680
rect 26697 18683 26755 18689
rect 26697 18649 26709 18683
rect 26743 18680 26755 18683
rect 26970 18680 26976 18692
rect 26743 18652 26976 18680
rect 26743 18649 26755 18652
rect 26697 18643 26755 18649
rect 26970 18640 26976 18652
rect 27028 18640 27034 18692
rect 30558 18640 30564 18692
rect 30616 18680 30622 18692
rect 31496 18689 31524 18720
rect 34054 18708 34060 18720
rect 34112 18708 34118 18760
rect 34330 18748 34336 18760
rect 34291 18720 34336 18748
rect 34330 18708 34336 18720
rect 34388 18708 34394 18760
rect 31481 18683 31539 18689
rect 31481 18680 31493 18683
rect 30616 18652 31493 18680
rect 30616 18640 30622 18652
rect 31481 18649 31493 18652
rect 31527 18649 31539 18683
rect 31481 18643 31539 18649
rect 16298 18572 16304 18624
rect 16356 18612 16362 18624
rect 17681 18615 17739 18621
rect 17681 18612 17693 18615
rect 16356 18584 17693 18612
rect 16356 18572 16362 18584
rect 17681 18581 17693 18584
rect 17727 18612 17739 18615
rect 18046 18612 18052 18624
rect 17727 18584 18052 18612
rect 17727 18581 17739 18584
rect 17681 18575 17739 18581
rect 18046 18572 18052 18584
rect 18104 18572 18110 18624
rect 21913 18615 21971 18621
rect 21913 18581 21925 18615
rect 21959 18612 21971 18615
rect 23382 18612 23388 18624
rect 21959 18584 23388 18612
rect 21959 18581 21971 18584
rect 21913 18575 21971 18581
rect 23382 18572 23388 18584
rect 23440 18572 23446 18624
rect 27985 18615 28043 18621
rect 27985 18581 27997 18615
rect 28031 18612 28043 18615
rect 28810 18612 28816 18624
rect 28031 18584 28816 18612
rect 28031 18581 28043 18584
rect 27985 18575 28043 18581
rect 28810 18572 28816 18584
rect 28868 18572 28874 18624
rect 32122 18572 32128 18624
rect 32180 18612 32186 18624
rect 32585 18615 32643 18621
rect 32585 18612 32597 18615
rect 32180 18584 32597 18612
rect 32180 18572 32186 18584
rect 32585 18581 32597 18584
rect 32631 18612 32643 18615
rect 32766 18612 32772 18624
rect 32631 18584 32772 18612
rect 32631 18581 32643 18584
rect 32585 18575 32643 18581
rect 32766 18572 32772 18584
rect 32824 18572 32830 18624
rect 35710 18612 35716 18624
rect 35671 18584 35716 18612
rect 35710 18572 35716 18584
rect 35768 18572 35774 18624
rect 1104 18522 38824 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 34966 18522
rect 35018 18470 35030 18522
rect 35082 18470 35094 18522
rect 35146 18470 35158 18522
rect 35210 18470 38824 18522
rect 1104 18448 38824 18470
rect 15381 18411 15439 18417
rect 15381 18377 15393 18411
rect 15427 18408 15439 18411
rect 15838 18408 15844 18420
rect 15427 18380 15844 18408
rect 15427 18377 15439 18380
rect 15381 18371 15439 18377
rect 15838 18368 15844 18380
rect 15896 18408 15902 18420
rect 15933 18411 15991 18417
rect 15933 18408 15945 18411
rect 15896 18380 15945 18408
rect 15896 18368 15902 18380
rect 15933 18377 15945 18380
rect 15979 18377 15991 18411
rect 17862 18408 17868 18420
rect 17823 18380 17868 18408
rect 15933 18371 15991 18377
rect 17862 18368 17868 18380
rect 17920 18368 17926 18420
rect 19797 18411 19855 18417
rect 19797 18377 19809 18411
rect 19843 18408 19855 18411
rect 22370 18408 22376 18420
rect 19843 18380 22376 18408
rect 19843 18377 19855 18380
rect 19797 18371 19855 18377
rect 22370 18368 22376 18380
rect 22428 18408 22434 18420
rect 22557 18411 22615 18417
rect 22557 18408 22569 18411
rect 22428 18380 22569 18408
rect 22428 18368 22434 18380
rect 22557 18377 22569 18380
rect 22603 18377 22615 18411
rect 22922 18408 22928 18420
rect 22883 18380 22928 18408
rect 22557 18371 22615 18377
rect 22922 18368 22928 18380
rect 22980 18368 22986 18420
rect 23477 18411 23535 18417
rect 23477 18377 23489 18411
rect 23523 18408 23535 18411
rect 23658 18408 23664 18420
rect 23523 18380 23664 18408
rect 23523 18377 23535 18380
rect 23477 18371 23535 18377
rect 23658 18368 23664 18380
rect 23716 18368 23722 18420
rect 24394 18408 24400 18420
rect 24355 18380 24400 18408
rect 24394 18368 24400 18380
rect 24452 18368 24458 18420
rect 25498 18408 25504 18420
rect 25459 18380 25504 18408
rect 25498 18368 25504 18380
rect 25556 18368 25562 18420
rect 25774 18408 25780 18420
rect 25735 18380 25780 18408
rect 25774 18368 25780 18380
rect 25832 18368 25838 18420
rect 28442 18408 28448 18420
rect 28403 18380 28448 18408
rect 28442 18368 28448 18380
rect 28500 18368 28506 18420
rect 28718 18408 28724 18420
rect 28679 18380 28724 18408
rect 28718 18368 28724 18380
rect 28776 18368 28782 18420
rect 30374 18408 30380 18420
rect 30335 18380 30380 18408
rect 30374 18368 30380 18380
rect 30432 18368 30438 18420
rect 35802 18408 35808 18420
rect 33796 18380 35808 18408
rect 13909 18275 13967 18281
rect 13909 18241 13921 18275
rect 13955 18272 13967 18275
rect 17880 18272 17908 18368
rect 19429 18343 19487 18349
rect 19429 18309 19441 18343
rect 19475 18340 19487 18343
rect 19978 18340 19984 18352
rect 19475 18312 19984 18340
rect 19475 18309 19487 18312
rect 19429 18303 19487 18309
rect 19978 18300 19984 18312
rect 20036 18300 20042 18352
rect 20530 18340 20536 18352
rect 20456 18312 20536 18340
rect 20456 18281 20484 18312
rect 20530 18300 20536 18312
rect 20588 18300 20594 18352
rect 23842 18300 23848 18352
rect 23900 18340 23906 18352
rect 24305 18343 24363 18349
rect 24305 18340 24317 18343
rect 23900 18312 24317 18340
rect 23900 18300 23906 18312
rect 24305 18309 24317 18312
rect 24351 18340 24363 18343
rect 25222 18340 25228 18352
rect 24351 18312 25228 18340
rect 24351 18309 24363 18312
rect 24305 18303 24363 18309
rect 25222 18300 25228 18312
rect 25280 18300 25286 18352
rect 27985 18343 28043 18349
rect 27985 18309 27997 18343
rect 28031 18340 28043 18343
rect 30009 18343 30067 18349
rect 30009 18340 30021 18343
rect 28031 18312 30021 18340
rect 28031 18309 28043 18312
rect 27985 18303 28043 18309
rect 30009 18309 30021 18312
rect 30055 18309 30067 18343
rect 30009 18303 30067 18309
rect 20441 18275 20499 18281
rect 13955 18244 14136 18272
rect 17880 18244 18184 18272
rect 13955 18241 13967 18244
rect 13909 18235 13967 18241
rect 13446 18164 13452 18216
rect 13504 18204 13510 18216
rect 13998 18204 14004 18216
rect 13504 18176 14004 18204
rect 13504 18164 13510 18176
rect 13998 18164 14004 18176
rect 14056 18164 14062 18216
rect 14108 18204 14136 18244
rect 14268 18207 14326 18213
rect 14268 18204 14280 18207
rect 14108 18176 14280 18204
rect 14268 18173 14280 18176
rect 14314 18204 14326 18207
rect 14826 18204 14832 18216
rect 14314 18176 14832 18204
rect 14314 18173 14326 18176
rect 14268 18167 14326 18173
rect 14826 18164 14832 18176
rect 14884 18164 14890 18216
rect 18046 18204 18052 18216
rect 18007 18176 18052 18204
rect 18046 18164 18052 18176
rect 18104 18164 18110 18216
rect 18156 18204 18184 18244
rect 20441 18241 20453 18275
rect 20487 18241 20499 18275
rect 20622 18272 20628 18284
rect 20583 18244 20628 18272
rect 20441 18235 20499 18241
rect 20622 18232 20628 18244
rect 20680 18232 20686 18284
rect 24486 18232 24492 18284
rect 24544 18272 24550 18284
rect 24949 18275 25007 18281
rect 24949 18272 24961 18275
rect 24544 18244 24961 18272
rect 24544 18232 24550 18244
rect 24949 18241 24961 18244
rect 24995 18241 25007 18275
rect 24949 18235 25007 18241
rect 27709 18275 27767 18281
rect 27709 18241 27721 18275
rect 27755 18272 27767 18275
rect 28626 18272 28632 18284
rect 27755 18244 28632 18272
rect 27755 18241 27767 18244
rect 27709 18235 27767 18241
rect 28626 18232 28632 18244
rect 28684 18232 28690 18284
rect 30024 18272 30052 18303
rect 33796 18281 33824 18380
rect 35802 18368 35808 18380
rect 35860 18408 35866 18420
rect 36449 18411 36507 18417
rect 36449 18408 36461 18411
rect 35860 18380 36461 18408
rect 35860 18368 35866 18380
rect 36449 18377 36461 18380
rect 36495 18377 36507 18411
rect 36449 18371 36507 18377
rect 33870 18300 33876 18352
rect 33928 18340 33934 18352
rect 34241 18343 34299 18349
rect 34241 18340 34253 18343
rect 33928 18312 34253 18340
rect 33928 18300 33934 18312
rect 34241 18309 34253 18312
rect 34287 18309 34299 18343
rect 34241 18303 34299 18309
rect 31024 18275 31082 18281
rect 31024 18272 31036 18275
rect 30024 18244 31036 18272
rect 31024 18241 31036 18244
rect 31070 18272 31082 18275
rect 32769 18275 32827 18281
rect 31070 18244 31708 18272
rect 31070 18241 31082 18244
rect 31024 18235 31082 18241
rect 18305 18207 18363 18213
rect 18305 18204 18317 18207
rect 18156 18176 18317 18204
rect 18305 18173 18317 18176
rect 18351 18173 18363 18207
rect 25958 18204 25964 18216
rect 25919 18176 25964 18204
rect 18305 18167 18363 18173
rect 25958 18164 25964 18176
rect 26016 18164 26022 18216
rect 27798 18204 27804 18216
rect 27759 18176 27804 18204
rect 27798 18164 27804 18176
rect 27856 18164 27862 18216
rect 28644 18204 28672 18232
rect 30558 18204 30564 18216
rect 28644 18176 30564 18204
rect 30558 18164 30564 18176
rect 30616 18164 30622 18216
rect 30884 18207 30942 18213
rect 30884 18204 30896 18207
rect 30668 18176 30896 18204
rect 20257 18139 20315 18145
rect 20257 18105 20269 18139
rect 20303 18136 20315 18139
rect 20714 18136 20720 18148
rect 20303 18108 20720 18136
rect 20303 18105 20315 18108
rect 20257 18099 20315 18105
rect 20714 18096 20720 18108
rect 20772 18136 20778 18148
rect 20870 18139 20928 18145
rect 20870 18136 20882 18139
rect 20772 18108 20882 18136
rect 20772 18096 20778 18108
rect 20870 18105 20882 18108
rect 20916 18105 20928 18139
rect 20870 18099 20928 18105
rect 23937 18139 23995 18145
rect 23937 18105 23949 18139
rect 23983 18136 23995 18139
rect 24854 18136 24860 18148
rect 23983 18108 24860 18136
rect 23983 18105 23995 18108
rect 23937 18099 23995 18105
rect 24854 18096 24860 18108
rect 24912 18096 24918 18148
rect 30374 18096 30380 18148
rect 30432 18136 30438 18148
rect 30668 18136 30696 18176
rect 30884 18173 30896 18176
rect 30930 18173 30942 18207
rect 31294 18204 31300 18216
rect 31255 18176 31300 18204
rect 30884 18167 30942 18173
rect 31294 18164 31300 18176
rect 31352 18164 31358 18216
rect 31680 18204 31708 18244
rect 32769 18241 32781 18275
rect 32815 18272 32827 18275
rect 33781 18275 33839 18281
rect 33781 18272 33793 18275
rect 32815 18244 33793 18272
rect 32815 18241 32827 18244
rect 32769 18235 32827 18241
rect 33781 18241 33793 18244
rect 33827 18241 33839 18275
rect 33781 18235 33839 18241
rect 31754 18204 31760 18216
rect 31680 18176 31760 18204
rect 31754 18164 31760 18176
rect 31812 18164 31818 18216
rect 33137 18207 33195 18213
rect 33137 18173 33149 18207
rect 33183 18204 33195 18207
rect 33594 18204 33600 18216
rect 33183 18176 33600 18204
rect 33183 18173 33195 18176
rect 33137 18167 33195 18173
rect 33594 18164 33600 18176
rect 33652 18204 33658 18216
rect 34330 18204 34336 18216
rect 33652 18176 34336 18204
rect 33652 18164 33658 18176
rect 34330 18164 34336 18176
rect 34388 18164 34394 18216
rect 35069 18207 35127 18213
rect 35069 18173 35081 18207
rect 35115 18204 35127 18207
rect 35894 18204 35900 18216
rect 35115 18176 35900 18204
rect 35115 18173 35127 18176
rect 35069 18167 35127 18173
rect 35894 18164 35900 18176
rect 35952 18164 35958 18216
rect 30432 18108 30696 18136
rect 30432 18096 30438 18108
rect 33410 18096 33416 18148
rect 33468 18136 33474 18148
rect 33689 18139 33747 18145
rect 33689 18136 33701 18139
rect 33468 18108 33701 18136
rect 33468 18096 33474 18108
rect 33689 18105 33701 18108
rect 33735 18105 33747 18139
rect 33689 18099 33747 18105
rect 34701 18139 34759 18145
rect 34701 18105 34713 18139
rect 34747 18136 34759 18139
rect 35314 18139 35372 18145
rect 35314 18136 35326 18139
rect 34747 18108 35326 18136
rect 34747 18105 34759 18108
rect 34701 18099 34759 18105
rect 35314 18105 35326 18108
rect 35360 18136 35372 18139
rect 35710 18136 35716 18148
rect 35360 18108 35716 18136
rect 35360 18105 35372 18108
rect 35314 18099 35372 18105
rect 35710 18096 35716 18108
rect 35768 18096 35774 18148
rect 16298 18068 16304 18080
rect 16259 18040 16304 18068
rect 16298 18028 16304 18040
rect 16356 18028 16362 18080
rect 20162 18068 20168 18080
rect 20123 18040 20168 18068
rect 20162 18028 20168 18040
rect 20220 18068 20226 18080
rect 22005 18071 22063 18077
rect 22005 18068 22017 18071
rect 20220 18040 22017 18068
rect 20220 18028 20226 18040
rect 22005 18037 22017 18040
rect 22051 18037 22063 18071
rect 24762 18068 24768 18080
rect 24723 18040 24768 18068
rect 22005 18031 22063 18037
rect 24762 18028 24768 18040
rect 24820 18028 24826 18080
rect 29546 18068 29552 18080
rect 29507 18040 29552 18068
rect 29546 18028 29552 18040
rect 29604 18028 29610 18080
rect 32401 18071 32459 18077
rect 32401 18037 32413 18071
rect 32447 18068 32459 18071
rect 32582 18068 32588 18080
rect 32447 18040 32588 18068
rect 32447 18037 32459 18040
rect 32401 18031 32459 18037
rect 32582 18028 32588 18040
rect 32640 18028 32646 18080
rect 33226 18068 33232 18080
rect 33187 18040 33232 18068
rect 33226 18028 33232 18040
rect 33284 18028 33290 18080
rect 1104 17978 38824 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 38824 17978
rect 1104 17904 38824 17926
rect 13998 17864 14004 17876
rect 13959 17836 14004 17864
rect 13998 17824 14004 17836
rect 14056 17864 14062 17876
rect 15473 17867 15531 17873
rect 15473 17864 15485 17867
rect 14056 17836 15485 17864
rect 14056 17824 14062 17836
rect 15473 17833 15485 17836
rect 15519 17864 15531 17867
rect 16298 17864 16304 17876
rect 15519 17836 16304 17864
rect 15519 17833 15531 17836
rect 15473 17827 15531 17833
rect 16298 17824 16304 17836
rect 16356 17824 16362 17876
rect 18046 17864 18052 17876
rect 18007 17836 18052 17864
rect 18046 17824 18052 17836
rect 18104 17824 18110 17876
rect 20162 17864 20168 17876
rect 20123 17836 20168 17864
rect 20162 17824 20168 17836
rect 20220 17824 20226 17876
rect 20806 17824 20812 17876
rect 20864 17864 20870 17876
rect 21085 17867 21143 17873
rect 21085 17864 21097 17867
rect 20864 17836 21097 17864
rect 20864 17824 20870 17836
rect 21085 17833 21097 17836
rect 21131 17833 21143 17867
rect 21085 17827 21143 17833
rect 23569 17867 23627 17873
rect 23569 17833 23581 17867
rect 23615 17864 23627 17867
rect 24302 17864 24308 17876
rect 23615 17836 24308 17864
rect 23615 17833 23627 17836
rect 23569 17827 23627 17833
rect 24302 17824 24308 17836
rect 24360 17824 24366 17876
rect 24854 17864 24860 17876
rect 24815 17836 24860 17864
rect 24854 17824 24860 17836
rect 24912 17824 24918 17876
rect 25406 17824 25412 17876
rect 25464 17864 25470 17876
rect 25869 17867 25927 17873
rect 25869 17864 25881 17867
rect 25464 17836 25881 17864
rect 25464 17824 25470 17836
rect 25869 17833 25881 17836
rect 25915 17833 25927 17867
rect 26510 17864 26516 17876
rect 26471 17836 26516 17864
rect 25869 17827 25927 17833
rect 26510 17824 26516 17836
rect 26568 17824 26574 17876
rect 27798 17864 27804 17876
rect 27759 17836 27804 17864
rect 27798 17824 27804 17836
rect 27856 17824 27862 17876
rect 31294 17864 31300 17876
rect 31255 17836 31300 17864
rect 31294 17824 31300 17836
rect 31352 17824 31358 17876
rect 31754 17824 31760 17876
rect 31812 17864 31818 17876
rect 32490 17864 32496 17876
rect 31812 17836 32496 17864
rect 31812 17824 31818 17836
rect 32490 17824 32496 17836
rect 32548 17824 32554 17876
rect 32582 17824 32588 17876
rect 32640 17864 32646 17876
rect 33594 17864 33600 17876
rect 32640 17836 33600 17864
rect 32640 17824 32646 17836
rect 33594 17824 33600 17836
rect 33652 17824 33658 17876
rect 34054 17864 34060 17876
rect 34015 17836 34060 17864
rect 34054 17824 34060 17836
rect 34112 17864 34118 17876
rect 34425 17867 34483 17873
rect 34425 17864 34437 17867
rect 34112 17836 34437 17864
rect 34112 17824 34118 17836
rect 34425 17833 34437 17836
rect 34471 17833 34483 17867
rect 35894 17864 35900 17876
rect 35855 17836 35900 17864
rect 34425 17827 34483 17833
rect 35894 17824 35900 17836
rect 35952 17824 35958 17876
rect 19061 17799 19119 17805
rect 19061 17765 19073 17799
rect 19107 17796 19119 17799
rect 19610 17796 19616 17808
rect 19107 17768 19616 17796
rect 19107 17765 19119 17768
rect 19061 17759 19119 17765
rect 19610 17756 19616 17768
rect 19668 17796 19674 17808
rect 20530 17796 20536 17808
rect 19668 17768 20536 17796
rect 19668 17756 19674 17768
rect 20530 17756 20536 17768
rect 20588 17756 20594 17808
rect 24397 17799 24455 17805
rect 24397 17765 24409 17799
rect 24443 17796 24455 17799
rect 24762 17796 24768 17808
rect 24443 17768 24768 17796
rect 24443 17765 24455 17768
rect 24397 17759 24455 17765
rect 24762 17756 24768 17768
rect 24820 17756 24826 17808
rect 28261 17799 28319 17805
rect 28261 17765 28273 17799
rect 28307 17796 28319 17799
rect 28902 17796 28908 17808
rect 28307 17768 28908 17796
rect 28307 17765 28319 17768
rect 28261 17759 28319 17765
rect 28902 17756 28908 17768
rect 28960 17796 28966 17808
rect 29454 17796 29460 17808
rect 28960 17768 29460 17796
rect 28960 17756 28966 17768
rect 29454 17756 29460 17768
rect 29512 17805 29518 17808
rect 29512 17799 29576 17805
rect 29512 17765 29530 17799
rect 29564 17765 29576 17799
rect 29512 17759 29576 17765
rect 33321 17799 33379 17805
rect 33321 17765 33333 17799
rect 33367 17796 33379 17799
rect 33410 17796 33416 17808
rect 33367 17768 33416 17796
rect 33367 17765 33379 17768
rect 33321 17759 33379 17765
rect 29512 17756 29518 17759
rect 33410 17756 33416 17768
rect 33468 17756 33474 17808
rect 35342 17756 35348 17808
rect 35400 17796 35406 17808
rect 36262 17796 36268 17808
rect 35400 17768 36268 17796
rect 35400 17756 35406 17768
rect 36262 17756 36268 17768
rect 36320 17756 36326 17808
rect 22186 17728 22192 17740
rect 22147 17700 22192 17728
rect 22186 17688 22192 17700
rect 22244 17688 22250 17740
rect 22281 17731 22339 17737
rect 22281 17697 22293 17731
rect 22327 17728 22339 17731
rect 22462 17728 22468 17740
rect 22327 17700 22468 17728
rect 22327 17697 22339 17700
rect 22281 17691 22339 17697
rect 22462 17688 22468 17700
rect 22520 17688 22526 17740
rect 23382 17728 23388 17740
rect 23343 17700 23388 17728
rect 23382 17688 23388 17700
rect 23440 17688 23446 17740
rect 24029 17731 24087 17737
rect 24029 17697 24041 17731
rect 24075 17728 24087 17731
rect 24486 17728 24492 17740
rect 24075 17700 24492 17728
rect 24075 17697 24087 17700
rect 24029 17691 24087 17697
rect 21729 17663 21787 17669
rect 21729 17629 21741 17663
rect 21775 17660 21787 17663
rect 22373 17663 22431 17669
rect 22373 17660 22385 17663
rect 21775 17632 22385 17660
rect 21775 17629 21787 17632
rect 21729 17623 21787 17629
rect 22373 17629 22385 17632
rect 22419 17660 22431 17663
rect 24044 17660 24072 17691
rect 24486 17688 24492 17700
rect 24544 17688 24550 17740
rect 25222 17728 25228 17740
rect 25183 17700 25228 17728
rect 25222 17688 25228 17700
rect 25280 17688 25286 17740
rect 26878 17728 26884 17740
rect 26839 17700 26884 17728
rect 26878 17688 26884 17700
rect 26936 17688 26942 17740
rect 34793 17731 34851 17737
rect 34793 17697 34805 17731
rect 34839 17728 34851 17731
rect 35250 17728 35256 17740
rect 34839 17700 35256 17728
rect 34839 17697 34851 17700
rect 34793 17691 34851 17697
rect 35250 17688 35256 17700
rect 35308 17728 35314 17740
rect 35989 17731 36047 17737
rect 35989 17728 36001 17731
rect 35308 17700 36001 17728
rect 35308 17688 35314 17700
rect 35989 17697 36001 17700
rect 36035 17697 36047 17731
rect 35989 17691 36047 17697
rect 25314 17660 25320 17672
rect 22419 17632 24072 17660
rect 25275 17632 25320 17660
rect 22419 17629 22431 17632
rect 22373 17623 22431 17629
rect 25314 17620 25320 17632
rect 25372 17620 25378 17672
rect 25409 17663 25467 17669
rect 25409 17629 25421 17663
rect 25455 17629 25467 17663
rect 26970 17660 26976 17672
rect 26931 17632 26976 17660
rect 25409 17623 25467 17629
rect 19889 17595 19947 17601
rect 19889 17561 19901 17595
rect 19935 17592 19947 17595
rect 19935 17564 20760 17592
rect 19935 17561 19947 17564
rect 19889 17555 19947 17561
rect 20732 17536 20760 17564
rect 25130 17552 25136 17604
rect 25188 17592 25194 17604
rect 25424 17592 25452 17623
rect 26970 17620 26976 17632
rect 27028 17620 27034 17672
rect 27065 17663 27123 17669
rect 27065 17629 27077 17663
rect 27111 17629 27123 17663
rect 29273 17663 29331 17669
rect 29273 17660 29285 17663
rect 27065 17623 27123 17629
rect 29104 17632 29285 17660
rect 25188 17564 25452 17592
rect 25188 17552 25194 17564
rect 18414 17524 18420 17536
rect 18375 17496 18420 17524
rect 18414 17484 18420 17496
rect 18472 17484 18478 17536
rect 20714 17524 20720 17536
rect 20675 17496 20720 17524
rect 20714 17484 20720 17496
rect 20772 17484 20778 17536
rect 21818 17524 21824 17536
rect 21779 17496 21824 17524
rect 21818 17484 21824 17496
rect 21876 17484 21882 17536
rect 24765 17527 24823 17533
rect 24765 17493 24777 17527
rect 24811 17524 24823 17527
rect 24946 17524 24952 17536
rect 24811 17496 24952 17524
rect 24811 17493 24823 17496
rect 24765 17487 24823 17493
rect 24946 17484 24952 17496
rect 25004 17484 25010 17536
rect 25424 17524 25452 17564
rect 25866 17524 25872 17536
rect 25424 17496 25872 17524
rect 25866 17484 25872 17496
rect 25924 17524 25930 17536
rect 27080 17524 27108 17623
rect 29104 17536 29132 17632
rect 29273 17629 29285 17632
rect 29319 17629 29331 17663
rect 32766 17660 32772 17672
rect 32727 17632 32772 17660
rect 29273 17623 29331 17629
rect 32766 17620 32772 17632
rect 32824 17620 32830 17672
rect 34054 17620 34060 17672
rect 34112 17660 34118 17672
rect 34885 17663 34943 17669
rect 34885 17660 34897 17663
rect 34112 17632 34897 17660
rect 34112 17620 34118 17632
rect 34885 17629 34897 17632
rect 34931 17629 34943 17663
rect 34885 17623 34943 17629
rect 35069 17663 35127 17669
rect 35069 17629 35081 17663
rect 35115 17660 35127 17663
rect 35342 17660 35348 17672
rect 35115 17632 35348 17660
rect 35115 17629 35127 17632
rect 35069 17623 35127 17629
rect 35342 17620 35348 17632
rect 35400 17620 35406 17672
rect 32122 17592 32128 17604
rect 32083 17564 32128 17592
rect 32122 17552 32128 17564
rect 32180 17552 32186 17604
rect 34238 17552 34244 17604
rect 34296 17592 34302 17604
rect 34514 17592 34520 17604
rect 34296 17564 34520 17592
rect 34296 17552 34302 17564
rect 34514 17552 34520 17564
rect 34572 17552 34578 17604
rect 35618 17552 35624 17604
rect 35676 17592 35682 17604
rect 35894 17592 35900 17604
rect 35676 17564 35900 17592
rect 35676 17552 35682 17564
rect 35894 17552 35900 17564
rect 35952 17552 35958 17604
rect 27890 17524 27896 17536
rect 25924 17496 27896 17524
rect 25924 17484 25930 17496
rect 27890 17484 27896 17496
rect 27948 17484 27954 17536
rect 29086 17524 29092 17536
rect 29047 17496 29092 17524
rect 29086 17484 29092 17496
rect 29144 17484 29150 17536
rect 30466 17484 30472 17536
rect 30524 17524 30530 17536
rect 30653 17527 30711 17533
rect 30653 17524 30665 17527
rect 30524 17496 30665 17524
rect 30524 17484 30530 17496
rect 30653 17493 30665 17496
rect 30699 17493 30711 17527
rect 30653 17487 30711 17493
rect 35529 17527 35587 17533
rect 35529 17493 35541 17527
rect 35575 17524 35587 17527
rect 35710 17524 35716 17536
rect 35575 17496 35716 17524
rect 35575 17493 35587 17496
rect 35529 17487 35587 17493
rect 35710 17484 35716 17496
rect 35768 17484 35774 17536
rect 1104 17434 38824 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 34966 17434
rect 35018 17382 35030 17434
rect 35082 17382 35094 17434
rect 35146 17382 35158 17434
rect 35210 17382 38824 17434
rect 1104 17360 38824 17382
rect 18966 17320 18972 17332
rect 18927 17292 18972 17320
rect 18966 17280 18972 17292
rect 19024 17280 19030 17332
rect 20714 17280 20720 17332
rect 20772 17320 20778 17332
rect 21913 17323 21971 17329
rect 21913 17320 21925 17323
rect 20772 17292 21925 17320
rect 20772 17280 20778 17292
rect 21913 17289 21925 17292
rect 21959 17289 21971 17323
rect 21913 17283 21971 17289
rect 22186 17280 22192 17332
rect 22244 17320 22250 17332
rect 22833 17323 22891 17329
rect 22833 17320 22845 17323
rect 22244 17292 22845 17320
rect 22244 17280 22250 17292
rect 22833 17289 22845 17292
rect 22879 17289 22891 17323
rect 23382 17320 23388 17332
rect 23343 17292 23388 17320
rect 22833 17283 22891 17289
rect 23382 17280 23388 17292
rect 23440 17280 23446 17332
rect 23842 17320 23848 17332
rect 23803 17292 23848 17320
rect 23842 17280 23848 17292
rect 23900 17280 23906 17332
rect 27430 17320 27436 17332
rect 27391 17292 27436 17320
rect 27430 17280 27436 17292
rect 27488 17280 27494 17332
rect 27890 17320 27896 17332
rect 27851 17292 27896 17320
rect 27890 17280 27896 17292
rect 27948 17280 27954 17332
rect 29086 17320 29092 17332
rect 29047 17292 29092 17320
rect 29086 17280 29092 17292
rect 29144 17280 29150 17332
rect 29454 17320 29460 17332
rect 29415 17292 29460 17320
rect 29454 17280 29460 17292
rect 29512 17280 29518 17332
rect 30374 17280 30380 17332
rect 30432 17320 30438 17332
rect 31573 17323 31631 17329
rect 31573 17320 31585 17323
rect 30432 17292 31585 17320
rect 30432 17280 30438 17292
rect 31573 17289 31585 17292
rect 31619 17320 31631 17323
rect 32766 17320 32772 17332
rect 31619 17292 32772 17320
rect 31619 17289 31631 17292
rect 31573 17283 31631 17289
rect 32766 17280 32772 17292
rect 32824 17320 32830 17332
rect 32861 17323 32919 17329
rect 32861 17320 32873 17323
rect 32824 17292 32873 17320
rect 32824 17280 32830 17292
rect 32861 17289 32873 17292
rect 32907 17289 32919 17323
rect 32861 17283 32919 17289
rect 33226 17280 33232 17332
rect 33284 17320 33290 17332
rect 34054 17320 34060 17332
rect 33284 17292 34060 17320
rect 33284 17280 33290 17292
rect 34054 17280 34060 17292
rect 34112 17280 34118 17332
rect 35161 17323 35219 17329
rect 35161 17289 35173 17323
rect 35207 17320 35219 17323
rect 35250 17320 35256 17332
rect 35207 17292 35256 17320
rect 35207 17289 35219 17292
rect 35161 17283 35219 17289
rect 35250 17280 35256 17292
rect 35308 17280 35314 17332
rect 35710 17320 35716 17332
rect 35452 17292 35716 17320
rect 32490 17252 32496 17264
rect 32451 17224 32496 17252
rect 32490 17212 32496 17224
rect 32548 17212 32554 17264
rect 33686 17252 33692 17264
rect 33647 17224 33692 17252
rect 33686 17212 33692 17224
rect 33744 17212 33750 17264
rect 19610 17184 19616 17196
rect 19571 17156 19616 17184
rect 19610 17144 19616 17156
rect 19668 17184 19674 17196
rect 19886 17184 19892 17196
rect 19668 17156 19892 17184
rect 19668 17144 19674 17156
rect 19886 17144 19892 17156
rect 19944 17144 19950 17196
rect 32217 17187 32275 17193
rect 32217 17153 32229 17187
rect 32263 17184 32275 17187
rect 32582 17184 32588 17196
rect 32263 17156 32588 17184
rect 32263 17153 32275 17156
rect 32217 17147 32275 17153
rect 32582 17144 32588 17156
rect 32640 17144 32646 17196
rect 35452 17193 35480 17292
rect 35710 17280 35716 17292
rect 35768 17280 35774 17332
rect 35437 17187 35495 17193
rect 35437 17153 35449 17187
rect 35483 17153 35495 17187
rect 35437 17147 35495 17153
rect 20533 17119 20591 17125
rect 20533 17085 20545 17119
rect 20579 17116 20591 17119
rect 20622 17116 20628 17128
rect 20579 17088 20628 17116
rect 20579 17085 20591 17088
rect 20533 17079 20591 17085
rect 20622 17076 20628 17088
rect 20680 17076 20686 17128
rect 22462 17116 22468 17128
rect 22423 17088 22468 17116
rect 22462 17076 22468 17088
rect 22520 17076 22526 17128
rect 23658 17116 23664 17128
rect 23619 17088 23664 17116
rect 23658 17076 23664 17088
rect 23716 17076 23722 17128
rect 24854 17116 24860 17128
rect 24815 17088 24860 17116
rect 24854 17076 24860 17088
rect 24912 17076 24918 17128
rect 24946 17076 24952 17128
rect 25004 17116 25010 17128
rect 25113 17119 25171 17125
rect 25113 17116 25125 17119
rect 25004 17088 25125 17116
rect 25004 17076 25010 17088
rect 25113 17085 25125 17088
rect 25159 17116 25171 17119
rect 26789 17119 26847 17125
rect 26789 17116 26801 17119
rect 25159 17088 26801 17116
rect 25159 17085 25171 17088
rect 25113 17079 25171 17085
rect 26789 17085 26801 17088
rect 26835 17116 26847 17119
rect 26970 17116 26976 17128
rect 26835 17088 26976 17116
rect 26835 17085 26847 17088
rect 26789 17079 26847 17085
rect 26970 17076 26976 17088
rect 27028 17076 27034 17128
rect 27614 17116 27620 17128
rect 27575 17088 27620 17116
rect 27614 17076 27620 17088
rect 27672 17116 27678 17128
rect 28261 17119 28319 17125
rect 28261 17116 28273 17119
rect 27672 17088 28273 17116
rect 27672 17076 27678 17088
rect 28261 17085 28273 17088
rect 28307 17085 28319 17119
rect 28261 17079 28319 17085
rect 30193 17119 30251 17125
rect 30193 17085 30205 17119
rect 30239 17116 30251 17119
rect 30282 17116 30288 17128
rect 30239 17088 30288 17116
rect 30239 17085 30251 17088
rect 30193 17079 30251 17085
rect 30282 17076 30288 17088
rect 30340 17076 30346 17128
rect 30466 17125 30472 17128
rect 30460 17116 30472 17125
rect 30392 17088 30472 17116
rect 19058 17008 19064 17060
rect 19116 17048 19122 17060
rect 19337 17051 19395 17057
rect 19337 17048 19349 17051
rect 19116 17020 19349 17048
rect 19116 17008 19122 17020
rect 19337 17017 19349 17020
rect 19383 17048 19395 17051
rect 20441 17051 20499 17057
rect 20441 17048 20453 17051
rect 19383 17020 20453 17048
rect 19383 17017 19395 17020
rect 19337 17011 19395 17017
rect 20441 17017 20453 17020
rect 20487 17048 20499 17051
rect 20800 17051 20858 17057
rect 20800 17048 20812 17051
rect 20487 17020 20812 17048
rect 20487 17017 20499 17020
rect 20441 17011 20499 17017
rect 20800 17017 20812 17020
rect 20846 17048 20858 17051
rect 22278 17048 22284 17060
rect 20846 17020 22284 17048
rect 20846 17017 20858 17020
rect 20800 17011 20858 17017
rect 22278 17008 22284 17020
rect 22336 17008 22342 17060
rect 24118 17008 24124 17060
rect 24176 17048 24182 17060
rect 24673 17051 24731 17057
rect 24673 17048 24685 17051
rect 24176 17020 24685 17048
rect 24176 17008 24182 17020
rect 24673 17017 24685 17020
rect 24719 17048 24731 17051
rect 25314 17048 25320 17060
rect 24719 17020 25320 17048
rect 24719 17017 24731 17020
rect 24673 17011 24731 17017
rect 25314 17008 25320 17020
rect 25372 17008 25378 17060
rect 30101 17051 30159 17057
rect 30101 17017 30113 17051
rect 30147 17048 30159 17051
rect 30392 17048 30420 17088
rect 30460 17079 30472 17088
rect 30466 17076 30472 17079
rect 30524 17076 30530 17128
rect 30147 17020 30420 17048
rect 35704 17051 35762 17057
rect 30147 17017 30159 17020
rect 30101 17011 30159 17017
rect 35704 17017 35716 17051
rect 35750 17048 35762 17051
rect 35802 17048 35808 17060
rect 35750 17020 35808 17048
rect 35750 17017 35762 17020
rect 35704 17011 35762 17017
rect 35802 17008 35808 17020
rect 35860 17008 35866 17060
rect 18877 16983 18935 16989
rect 18877 16949 18889 16983
rect 18923 16980 18935 16983
rect 19429 16983 19487 16989
rect 19429 16980 19441 16983
rect 18923 16952 19441 16980
rect 18923 16949 18935 16952
rect 18877 16943 18935 16949
rect 19429 16949 19441 16952
rect 19475 16980 19487 16983
rect 20162 16980 20168 16992
rect 19475 16952 20168 16980
rect 19475 16949 19487 16952
rect 19429 16943 19487 16949
rect 20162 16940 20168 16952
rect 20220 16940 20226 16992
rect 24397 16983 24455 16989
rect 24397 16949 24409 16983
rect 24443 16980 24455 16983
rect 25222 16980 25228 16992
rect 24443 16952 25228 16980
rect 24443 16949 24455 16952
rect 24397 16943 24455 16949
rect 25222 16940 25228 16952
rect 25280 16940 25286 16992
rect 26234 16980 26240 16992
rect 26195 16952 26240 16980
rect 26234 16940 26240 16952
rect 26292 16980 26298 16992
rect 26878 16980 26884 16992
rect 26292 16952 26884 16980
rect 26292 16940 26298 16952
rect 26878 16940 26884 16952
rect 26936 16980 26942 16992
rect 27157 16983 27215 16989
rect 27157 16980 27169 16983
rect 26936 16952 27169 16980
rect 26936 16940 26942 16952
rect 27157 16949 27169 16952
rect 27203 16949 27215 16983
rect 27157 16943 27215 16949
rect 34517 16983 34575 16989
rect 34517 16949 34529 16983
rect 34563 16980 34575 16983
rect 35342 16980 35348 16992
rect 34563 16952 35348 16980
rect 34563 16949 34575 16952
rect 34517 16943 34575 16949
rect 35342 16940 35348 16952
rect 35400 16980 35406 16992
rect 36817 16983 36875 16989
rect 36817 16980 36829 16983
rect 35400 16952 36829 16980
rect 35400 16940 35406 16952
rect 36817 16949 36829 16952
rect 36863 16980 36875 16983
rect 36906 16980 36912 16992
rect 36863 16952 36912 16980
rect 36863 16949 36875 16952
rect 36817 16943 36875 16949
rect 36906 16940 36912 16952
rect 36964 16940 36970 16992
rect 1104 16890 38824 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 38824 16890
rect 1104 16816 38824 16838
rect 19058 16776 19064 16788
rect 19019 16748 19064 16776
rect 19058 16736 19064 16748
rect 19116 16736 19122 16788
rect 19242 16776 19248 16788
rect 19203 16748 19248 16776
rect 19242 16736 19248 16748
rect 19300 16736 19306 16788
rect 22278 16776 22284 16788
rect 22239 16748 22284 16776
rect 22278 16736 22284 16748
rect 22336 16736 22342 16788
rect 23658 16776 23664 16788
rect 23619 16748 23664 16776
rect 23658 16736 23664 16748
rect 23716 16736 23722 16788
rect 25222 16736 25228 16788
rect 25280 16776 25286 16788
rect 25317 16779 25375 16785
rect 25317 16776 25329 16779
rect 25280 16748 25329 16776
rect 25280 16736 25286 16748
rect 25317 16745 25329 16748
rect 25363 16776 25375 16779
rect 25363 16748 26823 16776
rect 25363 16745 25375 16748
rect 25317 16739 25375 16745
rect 20162 16668 20168 16720
rect 20220 16708 20226 16720
rect 21146 16711 21204 16717
rect 21146 16708 21158 16711
rect 20220 16680 21158 16708
rect 20220 16668 20226 16680
rect 21146 16677 21158 16680
rect 21192 16708 21204 16711
rect 22094 16708 22100 16720
rect 21192 16680 22100 16708
rect 21192 16677 21204 16680
rect 21146 16671 21204 16677
rect 22094 16668 22100 16680
rect 22152 16668 22158 16720
rect 24118 16668 24124 16720
rect 24176 16717 24182 16720
rect 24176 16711 24240 16717
rect 24176 16677 24194 16711
rect 24228 16677 24240 16711
rect 24176 16671 24240 16677
rect 24176 16668 24182 16671
rect 24854 16668 24860 16720
rect 24912 16668 24918 16720
rect 19610 16640 19616 16652
rect 19571 16612 19616 16640
rect 19610 16600 19616 16612
rect 19668 16600 19674 16652
rect 20625 16643 20683 16649
rect 20625 16609 20637 16643
rect 20671 16640 20683 16643
rect 20714 16640 20720 16652
rect 20671 16612 20720 16640
rect 20671 16609 20683 16612
rect 20625 16603 20683 16609
rect 20714 16600 20720 16612
rect 20772 16640 20778 16652
rect 20901 16643 20959 16649
rect 20901 16640 20913 16643
rect 20772 16612 20913 16640
rect 20772 16600 20778 16612
rect 20901 16609 20913 16612
rect 20947 16609 20959 16643
rect 20901 16603 20959 16609
rect 23937 16643 23995 16649
rect 23937 16609 23949 16643
rect 23983 16640 23995 16643
rect 24872 16640 24900 16668
rect 26795 16649 26823 16748
rect 26970 16736 26976 16788
rect 27028 16776 27034 16788
rect 27893 16779 27951 16785
rect 27893 16776 27905 16779
rect 27028 16748 27905 16776
rect 27028 16736 27034 16748
rect 27893 16745 27905 16748
rect 27939 16745 27951 16779
rect 29914 16776 29920 16788
rect 29875 16748 29920 16776
rect 27893 16739 27951 16745
rect 29914 16736 29920 16748
rect 29972 16736 29978 16788
rect 30374 16736 30380 16788
rect 30432 16776 30438 16788
rect 30929 16779 30987 16785
rect 30929 16776 30941 16779
rect 30432 16748 30941 16776
rect 30432 16736 30438 16748
rect 30929 16745 30941 16748
rect 30975 16745 30987 16779
rect 30929 16739 30987 16745
rect 35529 16779 35587 16785
rect 35529 16745 35541 16779
rect 35575 16776 35587 16779
rect 35802 16776 35808 16788
rect 35575 16748 35808 16776
rect 35575 16745 35587 16748
rect 35529 16739 35587 16745
rect 35802 16736 35808 16748
rect 35860 16736 35866 16788
rect 29546 16668 29552 16720
rect 29604 16708 29610 16720
rect 30190 16708 30196 16720
rect 29604 16680 30196 16708
rect 29604 16668 29610 16680
rect 30190 16668 30196 16680
rect 30248 16708 30254 16720
rect 30285 16711 30343 16717
rect 30285 16708 30297 16711
rect 30248 16680 30297 16708
rect 30248 16668 30254 16680
rect 30285 16677 30297 16680
rect 30331 16677 30343 16711
rect 30285 16671 30343 16677
rect 23983 16612 24900 16640
rect 26780 16643 26838 16649
rect 23983 16609 23995 16612
rect 23937 16603 23995 16609
rect 26780 16609 26792 16643
rect 26826 16640 26838 16643
rect 27062 16640 27068 16652
rect 26826 16612 27068 16640
rect 26826 16609 26838 16612
rect 26780 16603 26838 16609
rect 27062 16600 27068 16612
rect 27120 16600 27126 16652
rect 28994 16600 29000 16652
rect 29052 16640 29058 16652
rect 29052 16612 30328 16640
rect 29052 16600 29058 16612
rect 19702 16572 19708 16584
rect 19663 16544 19708 16572
rect 19702 16532 19708 16544
rect 19760 16532 19766 16584
rect 19886 16572 19892 16584
rect 19847 16544 19892 16572
rect 19886 16532 19892 16544
rect 19944 16532 19950 16584
rect 25961 16575 26019 16581
rect 25961 16541 25973 16575
rect 26007 16572 26019 16575
rect 26510 16572 26516 16584
rect 26007 16544 26516 16572
rect 26007 16541 26019 16544
rect 25961 16535 26019 16541
rect 26510 16532 26516 16544
rect 26568 16532 26574 16584
rect 30300 16572 30328 16612
rect 30374 16572 30380 16584
rect 30287 16544 30380 16572
rect 30374 16532 30380 16544
rect 30432 16532 30438 16584
rect 30466 16532 30472 16584
rect 30524 16572 30530 16584
rect 30524 16544 30569 16572
rect 30524 16532 30530 16544
rect 35434 16532 35440 16584
rect 35492 16572 35498 16584
rect 36630 16572 36636 16584
rect 35492 16544 36636 16572
rect 35492 16532 35498 16544
rect 36630 16532 36636 16544
rect 36688 16532 36694 16584
rect 1104 16346 38824 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 34966 16346
rect 35018 16294 35030 16346
rect 35082 16294 35094 16346
rect 35146 16294 35158 16346
rect 35210 16294 38824 16346
rect 1104 16272 38824 16294
rect 18969 16235 19027 16241
rect 18969 16201 18981 16235
rect 19015 16232 19027 16235
rect 19886 16232 19892 16244
rect 19015 16204 19892 16232
rect 19015 16201 19027 16204
rect 18969 16195 19027 16201
rect 19886 16192 19892 16204
rect 19944 16192 19950 16244
rect 20162 16232 20168 16244
rect 20123 16204 20168 16232
rect 20162 16192 20168 16204
rect 20220 16192 20226 16244
rect 22094 16192 22100 16244
rect 22152 16232 22158 16244
rect 24029 16235 24087 16241
rect 22152 16204 22197 16232
rect 22152 16192 22158 16204
rect 24029 16201 24041 16235
rect 24075 16232 24087 16235
rect 24118 16232 24124 16244
rect 24075 16204 24124 16232
rect 24075 16201 24087 16204
rect 24029 16195 24087 16201
rect 24118 16192 24124 16204
rect 24176 16232 24182 16244
rect 26881 16235 26939 16241
rect 26881 16232 26893 16235
rect 24176 16204 26893 16232
rect 24176 16192 24182 16204
rect 26881 16201 26893 16204
rect 26927 16201 26939 16235
rect 26881 16195 26939 16201
rect 27062 16192 27068 16244
rect 27120 16232 27126 16244
rect 27433 16235 27491 16241
rect 27433 16232 27445 16235
rect 27120 16204 27445 16232
rect 27120 16192 27126 16204
rect 27433 16201 27445 16204
rect 27479 16201 27491 16235
rect 29914 16232 29920 16244
rect 29875 16204 29920 16232
rect 27433 16195 27491 16201
rect 29914 16192 29920 16204
rect 29972 16192 29978 16244
rect 30190 16232 30196 16244
rect 30151 16204 30196 16232
rect 30190 16192 30196 16204
rect 30248 16192 30254 16244
rect 30466 16192 30472 16244
rect 30524 16232 30530 16244
rect 30561 16235 30619 16241
rect 30561 16232 30573 16235
rect 30524 16204 30573 16232
rect 30524 16192 30530 16204
rect 30561 16201 30573 16204
rect 30607 16201 30619 16235
rect 30561 16195 30619 16201
rect 24949 16167 25007 16173
rect 24949 16133 24961 16167
rect 24995 16164 25007 16167
rect 25130 16164 25136 16176
rect 24995 16136 25136 16164
rect 24995 16133 25007 16136
rect 24949 16127 25007 16133
rect 25130 16124 25136 16136
rect 25188 16124 25194 16176
rect 33042 16124 33048 16176
rect 33100 16164 33106 16176
rect 34606 16164 34612 16176
rect 33100 16136 34612 16164
rect 33100 16124 33106 16136
rect 34606 16124 34612 16136
rect 34664 16124 34670 16176
rect 19337 16099 19395 16105
rect 19337 16065 19349 16099
rect 19383 16096 19395 16099
rect 19702 16096 19708 16108
rect 19383 16068 19708 16096
rect 19383 16065 19395 16068
rect 19337 16059 19395 16065
rect 19702 16056 19708 16068
rect 19760 16096 19766 16108
rect 20622 16096 20628 16108
rect 19760 16068 20628 16096
rect 19760 16056 19766 16068
rect 20622 16056 20628 16068
rect 20680 16056 20686 16108
rect 28626 16096 28632 16108
rect 28000 16068 28632 16096
rect 20714 16028 20720 16040
rect 20675 16000 20720 16028
rect 20714 15988 20720 16000
rect 20772 15988 20778 16040
rect 22741 16031 22799 16037
rect 22741 15997 22753 16031
rect 22787 16028 22799 16031
rect 24397 16031 24455 16037
rect 24397 16028 24409 16031
rect 22787 16000 24409 16028
rect 22787 15997 22799 16000
rect 22741 15991 22799 15997
rect 24397 15997 24409 16000
rect 24443 16028 24455 16031
rect 24578 16028 24584 16040
rect 24443 16000 24584 16028
rect 24443 15997 24455 16000
rect 24397 15991 24455 15997
rect 24578 15988 24584 16000
rect 24636 16028 24642 16040
rect 24854 16028 24860 16040
rect 24636 16000 24860 16028
rect 24636 15988 24642 16000
rect 24854 15988 24860 16000
rect 24912 16028 24918 16040
rect 25501 16031 25559 16037
rect 25501 16028 25513 16031
rect 24912 16000 25513 16028
rect 24912 15988 24918 16000
rect 25501 15997 25513 16000
rect 25547 16028 25559 16031
rect 26510 16028 26516 16040
rect 25547 16000 26516 16028
rect 25547 15997 25559 16000
rect 25501 15991 25559 15997
rect 26510 15988 26516 16000
rect 26568 15988 26574 16040
rect 28000 16037 28028 16068
rect 28626 16056 28632 16068
rect 28684 16056 28690 16108
rect 27985 16031 28043 16037
rect 27985 15997 27997 16031
rect 28031 15997 28043 16031
rect 27985 15991 28043 15997
rect 29273 16031 29331 16037
rect 29273 15997 29285 16031
rect 29319 16028 29331 16031
rect 29914 16028 29920 16040
rect 29319 16000 29920 16028
rect 29319 15997 29331 16000
rect 29273 15991 29331 15997
rect 29914 15988 29920 16000
rect 29972 15988 29978 16040
rect 19610 15920 19616 15972
rect 19668 15960 19674 15972
rect 19705 15963 19763 15969
rect 19705 15960 19717 15963
rect 19668 15932 19717 15960
rect 19668 15920 19674 15932
rect 19705 15929 19717 15932
rect 19751 15960 19763 15963
rect 20625 15963 20683 15969
rect 20625 15960 20637 15963
rect 19751 15932 20637 15960
rect 19751 15929 19763 15932
rect 19705 15923 19763 15929
rect 20625 15929 20637 15932
rect 20671 15960 20683 15963
rect 20984 15963 21042 15969
rect 20984 15960 20996 15963
rect 20671 15932 20996 15960
rect 20671 15929 20683 15932
rect 20625 15923 20683 15929
rect 20984 15929 20996 15932
rect 21030 15960 21042 15963
rect 22278 15960 22284 15972
rect 21030 15932 22284 15960
rect 21030 15929 21042 15932
rect 20984 15923 21042 15929
rect 22278 15920 22284 15932
rect 22336 15920 22342 15972
rect 25774 15969 25780 15972
rect 25409 15963 25467 15969
rect 25409 15929 25421 15963
rect 25455 15960 25467 15963
rect 25768 15960 25780 15969
rect 25455 15932 25780 15960
rect 25455 15929 25467 15932
rect 25409 15923 25467 15929
rect 25768 15923 25780 15932
rect 25774 15920 25780 15923
rect 25832 15920 25838 15972
rect 27154 15852 27160 15904
rect 27212 15892 27218 15904
rect 28169 15895 28227 15901
rect 28169 15892 28181 15895
rect 27212 15864 28181 15892
rect 27212 15852 27218 15864
rect 28169 15861 28181 15864
rect 28215 15861 28227 15895
rect 29454 15892 29460 15904
rect 29415 15864 29460 15892
rect 28169 15855 28227 15861
rect 29454 15852 29460 15864
rect 29512 15852 29518 15904
rect 32493 15895 32551 15901
rect 32493 15861 32505 15895
rect 32539 15892 32551 15895
rect 33042 15892 33048 15904
rect 32539 15864 33048 15892
rect 32539 15861 32551 15864
rect 32493 15855 32551 15861
rect 33042 15852 33048 15864
rect 33100 15852 33106 15904
rect 35437 15895 35495 15901
rect 35437 15861 35449 15895
rect 35483 15892 35495 15895
rect 35802 15892 35808 15904
rect 35483 15864 35808 15892
rect 35483 15861 35495 15864
rect 35437 15855 35495 15861
rect 35802 15852 35808 15864
rect 35860 15852 35866 15904
rect 1104 15802 38824 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 38824 15802
rect 1104 15728 38824 15750
rect 22278 15688 22284 15700
rect 22239 15660 22284 15688
rect 22278 15648 22284 15660
rect 22336 15648 22342 15700
rect 30374 15688 30380 15700
rect 30335 15660 30380 15688
rect 30374 15648 30380 15660
rect 30432 15648 30438 15700
rect 35710 15648 35716 15700
rect 35768 15688 35774 15700
rect 35986 15688 35992 15700
rect 35768 15660 35992 15688
rect 35768 15648 35774 15660
rect 35986 15648 35992 15660
rect 36044 15648 36050 15700
rect 20622 15512 20628 15564
rect 20680 15552 20686 15564
rect 21168 15555 21226 15561
rect 21168 15552 21180 15555
rect 20680 15524 21180 15552
rect 20680 15512 20686 15524
rect 21168 15521 21180 15524
rect 21214 15552 21226 15555
rect 22002 15552 22008 15564
rect 21214 15524 22008 15552
rect 21214 15521 21226 15524
rect 21168 15515 21226 15521
rect 22002 15512 22008 15524
rect 22060 15512 22066 15564
rect 27709 15555 27767 15561
rect 27709 15521 27721 15555
rect 27755 15552 27767 15555
rect 27982 15552 27988 15564
rect 27755 15524 27988 15552
rect 27755 15521 27767 15524
rect 27709 15515 27767 15521
rect 27982 15512 27988 15524
rect 28040 15512 28046 15564
rect 29730 15552 29736 15564
rect 29691 15524 29736 15552
rect 29730 15512 29736 15524
rect 29788 15512 29794 15564
rect 32214 15512 32220 15564
rect 32272 15552 32278 15564
rect 32769 15555 32827 15561
rect 32769 15552 32781 15555
rect 32272 15524 32781 15552
rect 32272 15512 32278 15524
rect 32769 15521 32781 15524
rect 32815 15521 32827 15555
rect 32769 15515 32827 15521
rect 32861 15555 32919 15561
rect 32861 15521 32873 15555
rect 32907 15552 32919 15555
rect 33042 15552 33048 15564
rect 32907 15524 33048 15552
rect 32907 15521 32919 15524
rect 32861 15515 32919 15521
rect 33042 15512 33048 15524
rect 33100 15512 33106 15564
rect 35434 15552 35440 15564
rect 35395 15524 35440 15552
rect 35434 15512 35440 15524
rect 35492 15512 35498 15564
rect 20714 15484 20720 15496
rect 20627 15456 20720 15484
rect 20714 15444 20720 15456
rect 20772 15484 20778 15496
rect 20898 15484 20904 15496
rect 20772 15456 20904 15484
rect 20772 15444 20778 15456
rect 20898 15444 20904 15456
rect 20956 15444 20962 15496
rect 27798 15484 27804 15496
rect 27759 15456 27804 15484
rect 27798 15444 27804 15456
rect 27856 15444 27862 15496
rect 27890 15444 27896 15496
rect 27948 15484 27954 15496
rect 29454 15484 29460 15496
rect 27948 15456 29460 15484
rect 27948 15444 27954 15456
rect 29454 15444 29460 15456
rect 29512 15444 29518 15496
rect 31754 15444 31760 15496
rect 31812 15484 31818 15496
rect 32950 15484 32956 15496
rect 31812 15456 32956 15484
rect 31812 15444 31818 15456
rect 32950 15444 32956 15456
rect 33008 15444 33014 15496
rect 26789 15419 26847 15425
rect 26789 15385 26801 15419
rect 26835 15416 26847 15419
rect 27154 15416 27160 15428
rect 26835 15388 27160 15416
rect 26835 15385 26847 15388
rect 26789 15379 26847 15385
rect 27154 15376 27160 15388
rect 27212 15376 27218 15428
rect 25593 15351 25651 15357
rect 25593 15317 25605 15351
rect 25639 15348 25651 15351
rect 26510 15348 26516 15360
rect 25639 15320 26516 15348
rect 25639 15317 25651 15320
rect 25593 15311 25651 15317
rect 26510 15308 26516 15320
rect 26568 15348 26574 15360
rect 27062 15348 27068 15360
rect 26568 15320 27068 15348
rect 26568 15308 26574 15320
rect 27062 15308 27068 15320
rect 27120 15308 27126 15360
rect 27338 15348 27344 15360
rect 27299 15320 27344 15348
rect 27338 15308 27344 15320
rect 27396 15308 27402 15360
rect 29917 15351 29975 15357
rect 29917 15317 29929 15351
rect 29963 15348 29975 15351
rect 30190 15348 30196 15360
rect 29963 15320 30196 15348
rect 29963 15317 29975 15320
rect 29917 15311 29975 15317
rect 30190 15308 30196 15320
rect 30248 15308 30254 15360
rect 32398 15348 32404 15360
rect 32359 15320 32404 15348
rect 32398 15308 32404 15320
rect 32456 15308 32462 15360
rect 34514 15308 34520 15360
rect 34572 15348 34578 15360
rect 35621 15351 35679 15357
rect 35621 15348 35633 15351
rect 34572 15320 35633 15348
rect 34572 15308 34578 15320
rect 35621 15317 35633 15320
rect 35667 15317 35679 15351
rect 35621 15311 35679 15317
rect 1104 15258 38824 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 34966 15258
rect 35018 15206 35030 15258
rect 35082 15206 35094 15258
rect 35146 15206 35158 15258
rect 35210 15206 38824 15258
rect 1104 15184 38824 15206
rect 20622 15144 20628 15156
rect 20583 15116 20628 15144
rect 20622 15104 20628 15116
rect 20680 15104 20686 15156
rect 22094 15104 22100 15156
rect 22152 15144 22158 15156
rect 22465 15147 22523 15153
rect 22465 15144 22477 15147
rect 22152 15116 22477 15144
rect 22152 15104 22158 15116
rect 22465 15113 22477 15116
rect 22511 15113 22523 15147
rect 22465 15107 22523 15113
rect 27709 15147 27767 15153
rect 27709 15113 27721 15147
rect 27755 15144 27767 15147
rect 27798 15144 27804 15156
rect 27755 15116 27804 15144
rect 27755 15113 27767 15116
rect 27709 15107 27767 15113
rect 27798 15104 27804 15116
rect 27856 15104 27862 15156
rect 27982 15144 27988 15156
rect 27943 15116 27988 15144
rect 27982 15104 27988 15116
rect 28040 15104 28046 15156
rect 29089 15147 29147 15153
rect 29089 15113 29101 15147
rect 29135 15144 29147 15147
rect 29730 15144 29736 15156
rect 29135 15116 29736 15144
rect 29135 15113 29147 15116
rect 29089 15107 29147 15113
rect 29730 15104 29736 15116
rect 29788 15144 29794 15156
rect 30193 15147 30251 15153
rect 30193 15144 30205 15147
rect 29788 15116 30205 15144
rect 29788 15104 29794 15116
rect 30193 15113 30205 15116
rect 30239 15113 30251 15147
rect 30193 15107 30251 15113
rect 31754 15104 31760 15156
rect 31812 15144 31818 15156
rect 32214 15144 32220 15156
rect 31812 15116 31857 15144
rect 32175 15116 32220 15144
rect 31812 15104 31818 15116
rect 32214 15104 32220 15116
rect 32272 15104 32278 15156
rect 32950 15104 32956 15156
rect 33008 15144 33014 15156
rect 33689 15147 33747 15153
rect 33689 15144 33701 15147
rect 33008 15116 33701 15144
rect 33008 15104 33014 15116
rect 33689 15113 33701 15116
rect 33735 15113 33747 15147
rect 33689 15107 33747 15113
rect 35345 15147 35403 15153
rect 35345 15113 35357 15147
rect 35391 15144 35403 15147
rect 35434 15144 35440 15156
rect 35391 15116 35440 15144
rect 35391 15113 35403 15116
rect 35345 15107 35403 15113
rect 35434 15104 35440 15116
rect 35492 15104 35498 15156
rect 27062 15036 27068 15088
rect 27120 15076 27126 15088
rect 28074 15076 28080 15088
rect 27120 15048 28080 15076
rect 27120 15036 27126 15048
rect 28074 15036 28080 15048
rect 28132 15036 28138 15088
rect 20993 15011 21051 15017
rect 20993 14977 21005 15011
rect 21039 15008 21051 15011
rect 27154 15008 27160 15020
rect 21039 14980 21220 15008
rect 27115 14980 27160 15008
rect 21039 14977 21051 14980
rect 20993 14971 21051 14977
rect 20257 14943 20315 14949
rect 20257 14909 20269 14943
rect 20303 14940 20315 14943
rect 20898 14940 20904 14952
rect 20303 14912 20904 14940
rect 20303 14909 20315 14912
rect 20257 14903 20315 14909
rect 20898 14900 20904 14912
rect 20956 14940 20962 14952
rect 21085 14943 21143 14949
rect 21085 14940 21097 14943
rect 20956 14912 21097 14940
rect 20956 14900 20962 14912
rect 21085 14909 21097 14912
rect 21131 14909 21143 14943
rect 21192 14940 21220 14980
rect 27154 14968 27160 14980
rect 27212 14968 27218 15020
rect 30558 15008 30564 15020
rect 30519 14980 30564 15008
rect 30558 14968 30564 14980
rect 30616 14968 30622 15020
rect 21358 14949 21364 14952
rect 21352 14940 21364 14949
rect 21192 14912 21364 14940
rect 21085 14903 21143 14909
rect 21352 14903 21364 14912
rect 21100 14872 21128 14903
rect 21358 14900 21364 14903
rect 21416 14900 21422 14952
rect 26145 14943 26203 14949
rect 26145 14909 26157 14943
rect 26191 14940 26203 14943
rect 26973 14943 27031 14949
rect 26973 14940 26985 14943
rect 26191 14912 26985 14940
rect 26191 14909 26203 14912
rect 26145 14903 26203 14909
rect 26973 14909 26985 14912
rect 27019 14940 27031 14943
rect 27338 14940 27344 14952
rect 27019 14912 27344 14940
rect 27019 14909 27031 14912
rect 26973 14903 27031 14909
rect 27338 14900 27344 14912
rect 27396 14900 27402 14952
rect 29733 14943 29791 14949
rect 29733 14909 29745 14943
rect 29779 14940 29791 14943
rect 30006 14940 30012 14952
rect 29779 14912 30012 14940
rect 29779 14909 29791 14912
rect 29733 14903 29791 14909
rect 30006 14900 30012 14912
rect 30064 14900 30070 14952
rect 21174 14872 21180 14884
rect 21100 14844 21180 14872
rect 21174 14832 21180 14844
rect 21232 14832 21238 14884
rect 26510 14872 26516 14884
rect 26423 14844 26516 14872
rect 26510 14832 26516 14844
rect 26568 14872 26574 14884
rect 27065 14875 27123 14881
rect 27065 14872 27077 14875
rect 26568 14844 27077 14872
rect 26568 14832 26574 14844
rect 27065 14841 27077 14844
rect 27111 14841 27123 14875
rect 27065 14835 27123 14841
rect 29825 14875 29883 14881
rect 29825 14841 29837 14875
rect 29871 14872 29883 14875
rect 30576 14872 30604 14968
rect 30742 14900 30748 14952
rect 30800 14940 30806 14952
rect 30929 14943 30987 14949
rect 30929 14940 30941 14943
rect 30800 14912 30941 14940
rect 30800 14900 30806 14912
rect 30929 14909 30941 14912
rect 30975 14940 30987 14943
rect 31021 14943 31079 14949
rect 31021 14940 31033 14943
rect 30975 14912 31033 14940
rect 30975 14909 30987 14912
rect 30929 14903 30987 14909
rect 31021 14909 31033 14912
rect 31067 14909 31079 14943
rect 32306 14940 32312 14952
rect 32267 14912 32312 14940
rect 31021 14903 31079 14909
rect 32306 14900 32312 14912
rect 32364 14900 32370 14952
rect 35250 14900 35256 14952
rect 35308 14940 35314 14952
rect 35437 14943 35495 14949
rect 35437 14940 35449 14943
rect 35308 14912 35449 14940
rect 35308 14900 35314 14912
rect 35437 14909 35449 14912
rect 35483 14940 35495 14943
rect 35986 14940 35992 14952
rect 35483 14912 35992 14940
rect 35483 14909 35495 14912
rect 35437 14903 35495 14909
rect 35986 14900 35992 14912
rect 36044 14900 36050 14952
rect 29871 14844 30604 14872
rect 32576 14875 32634 14881
rect 29871 14841 29883 14844
rect 29825 14835 29883 14841
rect 32576 14841 32588 14875
rect 32622 14872 32634 14875
rect 32766 14872 32772 14884
rect 32622 14844 32772 14872
rect 32622 14841 32634 14844
rect 32576 14835 32634 14841
rect 32766 14832 32772 14844
rect 32824 14832 32830 14884
rect 34701 14875 34759 14881
rect 34701 14841 34713 14875
rect 34747 14872 34759 14875
rect 35682 14875 35740 14881
rect 35682 14872 35694 14875
rect 34747 14844 35694 14872
rect 34747 14841 34759 14844
rect 34701 14835 34759 14841
rect 35682 14841 35694 14844
rect 35728 14872 35740 14875
rect 36446 14872 36452 14884
rect 35728 14844 36452 14872
rect 35728 14841 35740 14844
rect 35682 14835 35740 14841
rect 36446 14832 36452 14844
rect 36504 14832 36510 14884
rect 26602 14804 26608 14816
rect 26563 14776 26608 14804
rect 26602 14764 26608 14776
rect 26660 14764 26666 14816
rect 31205 14807 31263 14813
rect 31205 14773 31217 14807
rect 31251 14804 31263 14807
rect 33778 14804 33784 14816
rect 31251 14776 33784 14804
rect 31251 14773 31263 14776
rect 31205 14767 31263 14773
rect 33778 14764 33784 14776
rect 33836 14764 33842 14816
rect 35526 14764 35532 14816
rect 35584 14804 35590 14816
rect 36817 14807 36875 14813
rect 36817 14804 36829 14807
rect 35584 14776 36829 14804
rect 35584 14764 35590 14776
rect 36817 14773 36829 14776
rect 36863 14773 36875 14807
rect 36817 14767 36875 14773
rect 1104 14714 38824 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 38824 14714
rect 1104 14640 38824 14662
rect 24578 14600 24584 14612
rect 24539 14572 24584 14600
rect 24578 14560 24584 14572
rect 24636 14560 24642 14612
rect 26510 14600 26516 14612
rect 26471 14572 26516 14600
rect 26510 14560 26516 14572
rect 26568 14560 26574 14612
rect 27617 14603 27675 14609
rect 27617 14569 27629 14603
rect 27663 14600 27675 14603
rect 27890 14600 27896 14612
rect 27663 14572 27896 14600
rect 27663 14569 27675 14572
rect 27617 14563 27675 14569
rect 26881 14535 26939 14541
rect 26881 14501 26893 14535
rect 26927 14532 26939 14535
rect 27062 14532 27068 14544
rect 26927 14504 27068 14532
rect 26927 14501 26939 14504
rect 26881 14495 26939 14501
rect 27062 14492 27068 14504
rect 27120 14492 27126 14544
rect 23842 14464 23848 14476
rect 23803 14436 23848 14464
rect 23842 14424 23848 14436
rect 23900 14424 23906 14476
rect 23934 14396 23940 14408
rect 23895 14368 23940 14396
rect 23934 14356 23940 14368
rect 23992 14356 23998 14408
rect 24121 14399 24179 14405
rect 24121 14365 24133 14399
rect 24167 14365 24179 14399
rect 26970 14396 26976 14408
rect 26931 14368 26976 14396
rect 24121 14359 24179 14365
rect 23106 14288 23112 14340
rect 23164 14328 23170 14340
rect 24136 14328 24164 14359
rect 26970 14356 26976 14368
rect 27028 14356 27034 14408
rect 27157 14399 27215 14405
rect 27157 14365 27169 14399
rect 27203 14396 27215 14399
rect 27338 14396 27344 14408
rect 27203 14368 27344 14396
rect 27203 14365 27215 14368
rect 27157 14359 27215 14365
rect 27172 14328 27200 14359
rect 27338 14356 27344 14368
rect 27396 14396 27402 14408
rect 27632 14396 27660 14563
rect 27890 14560 27896 14572
rect 27948 14560 27954 14612
rect 30006 14560 30012 14612
rect 30064 14600 30070 14612
rect 30101 14603 30159 14609
rect 30101 14600 30113 14603
rect 30064 14572 30113 14600
rect 30064 14560 30070 14572
rect 30101 14569 30113 14572
rect 30147 14569 30159 14603
rect 32214 14600 32220 14612
rect 32175 14572 32220 14600
rect 30101 14563 30159 14569
rect 32214 14560 32220 14572
rect 32272 14560 32278 14612
rect 33695 14603 33753 14609
rect 33695 14569 33707 14603
rect 33741 14600 33753 14603
rect 33870 14600 33876 14612
rect 33741 14572 33876 14600
rect 33741 14569 33753 14572
rect 33695 14563 33753 14569
rect 33870 14560 33876 14572
rect 33928 14560 33934 14612
rect 34606 14560 34612 14612
rect 34664 14600 34670 14612
rect 35069 14603 35127 14609
rect 35069 14600 35081 14603
rect 34664 14572 35081 14600
rect 34664 14560 34670 14572
rect 35069 14569 35081 14572
rect 35115 14600 35127 14603
rect 35526 14600 35532 14612
rect 35115 14572 35388 14600
rect 35487 14572 35532 14600
rect 35115 14569 35127 14572
rect 35069 14563 35127 14569
rect 27982 14492 27988 14544
rect 28040 14532 28046 14544
rect 28718 14532 28724 14544
rect 28040 14504 28724 14532
rect 28040 14492 28046 14504
rect 28718 14492 28724 14504
rect 28776 14532 28782 14544
rect 28966 14535 29024 14541
rect 28966 14532 28978 14535
rect 28776 14504 28978 14532
rect 28776 14492 28782 14504
rect 28966 14501 28978 14504
rect 29012 14501 29024 14535
rect 35360 14532 35388 14572
rect 35526 14560 35532 14572
rect 35584 14560 35590 14612
rect 36170 14560 36176 14612
rect 36228 14600 36234 14612
rect 36265 14603 36323 14609
rect 36265 14600 36277 14603
rect 36228 14572 36277 14600
rect 36228 14560 36234 14572
rect 36265 14569 36277 14572
rect 36311 14569 36323 14603
rect 36265 14563 36323 14569
rect 36078 14532 36084 14544
rect 35360 14504 36084 14532
rect 28966 14495 29024 14501
rect 36078 14492 36084 14504
rect 36136 14532 36142 14544
rect 36357 14535 36415 14541
rect 36357 14532 36369 14535
rect 36136 14504 36369 14532
rect 36136 14492 36142 14504
rect 36357 14501 36369 14504
rect 36403 14501 36415 14535
rect 36357 14495 36415 14501
rect 30282 14464 30288 14476
rect 28736 14436 30288 14464
rect 27396 14368 27660 14396
rect 27396 14356 27402 14368
rect 28074 14356 28080 14408
rect 28132 14396 28138 14408
rect 28736 14405 28764 14436
rect 30282 14424 30288 14436
rect 30340 14424 30346 14476
rect 33965 14467 34023 14473
rect 33965 14464 33977 14467
rect 33152 14436 33977 14464
rect 28721 14399 28779 14405
rect 28721 14396 28733 14399
rect 28132 14368 28733 14396
rect 28132 14356 28138 14368
rect 28721 14365 28733 14368
rect 28767 14365 28779 14399
rect 28721 14359 28779 14365
rect 23164 14300 27200 14328
rect 23164 14288 23170 14300
rect 21174 14260 21180 14272
rect 21135 14232 21180 14260
rect 21174 14220 21180 14232
rect 21232 14220 21238 14272
rect 23477 14263 23535 14269
rect 23477 14229 23489 14263
rect 23523 14260 23535 14263
rect 24026 14260 24032 14272
rect 23523 14232 24032 14260
rect 23523 14229 23535 14232
rect 23477 14223 23535 14229
rect 24026 14220 24032 14232
rect 24084 14220 24090 14272
rect 31941 14263 31999 14269
rect 31941 14229 31953 14263
rect 31987 14260 31999 14263
rect 32306 14260 32312 14272
rect 31987 14232 32312 14260
rect 31987 14229 31999 14232
rect 31941 14223 31999 14229
rect 32306 14220 32312 14232
rect 32364 14220 32370 14272
rect 32766 14260 32772 14272
rect 32727 14232 32772 14260
rect 32766 14220 32772 14232
rect 32824 14220 32830 14272
rect 33152 14269 33180 14436
rect 33965 14433 33977 14436
rect 34011 14464 34023 14467
rect 34422 14464 34428 14476
rect 34011 14436 34428 14464
rect 34011 14433 34023 14436
rect 33965 14427 34023 14433
rect 34422 14424 34428 14436
rect 34480 14424 34486 14476
rect 33229 14399 33287 14405
rect 33229 14365 33241 14399
rect 33275 14396 33287 14399
rect 33594 14396 33600 14408
rect 33275 14368 33600 14396
rect 33275 14365 33287 14368
rect 33229 14359 33287 14365
rect 33594 14356 33600 14368
rect 33652 14356 33658 14408
rect 33778 14405 33784 14408
rect 33735 14399 33784 14405
rect 33735 14365 33747 14399
rect 33781 14365 33784 14399
rect 33735 14359 33784 14365
rect 33778 14356 33784 14359
rect 33836 14396 33842 14408
rect 36170 14396 36176 14408
rect 33836 14368 36176 14396
rect 33836 14356 33842 14368
rect 36170 14356 36176 14368
rect 36228 14356 36234 14408
rect 36446 14396 36452 14408
rect 36407 14368 36452 14396
rect 36446 14356 36452 14368
rect 36504 14356 36510 14408
rect 33137 14263 33195 14269
rect 33137 14229 33149 14263
rect 33183 14260 33195 14263
rect 33226 14260 33232 14272
rect 33183 14232 33232 14260
rect 33183 14229 33195 14232
rect 33137 14223 33195 14229
rect 33226 14220 33232 14232
rect 33284 14220 33290 14272
rect 35894 14260 35900 14272
rect 35855 14232 35900 14260
rect 35894 14220 35900 14232
rect 35952 14220 35958 14272
rect 1104 14170 38824 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 34966 14170
rect 35018 14118 35030 14170
rect 35082 14118 35094 14170
rect 35146 14118 35158 14170
rect 35210 14118 38824 14170
rect 1104 14096 38824 14118
rect 22741 14059 22799 14065
rect 22741 14025 22753 14059
rect 22787 14056 22799 14059
rect 23106 14056 23112 14068
rect 22787 14028 23112 14056
rect 22787 14025 22799 14028
rect 22741 14019 22799 14025
rect 23106 14016 23112 14028
rect 23164 14016 23170 14068
rect 23842 14016 23848 14068
rect 23900 14056 23906 14068
rect 25041 14059 25099 14065
rect 25041 14056 25053 14059
rect 23900 14028 25053 14056
rect 23900 14016 23906 14028
rect 25041 14025 25053 14028
rect 25087 14025 25099 14059
rect 25041 14019 25099 14025
rect 26142 14016 26148 14068
rect 26200 14056 26206 14068
rect 26605 14059 26663 14065
rect 26605 14056 26617 14059
rect 26200 14028 26617 14056
rect 26200 14016 26206 14028
rect 26605 14025 26617 14028
rect 26651 14056 26663 14059
rect 26970 14056 26976 14068
rect 26651 14028 26976 14056
rect 26651 14025 26663 14028
rect 26605 14019 26663 14025
rect 26970 14016 26976 14028
rect 27028 14016 27034 14068
rect 27798 14016 27804 14068
rect 27856 14056 27862 14068
rect 28077 14059 28135 14065
rect 28077 14056 28089 14059
rect 27856 14028 28089 14056
rect 27856 14016 27862 14028
rect 28077 14025 28089 14028
rect 28123 14025 28135 14059
rect 28718 14056 28724 14068
rect 28679 14028 28724 14056
rect 28077 14019 28135 14025
rect 28718 14016 28724 14028
rect 28776 14056 28782 14068
rect 28994 14056 29000 14068
rect 28776 14028 29000 14056
rect 28776 14016 28782 14028
rect 28994 14016 29000 14028
rect 29052 14016 29058 14068
rect 29641 14059 29699 14065
rect 29641 14025 29653 14059
rect 29687 14056 29699 14059
rect 30006 14056 30012 14068
rect 29687 14028 30012 14056
rect 29687 14025 29699 14028
rect 29641 14019 29699 14025
rect 30006 14016 30012 14028
rect 30064 14016 30070 14068
rect 31849 14059 31907 14065
rect 31849 14025 31861 14059
rect 31895 14056 31907 14059
rect 32674 14056 32680 14068
rect 31895 14028 32680 14056
rect 31895 14025 31907 14028
rect 31849 14019 31907 14025
rect 32674 14016 32680 14028
rect 32732 14056 32738 14068
rect 33594 14056 33600 14068
rect 32732 14028 33600 14056
rect 32732 14016 32738 14028
rect 33594 14016 33600 14028
rect 33652 14016 33658 14068
rect 33870 14016 33876 14068
rect 33928 14056 33934 14068
rect 34241 14059 34299 14065
rect 34241 14056 34253 14059
rect 33928 14028 34253 14056
rect 33928 14016 33934 14028
rect 34241 14025 34253 14028
rect 34287 14025 34299 14059
rect 34241 14019 34299 14025
rect 35345 14059 35403 14065
rect 35345 14025 35357 14059
rect 35391 14056 35403 14059
rect 36078 14056 36084 14068
rect 35391 14028 36084 14056
rect 35391 14025 35403 14028
rect 35345 14019 35403 14025
rect 36078 14016 36084 14028
rect 36136 14016 36142 14068
rect 36446 14016 36452 14068
rect 36504 14056 36510 14068
rect 37369 14059 37427 14065
rect 37369 14056 37381 14059
rect 36504 14028 37381 14056
rect 36504 14016 36510 14028
rect 37369 14025 37381 14028
rect 37415 14025 37427 14059
rect 37369 14019 37427 14025
rect 36814 13988 36820 14000
rect 36775 13960 36820 13988
rect 36814 13948 36820 13960
rect 36872 13948 36878 14000
rect 33778 13880 33784 13932
rect 33836 13920 33842 13932
rect 34609 13923 34667 13929
rect 34609 13920 34621 13923
rect 33836 13892 34621 13920
rect 33836 13880 33842 13892
rect 34609 13889 34621 13892
rect 34655 13889 34667 13923
rect 34609 13883 34667 13889
rect 23658 13852 23664 13864
rect 23619 13824 23664 13852
rect 23658 13812 23664 13824
rect 23716 13812 23722 13864
rect 23934 13861 23940 13864
rect 23917 13855 23940 13861
rect 23917 13852 23929 13855
rect 23768 13824 23929 13852
rect 23768 13784 23796 13824
rect 23917 13821 23929 13824
rect 23992 13852 23998 13864
rect 25869 13855 25927 13861
rect 23992 13824 24065 13852
rect 23917 13815 23940 13821
rect 23934 13812 23940 13815
rect 23992 13812 23998 13824
rect 25869 13821 25881 13855
rect 25915 13852 25927 13855
rect 26694 13852 26700 13864
rect 25915 13824 26280 13852
rect 26607 13824 26700 13852
rect 25915 13821 25927 13824
rect 25869 13815 25927 13821
rect 26252 13793 26280 13824
rect 26694 13812 26700 13824
rect 26752 13852 26758 13864
rect 28074 13852 28080 13864
rect 26752 13824 28080 13852
rect 26752 13812 26758 13824
rect 28074 13812 28080 13824
rect 28132 13812 28138 13864
rect 30006 13861 30012 13864
rect 29733 13855 29791 13861
rect 29733 13821 29745 13855
rect 29779 13821 29791 13855
rect 30000 13852 30012 13861
rect 29967 13824 30012 13852
rect 29733 13815 29791 13821
rect 30000 13815 30012 13824
rect 23400 13756 23796 13784
rect 26237 13787 26295 13793
rect 23014 13716 23020 13728
rect 22975 13688 23020 13716
rect 23014 13676 23020 13688
rect 23072 13716 23078 13728
rect 23400 13725 23428 13756
rect 26237 13753 26249 13787
rect 26283 13784 26295 13787
rect 26964 13787 27022 13793
rect 26964 13784 26976 13787
rect 26283 13756 26976 13784
rect 26283 13753 26295 13756
rect 26237 13747 26295 13753
rect 26964 13753 26976 13756
rect 27010 13784 27022 13787
rect 27062 13784 27068 13796
rect 27010 13756 27068 13784
rect 27010 13753 27022 13756
rect 26964 13747 27022 13753
rect 27062 13744 27068 13756
rect 27120 13744 27126 13796
rect 29748 13784 29776 13815
rect 30006 13812 30012 13815
rect 30064 13812 30070 13864
rect 32306 13852 32312 13864
rect 32219 13824 32312 13852
rect 32306 13812 32312 13824
rect 32364 13852 32370 13864
rect 35250 13852 35256 13864
rect 32364 13824 35256 13852
rect 32364 13812 32370 13824
rect 35250 13812 35256 13824
rect 35308 13852 35314 13864
rect 35437 13855 35495 13861
rect 35437 13852 35449 13855
rect 35308 13824 35449 13852
rect 35308 13812 35314 13824
rect 35437 13821 35449 13824
rect 35483 13821 35495 13855
rect 35437 13815 35495 13821
rect 35526 13812 35532 13864
rect 35584 13852 35590 13864
rect 35693 13855 35751 13861
rect 35693 13852 35705 13855
rect 35584 13824 35705 13852
rect 35584 13812 35590 13824
rect 35693 13821 35705 13824
rect 35739 13821 35751 13855
rect 35693 13815 35751 13821
rect 30282 13784 30288 13796
rect 29748 13756 30288 13784
rect 30282 13744 30288 13756
rect 30340 13744 30346 13796
rect 32554 13787 32612 13793
rect 32554 13784 32566 13787
rect 32140 13756 32566 13784
rect 32140 13728 32168 13756
rect 32554 13753 32566 13756
rect 32600 13753 32612 13787
rect 32554 13747 32612 13753
rect 23385 13719 23443 13725
rect 23385 13716 23397 13719
rect 23072 13688 23397 13716
rect 23072 13676 23078 13688
rect 23385 13685 23397 13688
rect 23431 13685 23443 13719
rect 23385 13679 23443 13685
rect 30926 13676 30932 13728
rect 30984 13716 30990 13728
rect 31113 13719 31171 13725
rect 31113 13716 31125 13719
rect 30984 13688 31125 13716
rect 30984 13676 30990 13688
rect 31113 13685 31125 13688
rect 31159 13685 31171 13719
rect 32122 13716 32128 13728
rect 32083 13688 32128 13716
rect 31113 13679 31171 13685
rect 32122 13676 32128 13688
rect 32180 13676 32186 13728
rect 33686 13716 33692 13728
rect 33647 13688 33692 13716
rect 33686 13676 33692 13688
rect 33744 13676 33750 13728
rect 34790 13676 34796 13728
rect 34848 13716 34854 13728
rect 35342 13716 35348 13728
rect 34848 13688 35348 13716
rect 34848 13676 34854 13688
rect 35342 13676 35348 13688
rect 35400 13676 35406 13728
rect 1104 13626 38824 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 38824 13626
rect 1104 13552 38824 13574
rect 23569 13515 23627 13521
rect 23569 13481 23581 13515
rect 23615 13512 23627 13515
rect 23842 13512 23848 13524
rect 23615 13484 23848 13512
rect 23615 13481 23627 13484
rect 23569 13475 23627 13481
rect 23842 13472 23848 13484
rect 23900 13472 23906 13524
rect 25317 13515 25375 13521
rect 25317 13481 25329 13515
rect 25363 13512 25375 13515
rect 25590 13512 25596 13524
rect 25363 13484 25596 13512
rect 25363 13481 25375 13484
rect 25317 13475 25375 13481
rect 25590 13472 25596 13484
rect 25648 13512 25654 13524
rect 26142 13512 26148 13524
rect 25648 13484 26148 13512
rect 25648 13472 25654 13484
rect 26142 13472 26148 13484
rect 26200 13472 26206 13524
rect 27157 13515 27215 13521
rect 27157 13481 27169 13515
rect 27203 13512 27215 13515
rect 27338 13512 27344 13524
rect 27203 13484 27344 13512
rect 27203 13481 27215 13484
rect 27157 13475 27215 13481
rect 27338 13472 27344 13484
rect 27396 13472 27402 13524
rect 28994 13512 29000 13524
rect 28955 13484 29000 13512
rect 28994 13472 29000 13484
rect 29052 13472 29058 13524
rect 29641 13515 29699 13521
rect 29641 13481 29653 13515
rect 29687 13512 29699 13515
rect 30009 13515 30067 13521
rect 30009 13512 30021 13515
rect 29687 13484 30021 13512
rect 29687 13481 29699 13484
rect 29641 13475 29699 13481
rect 30009 13481 30021 13484
rect 30055 13512 30067 13515
rect 30282 13512 30288 13524
rect 30055 13484 30288 13512
rect 30055 13481 30067 13484
rect 30009 13475 30067 13481
rect 30282 13472 30288 13484
rect 30340 13472 30346 13524
rect 30466 13512 30472 13524
rect 30379 13484 30472 13512
rect 30466 13472 30472 13484
rect 30524 13512 30530 13524
rect 30742 13512 30748 13524
rect 30524 13484 30748 13512
rect 30524 13472 30530 13484
rect 30742 13472 30748 13484
rect 30800 13472 30806 13524
rect 31205 13515 31263 13521
rect 31205 13481 31217 13515
rect 31251 13512 31263 13515
rect 31941 13515 31999 13521
rect 31941 13512 31953 13515
rect 31251 13484 31953 13512
rect 31251 13481 31263 13484
rect 31205 13475 31263 13481
rect 31941 13481 31953 13484
rect 31987 13512 31999 13515
rect 32306 13512 32312 13524
rect 31987 13484 32312 13512
rect 31987 13481 31999 13484
rect 31941 13475 31999 13481
rect 23860 13444 23888 13472
rect 24182 13447 24240 13453
rect 24182 13444 24194 13447
rect 23860 13416 24194 13444
rect 24182 13413 24194 13416
rect 24228 13444 24240 13447
rect 24670 13444 24676 13456
rect 24228 13416 24676 13444
rect 24228 13413 24240 13416
rect 24182 13407 24240 13413
rect 24670 13404 24676 13416
rect 24728 13404 24734 13456
rect 27798 13404 27804 13456
rect 27856 13453 27862 13456
rect 27856 13447 27920 13453
rect 27856 13413 27874 13447
rect 27908 13413 27920 13447
rect 27856 13407 27920 13413
rect 27856 13404 27862 13407
rect 28074 13404 28080 13456
rect 28132 13404 28138 13456
rect 30650 13404 30656 13456
rect 30708 13444 30714 13456
rect 31220 13444 31248 13475
rect 32306 13472 32312 13484
rect 32364 13472 32370 13524
rect 32398 13472 32404 13524
rect 32456 13512 32462 13524
rect 32493 13515 32551 13521
rect 32493 13512 32505 13515
rect 32456 13484 32505 13512
rect 32456 13472 32462 13484
rect 32493 13481 32505 13484
rect 32539 13481 32551 13515
rect 32493 13475 32551 13481
rect 30708 13416 31248 13444
rect 30708 13404 30714 13416
rect 22741 13379 22799 13385
rect 22741 13345 22753 13379
rect 22787 13376 22799 13379
rect 23658 13376 23664 13388
rect 22787 13348 23664 13376
rect 22787 13345 22799 13348
rect 22741 13339 22799 13345
rect 23658 13336 23664 13348
rect 23716 13336 23722 13388
rect 23750 13336 23756 13388
rect 23808 13376 23814 13388
rect 23937 13379 23995 13385
rect 23937 13376 23949 13379
rect 23808 13348 23949 13376
rect 23808 13336 23814 13348
rect 23937 13345 23949 13348
rect 23983 13376 23995 13379
rect 24578 13376 24584 13388
rect 23983 13348 24584 13376
rect 23983 13345 23995 13348
rect 23937 13339 23995 13345
rect 24578 13336 24584 13348
rect 24636 13336 24642 13388
rect 26513 13379 26571 13385
rect 26513 13345 26525 13379
rect 26559 13376 26571 13379
rect 26602 13376 26608 13388
rect 26559 13348 26608 13376
rect 26559 13345 26571 13348
rect 26513 13339 26571 13345
rect 26602 13336 26608 13348
rect 26660 13336 26666 13388
rect 27525 13379 27583 13385
rect 27525 13345 27537 13379
rect 27571 13376 27583 13379
rect 27617 13379 27675 13385
rect 27617 13376 27629 13379
rect 27571 13348 27629 13376
rect 27571 13345 27583 13348
rect 27525 13339 27583 13345
rect 27617 13345 27629 13348
rect 27663 13376 27675 13379
rect 28092 13376 28120 13404
rect 27663 13348 28120 13376
rect 27663 13345 27675 13348
rect 27617 13339 27675 13345
rect 30374 13336 30380 13388
rect 30432 13376 30438 13388
rect 32508 13376 32536 13475
rect 32766 13472 32772 13524
rect 32824 13512 32830 13524
rect 33143 13515 33201 13521
rect 33143 13512 33155 13515
rect 32824 13484 33155 13512
rect 32824 13472 32830 13484
rect 33143 13481 33155 13484
rect 33189 13512 33201 13515
rect 33870 13512 33876 13524
rect 33189 13484 33876 13512
rect 33189 13481 33201 13484
rect 33143 13475 33201 13481
rect 33870 13472 33876 13484
rect 33928 13472 33934 13524
rect 34422 13472 34428 13524
rect 34480 13512 34486 13524
rect 34517 13515 34575 13521
rect 34517 13512 34529 13515
rect 34480 13484 34529 13512
rect 34480 13472 34486 13484
rect 34517 13481 34529 13484
rect 34563 13481 34575 13515
rect 34517 13475 34575 13481
rect 34790 13472 34796 13524
rect 34848 13512 34854 13524
rect 34885 13515 34943 13521
rect 34885 13512 34897 13515
rect 34848 13484 34897 13512
rect 34848 13472 34854 13484
rect 34885 13481 34897 13484
rect 34931 13512 34943 13515
rect 35250 13512 35256 13524
rect 34931 13484 35256 13512
rect 34931 13481 34943 13484
rect 34885 13475 34943 13481
rect 35250 13472 35256 13484
rect 35308 13472 35314 13524
rect 35802 13512 35808 13524
rect 35763 13484 35808 13512
rect 35802 13472 35808 13484
rect 35860 13472 35866 13524
rect 36170 13472 36176 13524
rect 36228 13512 36234 13524
rect 36449 13515 36507 13521
rect 36449 13512 36461 13515
rect 36228 13484 36461 13512
rect 36228 13472 36234 13484
rect 36449 13481 36461 13484
rect 36495 13481 36507 13515
rect 36449 13475 36507 13481
rect 35268 13444 35296 13472
rect 36817 13447 36875 13453
rect 36817 13444 36829 13447
rect 35268 13416 36829 13444
rect 36817 13413 36829 13416
rect 36863 13413 36875 13447
rect 36817 13407 36875 13413
rect 30432 13348 30696 13376
rect 32508 13348 33180 13376
rect 30432 13336 30438 13348
rect 22830 13308 22836 13320
rect 22791 13280 22836 13308
rect 22830 13268 22836 13280
rect 22888 13268 22894 13320
rect 23017 13311 23075 13317
rect 23017 13277 23029 13311
rect 23063 13308 23075 13311
rect 23106 13308 23112 13320
rect 23063 13280 23112 13308
rect 23063 13277 23075 13280
rect 23017 13271 23075 13277
rect 22281 13243 22339 13249
rect 22281 13209 22293 13243
rect 22327 13240 22339 13243
rect 23032 13240 23060 13271
rect 23106 13268 23112 13280
rect 23164 13268 23170 13320
rect 30558 13308 30564 13320
rect 30519 13280 30564 13308
rect 30558 13268 30564 13280
rect 30616 13268 30622 13320
rect 30668 13317 30696 13348
rect 30653 13311 30711 13317
rect 30653 13277 30665 13311
rect 30699 13277 30711 13311
rect 32674 13308 32680 13320
rect 32635 13280 32680 13308
rect 30653 13271 30711 13277
rect 32674 13268 32680 13280
rect 32732 13268 32738 13320
rect 33152 13317 33180 13348
rect 35526 13336 35532 13388
rect 35584 13376 35590 13388
rect 35584 13348 36032 13376
rect 35584 13336 35590 13348
rect 33140 13311 33198 13317
rect 33140 13277 33152 13311
rect 33186 13277 33198 13311
rect 33410 13308 33416 13320
rect 33371 13280 33416 13308
rect 33140 13271 33198 13277
rect 33410 13268 33416 13280
rect 33468 13268 33474 13320
rect 35894 13308 35900 13320
rect 35855 13280 35900 13308
rect 35894 13268 35900 13280
rect 35952 13268 35958 13320
rect 36004 13317 36032 13348
rect 35989 13311 36047 13317
rect 35989 13277 36001 13311
rect 36035 13308 36047 13311
rect 36078 13308 36084 13320
rect 36035 13280 36084 13308
rect 36035 13277 36047 13280
rect 35989 13271 36047 13277
rect 36078 13268 36084 13280
rect 36136 13268 36142 13320
rect 22327 13212 23060 13240
rect 22327 13209 22339 13212
rect 22281 13203 22339 13209
rect 34238 13200 34244 13252
rect 34296 13240 34302 13252
rect 35526 13240 35532 13252
rect 34296 13212 35532 13240
rect 34296 13200 34302 13212
rect 35526 13200 35532 13212
rect 35584 13200 35590 13252
rect 22370 13172 22376 13184
rect 22331 13144 22376 13172
rect 22370 13132 22376 13144
rect 22428 13132 22434 13184
rect 26697 13175 26755 13181
rect 26697 13141 26709 13175
rect 26743 13172 26755 13175
rect 27614 13172 27620 13184
rect 26743 13144 27620 13172
rect 26743 13141 26755 13144
rect 26697 13135 26755 13141
rect 27614 13132 27620 13144
rect 27672 13132 27678 13184
rect 30006 13132 30012 13184
rect 30064 13172 30070 13184
rect 30101 13175 30159 13181
rect 30101 13172 30113 13175
rect 30064 13144 30113 13172
rect 30064 13132 30070 13144
rect 30101 13141 30113 13144
rect 30147 13141 30159 13175
rect 35250 13172 35256 13184
rect 35211 13144 35256 13172
rect 30101 13135 30159 13141
rect 35250 13132 35256 13144
rect 35308 13132 35314 13184
rect 35437 13175 35495 13181
rect 35437 13141 35449 13175
rect 35483 13172 35495 13175
rect 35986 13172 35992 13184
rect 35483 13144 35992 13172
rect 35483 13141 35495 13144
rect 35437 13135 35495 13141
rect 35986 13132 35992 13144
rect 36044 13132 36050 13184
rect 1104 13082 38824 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 34966 13082
rect 35018 13030 35030 13082
rect 35082 13030 35094 13082
rect 35146 13030 35158 13082
rect 35210 13030 38824 13082
rect 1104 13008 38824 13030
rect 22465 12971 22523 12977
rect 22465 12937 22477 12971
rect 22511 12968 22523 12971
rect 23014 12968 23020 12980
rect 22511 12940 23020 12968
rect 22511 12937 22523 12940
rect 22465 12931 22523 12937
rect 23014 12928 23020 12940
rect 23072 12928 23078 12980
rect 24670 12968 24676 12980
rect 24631 12940 24676 12968
rect 24670 12928 24676 12940
rect 24728 12928 24734 12980
rect 25590 12968 25596 12980
rect 25551 12940 25596 12968
rect 25590 12928 25596 12940
rect 25648 12928 25654 12980
rect 27062 12968 27068 12980
rect 27023 12940 27068 12968
rect 27062 12928 27068 12940
rect 27120 12928 27126 12980
rect 27709 12971 27767 12977
rect 27709 12937 27721 12971
rect 27755 12968 27767 12971
rect 27798 12968 27804 12980
rect 27755 12940 27804 12968
rect 27755 12937 27767 12940
rect 27709 12931 27767 12937
rect 27798 12928 27804 12940
rect 27856 12928 27862 12980
rect 28074 12968 28080 12980
rect 28035 12940 28080 12968
rect 28074 12928 28080 12940
rect 28132 12928 28138 12980
rect 30190 12968 30196 12980
rect 30103 12940 30196 12968
rect 30190 12928 30196 12940
rect 30248 12968 30254 12980
rect 30558 12968 30564 12980
rect 30248 12940 30564 12968
rect 30248 12928 30254 12940
rect 30558 12928 30564 12940
rect 30616 12928 30622 12980
rect 32766 12968 32772 12980
rect 32727 12940 32772 12968
rect 32766 12928 32772 12940
rect 32824 12928 32830 12980
rect 33042 12928 33048 12980
rect 33100 12968 33106 12980
rect 33137 12971 33195 12977
rect 33137 12968 33149 12971
rect 33100 12940 33149 12968
rect 33100 12928 33106 12940
rect 33137 12937 33149 12940
rect 33183 12937 33195 12971
rect 33137 12931 33195 12937
rect 34701 12971 34759 12977
rect 34701 12937 34713 12971
rect 34747 12968 34759 12971
rect 35802 12968 35808 12980
rect 34747 12940 35808 12968
rect 34747 12937 34759 12940
rect 34701 12931 34759 12937
rect 35802 12928 35808 12940
rect 35860 12928 35866 12980
rect 35894 12928 35900 12980
rect 35952 12968 35958 12980
rect 37093 12971 37151 12977
rect 37093 12968 37105 12971
rect 35952 12940 37105 12968
rect 35952 12928 35958 12940
rect 37093 12937 37105 12940
rect 37139 12937 37151 12971
rect 37093 12931 37151 12937
rect 23661 12903 23719 12909
rect 23661 12869 23673 12903
rect 23707 12900 23719 12903
rect 24854 12900 24860 12912
rect 23707 12872 24860 12900
rect 23707 12869 23719 12872
rect 23661 12863 23719 12869
rect 24854 12860 24860 12872
rect 24912 12860 24918 12912
rect 22370 12792 22376 12844
rect 22428 12832 22434 12844
rect 24118 12832 24124 12844
rect 22428 12804 24124 12832
rect 22428 12792 22434 12804
rect 24118 12792 24124 12804
rect 24176 12792 24182 12844
rect 24305 12835 24363 12841
rect 24305 12801 24317 12835
rect 24351 12832 24363 12835
rect 24578 12832 24584 12844
rect 24351 12804 24584 12832
rect 24351 12801 24363 12804
rect 24305 12795 24363 12801
rect 24578 12792 24584 12804
rect 24636 12792 24642 12844
rect 25608 12832 25636 12928
rect 29733 12903 29791 12909
rect 29733 12869 29745 12903
rect 29779 12900 29791 12903
rect 30374 12900 30380 12912
rect 29779 12872 30380 12900
rect 29779 12869 29791 12872
rect 29733 12863 29791 12869
rect 30374 12860 30380 12872
rect 30432 12860 30438 12912
rect 30466 12860 30472 12912
rect 30524 12900 30530 12912
rect 30524 12872 30569 12900
rect 30524 12860 30530 12872
rect 33870 12860 33876 12912
rect 33928 12900 33934 12912
rect 33928 12872 34836 12900
rect 33928 12860 33934 12872
rect 34808 12844 34836 12872
rect 36446 12860 36452 12912
rect 36504 12900 36510 12912
rect 36541 12903 36599 12909
rect 36541 12900 36553 12903
rect 36504 12872 36553 12900
rect 36504 12860 36510 12872
rect 36541 12869 36553 12872
rect 36587 12869 36599 12903
rect 36541 12863 36599 12869
rect 30650 12832 30656 12844
rect 25608 12804 25820 12832
rect 30611 12804 30656 12832
rect 21085 12767 21143 12773
rect 21085 12733 21097 12767
rect 21131 12764 21143 12767
rect 21174 12764 21180 12776
rect 21131 12736 21180 12764
rect 21131 12733 21143 12736
rect 21085 12727 21143 12733
rect 21174 12724 21180 12736
rect 21232 12724 21238 12776
rect 24026 12764 24032 12776
rect 23987 12736 24032 12764
rect 24026 12724 24032 12736
rect 24084 12764 24090 12776
rect 25041 12767 25099 12773
rect 25041 12764 25053 12767
rect 24084 12736 25053 12764
rect 24084 12724 24090 12736
rect 25041 12733 25053 12736
rect 25087 12733 25099 12767
rect 25682 12764 25688 12776
rect 25643 12736 25688 12764
rect 25041 12727 25099 12733
rect 25682 12724 25688 12736
rect 25740 12724 25746 12776
rect 25792 12764 25820 12804
rect 30650 12792 30656 12804
rect 30708 12792 30714 12844
rect 33778 12832 33784 12844
rect 33739 12804 33784 12832
rect 33778 12792 33784 12804
rect 33836 12792 33842 12844
rect 34330 12792 34336 12844
rect 34388 12832 34394 12844
rect 34388 12804 34560 12832
rect 34388 12792 34394 12804
rect 25941 12767 25999 12773
rect 25941 12764 25953 12767
rect 25792 12736 25953 12764
rect 25941 12733 25953 12736
rect 25987 12733 25999 12767
rect 25941 12727 25999 12733
rect 29549 12767 29607 12773
rect 29549 12733 29561 12767
rect 29595 12764 29607 12767
rect 29638 12764 29644 12776
rect 29595 12736 29644 12764
rect 29595 12733 29607 12736
rect 29549 12727 29607 12733
rect 29638 12724 29644 12736
rect 29696 12764 29702 12776
rect 30006 12764 30012 12776
rect 29696 12736 30012 12764
rect 29696 12724 29702 12736
rect 30006 12724 30012 12736
rect 30064 12724 30070 12776
rect 30926 12773 30932 12776
rect 30920 12764 30932 12773
rect 30887 12736 30932 12764
rect 30920 12727 30932 12736
rect 30926 12724 30932 12727
rect 30984 12724 30990 12776
rect 20993 12699 21051 12705
rect 20993 12665 21005 12699
rect 21039 12696 21051 12699
rect 21330 12699 21388 12705
rect 21330 12696 21342 12699
rect 21039 12668 21342 12696
rect 21039 12665 21051 12668
rect 20993 12659 21051 12665
rect 21330 12665 21342 12668
rect 21376 12696 21388 12699
rect 21376 12668 22140 12696
rect 21376 12665 21388 12668
rect 21330 12659 21388 12665
rect 22112 12628 22140 12668
rect 22370 12656 22376 12708
rect 22428 12696 22434 12708
rect 22830 12696 22836 12708
rect 22428 12668 22836 12696
rect 22428 12656 22434 12668
rect 22830 12656 22836 12668
rect 22888 12696 22894 12708
rect 23017 12699 23075 12705
rect 23017 12696 23029 12699
rect 22888 12668 23029 12696
rect 22888 12656 22894 12668
rect 23017 12665 23029 12668
rect 23063 12665 23075 12699
rect 23017 12659 23075 12665
rect 33134 12656 33140 12708
rect 33192 12696 33198 12708
rect 33410 12696 33416 12708
rect 33192 12668 33416 12696
rect 33192 12656 33198 12668
rect 33410 12656 33416 12668
rect 33468 12696 33474 12708
rect 33505 12699 33563 12705
rect 33505 12696 33517 12699
rect 33468 12668 33517 12696
rect 33468 12656 33474 12668
rect 33505 12665 33517 12668
rect 33551 12696 33563 12699
rect 33551 12668 34284 12696
rect 33551 12665 33563 12668
rect 33505 12659 33563 12665
rect 23477 12631 23535 12637
rect 23477 12628 23489 12631
rect 22112 12600 23489 12628
rect 23477 12597 23489 12600
rect 23523 12628 23535 12631
rect 23658 12628 23664 12640
rect 23523 12600 23664 12628
rect 23523 12597 23535 12600
rect 23477 12591 23535 12597
rect 23658 12588 23664 12600
rect 23716 12588 23722 12640
rect 31754 12588 31760 12640
rect 31812 12628 31818 12640
rect 32033 12631 32091 12637
rect 32033 12628 32045 12631
rect 31812 12600 32045 12628
rect 31812 12588 31818 12600
rect 32033 12597 32045 12600
rect 32079 12628 32091 12631
rect 32122 12628 32128 12640
rect 32079 12600 32128 12628
rect 32079 12597 32091 12600
rect 32033 12591 32091 12597
rect 32122 12588 32128 12600
rect 32180 12588 32186 12640
rect 33594 12588 33600 12640
rect 33652 12628 33658 12640
rect 33652 12600 33697 12628
rect 33652 12588 33658 12600
rect 33778 12588 33784 12640
rect 33836 12628 33842 12640
rect 34146 12628 34152 12640
rect 33836 12600 34152 12628
rect 33836 12588 33842 12600
rect 34146 12588 34152 12600
rect 34204 12588 34210 12640
rect 34256 12637 34284 12668
rect 34532 12640 34560 12804
rect 34790 12792 34796 12844
rect 34848 12832 34854 12844
rect 35161 12835 35219 12841
rect 35161 12832 35173 12835
rect 34848 12804 35173 12832
rect 34848 12792 34854 12804
rect 35161 12801 35173 12804
rect 35207 12801 35219 12835
rect 35161 12795 35219 12801
rect 35250 12724 35256 12776
rect 35308 12764 35314 12776
rect 35417 12767 35475 12773
rect 35417 12764 35429 12767
rect 35308 12736 35429 12764
rect 35308 12724 35314 12736
rect 35417 12733 35429 12736
rect 35463 12764 35475 12767
rect 35710 12764 35716 12776
rect 35463 12736 35716 12764
rect 35463 12733 35475 12736
rect 35417 12727 35475 12733
rect 35710 12724 35716 12736
rect 35768 12724 35774 12776
rect 34241 12631 34299 12637
rect 34241 12597 34253 12631
rect 34287 12628 34299 12631
rect 34422 12628 34428 12640
rect 34287 12600 34428 12628
rect 34287 12597 34299 12600
rect 34241 12591 34299 12597
rect 34422 12588 34428 12600
rect 34480 12588 34486 12640
rect 34514 12588 34520 12640
rect 34572 12588 34578 12640
rect 1104 12538 38824 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 38824 12538
rect 1104 12464 38824 12486
rect 23658 12424 23664 12436
rect 23619 12396 23664 12424
rect 23658 12384 23664 12396
rect 23716 12384 23722 12436
rect 24118 12384 24124 12436
rect 24176 12424 24182 12436
rect 24213 12427 24271 12433
rect 24213 12424 24225 12427
rect 24176 12396 24225 12424
rect 24176 12384 24182 12396
rect 24213 12393 24225 12396
rect 24259 12393 24271 12427
rect 24213 12387 24271 12393
rect 26602 12384 26608 12436
rect 26660 12424 26666 12436
rect 26697 12427 26755 12433
rect 26697 12424 26709 12427
rect 26660 12396 26709 12424
rect 26660 12384 26666 12396
rect 26697 12393 26709 12396
rect 26743 12393 26755 12427
rect 27430 12424 27436 12436
rect 27391 12396 27436 12424
rect 26697 12387 26755 12393
rect 27430 12384 27436 12396
rect 27488 12384 27494 12436
rect 29638 12424 29644 12436
rect 29599 12396 29644 12424
rect 29638 12384 29644 12396
rect 29696 12384 29702 12436
rect 30009 12427 30067 12433
rect 30009 12393 30021 12427
rect 30055 12424 30067 12427
rect 30282 12424 30288 12436
rect 30055 12396 30288 12424
rect 30055 12393 30067 12396
rect 30009 12387 30067 12393
rect 30282 12384 30288 12396
rect 30340 12384 30346 12436
rect 30374 12384 30380 12436
rect 30432 12424 30438 12436
rect 30561 12427 30619 12433
rect 30561 12424 30573 12427
rect 30432 12396 30573 12424
rect 30432 12384 30438 12396
rect 30561 12393 30573 12396
rect 30607 12393 30619 12427
rect 30561 12387 30619 12393
rect 32677 12427 32735 12433
rect 32677 12393 32689 12427
rect 32723 12424 32735 12427
rect 33134 12424 33140 12436
rect 32723 12396 33140 12424
rect 32723 12393 32735 12396
rect 32677 12387 32735 12393
rect 33134 12384 33140 12396
rect 33192 12384 33198 12436
rect 33318 12384 33324 12436
rect 33376 12424 33382 12436
rect 34238 12424 34244 12436
rect 33376 12396 34008 12424
rect 34199 12396 34244 12424
rect 33376 12384 33382 12396
rect 22370 12316 22376 12368
rect 22428 12356 22434 12368
rect 22526 12359 22584 12365
rect 22526 12356 22538 12359
rect 22428 12328 22538 12356
rect 22428 12316 22434 12328
rect 22526 12325 22538 12328
rect 22572 12325 22584 12359
rect 30190 12356 30196 12368
rect 22526 12319 22584 12325
rect 29012 12328 30196 12356
rect 29012 12300 29040 12328
rect 30190 12316 30196 12328
rect 30248 12316 30254 12368
rect 33781 12359 33839 12365
rect 33781 12356 33793 12359
rect 33612 12328 33793 12356
rect 33612 12300 33640 12328
rect 33781 12325 33793 12328
rect 33827 12325 33839 12359
rect 33980 12356 34008 12396
rect 34238 12384 34244 12396
rect 34296 12384 34302 12436
rect 34330 12384 34336 12436
rect 34388 12384 34394 12436
rect 36078 12384 36084 12436
rect 36136 12424 36142 12436
rect 36265 12427 36323 12433
rect 36265 12424 36277 12427
rect 36136 12396 36277 12424
rect 36136 12384 36142 12396
rect 36265 12393 36277 12396
rect 36311 12393 36323 12427
rect 36265 12387 36323 12393
rect 34348 12356 34376 12384
rect 33980 12328 34376 12356
rect 33781 12319 33839 12325
rect 24854 12248 24860 12300
rect 24912 12288 24918 12300
rect 25133 12291 25191 12297
rect 25133 12288 25145 12291
rect 24912 12260 25145 12288
rect 24912 12248 24918 12260
rect 25133 12257 25145 12260
rect 25179 12257 25191 12291
rect 25133 12251 25191 12257
rect 27614 12248 27620 12300
rect 27672 12288 27678 12300
rect 27798 12288 27804 12300
rect 27672 12260 27804 12288
rect 27672 12248 27678 12260
rect 27798 12248 27804 12260
rect 27856 12248 27862 12300
rect 28994 12288 29000 12300
rect 28907 12260 29000 12288
rect 28994 12248 29000 12260
rect 29052 12248 29058 12300
rect 30098 12248 30104 12300
rect 30156 12288 30162 12300
rect 30469 12291 30527 12297
rect 30469 12288 30481 12291
rect 30156 12260 30481 12288
rect 30156 12248 30162 12260
rect 30469 12257 30481 12260
rect 30515 12257 30527 12291
rect 33134 12288 33140 12300
rect 33095 12260 33140 12288
rect 30469 12251 30527 12257
rect 33134 12248 33140 12260
rect 33192 12288 33198 12300
rect 33594 12288 33600 12300
rect 33192 12260 33600 12288
rect 33192 12248 33198 12260
rect 33594 12248 33600 12260
rect 33652 12248 33658 12300
rect 33870 12248 33876 12300
rect 33928 12288 33934 12300
rect 34606 12297 34612 12300
rect 34333 12291 34391 12297
rect 34333 12288 34345 12291
rect 33928 12260 34345 12288
rect 33928 12248 33934 12260
rect 34333 12257 34345 12260
rect 34379 12257 34391 12291
rect 34333 12251 34391 12257
rect 34600 12251 34612 12297
rect 34664 12288 34670 12300
rect 34664 12260 34700 12288
rect 34606 12248 34612 12251
rect 34664 12248 34670 12260
rect 21174 12220 21180 12232
rect 21087 12192 21180 12220
rect 21174 12180 21180 12192
rect 21232 12220 21238 12232
rect 22278 12220 22284 12232
rect 21232 12192 22284 12220
rect 21232 12180 21238 12192
rect 22278 12180 22284 12192
rect 22336 12180 22342 12232
rect 26602 12220 26608 12232
rect 25332 12192 26608 12220
rect 25332 12161 25360 12192
rect 26602 12180 26608 12192
rect 26660 12220 26666 12232
rect 27893 12223 27951 12229
rect 27893 12220 27905 12223
rect 26660 12192 27905 12220
rect 26660 12180 26666 12192
rect 27893 12189 27905 12192
rect 27939 12189 27951 12223
rect 28074 12220 28080 12232
rect 28035 12192 28080 12220
rect 27893 12183 27951 12189
rect 28074 12180 28080 12192
rect 28132 12180 28138 12232
rect 30650 12220 30656 12232
rect 30611 12192 30656 12220
rect 30650 12180 30656 12192
rect 30708 12220 30714 12232
rect 30926 12220 30932 12232
rect 30708 12192 30932 12220
rect 30708 12180 30714 12192
rect 30926 12180 30932 12192
rect 30984 12220 30990 12232
rect 31113 12223 31171 12229
rect 31113 12220 31125 12223
rect 30984 12192 31125 12220
rect 30984 12180 30990 12192
rect 31113 12189 31125 12192
rect 31159 12189 31171 12223
rect 33226 12220 33232 12232
rect 33187 12192 33232 12220
rect 31113 12183 31171 12189
rect 33226 12180 33232 12192
rect 33284 12180 33290 12232
rect 33413 12223 33471 12229
rect 33413 12189 33425 12223
rect 33459 12220 33471 12223
rect 33686 12220 33692 12232
rect 33459 12192 33692 12220
rect 33459 12189 33471 12192
rect 33413 12183 33471 12189
rect 33686 12180 33692 12192
rect 33744 12180 33750 12232
rect 25317 12155 25375 12161
rect 25317 12121 25329 12155
rect 25363 12121 25375 12155
rect 25317 12115 25375 12121
rect 27341 12155 27399 12161
rect 27341 12121 27353 12155
rect 27387 12152 27399 12155
rect 28092 12152 28120 12180
rect 27387 12124 28120 12152
rect 30101 12155 30159 12161
rect 27387 12121 27399 12124
rect 27341 12115 27399 12121
rect 30101 12121 30113 12155
rect 30147 12152 30159 12155
rect 31478 12152 31484 12164
rect 30147 12124 31484 12152
rect 30147 12121 30159 12124
rect 30101 12115 30159 12121
rect 31478 12112 31484 12124
rect 31536 12112 31542 12164
rect 32674 12152 32680 12164
rect 31956 12124 32680 12152
rect 31956 12096 31984 12124
rect 32674 12112 32680 12124
rect 32732 12112 32738 12164
rect 24578 12084 24584 12096
rect 24539 12056 24584 12084
rect 24578 12044 24584 12056
rect 24636 12044 24642 12096
rect 25041 12087 25099 12093
rect 25041 12053 25053 12087
rect 25087 12084 25099 12087
rect 25498 12084 25504 12096
rect 25087 12056 25504 12084
rect 25087 12053 25099 12056
rect 25041 12047 25099 12053
rect 25498 12044 25504 12056
rect 25556 12044 25562 12096
rect 25682 12084 25688 12096
rect 25643 12056 25688 12084
rect 25682 12044 25688 12056
rect 25740 12044 25746 12096
rect 29178 12084 29184 12096
rect 29139 12056 29184 12084
rect 29178 12044 29184 12056
rect 29236 12044 29242 12096
rect 31938 12084 31944 12096
rect 31899 12056 31944 12084
rect 31938 12044 31944 12056
rect 31996 12044 32002 12096
rect 32766 12084 32772 12096
rect 32727 12056 32772 12084
rect 32766 12044 32772 12056
rect 32824 12044 32830 12096
rect 33686 12044 33692 12096
rect 33744 12084 33750 12096
rect 34330 12084 34336 12096
rect 33744 12056 34336 12084
rect 33744 12044 33750 12056
rect 34330 12044 34336 12056
rect 34388 12084 34394 12096
rect 34606 12084 34612 12096
rect 34388 12056 34612 12084
rect 34388 12044 34394 12056
rect 34606 12044 34612 12056
rect 34664 12044 34670 12096
rect 35434 12044 35440 12096
rect 35492 12084 35498 12096
rect 35710 12084 35716 12096
rect 35492 12056 35716 12084
rect 35492 12044 35498 12056
rect 35710 12044 35716 12056
rect 35768 12044 35774 12096
rect 1104 11994 38824 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 34966 11994
rect 35018 11942 35030 11994
rect 35082 11942 35094 11994
rect 35146 11942 35158 11994
rect 35210 11942 38824 11994
rect 1104 11920 38824 11942
rect 24854 11840 24860 11892
rect 24912 11880 24918 11892
rect 25133 11883 25191 11889
rect 25133 11880 25145 11883
rect 24912 11852 25145 11880
rect 24912 11840 24918 11852
rect 25133 11849 25145 11852
rect 25179 11849 25191 11883
rect 25133 11843 25191 11849
rect 25498 11840 25504 11892
rect 25556 11880 25562 11892
rect 26694 11880 26700 11892
rect 25556 11852 26700 11880
rect 25556 11840 25562 11852
rect 26694 11840 26700 11852
rect 26752 11840 26758 11892
rect 27798 11840 27804 11892
rect 27856 11880 27862 11892
rect 28537 11883 28595 11889
rect 28537 11880 28549 11883
rect 27856 11852 28549 11880
rect 27856 11840 27862 11852
rect 28537 11849 28549 11852
rect 28583 11849 28595 11883
rect 28994 11880 29000 11892
rect 28955 11852 29000 11880
rect 28537 11843 28595 11849
rect 28994 11840 29000 11852
rect 29052 11840 29058 11892
rect 29178 11840 29184 11892
rect 29236 11880 29242 11892
rect 30098 11880 30104 11892
rect 29236 11852 30104 11880
rect 29236 11840 29242 11852
rect 30098 11840 30104 11852
rect 30156 11840 30162 11892
rect 30374 11840 30380 11892
rect 30432 11880 30438 11892
rect 30469 11883 30527 11889
rect 30469 11880 30481 11883
rect 30432 11852 30481 11880
rect 30432 11840 30438 11852
rect 30469 11849 30481 11852
rect 30515 11849 30527 11883
rect 30469 11843 30527 11849
rect 31297 11883 31355 11889
rect 31297 11849 31309 11883
rect 31343 11880 31355 11883
rect 32861 11883 32919 11889
rect 31343 11852 31984 11880
rect 31343 11849 31355 11852
rect 31297 11843 31355 11849
rect 22278 11772 22284 11824
rect 22336 11812 22342 11824
rect 22741 11815 22799 11821
rect 22741 11812 22753 11815
rect 22336 11784 22753 11812
rect 22336 11772 22342 11784
rect 22741 11781 22753 11784
rect 22787 11812 22799 11815
rect 23382 11812 23388 11824
rect 22787 11784 23388 11812
rect 22787 11781 22799 11784
rect 22741 11775 22799 11781
rect 23382 11772 23388 11784
rect 23440 11772 23446 11824
rect 26602 11812 26608 11824
rect 26563 11784 26608 11812
rect 26602 11772 26608 11784
rect 26660 11772 26666 11824
rect 27525 11815 27583 11821
rect 27525 11781 27537 11815
rect 27571 11812 27583 11815
rect 29012 11812 29040 11840
rect 27571 11784 29040 11812
rect 29825 11815 29883 11821
rect 27571 11781 27583 11784
rect 27525 11775 27583 11781
rect 29825 11781 29837 11815
rect 29871 11812 29883 11815
rect 30650 11812 30656 11824
rect 29871 11784 30656 11812
rect 29871 11781 29883 11784
rect 29825 11775 29883 11781
rect 30650 11772 30656 11784
rect 30708 11772 30714 11824
rect 23477 11747 23535 11753
rect 23477 11713 23489 11747
rect 23523 11744 23535 11747
rect 23658 11744 23664 11756
rect 23523 11716 23664 11744
rect 23523 11713 23535 11716
rect 23477 11707 23535 11713
rect 23658 11704 23664 11716
rect 23716 11744 23722 11756
rect 24213 11747 24271 11753
rect 24213 11744 24225 11747
rect 23716 11716 24225 11744
rect 23716 11704 23722 11716
rect 24213 11713 24225 11716
rect 24259 11713 24271 11747
rect 24213 11707 24271 11713
rect 24397 11747 24455 11753
rect 24397 11713 24409 11747
rect 24443 11744 24455 11747
rect 24857 11747 24915 11753
rect 24857 11744 24869 11747
rect 24443 11716 24869 11744
rect 24443 11713 24455 11716
rect 24397 11707 24455 11713
rect 24857 11713 24869 11716
rect 24903 11744 24915 11747
rect 27430 11744 27436 11756
rect 24903 11716 27436 11744
rect 24903 11713 24915 11716
rect 24857 11707 24915 11713
rect 22554 11636 22560 11688
rect 22612 11676 22618 11688
rect 24412 11676 24440 11707
rect 27430 11704 27436 11716
rect 27488 11704 27494 11756
rect 28074 11744 28080 11756
rect 28035 11716 28080 11744
rect 28074 11704 28080 11716
rect 28132 11704 28138 11756
rect 31478 11704 31484 11756
rect 31536 11744 31542 11756
rect 31757 11747 31815 11753
rect 31757 11744 31769 11747
rect 31536 11716 31769 11744
rect 31536 11704 31542 11716
rect 31757 11713 31769 11716
rect 31803 11713 31815 11747
rect 31757 11707 31815 11713
rect 31849 11747 31907 11753
rect 31849 11713 31861 11747
rect 31895 11713 31907 11747
rect 31956 11744 31984 11852
rect 32861 11849 32873 11883
rect 32907 11880 32919 11883
rect 33226 11880 33232 11892
rect 32907 11852 33232 11880
rect 32907 11849 32919 11852
rect 32861 11843 32919 11849
rect 33226 11840 33232 11852
rect 33284 11840 33290 11892
rect 33597 11883 33655 11889
rect 33597 11849 33609 11883
rect 33643 11880 33655 11883
rect 33686 11880 33692 11892
rect 33643 11852 33692 11880
rect 33643 11849 33655 11852
rect 33597 11843 33655 11849
rect 33686 11840 33692 11852
rect 33744 11840 33750 11892
rect 33870 11880 33876 11892
rect 33831 11852 33876 11880
rect 33870 11840 33876 11852
rect 33928 11840 33934 11892
rect 34330 11880 34336 11892
rect 34291 11852 34336 11880
rect 34330 11840 34336 11852
rect 34388 11840 34394 11892
rect 34606 11840 34612 11892
rect 34664 11880 34670 11892
rect 35342 11880 35348 11892
rect 34664 11852 35348 11880
rect 34664 11840 34670 11852
rect 35342 11840 35348 11852
rect 35400 11840 35406 11892
rect 35710 11840 35716 11892
rect 35768 11880 35774 11892
rect 36262 11880 36268 11892
rect 35768 11852 36268 11880
rect 35768 11840 35774 11852
rect 36262 11840 36268 11852
rect 36320 11840 36326 11892
rect 34885 11815 34943 11821
rect 34885 11781 34897 11815
rect 34931 11812 34943 11815
rect 35250 11812 35256 11824
rect 34931 11784 35256 11812
rect 34931 11781 34943 11784
rect 34885 11775 34943 11781
rect 35250 11772 35256 11784
rect 35308 11812 35314 11824
rect 36078 11812 36084 11824
rect 35308 11784 36084 11812
rect 35308 11772 35314 11784
rect 36078 11772 36084 11784
rect 36136 11772 36142 11824
rect 33134 11744 33140 11756
rect 31956 11716 33140 11744
rect 31849 11707 31907 11713
rect 26881 11679 26939 11685
rect 26881 11676 26893 11679
rect 22612 11648 24440 11676
rect 26252 11648 26893 11676
rect 22612 11636 22618 11648
rect 23109 11611 23167 11617
rect 23109 11577 23121 11611
rect 23155 11608 23167 11611
rect 23474 11608 23480 11620
rect 23155 11580 23480 11608
rect 23155 11577 23167 11580
rect 23109 11571 23167 11577
rect 23474 11568 23480 11580
rect 23532 11608 23538 11620
rect 24121 11611 24179 11617
rect 24121 11608 24133 11611
rect 23532 11580 24133 11608
rect 23532 11568 23538 11580
rect 24121 11577 24133 11580
rect 24167 11577 24179 11611
rect 24121 11571 24179 11577
rect 26252 11552 26280 11648
rect 26881 11645 26893 11648
rect 26927 11676 26939 11679
rect 27338 11676 27344 11688
rect 26927 11648 27344 11676
rect 26927 11645 26939 11648
rect 26881 11639 26939 11645
rect 27338 11636 27344 11648
rect 27396 11636 27402 11688
rect 31386 11636 31392 11688
rect 31444 11676 31450 11688
rect 31570 11676 31576 11688
rect 31444 11648 31576 11676
rect 31444 11636 31450 11648
rect 31570 11636 31576 11648
rect 31628 11676 31634 11688
rect 31864 11676 31892 11707
rect 33134 11704 33140 11716
rect 33192 11704 33198 11756
rect 35434 11744 35440 11756
rect 35395 11716 35440 11744
rect 35434 11704 35440 11716
rect 35492 11704 35498 11756
rect 35342 11676 35348 11688
rect 31628 11648 31892 11676
rect 35303 11648 35348 11676
rect 31628 11636 31634 11648
rect 35342 11636 35348 11648
rect 35400 11676 35406 11688
rect 35897 11679 35955 11685
rect 35897 11676 35909 11679
rect 35400 11648 35909 11676
rect 35400 11636 35406 11648
rect 35897 11645 35909 11648
rect 35943 11645 35955 11679
rect 35897 11639 35955 11645
rect 27433 11611 27491 11617
rect 27433 11577 27445 11611
rect 27479 11608 27491 11611
rect 27985 11611 28043 11617
rect 27985 11608 27997 11611
rect 27479 11580 27997 11608
rect 27479 11577 27491 11580
rect 27433 11571 27491 11577
rect 27985 11577 27997 11580
rect 28031 11608 28043 11611
rect 28718 11608 28724 11620
rect 28031 11580 28724 11608
rect 28031 11577 28043 11580
rect 27985 11571 28043 11577
rect 28718 11568 28724 11580
rect 28776 11568 28782 11620
rect 31205 11611 31263 11617
rect 31205 11577 31217 11611
rect 31251 11608 31263 11611
rect 31665 11611 31723 11617
rect 31665 11608 31677 11611
rect 31251 11580 31677 11608
rect 31251 11577 31263 11580
rect 31205 11571 31263 11577
rect 31665 11577 31677 11580
rect 31711 11608 31723 11611
rect 32122 11608 32128 11620
rect 31711 11580 32128 11608
rect 31711 11577 31723 11580
rect 31665 11571 31723 11577
rect 32122 11568 32128 11580
rect 32180 11568 32186 11620
rect 34701 11611 34759 11617
rect 34701 11577 34713 11611
rect 34747 11608 34759 11611
rect 35066 11608 35072 11620
rect 34747 11580 35072 11608
rect 34747 11577 34759 11580
rect 34701 11571 34759 11577
rect 35066 11568 35072 11580
rect 35124 11608 35130 11620
rect 35253 11611 35311 11617
rect 35253 11608 35265 11611
rect 35124 11580 35265 11608
rect 35124 11568 35130 11580
rect 35253 11577 35265 11580
rect 35299 11577 35311 11611
rect 35253 11571 35311 11577
rect 22370 11540 22376 11552
rect 22331 11512 22376 11540
rect 22370 11500 22376 11512
rect 22428 11500 22434 11552
rect 23750 11540 23756 11552
rect 23711 11512 23756 11540
rect 23750 11500 23756 11512
rect 23808 11500 23814 11552
rect 26234 11540 26240 11552
rect 26195 11512 26240 11540
rect 26234 11500 26240 11512
rect 26292 11500 26298 11552
rect 27890 11540 27896 11552
rect 27851 11512 27896 11540
rect 27890 11500 27896 11512
rect 27948 11500 27954 11552
rect 1104 11450 38824 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 38824 11450
rect 1104 11376 38824 11398
rect 22370 11296 22376 11348
rect 22428 11336 22434 11348
rect 23753 11339 23811 11345
rect 23753 11336 23765 11339
rect 22428 11308 23765 11336
rect 22428 11296 22434 11308
rect 23753 11305 23765 11308
rect 23799 11305 23811 11339
rect 23753 11299 23811 11305
rect 26789 11339 26847 11345
rect 26789 11305 26801 11339
rect 26835 11336 26847 11339
rect 27154 11336 27160 11348
rect 26835 11308 27160 11336
rect 26835 11305 26847 11308
rect 26789 11299 26847 11305
rect 27154 11296 27160 11308
rect 27212 11296 27218 11348
rect 28074 11296 28080 11348
rect 28132 11336 28138 11348
rect 28353 11339 28411 11345
rect 28353 11336 28365 11339
rect 28132 11308 28365 11336
rect 28132 11296 28138 11308
rect 28353 11305 28365 11308
rect 28399 11305 28411 11339
rect 28718 11336 28724 11348
rect 28679 11308 28724 11336
rect 28353 11299 28411 11305
rect 28718 11296 28724 11308
rect 28776 11296 28782 11348
rect 31386 11336 31392 11348
rect 31347 11308 31392 11336
rect 31386 11296 31392 11308
rect 31444 11296 31450 11348
rect 32122 11336 32128 11348
rect 32083 11308 32128 11336
rect 32122 11296 32128 11308
rect 32180 11296 32186 11348
rect 35066 11336 35072 11348
rect 35027 11308 35072 11336
rect 35066 11296 35072 11308
rect 35124 11296 35130 11348
rect 27433 11271 27491 11277
rect 27433 11237 27445 11271
rect 27479 11268 27491 11271
rect 27522 11268 27528 11280
rect 27479 11240 27528 11268
rect 27479 11237 27491 11240
rect 27433 11231 27491 11237
rect 27522 11228 27528 11240
rect 27580 11228 27586 11280
rect 34977 11271 35035 11277
rect 34977 11237 34989 11271
rect 35023 11268 35035 11271
rect 35434 11268 35440 11280
rect 35023 11240 35440 11268
rect 35023 11237 35035 11240
rect 34977 11231 35035 11237
rect 35434 11228 35440 11240
rect 35492 11228 35498 11280
rect 22373 11203 22431 11209
rect 22373 11169 22385 11203
rect 22419 11200 22431 11203
rect 22462 11200 22468 11212
rect 22419 11172 22468 11200
rect 22419 11169 22431 11172
rect 22373 11163 22431 11169
rect 22462 11160 22468 11172
rect 22520 11160 22526 11212
rect 22646 11209 22652 11212
rect 22640 11200 22652 11209
rect 22607 11172 22652 11200
rect 22640 11163 22652 11172
rect 22646 11160 22652 11163
rect 22704 11160 22710 11212
rect 25314 11200 25320 11212
rect 25275 11172 25320 11200
rect 25314 11160 25320 11172
rect 25372 11160 25378 11212
rect 26418 11160 26424 11212
rect 26476 11200 26482 11212
rect 27341 11203 27399 11209
rect 27341 11200 27353 11203
rect 26476 11172 27353 11200
rect 26476 11160 26482 11172
rect 27341 11169 27353 11172
rect 27387 11169 27399 11203
rect 28534 11200 28540 11212
rect 28495 11172 28540 11200
rect 27341 11163 27399 11169
rect 28534 11160 28540 11172
rect 28592 11160 28598 11212
rect 33870 11160 33876 11212
rect 33928 11200 33934 11212
rect 35529 11203 35587 11209
rect 35529 11200 35541 11203
rect 33928 11172 35541 11200
rect 33928 11160 33934 11172
rect 35452 11144 35480 11172
rect 35529 11169 35541 11172
rect 35575 11169 35587 11203
rect 35529 11163 35587 11169
rect 27430 11092 27436 11144
rect 27488 11132 27494 11144
rect 27525 11135 27583 11141
rect 27525 11132 27537 11135
rect 27488 11104 27537 11132
rect 27488 11092 27494 11104
rect 27525 11101 27537 11104
rect 27571 11101 27583 11135
rect 27525 11095 27583 11101
rect 35434 11092 35440 11144
rect 35492 11092 35498 11144
rect 25501 11067 25559 11073
rect 25501 11033 25513 11067
rect 25547 11064 25559 11067
rect 27890 11064 27896 11076
rect 25547 11036 27896 11064
rect 25547 11033 25559 11036
rect 25501 11027 25559 11033
rect 27890 11024 27896 11036
rect 27948 11064 27954 11076
rect 27985 11067 28043 11073
rect 27985 11064 27997 11067
rect 27948 11036 27997 11064
rect 27948 11024 27954 11036
rect 27985 11033 27997 11036
rect 28031 11033 28043 11067
rect 29178 11064 29184 11076
rect 29139 11036 29184 11064
rect 27985 11027 28043 11033
rect 29178 11024 29184 11036
rect 29236 11024 29242 11076
rect 22097 10999 22155 11005
rect 22097 10965 22109 10999
rect 22143 10996 22155 10999
rect 22554 10996 22560 11008
rect 22143 10968 22560 10996
rect 22143 10965 22155 10968
rect 22097 10959 22155 10965
rect 22554 10956 22560 10968
rect 22612 10956 22618 11008
rect 24302 10996 24308 11008
rect 24263 10968 24308 10996
rect 24302 10956 24308 10968
rect 24360 10956 24366 11008
rect 26970 10996 26976 11008
rect 26931 10968 26976 10996
rect 26970 10956 26976 10968
rect 27028 10956 27034 11008
rect 29917 10999 29975 11005
rect 29917 10965 29929 10999
rect 29963 10996 29975 10999
rect 30282 10996 30288 11008
rect 29963 10968 30288 10996
rect 29963 10965 29975 10968
rect 29917 10959 29975 10965
rect 30282 10956 30288 10968
rect 30340 10956 30346 11008
rect 1104 10906 38824 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 34966 10906
rect 35018 10854 35030 10906
rect 35082 10854 35094 10906
rect 35146 10854 35158 10906
rect 35210 10854 38824 10906
rect 1104 10832 38824 10854
rect 23477 10795 23535 10801
rect 23477 10761 23489 10795
rect 23523 10792 23535 10795
rect 23750 10792 23756 10804
rect 23523 10764 23756 10792
rect 23523 10761 23535 10764
rect 23477 10755 23535 10761
rect 23750 10752 23756 10764
rect 23808 10752 23814 10804
rect 27338 10752 27344 10804
rect 27396 10792 27402 10804
rect 28077 10795 28135 10801
rect 28077 10792 28089 10795
rect 27396 10764 28089 10792
rect 27396 10752 27402 10764
rect 28077 10761 28089 10764
rect 28123 10761 28135 10795
rect 28077 10755 28135 10761
rect 28258 10752 28264 10804
rect 28316 10792 28322 10804
rect 29641 10795 29699 10801
rect 29641 10792 29653 10795
rect 28316 10764 29653 10792
rect 28316 10752 28322 10764
rect 29641 10761 29653 10764
rect 29687 10792 29699 10795
rect 30098 10792 30104 10804
rect 29687 10764 30104 10792
rect 29687 10761 29699 10764
rect 29641 10755 29699 10761
rect 30098 10752 30104 10764
rect 30156 10752 30162 10804
rect 22554 10656 22560 10668
rect 22515 10628 22560 10656
rect 22554 10616 22560 10628
rect 22612 10616 22618 10668
rect 23768 10656 23796 10752
rect 23937 10727 23995 10733
rect 23937 10693 23949 10727
rect 23983 10724 23995 10727
rect 25314 10724 25320 10736
rect 23983 10696 25320 10724
rect 23983 10693 23995 10696
rect 23937 10687 23995 10693
rect 25314 10684 25320 10696
rect 25372 10684 25378 10736
rect 26513 10727 26571 10733
rect 26513 10693 26525 10727
rect 26559 10724 26571 10727
rect 28534 10724 28540 10736
rect 26559 10696 28540 10724
rect 26559 10693 26571 10696
rect 26513 10687 26571 10693
rect 28534 10684 28540 10696
rect 28592 10684 28598 10736
rect 24397 10659 24455 10665
rect 24397 10656 24409 10659
rect 23768 10628 24409 10656
rect 24397 10625 24409 10628
rect 24443 10625 24455 10659
rect 24578 10656 24584 10668
rect 24491 10628 24584 10656
rect 24397 10619 24455 10625
rect 24578 10616 24584 10628
rect 24636 10616 24642 10668
rect 26053 10659 26111 10665
rect 26053 10625 26065 10659
rect 26099 10656 26111 10659
rect 26970 10656 26976 10668
rect 26099 10628 26976 10656
rect 26099 10625 26111 10628
rect 26053 10619 26111 10625
rect 26970 10616 26976 10628
rect 27028 10616 27034 10668
rect 27154 10656 27160 10668
rect 27115 10628 27160 10656
rect 27154 10616 27160 10628
rect 27212 10616 27218 10668
rect 29089 10659 29147 10665
rect 29089 10625 29101 10659
rect 29135 10656 29147 10659
rect 30190 10656 30196 10668
rect 29135 10628 30196 10656
rect 29135 10625 29147 10628
rect 29089 10619 29147 10625
rect 30190 10616 30196 10628
rect 30248 10656 30254 10668
rect 30377 10659 30435 10665
rect 30377 10656 30389 10659
rect 30248 10628 30389 10656
rect 30248 10616 30254 10628
rect 30377 10625 30389 10628
rect 30423 10625 30435 10659
rect 35434 10656 35440 10668
rect 35395 10628 35440 10656
rect 30377 10619 30435 10625
rect 35434 10616 35440 10628
rect 35492 10616 35498 10668
rect 21913 10591 21971 10597
rect 21913 10557 21925 10591
rect 21959 10588 21971 10591
rect 22278 10588 22284 10600
rect 21959 10560 22284 10588
rect 21959 10557 21971 10560
rect 21913 10551 21971 10557
rect 22278 10548 22284 10560
rect 22336 10548 22342 10600
rect 22373 10591 22431 10597
rect 22373 10557 22385 10591
rect 22419 10588 22431 10591
rect 22646 10588 22652 10600
rect 22419 10560 22652 10588
rect 22419 10557 22431 10560
rect 22373 10551 22431 10557
rect 22646 10548 22652 10560
rect 22704 10588 22710 10600
rect 23106 10588 23112 10600
rect 22704 10560 23112 10588
rect 22704 10548 22710 10560
rect 23106 10548 23112 10560
rect 23164 10548 23170 10600
rect 24596 10588 24624 10616
rect 25041 10591 25099 10597
rect 25041 10588 25053 10591
rect 24596 10560 25053 10588
rect 25041 10557 25053 10560
rect 25087 10588 25099 10591
rect 27172 10588 27200 10616
rect 25087 10560 27200 10588
rect 28261 10591 28319 10597
rect 25087 10557 25099 10560
rect 25041 10551 25099 10557
rect 28261 10557 28273 10591
rect 28307 10588 28319 10591
rect 28902 10588 28908 10600
rect 28307 10560 28908 10588
rect 28307 10557 28319 10560
rect 28261 10551 28319 10557
rect 28902 10548 28908 10560
rect 28960 10548 28966 10600
rect 24302 10520 24308 10532
rect 22020 10492 24308 10520
rect 22020 10461 22048 10492
rect 24302 10480 24308 10492
rect 24360 10480 24366 10532
rect 27154 10480 27160 10532
rect 27212 10520 27218 10532
rect 27430 10520 27436 10532
rect 27212 10492 27436 10520
rect 27212 10480 27218 10492
rect 27430 10480 27436 10492
rect 27488 10520 27494 10532
rect 27893 10523 27951 10529
rect 27893 10520 27905 10523
rect 27488 10492 27905 10520
rect 27488 10480 27494 10492
rect 27893 10489 27905 10492
rect 27939 10489 27951 10523
rect 27893 10483 27951 10489
rect 30098 10480 30104 10532
rect 30156 10520 30162 10532
rect 30193 10523 30251 10529
rect 30193 10520 30205 10523
rect 30156 10492 30205 10520
rect 30156 10480 30162 10492
rect 30193 10489 30205 10492
rect 30239 10489 30251 10523
rect 30193 10483 30251 10489
rect 35345 10523 35403 10529
rect 35345 10489 35357 10523
rect 35391 10520 35403 10523
rect 35682 10523 35740 10529
rect 35682 10520 35694 10523
rect 35391 10492 35694 10520
rect 35391 10489 35403 10492
rect 35345 10483 35403 10489
rect 35682 10489 35694 10492
rect 35728 10520 35740 10523
rect 35802 10520 35808 10532
rect 35728 10492 35808 10520
rect 35728 10489 35740 10492
rect 35682 10483 35740 10489
rect 35802 10480 35808 10492
rect 35860 10480 35866 10532
rect 22005 10455 22063 10461
rect 22005 10421 22017 10455
rect 22051 10421 22063 10455
rect 22005 10415 22063 10421
rect 22278 10412 22284 10464
rect 22336 10452 22342 10464
rect 22465 10455 22523 10461
rect 22465 10452 22477 10455
rect 22336 10424 22477 10452
rect 22336 10412 22342 10424
rect 22465 10421 22477 10424
rect 22511 10452 22523 10455
rect 22922 10452 22928 10464
rect 22511 10424 22928 10452
rect 22511 10421 22523 10424
rect 22465 10415 22523 10421
rect 22922 10412 22928 10424
rect 22980 10412 22986 10464
rect 23106 10452 23112 10464
rect 23067 10424 23112 10452
rect 23106 10412 23112 10424
rect 23164 10412 23170 10464
rect 26418 10452 26424 10464
rect 26379 10424 26424 10452
rect 26418 10412 26424 10424
rect 26476 10412 26482 10464
rect 26602 10412 26608 10464
rect 26660 10452 26666 10464
rect 26881 10455 26939 10461
rect 26881 10452 26893 10455
rect 26660 10424 26893 10452
rect 26660 10412 26666 10424
rect 26881 10421 26893 10424
rect 26927 10421 26939 10455
rect 27614 10452 27620 10464
rect 27575 10424 27620 10452
rect 26881 10415 26939 10421
rect 27614 10412 27620 10424
rect 27672 10412 27678 10464
rect 29825 10455 29883 10461
rect 29825 10421 29837 10455
rect 29871 10452 29883 10455
rect 29914 10452 29920 10464
rect 29871 10424 29920 10452
rect 29871 10421 29883 10424
rect 29825 10415 29883 10421
rect 29914 10412 29920 10424
rect 29972 10412 29978 10464
rect 30282 10412 30288 10464
rect 30340 10452 30346 10464
rect 33781 10455 33839 10461
rect 30340 10424 30385 10452
rect 30340 10412 30346 10424
rect 33781 10421 33793 10455
rect 33827 10452 33839 10455
rect 34514 10452 34520 10464
rect 33827 10424 34520 10452
rect 33827 10421 33839 10424
rect 33781 10415 33839 10421
rect 34514 10412 34520 10424
rect 34572 10412 34578 10464
rect 36814 10452 36820 10464
rect 36775 10424 36820 10452
rect 36814 10412 36820 10424
rect 36872 10412 36878 10464
rect 1104 10362 38824 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 38824 10362
rect 1104 10288 38824 10310
rect 22097 10251 22155 10257
rect 22097 10217 22109 10251
rect 22143 10248 22155 10251
rect 23106 10248 23112 10260
rect 22143 10220 23112 10248
rect 22143 10217 22155 10220
rect 22097 10211 22155 10217
rect 23106 10208 23112 10220
rect 23164 10248 23170 10260
rect 24121 10251 24179 10257
rect 24121 10248 24133 10251
rect 23164 10220 24133 10248
rect 23164 10208 23170 10220
rect 24121 10217 24133 10220
rect 24167 10217 24179 10251
rect 24121 10211 24179 10217
rect 26418 10208 26424 10260
rect 26476 10248 26482 10260
rect 28353 10251 28411 10257
rect 28353 10248 28365 10251
rect 26476 10220 28365 10248
rect 26476 10208 26482 10220
rect 28353 10217 28365 10220
rect 28399 10217 28411 10251
rect 28353 10211 28411 10217
rect 30098 10208 30104 10260
rect 30156 10248 30162 10260
rect 30469 10251 30527 10257
rect 30469 10248 30481 10251
rect 30156 10220 30481 10248
rect 30156 10208 30162 10220
rect 30469 10217 30481 10220
rect 30515 10248 30527 10251
rect 30558 10248 30564 10260
rect 30515 10220 30564 10248
rect 30515 10217 30527 10220
rect 30469 10211 30527 10217
rect 30558 10208 30564 10220
rect 30616 10208 30622 10260
rect 32490 10248 32496 10260
rect 32451 10220 32496 10248
rect 32490 10208 32496 10220
rect 32548 10208 32554 10260
rect 32861 10251 32919 10257
rect 32861 10217 32873 10251
rect 32907 10217 32919 10251
rect 35434 10248 35440 10260
rect 35395 10220 35440 10248
rect 32861 10211 32919 10217
rect 32876 10180 32904 10211
rect 35434 10208 35440 10220
rect 35492 10208 35498 10260
rect 35526 10208 35532 10260
rect 35584 10248 35590 10260
rect 35897 10251 35955 10257
rect 35897 10248 35909 10251
rect 35584 10220 35909 10248
rect 35584 10208 35590 10220
rect 35897 10217 35909 10220
rect 35943 10217 35955 10251
rect 35897 10211 35955 10217
rect 33134 10180 33140 10192
rect 32876 10152 33140 10180
rect 33134 10140 33140 10152
rect 33192 10180 33198 10192
rect 33870 10180 33876 10192
rect 33192 10152 33876 10180
rect 33192 10140 33198 10152
rect 23014 10121 23020 10124
rect 23008 10112 23020 10121
rect 22975 10084 23020 10112
rect 23008 10075 23020 10084
rect 23014 10072 23020 10075
rect 23072 10072 23078 10124
rect 27240 10115 27298 10121
rect 27240 10081 27252 10115
rect 27286 10112 27298 10115
rect 27614 10112 27620 10124
rect 27286 10084 27620 10112
rect 27286 10081 27298 10084
rect 27240 10075 27298 10081
rect 27614 10072 27620 10084
rect 27672 10072 27678 10124
rect 29086 10072 29092 10124
rect 29144 10112 29150 10124
rect 29825 10115 29883 10121
rect 29825 10112 29837 10115
rect 29144 10084 29837 10112
rect 29144 10072 29150 10084
rect 29825 10081 29837 10084
rect 29871 10081 29883 10115
rect 33042 10112 33048 10124
rect 33003 10084 33048 10112
rect 29825 10075 29883 10081
rect 33042 10072 33048 10084
rect 33100 10072 33106 10124
rect 33428 10121 33456 10152
rect 33870 10140 33876 10152
rect 33928 10140 33934 10192
rect 33413 10115 33471 10121
rect 33413 10081 33425 10115
rect 33459 10081 33471 10115
rect 33413 10075 33471 10081
rect 33502 10072 33508 10124
rect 33560 10112 33566 10124
rect 33669 10115 33727 10121
rect 33669 10112 33681 10115
rect 33560 10084 33681 10112
rect 33560 10072 33566 10084
rect 33669 10081 33681 10084
rect 33715 10081 33727 10115
rect 36262 10112 36268 10124
rect 36223 10084 36268 10112
rect 33669 10075 33727 10081
rect 36262 10072 36268 10084
rect 36320 10072 36326 10124
rect 22741 10047 22799 10053
rect 22741 10044 22753 10047
rect 22480 10016 22753 10044
rect 22480 9920 22508 10016
rect 22741 10013 22753 10016
rect 22787 10013 22799 10047
rect 26973 10047 27031 10053
rect 26973 10044 26985 10047
rect 22741 10007 22799 10013
rect 26344 10016 26985 10044
rect 26344 9920 26372 10016
rect 26973 10013 26985 10016
rect 27019 10013 27031 10047
rect 29914 10044 29920 10056
rect 29875 10016 29920 10044
rect 26973 10007 27031 10013
rect 29914 10004 29920 10016
rect 29972 10004 29978 10056
rect 30098 10044 30104 10056
rect 30059 10016 30104 10044
rect 30098 10004 30104 10016
rect 30156 10004 30162 10056
rect 36354 10044 36360 10056
rect 36315 10016 36360 10044
rect 36354 10004 36360 10016
rect 36412 10004 36418 10056
rect 36541 10047 36599 10053
rect 36541 10013 36553 10047
rect 36587 10044 36599 10047
rect 36814 10044 36820 10056
rect 36587 10016 36820 10044
rect 36587 10013 36599 10016
rect 36541 10007 36599 10013
rect 36814 10004 36820 10016
rect 36872 10004 36878 10056
rect 28997 9979 29055 9985
rect 28997 9945 29009 9979
rect 29043 9976 29055 9979
rect 29822 9976 29828 9988
rect 29043 9948 29828 9976
rect 29043 9945 29055 9948
rect 28997 9939 29055 9945
rect 29822 9936 29828 9948
rect 29880 9936 29886 9988
rect 22462 9908 22468 9920
rect 22423 9880 22468 9908
rect 22462 9868 22468 9880
rect 22520 9868 22526 9920
rect 26326 9908 26332 9920
rect 26287 9880 26332 9908
rect 26326 9868 26332 9880
rect 26384 9868 26390 9920
rect 26602 9868 26608 9920
rect 26660 9908 26666 9920
rect 26697 9911 26755 9917
rect 26697 9908 26709 9911
rect 26660 9880 26709 9908
rect 26660 9868 26666 9880
rect 26697 9877 26709 9880
rect 26743 9877 26755 9911
rect 26697 9871 26755 9877
rect 29365 9911 29423 9917
rect 29365 9877 29377 9911
rect 29411 9908 29423 9911
rect 29454 9908 29460 9920
rect 29411 9880 29460 9908
rect 29411 9877 29423 9880
rect 29365 9871 29423 9877
rect 29454 9868 29460 9880
rect 29512 9868 29518 9920
rect 34790 9908 34796 9920
rect 34751 9880 34796 9908
rect 34790 9868 34796 9880
rect 34848 9868 34854 9920
rect 1104 9818 38824 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 34966 9818
rect 35018 9766 35030 9818
rect 35082 9766 35094 9818
rect 35146 9766 35158 9818
rect 35210 9766 38824 9818
rect 1104 9744 38824 9766
rect 22833 9707 22891 9713
rect 22833 9673 22845 9707
rect 22879 9704 22891 9707
rect 23014 9704 23020 9716
rect 22879 9676 23020 9704
rect 22879 9673 22891 9676
rect 22833 9667 22891 9673
rect 23014 9664 23020 9676
rect 23072 9704 23078 9716
rect 29086 9704 29092 9716
rect 23072 9676 24624 9704
rect 29047 9676 29092 9704
rect 23072 9664 23078 9676
rect 23474 9636 23480 9648
rect 23435 9608 23480 9636
rect 23474 9596 23480 9608
rect 23532 9596 23538 9648
rect 24596 9636 24624 9676
rect 29086 9664 29092 9676
rect 29144 9664 29150 9716
rect 30098 9704 30104 9716
rect 29196 9676 30104 9704
rect 25041 9639 25099 9645
rect 25041 9636 25053 9639
rect 24596 9608 25053 9636
rect 25041 9605 25053 9608
rect 25087 9605 25099 9639
rect 28718 9636 28724 9648
rect 28631 9608 28724 9636
rect 25041 9599 25099 9605
rect 28718 9596 28724 9608
rect 28776 9636 28782 9648
rect 29196 9636 29224 9676
rect 30098 9664 30104 9676
rect 30156 9704 30162 9716
rect 30282 9704 30288 9716
rect 30156 9676 30288 9704
rect 30156 9664 30162 9676
rect 30282 9664 30288 9676
rect 30340 9664 30346 9716
rect 33042 9664 33048 9716
rect 33100 9664 33106 9716
rect 35802 9664 35808 9716
rect 35860 9664 35866 9716
rect 28776 9608 29224 9636
rect 28776 9596 28782 9608
rect 31846 9596 31852 9648
rect 31904 9636 31910 9648
rect 33060 9636 33088 9664
rect 33873 9639 33931 9645
rect 33873 9636 33885 9639
rect 31904 9608 33885 9636
rect 31904 9596 31910 9608
rect 33873 9605 33885 9608
rect 33919 9605 33931 9639
rect 35820 9636 35848 9664
rect 36265 9639 36323 9645
rect 36265 9636 36277 9639
rect 35820 9608 36277 9636
rect 33873 9599 33931 9605
rect 36265 9605 36277 9608
rect 36311 9605 36323 9639
rect 36265 9599 36323 9605
rect 23492 9568 23520 9596
rect 23492 9540 23796 9568
rect 23661 9503 23719 9509
rect 23661 9469 23673 9503
rect 23707 9469 23719 9503
rect 23768 9500 23796 9540
rect 29454 9528 29460 9580
rect 29512 9568 29518 9580
rect 30288 9571 30346 9577
rect 30288 9568 30300 9571
rect 29512 9540 30300 9568
rect 29512 9528 29518 9540
rect 30288 9537 30300 9540
rect 30334 9537 30346 9571
rect 30558 9568 30564 9580
rect 30519 9540 30564 9568
rect 30288 9531 30346 9537
rect 30558 9528 30564 9540
rect 30616 9528 30622 9580
rect 32033 9571 32091 9577
rect 32033 9537 32045 9571
rect 32079 9568 32091 9571
rect 33045 9571 33103 9577
rect 33045 9568 33057 9571
rect 32079 9540 33057 9568
rect 32079 9537 32091 9540
rect 32033 9531 32091 9537
rect 33045 9537 33057 9540
rect 33091 9568 33103 9571
rect 33502 9568 33508 9580
rect 33091 9540 33508 9568
rect 33091 9537 33103 9540
rect 33045 9531 33103 9537
rect 33502 9528 33508 9540
rect 33560 9528 33566 9580
rect 23917 9503 23975 9509
rect 23917 9500 23929 9503
rect 23768 9472 23929 9500
rect 23661 9463 23719 9469
rect 23917 9469 23929 9472
rect 23963 9500 23975 9503
rect 24854 9500 24860 9512
rect 23963 9472 24860 9500
rect 23963 9469 23975 9472
rect 23917 9463 23975 9469
rect 22462 9432 22468 9444
rect 22375 9404 22468 9432
rect 22462 9392 22468 9404
rect 22520 9432 22526 9444
rect 23474 9432 23480 9444
rect 22520 9404 23480 9432
rect 22520 9392 22526 9404
rect 23474 9392 23480 9404
rect 23532 9432 23538 9444
rect 23676 9432 23704 9463
rect 24854 9460 24860 9472
rect 24912 9460 24918 9512
rect 25682 9500 25688 9512
rect 25595 9472 25688 9500
rect 25682 9460 25688 9472
rect 25740 9500 25746 9512
rect 26145 9503 26203 9509
rect 26145 9500 26157 9503
rect 25740 9472 26157 9500
rect 25740 9460 25746 9472
rect 26145 9469 26157 9472
rect 26191 9500 26203 9503
rect 26234 9500 26240 9512
rect 26191 9472 26240 9500
rect 26191 9469 26203 9472
rect 26145 9463 26203 9469
rect 26234 9460 26240 9472
rect 26292 9460 26298 9512
rect 29822 9500 29828 9512
rect 29783 9472 29828 9500
rect 29822 9460 29828 9472
rect 29880 9460 29886 9512
rect 32490 9460 32496 9512
rect 32548 9500 32554 9512
rect 32861 9503 32919 9509
rect 32861 9500 32873 9503
rect 32548 9472 32873 9500
rect 32548 9460 32554 9472
rect 32861 9469 32873 9472
rect 32907 9469 32919 9503
rect 34885 9503 34943 9509
rect 34885 9500 34897 9503
rect 32861 9463 32919 9469
rect 34256 9472 34897 9500
rect 24486 9432 24492 9444
rect 23532 9404 24492 9432
rect 23532 9392 23538 9404
rect 24486 9392 24492 9404
rect 24544 9392 24550 9444
rect 26050 9432 26056 9444
rect 25963 9404 26056 9432
rect 26050 9392 26056 9404
rect 26108 9432 26114 9444
rect 26390 9435 26448 9441
rect 26390 9432 26402 9435
rect 26108 9404 26402 9432
rect 26108 9392 26114 9404
rect 26390 9401 26402 9404
rect 26436 9401 26448 9435
rect 32401 9435 32459 9441
rect 32401 9432 32413 9435
rect 26390 9395 26448 9401
rect 32324 9404 32413 9432
rect 27522 9364 27528 9376
rect 27483 9336 27528 9364
rect 27522 9324 27528 9336
rect 27580 9324 27586 9376
rect 27614 9324 27620 9376
rect 27672 9364 27678 9376
rect 28169 9367 28227 9373
rect 28169 9364 28181 9367
rect 27672 9336 28181 9364
rect 27672 9324 27678 9336
rect 28169 9333 28181 9336
rect 28215 9364 28227 9367
rect 28902 9364 28908 9376
rect 28215 9336 28908 9364
rect 28215 9333 28227 9336
rect 28169 9327 28227 9333
rect 28902 9324 28908 9336
rect 28960 9324 28966 9376
rect 29638 9364 29644 9376
rect 29599 9336 29644 9364
rect 29638 9324 29644 9336
rect 29696 9364 29702 9376
rect 30291 9367 30349 9373
rect 30291 9364 30303 9367
rect 29696 9336 30303 9364
rect 29696 9324 29702 9336
rect 30291 9333 30303 9336
rect 30337 9333 30349 9367
rect 30291 9327 30349 9333
rect 31665 9367 31723 9373
rect 31665 9333 31677 9367
rect 31711 9364 31723 9367
rect 32324 9364 32352 9404
rect 32401 9401 32413 9404
rect 32447 9432 32459 9435
rect 32447 9404 32720 9432
rect 32447 9401 32459 9404
rect 32401 9395 32459 9401
rect 32490 9364 32496 9376
rect 31711 9336 32352 9364
rect 32451 9336 32496 9364
rect 31711 9333 31723 9336
rect 31665 9327 31723 9333
rect 32490 9324 32496 9336
rect 32548 9324 32554 9376
rect 32692 9364 32720 9404
rect 33134 9392 33140 9444
rect 33192 9432 33198 9444
rect 34256 9441 34284 9472
rect 34885 9469 34897 9472
rect 34931 9469 34943 9503
rect 34885 9463 34943 9469
rect 36262 9460 36268 9512
rect 36320 9500 36326 9512
rect 37369 9503 37427 9509
rect 37369 9500 37381 9503
rect 36320 9472 37381 9500
rect 36320 9460 36326 9472
rect 37369 9469 37381 9472
rect 37415 9469 37427 9503
rect 37369 9463 37427 9469
rect 34241 9435 34299 9441
rect 34241 9432 34253 9435
rect 33192 9404 34253 9432
rect 33192 9392 33198 9404
rect 34241 9401 34253 9404
rect 34287 9401 34299 9435
rect 34241 9395 34299 9401
rect 34701 9435 34759 9441
rect 34701 9401 34713 9435
rect 34747 9432 34759 9435
rect 34790 9432 34796 9444
rect 34747 9404 34796 9432
rect 34747 9401 34759 9404
rect 34701 9395 34759 9401
rect 34790 9392 34796 9404
rect 34848 9432 34854 9444
rect 35152 9435 35210 9441
rect 35152 9432 35164 9435
rect 34848 9404 35164 9432
rect 34848 9392 34854 9404
rect 35152 9401 35164 9404
rect 35198 9432 35210 9435
rect 35434 9432 35440 9444
rect 35198 9404 35440 9432
rect 35198 9401 35210 9404
rect 35152 9395 35210 9401
rect 35434 9392 35440 9404
rect 35492 9392 35498 9444
rect 32953 9367 33011 9373
rect 32953 9364 32965 9367
rect 32692 9336 32965 9364
rect 32953 9333 32965 9336
rect 32999 9364 33011 9367
rect 33318 9364 33324 9376
rect 32999 9336 33324 9364
rect 32999 9333 33011 9336
rect 32953 9327 33011 9333
rect 33318 9324 33324 9336
rect 33376 9324 33382 9376
rect 34882 9324 34888 9376
rect 34940 9364 34946 9376
rect 35986 9364 35992 9376
rect 34940 9336 35992 9364
rect 34940 9324 34946 9336
rect 35986 9324 35992 9336
rect 36044 9324 36050 9376
rect 36814 9364 36820 9376
rect 36775 9336 36820 9364
rect 36814 9324 36820 9336
rect 36872 9324 36878 9376
rect 1104 9274 38824 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 38824 9274
rect 1104 9200 38824 9222
rect 24854 9160 24860 9172
rect 24815 9132 24860 9160
rect 24854 9120 24860 9132
rect 24912 9120 24918 9172
rect 28997 9163 29055 9169
rect 28997 9129 29009 9163
rect 29043 9160 29055 9163
rect 29914 9160 29920 9172
rect 29043 9132 29920 9160
rect 29043 9129 29055 9132
rect 28997 9123 29055 9129
rect 29914 9120 29920 9132
rect 29972 9120 29978 9172
rect 30190 9120 30196 9172
rect 30248 9160 30254 9172
rect 30929 9163 30987 9169
rect 30929 9160 30941 9163
rect 30248 9132 30941 9160
rect 30248 9120 30254 9132
rect 30929 9129 30941 9132
rect 30975 9129 30987 9163
rect 30929 9123 30987 9129
rect 32950 9120 32956 9172
rect 33008 9160 33014 9172
rect 33051 9163 33109 9169
rect 33051 9160 33063 9163
rect 33008 9132 33063 9160
rect 33008 9120 33014 9132
rect 33051 9129 33063 9132
rect 33097 9129 33109 9163
rect 33051 9123 33109 9129
rect 34238 9120 34244 9172
rect 34296 9160 34302 9172
rect 34425 9163 34483 9169
rect 34425 9160 34437 9163
rect 34296 9132 34437 9160
rect 34296 9120 34302 9132
rect 34425 9129 34437 9132
rect 34471 9160 34483 9163
rect 35161 9163 35219 9169
rect 35161 9160 35173 9163
rect 34471 9132 35173 9160
rect 34471 9129 34483 9132
rect 34425 9123 34483 9129
rect 35161 9129 35173 9132
rect 35207 9129 35219 9163
rect 35161 9123 35219 9129
rect 35253 9163 35311 9169
rect 35253 9129 35265 9163
rect 35299 9129 35311 9163
rect 36262 9160 36268 9172
rect 36223 9132 36268 9160
rect 35253 9123 35311 9129
rect 29822 9101 29828 9104
rect 29816 9092 29828 9101
rect 29783 9064 29828 9092
rect 29816 9055 29828 9064
rect 29822 9052 29828 9055
rect 29880 9052 29886 9104
rect 35268 9092 35296 9123
rect 36262 9120 36268 9132
rect 36320 9120 36326 9172
rect 36354 9120 36360 9172
rect 36412 9160 36418 9172
rect 36633 9163 36691 9169
rect 36633 9160 36645 9163
rect 36412 9132 36645 9160
rect 36412 9120 36418 9132
rect 36633 9129 36645 9132
rect 36679 9129 36691 9163
rect 36633 9123 36691 9129
rect 36372 9092 36400 9120
rect 35268 9064 36400 9092
rect 23385 9027 23443 9033
rect 23385 8993 23397 9027
rect 23431 9024 23443 9027
rect 23474 9024 23480 9036
rect 23431 8996 23480 9024
rect 23431 8993 23443 8996
rect 23385 8987 23443 8993
rect 23474 8984 23480 8996
rect 23532 8984 23538 9036
rect 23750 9033 23756 9036
rect 23744 9024 23756 9033
rect 23711 8996 23756 9024
rect 23744 8987 23756 8996
rect 23750 8984 23756 8987
rect 23808 8984 23814 9036
rect 26142 9024 26148 9036
rect 26103 8996 26148 9024
rect 26142 8984 26148 8996
rect 26200 8984 26206 9036
rect 26418 8984 26424 9036
rect 26476 9024 26482 9036
rect 26769 9027 26827 9033
rect 26769 9024 26781 9027
rect 26476 8996 26781 9024
rect 26476 8984 26482 8996
rect 26769 8993 26781 8996
rect 26815 8993 26827 9027
rect 26769 8987 26827 8993
rect 27706 8984 27712 9036
rect 27764 9024 27770 9036
rect 29273 9027 29331 9033
rect 29273 9024 29285 9027
rect 27764 8996 29285 9024
rect 27764 8984 27770 8996
rect 29273 8993 29285 8996
rect 29319 8993 29331 9027
rect 35342 9024 35348 9036
rect 29273 8987 29331 8993
rect 33060 8996 35348 9024
rect 33060 8968 33088 8996
rect 35342 8984 35348 8996
rect 35400 9024 35406 9036
rect 35621 9027 35679 9033
rect 35621 9024 35633 9027
rect 35400 8996 35633 9024
rect 35400 8984 35406 8996
rect 35621 8993 35633 8996
rect 35667 8993 35679 9027
rect 35621 8987 35679 8993
rect 26234 8956 26240 8968
rect 25976 8928 26240 8956
rect 24486 8848 24492 8900
rect 24544 8888 24550 8900
rect 25976 8897 26004 8928
rect 26234 8916 26240 8928
rect 26292 8956 26298 8968
rect 26510 8956 26516 8968
rect 26292 8928 26516 8956
rect 26292 8916 26298 8928
rect 26510 8916 26516 8928
rect 26568 8916 26574 8968
rect 28629 8959 28687 8965
rect 28629 8925 28641 8959
rect 28675 8956 28687 8959
rect 29362 8956 29368 8968
rect 28675 8928 29368 8956
rect 28675 8925 28687 8928
rect 28629 8919 28687 8925
rect 29362 8916 29368 8928
rect 29420 8956 29426 8968
rect 29549 8959 29607 8965
rect 29549 8956 29561 8959
rect 29420 8928 29561 8956
rect 29420 8916 29426 8928
rect 29549 8925 29561 8928
rect 29595 8925 29607 8959
rect 29549 8919 29607 8925
rect 31938 8916 31944 8968
rect 31996 8956 32002 8968
rect 32585 8959 32643 8965
rect 32585 8956 32597 8959
rect 31996 8928 32597 8956
rect 31996 8916 32002 8928
rect 32585 8925 32597 8928
rect 32631 8925 32643 8959
rect 32585 8919 32643 8925
rect 33042 8916 33048 8968
rect 33100 8956 33106 8968
rect 33318 8956 33324 8968
rect 33100 8928 33193 8956
rect 33279 8928 33324 8956
rect 33100 8916 33106 8928
rect 33318 8916 33324 8928
rect 33376 8916 33382 8968
rect 35161 8959 35219 8965
rect 35161 8925 35173 8959
rect 35207 8956 35219 8959
rect 35713 8959 35771 8965
rect 35713 8956 35725 8959
rect 35207 8928 35725 8956
rect 35207 8925 35219 8928
rect 35161 8919 35219 8925
rect 35713 8925 35725 8928
rect 35759 8925 35771 8959
rect 35713 8919 35771 8925
rect 25961 8891 26019 8897
rect 25961 8888 25973 8891
rect 24544 8860 25973 8888
rect 24544 8848 24550 8860
rect 25961 8857 25973 8860
rect 26007 8857 26019 8891
rect 25961 8851 26019 8857
rect 34977 8891 35035 8897
rect 34977 8857 34989 8891
rect 35023 8888 35035 8891
rect 35434 8888 35440 8900
rect 35023 8860 35440 8888
rect 35023 8857 35035 8860
rect 34977 8851 35035 8857
rect 35434 8848 35440 8860
rect 35492 8848 35498 8900
rect 35728 8888 35756 8919
rect 35802 8916 35808 8968
rect 35860 8956 35866 8968
rect 35860 8928 35905 8956
rect 35860 8916 35866 8928
rect 35894 8888 35900 8900
rect 35728 8860 35900 8888
rect 35894 8848 35900 8860
rect 35952 8848 35958 8900
rect 27890 8820 27896 8832
rect 27851 8792 27896 8820
rect 27890 8780 27896 8792
rect 27948 8780 27954 8832
rect 29089 8823 29147 8829
rect 29089 8789 29101 8823
rect 29135 8820 29147 8823
rect 29178 8820 29184 8832
rect 29135 8792 29184 8820
rect 29135 8789 29147 8792
rect 29089 8783 29147 8789
rect 29178 8780 29184 8792
rect 29236 8820 29242 8832
rect 31849 8823 31907 8829
rect 31849 8820 31861 8823
rect 29236 8792 31861 8820
rect 29236 8780 29242 8792
rect 31849 8789 31861 8792
rect 31895 8820 31907 8823
rect 32030 8820 32036 8832
rect 31895 8792 32036 8820
rect 31895 8789 31907 8792
rect 31849 8783 31907 8789
rect 32030 8780 32036 8792
rect 32088 8780 32094 8832
rect 32401 8823 32459 8829
rect 32401 8789 32413 8823
rect 32447 8820 32459 8823
rect 32858 8820 32864 8832
rect 32447 8792 32864 8820
rect 32447 8789 32459 8792
rect 32401 8783 32459 8789
rect 32858 8780 32864 8792
rect 32916 8780 32922 8832
rect 1104 8730 38824 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 34966 8730
rect 35018 8678 35030 8730
rect 35082 8678 35094 8730
rect 35146 8678 35158 8730
rect 35210 8678 38824 8730
rect 1104 8656 38824 8678
rect 23477 8619 23535 8625
rect 23477 8585 23489 8619
rect 23523 8616 23535 8619
rect 23750 8616 23756 8628
rect 23523 8588 23756 8616
rect 23523 8585 23535 8588
rect 23477 8579 23535 8585
rect 23750 8576 23756 8588
rect 23808 8616 23814 8628
rect 25501 8619 25559 8625
rect 25501 8616 25513 8619
rect 23808 8588 25513 8616
rect 23808 8576 23814 8588
rect 25501 8585 25513 8588
rect 25547 8585 25559 8619
rect 26050 8616 26056 8628
rect 26011 8588 26056 8616
rect 25501 8579 25559 8585
rect 26050 8576 26056 8588
rect 26108 8576 26114 8628
rect 26418 8616 26424 8628
rect 26379 8588 26424 8616
rect 26418 8576 26424 8588
rect 26476 8576 26482 8628
rect 26602 8616 26608 8628
rect 26563 8588 26608 8616
rect 26602 8576 26608 8588
rect 26660 8576 26666 8628
rect 27706 8576 27712 8628
rect 27764 8616 27770 8628
rect 28261 8619 28319 8625
rect 28261 8616 28273 8619
rect 27764 8588 28273 8616
rect 27764 8576 27770 8588
rect 28261 8585 28273 8588
rect 28307 8585 28319 8619
rect 28261 8579 28319 8585
rect 29089 8619 29147 8625
rect 29089 8585 29101 8619
rect 29135 8616 29147 8619
rect 29730 8616 29736 8628
rect 29135 8588 29736 8616
rect 29135 8585 29147 8588
rect 29089 8579 29147 8585
rect 29730 8576 29736 8588
rect 29788 8576 29794 8628
rect 30374 8576 30380 8628
rect 30432 8616 30438 8628
rect 30745 8619 30803 8625
rect 30745 8616 30757 8619
rect 30432 8588 30757 8616
rect 30432 8576 30438 8588
rect 30745 8585 30757 8588
rect 30791 8585 30803 8619
rect 31846 8616 31852 8628
rect 31807 8588 31852 8616
rect 30745 8579 30803 8585
rect 31846 8576 31852 8588
rect 31904 8576 31910 8628
rect 32490 8576 32496 8628
rect 32548 8616 32554 8628
rect 34241 8619 34299 8625
rect 34241 8616 34253 8619
rect 32548 8588 34253 8616
rect 32548 8576 32554 8588
rect 34241 8585 34253 8588
rect 34287 8585 34299 8619
rect 34241 8579 34299 8585
rect 26068 8480 26096 8576
rect 27890 8548 27896 8560
rect 27080 8520 27896 8548
rect 27080 8489 27108 8520
rect 27890 8508 27896 8520
rect 27948 8508 27954 8560
rect 33502 8508 33508 8560
rect 33560 8548 33566 8560
rect 33689 8551 33747 8557
rect 33689 8548 33701 8551
rect 33560 8520 33701 8548
rect 33560 8508 33566 8520
rect 33689 8517 33701 8520
rect 33735 8517 33747 8551
rect 33689 8511 33747 8517
rect 27065 8483 27123 8489
rect 27065 8480 27077 8483
rect 26068 8452 27077 8480
rect 27065 8449 27077 8452
rect 27111 8449 27123 8483
rect 27065 8443 27123 8449
rect 27154 8440 27160 8492
rect 27212 8480 27218 8492
rect 29362 8480 29368 8492
rect 27212 8452 27257 8480
rect 29323 8452 29368 8480
rect 27212 8440 27218 8452
rect 29362 8440 29368 8452
rect 29420 8480 29426 8492
rect 32309 8483 32367 8489
rect 32309 8480 32321 8483
rect 29420 8452 29500 8480
rect 29420 8440 29426 8452
rect 23109 8415 23167 8421
rect 23109 8381 23121 8415
rect 23155 8412 23167 8415
rect 24118 8412 24124 8424
rect 23155 8384 24124 8412
rect 23155 8381 23167 8384
rect 23109 8375 23167 8381
rect 24118 8372 24124 8384
rect 24176 8372 24182 8424
rect 24388 8415 24446 8421
rect 24388 8412 24400 8415
rect 24320 8384 24400 8412
rect 24029 8347 24087 8353
rect 24029 8313 24041 8347
rect 24075 8344 24087 8347
rect 24320 8344 24348 8384
rect 24388 8381 24400 8384
rect 24434 8412 24446 8415
rect 26878 8412 26884 8424
rect 24434 8384 26884 8412
rect 24434 8381 24446 8384
rect 24388 8375 24446 8381
rect 26878 8372 26884 8384
rect 26936 8412 26942 8424
rect 26973 8415 27031 8421
rect 26973 8412 26985 8415
rect 26936 8384 26985 8412
rect 26936 8372 26942 8384
rect 26973 8381 26985 8384
rect 27019 8412 27031 8415
rect 27522 8412 27528 8424
rect 27019 8384 27528 8412
rect 27019 8381 27031 8384
rect 26973 8375 27031 8381
rect 27522 8372 27528 8384
rect 27580 8372 27586 8424
rect 29472 8412 29500 8452
rect 31404 8452 32321 8480
rect 29472 8384 30328 8412
rect 24075 8316 24348 8344
rect 28721 8347 28779 8353
rect 24075 8313 24087 8316
rect 24029 8307 24087 8313
rect 28721 8313 28733 8347
rect 28767 8344 28779 8347
rect 29632 8347 29690 8353
rect 29632 8344 29644 8347
rect 28767 8316 29644 8344
rect 28767 8313 28779 8316
rect 28721 8307 28779 8313
rect 29632 8313 29644 8316
rect 29678 8344 29690 8347
rect 30190 8344 30196 8356
rect 29678 8316 30196 8344
rect 29678 8313 29690 8316
rect 29632 8307 29690 8313
rect 30190 8304 30196 8316
rect 30248 8304 30254 8356
rect 30300 8344 30328 8384
rect 30374 8344 30380 8356
rect 30300 8316 30380 8344
rect 30374 8304 30380 8316
rect 30432 8344 30438 8356
rect 31297 8347 31355 8353
rect 31297 8344 31309 8347
rect 30432 8316 31309 8344
rect 30432 8304 30438 8316
rect 31297 8313 31309 8316
rect 31343 8344 31355 8347
rect 31404 8344 31432 8452
rect 32309 8449 32321 8452
rect 32355 8449 32367 8483
rect 32309 8443 32367 8449
rect 32030 8412 32036 8424
rect 31991 8384 32036 8412
rect 32030 8372 32036 8384
rect 32088 8372 32094 8424
rect 32324 8412 32352 8443
rect 33134 8412 33140 8424
rect 32324 8384 33140 8412
rect 33134 8372 33140 8384
rect 33192 8372 33198 8424
rect 31343 8316 31432 8344
rect 32576 8347 32634 8353
rect 31343 8313 31355 8316
rect 31297 8307 31355 8313
rect 32576 8313 32588 8347
rect 32622 8344 32634 8347
rect 32858 8344 32864 8356
rect 32622 8316 32864 8344
rect 32622 8313 32634 8316
rect 32576 8307 32634 8313
rect 32858 8304 32864 8316
rect 32916 8304 32922 8356
rect 34256 8344 34284 8579
rect 34514 8576 34520 8628
rect 34572 8616 34578 8628
rect 34609 8619 34667 8625
rect 34609 8616 34621 8619
rect 34572 8588 34621 8616
rect 34572 8576 34578 8588
rect 34609 8585 34621 8588
rect 34655 8616 34667 8619
rect 34655 8588 35296 8616
rect 34655 8585 34667 8588
rect 34609 8579 34667 8585
rect 34698 8508 34704 8560
rect 34756 8548 34762 8560
rect 34885 8551 34943 8557
rect 34885 8548 34897 8551
rect 34756 8520 34897 8548
rect 34756 8508 34762 8520
rect 34885 8517 34897 8520
rect 34931 8548 34943 8551
rect 35158 8548 35164 8560
rect 34931 8520 35164 8548
rect 34931 8517 34943 8520
rect 34885 8511 34943 8517
rect 35158 8508 35164 8520
rect 35216 8508 35222 8560
rect 35268 8421 35296 8588
rect 35802 8576 35808 8628
rect 35860 8616 35866 8628
rect 36265 8619 36323 8625
rect 36265 8616 36277 8619
rect 35860 8588 36277 8616
rect 35860 8576 35866 8588
rect 36265 8585 36277 8588
rect 36311 8585 36323 8619
rect 37090 8616 37096 8628
rect 37051 8588 37096 8616
rect 36265 8579 36323 8585
rect 37090 8576 37096 8588
rect 37148 8576 37154 8628
rect 35894 8548 35900 8560
rect 35855 8520 35900 8548
rect 35894 8508 35900 8520
rect 35952 8508 35958 8560
rect 35434 8480 35440 8492
rect 35395 8452 35440 8480
rect 35434 8440 35440 8452
rect 35492 8440 35498 8492
rect 35253 8415 35311 8421
rect 35253 8381 35265 8415
rect 35299 8381 35311 8415
rect 35253 8375 35311 8381
rect 36449 8415 36507 8421
rect 36449 8381 36461 8415
rect 36495 8412 36507 8415
rect 37090 8412 37096 8424
rect 36495 8384 37096 8412
rect 36495 8381 36507 8384
rect 36449 8375 36507 8381
rect 37090 8372 37096 8384
rect 37148 8372 37154 8424
rect 35345 8347 35403 8353
rect 35345 8344 35357 8347
rect 34256 8316 35357 8344
rect 35345 8313 35357 8316
rect 35391 8313 35403 8347
rect 35345 8307 35403 8313
rect 35802 8304 35808 8356
rect 35860 8344 35866 8356
rect 36078 8344 36084 8356
rect 35860 8316 36084 8344
rect 35860 8304 35866 8316
rect 36078 8304 36084 8316
rect 36136 8304 36142 8356
rect 27709 8279 27767 8285
rect 27709 8245 27721 8279
rect 27755 8276 27767 8279
rect 28350 8276 28356 8288
rect 27755 8248 28356 8276
rect 27755 8245 27767 8248
rect 27709 8239 27767 8245
rect 28350 8236 28356 8248
rect 28408 8236 28414 8288
rect 31754 8236 31760 8288
rect 31812 8276 31818 8288
rect 36630 8276 36636 8288
rect 31812 8248 31857 8276
rect 36591 8248 36636 8276
rect 31812 8236 31818 8248
rect 36630 8236 36636 8248
rect 36688 8236 36694 8288
rect 1104 8186 38824 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 38824 8186
rect 1104 8112 38824 8134
rect 24118 8032 24124 8084
rect 24176 8072 24182 8084
rect 24213 8075 24271 8081
rect 24213 8072 24225 8075
rect 24176 8044 24225 8072
rect 24176 8032 24182 8044
rect 24213 8041 24225 8044
rect 24259 8072 24271 8075
rect 24486 8072 24492 8084
rect 24259 8044 24492 8072
rect 24259 8041 24271 8044
rect 24213 8035 24271 8041
rect 24486 8032 24492 8044
rect 24544 8032 24550 8084
rect 26053 8075 26111 8081
rect 26053 8041 26065 8075
rect 26099 8072 26111 8075
rect 26142 8072 26148 8084
rect 26099 8044 26148 8072
rect 26099 8041 26111 8044
rect 26053 8035 26111 8041
rect 26142 8032 26148 8044
rect 26200 8032 26206 8084
rect 26789 8075 26847 8081
rect 26789 8041 26801 8075
rect 26835 8072 26847 8075
rect 26878 8072 26884 8084
rect 26835 8044 26884 8072
rect 26835 8041 26847 8044
rect 26789 8035 26847 8041
rect 26878 8032 26884 8044
rect 26936 8032 26942 8084
rect 27154 8072 27160 8084
rect 27115 8044 27160 8072
rect 27154 8032 27160 8044
rect 27212 8032 27218 8084
rect 28994 8032 29000 8084
rect 29052 8072 29058 8084
rect 29733 8075 29791 8081
rect 29733 8072 29745 8075
rect 29052 8044 29745 8072
rect 29052 8032 29058 8044
rect 29733 8041 29745 8044
rect 29779 8041 29791 8075
rect 30374 8072 30380 8084
rect 30335 8044 30380 8072
rect 29733 8035 29791 8041
rect 30374 8032 30380 8044
rect 30432 8032 30438 8084
rect 31754 8032 31760 8084
rect 31812 8072 31818 8084
rect 32309 8075 32367 8081
rect 32309 8072 32321 8075
rect 31812 8044 32321 8072
rect 31812 8032 31818 8044
rect 32309 8041 32321 8044
rect 32355 8072 32367 8075
rect 33042 8072 33048 8084
rect 32355 8044 33048 8072
rect 32355 8041 32367 8044
rect 32309 8035 32367 8041
rect 33042 8032 33048 8044
rect 33100 8032 33106 8084
rect 33137 8075 33195 8081
rect 33137 8041 33149 8075
rect 33183 8072 33195 8075
rect 33318 8072 33324 8084
rect 33183 8044 33324 8072
rect 33183 8041 33195 8044
rect 33137 8035 33195 8041
rect 33318 8032 33324 8044
rect 33376 8032 33382 8084
rect 35342 8072 35348 8084
rect 35303 8044 35348 8072
rect 35342 8032 35348 8044
rect 35400 8032 35406 8084
rect 28620 8007 28678 8013
rect 28620 7973 28632 8007
rect 28666 8004 28678 8007
rect 28718 8004 28724 8016
rect 28666 7976 28724 8004
rect 28666 7973 28678 7976
rect 28620 7967 28678 7973
rect 28718 7964 28724 7976
rect 28776 7964 28782 8016
rect 31938 8004 31944 8016
rect 31899 7976 31944 8004
rect 31938 7964 31944 7976
rect 31996 7964 32002 8016
rect 32769 8007 32827 8013
rect 32769 7973 32781 8007
rect 32815 8004 32827 8007
rect 32950 8004 32956 8016
rect 32815 7976 32956 8004
rect 32815 7973 32827 7976
rect 32769 7967 32827 7973
rect 32950 7964 32956 7976
rect 33008 7964 33014 8016
rect 35618 7964 35624 8016
rect 35676 8004 35682 8016
rect 35713 8007 35771 8013
rect 35713 8004 35725 8007
rect 35676 7976 35725 8004
rect 35676 7964 35682 7976
rect 35713 7973 35725 7976
rect 35759 7973 35771 8007
rect 35713 7967 35771 7973
rect 32122 7936 32128 7948
rect 32083 7908 32128 7936
rect 32122 7896 32128 7908
rect 32180 7896 32186 7948
rect 33134 7896 33140 7948
rect 33192 7936 33198 7948
rect 33229 7939 33287 7945
rect 33229 7936 33241 7939
rect 33192 7908 33241 7936
rect 33192 7896 33198 7908
rect 33229 7905 33241 7908
rect 33275 7905 33287 7939
rect 33229 7899 33287 7905
rect 33318 7896 33324 7948
rect 33376 7936 33382 7948
rect 33485 7939 33543 7945
rect 33485 7936 33497 7939
rect 33376 7908 33497 7936
rect 33376 7896 33382 7908
rect 33485 7905 33497 7908
rect 33531 7905 33543 7939
rect 33485 7899 33543 7905
rect 35897 7939 35955 7945
rect 35897 7905 35909 7939
rect 35943 7936 35955 7939
rect 36170 7936 36176 7948
rect 35943 7908 36176 7936
rect 35943 7905 35955 7908
rect 35897 7899 35955 7905
rect 36170 7896 36176 7908
rect 36228 7896 36234 7948
rect 28350 7868 28356 7880
rect 28311 7840 28356 7868
rect 28350 7828 28356 7840
rect 28408 7828 28414 7880
rect 31021 7871 31079 7877
rect 31021 7837 31033 7871
rect 31067 7868 31079 7871
rect 32030 7868 32036 7880
rect 31067 7840 32036 7868
rect 31067 7837 31079 7840
rect 31021 7831 31079 7837
rect 32030 7828 32036 7840
rect 32088 7828 32094 7880
rect 35526 7760 35532 7812
rect 35584 7800 35590 7812
rect 36354 7800 36360 7812
rect 35584 7772 36360 7800
rect 35584 7760 35590 7772
rect 36354 7760 36360 7772
rect 36412 7760 36418 7812
rect 34606 7732 34612 7744
rect 34567 7704 34612 7732
rect 34606 7692 34612 7704
rect 34664 7692 34670 7744
rect 34790 7692 34796 7744
rect 34848 7732 34854 7744
rect 35710 7732 35716 7744
rect 34848 7704 35716 7732
rect 34848 7692 34854 7704
rect 35710 7692 35716 7704
rect 35768 7692 35774 7744
rect 36078 7732 36084 7744
rect 36039 7704 36084 7732
rect 36078 7692 36084 7704
rect 36136 7692 36142 7744
rect 1104 7642 38824 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 34966 7642
rect 35018 7590 35030 7642
rect 35082 7590 35094 7642
rect 35146 7590 35158 7642
rect 35210 7590 38824 7642
rect 1104 7568 38824 7590
rect 28445 7531 28503 7537
rect 28445 7497 28457 7531
rect 28491 7528 28503 7531
rect 28718 7528 28724 7540
rect 28491 7500 28724 7528
rect 28491 7497 28503 7500
rect 28445 7491 28503 7497
rect 28718 7488 28724 7500
rect 28776 7488 28782 7540
rect 32030 7528 32036 7540
rect 31991 7500 32036 7528
rect 32030 7488 32036 7500
rect 32088 7488 32094 7540
rect 32217 7531 32275 7537
rect 32217 7497 32229 7531
rect 32263 7528 32275 7531
rect 32398 7528 32404 7540
rect 32263 7500 32404 7528
rect 32263 7497 32275 7500
rect 32217 7491 32275 7497
rect 32398 7488 32404 7500
rect 32456 7488 32462 7540
rect 33134 7488 33140 7540
rect 33192 7528 33198 7540
rect 33965 7531 34023 7537
rect 33965 7528 33977 7531
rect 33192 7500 33977 7528
rect 33192 7488 33198 7500
rect 33965 7497 33977 7500
rect 34011 7497 34023 7531
rect 33965 7491 34023 7497
rect 35345 7531 35403 7537
rect 35345 7497 35357 7531
rect 35391 7528 35403 7531
rect 35618 7528 35624 7540
rect 35391 7500 35624 7528
rect 35391 7497 35403 7500
rect 35345 7491 35403 7497
rect 35618 7488 35624 7500
rect 35676 7488 35682 7540
rect 29086 7352 29092 7404
rect 29144 7392 29150 7404
rect 29457 7395 29515 7401
rect 29457 7392 29469 7395
rect 29144 7364 29469 7392
rect 29144 7352 29150 7364
rect 29457 7361 29469 7364
rect 29503 7361 29515 7395
rect 29457 7355 29515 7361
rect 31757 7395 31815 7401
rect 31757 7361 31769 7395
rect 31803 7392 31815 7395
rect 32858 7392 32864 7404
rect 31803 7364 32864 7392
rect 31803 7361 31815 7364
rect 31757 7355 31815 7361
rect 32858 7352 32864 7364
rect 32916 7352 32922 7404
rect 31113 7327 31171 7333
rect 31113 7293 31125 7327
rect 31159 7324 31171 7327
rect 31159 7296 31193 7324
rect 31159 7293 31171 7296
rect 31113 7287 31171 7293
rect 31021 7259 31079 7265
rect 31021 7225 31033 7259
rect 31067 7256 31079 7259
rect 31128 7256 31156 7287
rect 32030 7284 32036 7336
rect 32088 7324 32094 7336
rect 32585 7327 32643 7333
rect 32585 7324 32597 7327
rect 32088 7296 32597 7324
rect 32088 7284 32094 7296
rect 32585 7293 32597 7296
rect 32631 7293 32643 7327
rect 33318 7324 33324 7336
rect 33231 7296 33324 7324
rect 32585 7287 32643 7293
rect 33318 7284 33324 7296
rect 33376 7324 33382 7336
rect 35434 7324 35440 7336
rect 33376 7296 34100 7324
rect 35395 7296 35440 7324
rect 33376 7284 33382 7296
rect 31202 7256 31208 7268
rect 31067 7228 31208 7256
rect 31067 7225 31079 7228
rect 31021 7219 31079 7225
rect 31202 7216 31208 7228
rect 31260 7216 31266 7268
rect 32674 7256 32680 7268
rect 32587 7228 32680 7256
rect 32674 7216 32680 7228
rect 32732 7256 32738 7268
rect 33597 7259 33655 7265
rect 33597 7256 33609 7259
rect 32732 7228 33609 7256
rect 32732 7216 32738 7228
rect 33597 7225 33609 7228
rect 33643 7225 33655 7259
rect 33597 7219 33655 7225
rect 27614 7148 27620 7200
rect 27672 7188 27678 7200
rect 28350 7188 28356 7200
rect 27672 7160 28356 7188
rect 27672 7148 27678 7160
rect 28350 7148 28356 7160
rect 28408 7188 28414 7200
rect 28721 7191 28779 7197
rect 28721 7188 28733 7191
rect 28408 7160 28733 7188
rect 28408 7148 28414 7160
rect 28721 7157 28733 7160
rect 28767 7157 28779 7191
rect 31294 7188 31300 7200
rect 31255 7160 31300 7188
rect 28721 7151 28779 7157
rect 31294 7148 31300 7160
rect 31352 7148 31358 7200
rect 34072 7188 34100 7296
rect 35434 7284 35440 7296
rect 35492 7284 35498 7336
rect 34701 7259 34759 7265
rect 34701 7225 34713 7259
rect 34747 7256 34759 7259
rect 35704 7259 35762 7265
rect 35704 7256 35716 7259
rect 34747 7228 35716 7256
rect 34747 7225 34759 7228
rect 34701 7219 34759 7225
rect 35704 7225 35716 7228
rect 35750 7256 35762 7259
rect 36170 7256 36176 7268
rect 35750 7228 36176 7256
rect 35750 7225 35762 7228
rect 35704 7219 35762 7225
rect 36170 7216 36176 7228
rect 36228 7216 36234 7268
rect 36817 7191 36875 7197
rect 36817 7188 36829 7191
rect 34072 7160 36829 7188
rect 36817 7157 36829 7160
rect 36863 7157 36875 7191
rect 36817 7151 36875 7157
rect 1104 7098 38824 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 38824 7098
rect 1104 7024 38824 7046
rect 32122 6944 32128 6996
rect 32180 6984 32186 6996
rect 32309 6987 32367 6993
rect 32309 6984 32321 6987
rect 32180 6956 32321 6984
rect 32180 6944 32186 6956
rect 32309 6953 32321 6956
rect 32355 6953 32367 6987
rect 32674 6984 32680 6996
rect 32635 6956 32680 6984
rect 32309 6947 32367 6953
rect 32674 6944 32680 6956
rect 32732 6944 32738 6996
rect 34790 6944 34796 6996
rect 34848 6984 34854 6996
rect 35434 6984 35440 6996
rect 34848 6956 35440 6984
rect 34848 6944 34854 6956
rect 35434 6944 35440 6956
rect 35492 6984 35498 6996
rect 36265 6987 36323 6993
rect 36265 6984 36277 6987
rect 35492 6956 36277 6984
rect 35492 6944 35498 6956
rect 36265 6953 36277 6956
rect 36311 6953 36323 6987
rect 36265 6947 36323 6953
rect 31294 6876 31300 6928
rect 31352 6916 31358 6928
rect 32766 6916 32772 6928
rect 31352 6888 32772 6916
rect 31352 6876 31358 6888
rect 32766 6876 32772 6888
rect 32824 6916 32830 6928
rect 33045 6919 33103 6925
rect 33045 6916 33057 6919
rect 32824 6888 33057 6916
rect 32824 6876 32830 6888
rect 33045 6885 33057 6888
rect 33091 6885 33103 6919
rect 33045 6879 33103 6885
rect 33318 6876 33324 6928
rect 33376 6876 33382 6928
rect 26786 6857 26792 6860
rect 26780 6848 26792 6857
rect 26747 6820 26792 6848
rect 26780 6811 26792 6820
rect 26786 6808 26792 6811
rect 26844 6808 26850 6860
rect 30282 6848 30288 6860
rect 30243 6820 30288 6848
rect 30282 6808 30288 6820
rect 30340 6808 30346 6860
rect 31757 6851 31815 6857
rect 31757 6817 31769 6851
rect 31803 6848 31815 6851
rect 31846 6848 31852 6860
rect 31803 6820 31852 6848
rect 31803 6817 31815 6820
rect 31757 6811 31815 6817
rect 31846 6808 31852 6820
rect 31904 6808 31910 6860
rect 31938 6808 31944 6860
rect 31996 6848 32002 6860
rect 33336 6848 33364 6876
rect 34238 6848 34244 6860
rect 31996 6820 33364 6848
rect 34199 6820 34244 6848
rect 31996 6808 32002 6820
rect 26510 6780 26516 6792
rect 26471 6752 26516 6780
rect 26510 6740 26516 6752
rect 26568 6740 26574 6792
rect 33336 6789 33364 6820
rect 34238 6808 34244 6820
rect 34296 6808 34302 6860
rect 35345 6851 35403 6857
rect 35345 6817 35357 6851
rect 35391 6848 35403 6851
rect 35434 6848 35440 6860
rect 35391 6820 35440 6848
rect 35391 6817 35403 6820
rect 35345 6811 35403 6817
rect 35434 6808 35440 6820
rect 35492 6808 35498 6860
rect 36449 6851 36507 6857
rect 36449 6817 36461 6851
rect 36495 6848 36507 6851
rect 36998 6848 37004 6860
rect 36495 6820 37004 6848
rect 36495 6817 36507 6820
rect 36449 6811 36507 6817
rect 36998 6808 37004 6820
rect 37056 6808 37062 6860
rect 33137 6783 33195 6789
rect 33137 6749 33149 6783
rect 33183 6749 33195 6783
rect 33137 6743 33195 6749
rect 33321 6783 33379 6789
rect 33321 6749 33333 6783
rect 33367 6749 33379 6783
rect 33321 6743 33379 6749
rect 32398 6672 32404 6724
rect 32456 6712 32462 6724
rect 33152 6712 33180 6743
rect 34425 6715 34483 6721
rect 34425 6712 34437 6715
rect 32456 6684 34437 6712
rect 32456 6672 32462 6684
rect 34425 6681 34437 6684
rect 34471 6681 34483 6715
rect 34425 6675 34483 6681
rect 26510 6604 26516 6656
rect 26568 6644 26574 6656
rect 27522 6644 27528 6656
rect 26568 6616 27528 6644
rect 26568 6604 26574 6616
rect 27522 6604 27528 6616
rect 27580 6604 27586 6656
rect 27890 6644 27896 6656
rect 27851 6616 27896 6644
rect 27890 6604 27896 6616
rect 27948 6604 27954 6656
rect 29365 6647 29423 6653
rect 29365 6613 29377 6647
rect 29411 6644 29423 6647
rect 29822 6644 29828 6656
rect 29411 6616 29828 6644
rect 29411 6613 29423 6616
rect 29365 6607 29423 6613
rect 29822 6604 29828 6616
rect 29880 6604 29886 6656
rect 30469 6647 30527 6653
rect 30469 6613 30481 6647
rect 30515 6644 30527 6647
rect 30834 6644 30840 6656
rect 30515 6616 30840 6644
rect 30515 6613 30527 6616
rect 30469 6607 30527 6613
rect 30834 6604 30840 6616
rect 30892 6604 30898 6656
rect 31386 6644 31392 6656
rect 31347 6616 31392 6644
rect 31386 6604 31392 6616
rect 31444 6604 31450 6656
rect 33778 6644 33784 6656
rect 33739 6616 33784 6644
rect 33778 6604 33784 6616
rect 33836 6604 33842 6656
rect 35526 6644 35532 6656
rect 35487 6616 35532 6644
rect 35526 6604 35532 6616
rect 35584 6604 35590 6656
rect 35989 6647 36047 6653
rect 35989 6613 36001 6647
rect 36035 6644 36047 6647
rect 36170 6644 36176 6656
rect 36035 6616 36176 6644
rect 36035 6613 36047 6616
rect 35989 6607 36047 6613
rect 36170 6604 36176 6616
rect 36228 6604 36234 6656
rect 36446 6604 36452 6656
rect 36504 6644 36510 6656
rect 36633 6647 36691 6653
rect 36633 6644 36645 6647
rect 36504 6616 36645 6644
rect 36504 6604 36510 6616
rect 36633 6613 36645 6616
rect 36679 6613 36691 6647
rect 36633 6607 36691 6613
rect 1104 6554 38824 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 34966 6554
rect 35018 6502 35030 6554
rect 35082 6502 35094 6554
rect 35146 6502 35158 6554
rect 35210 6502 38824 6554
rect 1104 6480 38824 6502
rect 26605 6443 26663 6449
rect 26605 6409 26617 6443
rect 26651 6440 26663 6443
rect 26786 6440 26792 6452
rect 26651 6412 26792 6440
rect 26651 6409 26663 6412
rect 26605 6403 26663 6409
rect 26786 6400 26792 6412
rect 26844 6400 26850 6452
rect 30834 6440 30840 6452
rect 30795 6412 30840 6440
rect 30834 6400 30840 6412
rect 30892 6400 30898 6452
rect 32398 6440 32404 6452
rect 32359 6412 32404 6440
rect 32398 6400 32404 6412
rect 32456 6400 32462 6452
rect 32766 6440 32772 6452
rect 32727 6412 32772 6440
rect 32766 6400 32772 6412
rect 32824 6400 32830 6452
rect 36538 6440 36544 6452
rect 36499 6412 36544 6440
rect 36538 6400 36544 6412
rect 36596 6400 36602 6452
rect 36998 6440 37004 6452
rect 36959 6412 37004 6440
rect 36998 6400 37004 6412
rect 37056 6400 37062 6452
rect 27617 6375 27675 6381
rect 27617 6341 27629 6375
rect 27663 6372 27675 6375
rect 28997 6375 29055 6381
rect 28997 6372 29009 6375
rect 27663 6344 29009 6372
rect 27663 6341 27675 6344
rect 27617 6335 27675 6341
rect 28997 6341 29009 6344
rect 29043 6341 29055 6375
rect 28997 6335 29055 6341
rect 29273 6375 29331 6381
rect 29273 6341 29285 6375
rect 29319 6372 29331 6375
rect 30282 6372 30288 6384
rect 29319 6344 30288 6372
rect 29319 6341 29331 6344
rect 29273 6335 29331 6341
rect 27525 6307 27583 6313
rect 27525 6273 27537 6307
rect 27571 6304 27583 6307
rect 27890 6304 27896 6316
rect 27571 6276 27896 6304
rect 27571 6273 27583 6276
rect 27525 6267 27583 6273
rect 27890 6264 27896 6276
rect 27948 6304 27954 6316
rect 28077 6307 28135 6313
rect 28077 6304 28089 6307
rect 27948 6276 28089 6304
rect 27948 6264 27954 6276
rect 28077 6273 28089 6276
rect 28123 6273 28135 6307
rect 28077 6267 28135 6273
rect 28261 6307 28319 6313
rect 28261 6273 28273 6307
rect 28307 6304 28319 6307
rect 28718 6304 28724 6316
rect 28307 6276 28724 6304
rect 28307 6273 28319 6276
rect 28261 6267 28319 6273
rect 28718 6264 28724 6276
rect 28776 6264 28782 6316
rect 29012 6304 29040 6335
rect 30282 6332 30288 6344
rect 30340 6332 30346 6384
rect 29733 6307 29791 6313
rect 29733 6304 29745 6307
rect 29012 6276 29745 6304
rect 29733 6273 29745 6276
rect 29779 6273 29791 6307
rect 29733 6267 29791 6273
rect 29822 6264 29828 6316
rect 29880 6304 29886 6316
rect 29880 6276 29925 6304
rect 29880 6264 29886 6276
rect 30852 6168 30880 6400
rect 32861 6375 32919 6381
rect 32861 6341 32873 6375
rect 32907 6372 32919 6375
rect 34238 6372 34244 6384
rect 32907 6344 34244 6372
rect 32907 6341 32919 6344
rect 32861 6335 32919 6341
rect 34238 6332 34244 6344
rect 34296 6332 34302 6384
rect 31386 6264 31392 6316
rect 31444 6304 31450 6316
rect 31941 6307 31999 6313
rect 31941 6304 31953 6307
rect 31444 6276 31953 6304
rect 31444 6264 31450 6276
rect 31941 6273 31953 6276
rect 31987 6304 31999 6307
rect 33410 6304 33416 6316
rect 31987 6276 33416 6304
rect 31987 6273 31999 6276
rect 31941 6267 31999 6273
rect 33410 6264 33416 6276
rect 33468 6264 33474 6316
rect 33505 6307 33563 6313
rect 33505 6273 33517 6307
rect 33551 6304 33563 6307
rect 33778 6304 33784 6316
rect 33551 6276 33784 6304
rect 33551 6273 33563 6276
rect 33505 6267 33563 6273
rect 33778 6264 33784 6276
rect 33836 6264 33842 6316
rect 36556 6304 36584 6400
rect 37274 6372 37280 6384
rect 37235 6344 37280 6372
rect 37274 6332 37280 6344
rect 37332 6332 37338 6384
rect 36004 6276 36584 6304
rect 31205 6239 31263 6245
rect 31205 6205 31217 6239
rect 31251 6236 31263 6239
rect 31251 6208 31892 6236
rect 31251 6205 31263 6208
rect 31205 6199 31263 6205
rect 31864 6180 31892 6208
rect 32122 6196 32128 6248
rect 32180 6236 32186 6248
rect 33134 6236 33140 6248
rect 32180 6208 33140 6236
rect 32180 6196 32186 6208
rect 33134 6196 33140 6208
rect 33192 6236 33198 6248
rect 36004 6245 36032 6276
rect 33229 6239 33287 6245
rect 33229 6236 33241 6239
rect 33192 6208 33241 6236
rect 33192 6196 33198 6208
rect 33229 6205 33241 6208
rect 33275 6236 33287 6239
rect 33873 6239 33931 6245
rect 33873 6236 33885 6239
rect 33275 6208 33885 6236
rect 33275 6205 33287 6208
rect 33229 6199 33287 6205
rect 33873 6205 33885 6208
rect 33919 6205 33931 6239
rect 34885 6239 34943 6245
rect 34885 6236 34897 6239
rect 33873 6199 33931 6205
rect 34624 6208 34897 6236
rect 31757 6171 31815 6177
rect 31757 6168 31769 6171
rect 30852 6140 31769 6168
rect 31757 6137 31769 6140
rect 31803 6137 31815 6171
rect 31757 6131 31815 6137
rect 31846 6128 31852 6180
rect 31904 6128 31910 6180
rect 34624 6112 34652 6208
rect 34885 6205 34897 6208
rect 34931 6205 34943 6239
rect 34885 6199 34943 6205
rect 35989 6239 36047 6245
rect 35989 6205 36001 6239
rect 36035 6205 36047 6239
rect 35989 6199 36047 6205
rect 36078 6196 36084 6248
rect 36136 6236 36142 6248
rect 37093 6239 37151 6245
rect 37093 6236 37105 6239
rect 36136 6208 37105 6236
rect 36136 6196 36142 6208
rect 37093 6205 37105 6208
rect 37139 6236 37151 6239
rect 37645 6239 37703 6245
rect 37645 6236 37657 6239
rect 37139 6208 37657 6236
rect 37139 6205 37151 6208
rect 37093 6199 37151 6205
rect 37645 6205 37657 6208
rect 37691 6205 37703 6239
rect 37645 6199 37703 6205
rect 26237 6103 26295 6109
rect 26237 6069 26249 6103
rect 26283 6100 26295 6103
rect 26510 6100 26516 6112
rect 26283 6072 26516 6100
rect 26283 6069 26295 6072
rect 26237 6063 26295 6069
rect 26510 6060 26516 6072
rect 26568 6100 26574 6112
rect 26694 6100 26700 6112
rect 26568 6072 26700 6100
rect 26568 6060 26574 6072
rect 26694 6060 26700 6072
rect 26752 6060 26758 6112
rect 27157 6103 27215 6109
rect 27157 6069 27169 6103
rect 27203 6100 27215 6103
rect 27982 6100 27988 6112
rect 27203 6072 27988 6100
rect 27203 6069 27215 6072
rect 27157 6063 27215 6069
rect 27982 6060 27988 6072
rect 28040 6060 28046 6112
rect 28718 6100 28724 6112
rect 28679 6072 28724 6100
rect 28718 6060 28724 6072
rect 28776 6060 28782 6112
rect 28994 6060 29000 6112
rect 29052 6100 29058 6112
rect 29641 6103 29699 6109
rect 29641 6100 29653 6103
rect 29052 6072 29653 6100
rect 29052 6060 29058 6072
rect 29641 6069 29653 6072
rect 29687 6069 29699 6103
rect 29641 6063 29699 6069
rect 31021 6103 31079 6109
rect 31021 6069 31033 6103
rect 31067 6100 31079 6103
rect 31110 6100 31116 6112
rect 31067 6072 31116 6100
rect 31067 6069 31079 6072
rect 31021 6063 31079 6069
rect 31110 6060 31116 6072
rect 31168 6060 31174 6112
rect 31294 6100 31300 6112
rect 31255 6072 31300 6100
rect 31294 6060 31300 6072
rect 31352 6060 31358 6112
rect 31662 6100 31668 6112
rect 31623 6072 31668 6100
rect 31662 6060 31668 6072
rect 31720 6060 31726 6112
rect 32950 6060 32956 6112
rect 33008 6100 33014 6112
rect 33321 6103 33379 6109
rect 33321 6100 33333 6103
rect 33008 6072 33333 6100
rect 33008 6060 33014 6072
rect 33321 6069 33333 6072
rect 33367 6069 33379 6103
rect 34606 6100 34612 6112
rect 34567 6072 34612 6100
rect 33321 6063 33379 6069
rect 34606 6060 34612 6072
rect 34664 6060 34670 6112
rect 35066 6100 35072 6112
rect 35027 6072 35072 6100
rect 35066 6060 35072 6072
rect 35124 6060 35130 6112
rect 35434 6100 35440 6112
rect 35395 6072 35440 6100
rect 35434 6060 35440 6072
rect 35492 6060 35498 6112
rect 35894 6060 35900 6112
rect 35952 6100 35958 6112
rect 36173 6103 36231 6109
rect 36173 6100 36185 6103
rect 35952 6072 36185 6100
rect 35952 6060 35958 6072
rect 36173 6069 36185 6072
rect 36219 6069 36231 6103
rect 36173 6063 36231 6069
rect 1104 6010 38824 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 38824 6010
rect 1104 5936 38824 5958
rect 27982 5856 27988 5908
rect 28040 5896 28046 5908
rect 28721 5899 28779 5905
rect 28721 5896 28733 5899
rect 28040 5868 28733 5896
rect 28040 5856 28046 5868
rect 28721 5865 28733 5868
rect 28767 5865 28779 5899
rect 28721 5859 28779 5865
rect 31389 5899 31447 5905
rect 31389 5865 31401 5899
rect 31435 5896 31447 5899
rect 31662 5896 31668 5908
rect 31435 5868 31668 5896
rect 31435 5865 31447 5868
rect 31389 5859 31447 5865
rect 31662 5856 31668 5868
rect 31720 5856 31726 5908
rect 33505 5899 33563 5905
rect 33505 5865 33517 5899
rect 33551 5896 33563 5899
rect 33870 5896 33876 5908
rect 33551 5868 33876 5896
rect 33551 5865 33563 5868
rect 33505 5859 33563 5865
rect 33870 5856 33876 5868
rect 33928 5896 33934 5908
rect 35066 5896 35072 5908
rect 33928 5868 35072 5896
rect 33928 5856 33934 5868
rect 35066 5856 35072 5868
rect 35124 5856 35130 5908
rect 27430 5788 27436 5840
rect 27488 5828 27494 5840
rect 27608 5831 27666 5837
rect 27608 5828 27620 5831
rect 27488 5800 27620 5828
rect 27488 5788 27494 5800
rect 27608 5797 27620 5800
rect 27654 5828 27666 5831
rect 27890 5828 27896 5840
rect 27654 5800 27896 5828
rect 27654 5797 27666 5800
rect 27608 5791 27666 5797
rect 27890 5788 27896 5800
rect 27948 5788 27954 5840
rect 29822 5788 29828 5840
rect 29880 5828 29886 5840
rect 30282 5828 30288 5840
rect 29880 5800 30288 5828
rect 29880 5788 29886 5800
rect 30282 5788 30288 5800
rect 30340 5788 30346 5840
rect 31294 5788 31300 5840
rect 31352 5828 31358 5840
rect 31938 5828 31944 5840
rect 31352 5800 31800 5828
rect 31899 5800 31944 5828
rect 31352 5788 31358 5800
rect 30190 5760 30196 5772
rect 30151 5732 30196 5760
rect 30190 5720 30196 5732
rect 30248 5720 30254 5772
rect 30300 5760 30328 5788
rect 31772 5760 31800 5800
rect 31938 5788 31944 5800
rect 31996 5788 32002 5840
rect 32950 5828 32956 5840
rect 32911 5800 32956 5828
rect 32950 5788 32956 5800
rect 33008 5788 33014 5840
rect 33594 5828 33600 5840
rect 33507 5800 33600 5828
rect 33594 5788 33600 5800
rect 33652 5828 33658 5840
rect 35526 5828 35532 5840
rect 33652 5800 35532 5828
rect 33652 5788 33658 5800
rect 35526 5788 35532 5800
rect 35584 5788 35590 5840
rect 32968 5760 32996 5788
rect 30300 5732 30420 5760
rect 31772 5732 32996 5760
rect 26694 5652 26700 5704
rect 26752 5692 26758 5704
rect 27341 5695 27399 5701
rect 27341 5692 27353 5695
rect 26752 5664 27353 5692
rect 26752 5652 26758 5664
rect 27341 5661 27353 5664
rect 27387 5661 27399 5695
rect 27341 5655 27399 5661
rect 30098 5652 30104 5704
rect 30156 5692 30162 5704
rect 30392 5701 30420 5732
rect 34790 5720 34796 5772
rect 34848 5760 34854 5772
rect 35345 5763 35403 5769
rect 35345 5760 35357 5763
rect 34848 5732 35357 5760
rect 34848 5720 34854 5732
rect 35345 5729 35357 5732
rect 35391 5729 35403 5763
rect 35345 5723 35403 5729
rect 30285 5695 30343 5701
rect 30285 5692 30297 5695
rect 30156 5664 30297 5692
rect 30156 5652 30162 5664
rect 30285 5661 30297 5664
rect 30331 5661 30343 5695
rect 30285 5655 30343 5661
rect 30377 5695 30435 5701
rect 30377 5661 30389 5695
rect 30423 5661 30435 5695
rect 30377 5655 30435 5661
rect 33410 5652 33416 5704
rect 33468 5692 33474 5704
rect 33781 5695 33839 5701
rect 33781 5692 33793 5695
rect 33468 5664 33793 5692
rect 33468 5652 33474 5664
rect 33781 5661 33793 5664
rect 33827 5692 33839 5695
rect 34238 5692 34244 5704
rect 33827 5664 34244 5692
rect 33827 5661 33839 5664
rect 33781 5655 33839 5661
rect 34238 5652 34244 5664
rect 34296 5652 34302 5704
rect 34422 5652 34428 5704
rect 34480 5692 34486 5704
rect 34882 5692 34888 5704
rect 34480 5664 34888 5692
rect 34480 5652 34486 5664
rect 34882 5652 34888 5664
rect 34940 5652 34946 5704
rect 35250 5652 35256 5704
rect 35308 5692 35314 5704
rect 35437 5695 35495 5701
rect 35437 5692 35449 5695
rect 35308 5664 35449 5692
rect 35308 5652 35314 5664
rect 35437 5661 35449 5664
rect 35483 5661 35495 5695
rect 35437 5655 35495 5661
rect 35526 5652 35532 5704
rect 35584 5692 35590 5704
rect 35584 5664 35629 5692
rect 35584 5652 35590 5664
rect 29733 5627 29791 5633
rect 29733 5593 29745 5627
rect 29779 5624 29791 5627
rect 31110 5624 31116 5636
rect 29779 5596 31116 5624
rect 29779 5593 29791 5596
rect 29733 5587 29791 5593
rect 31110 5584 31116 5596
rect 31168 5584 31174 5636
rect 33134 5624 33140 5636
rect 33095 5596 33140 5624
rect 33134 5584 33140 5596
rect 33192 5584 33198 5636
rect 34514 5584 34520 5636
rect 34572 5624 34578 5636
rect 34977 5627 35035 5633
rect 34977 5624 34989 5627
rect 34572 5596 34989 5624
rect 34572 5584 34578 5596
rect 34977 5593 34989 5596
rect 35023 5593 35035 5627
rect 34977 5587 35035 5593
rect 28994 5516 29000 5568
rect 29052 5556 29058 5568
rect 29273 5559 29331 5565
rect 29273 5556 29285 5559
rect 29052 5528 29285 5556
rect 29052 5516 29058 5528
rect 29273 5525 29285 5528
rect 29319 5525 29331 5559
rect 29822 5556 29828 5568
rect 29783 5528 29828 5556
rect 29273 5519 29331 5525
rect 29822 5516 29828 5528
rect 29880 5516 29886 5568
rect 32493 5559 32551 5565
rect 32493 5525 32505 5559
rect 32539 5556 32551 5559
rect 32766 5556 32772 5568
rect 32539 5528 32772 5556
rect 32539 5525 32551 5528
rect 32493 5519 32551 5525
rect 32766 5516 32772 5528
rect 32824 5516 32830 5568
rect 36081 5559 36139 5565
rect 36081 5525 36093 5559
rect 36127 5556 36139 5559
rect 36262 5556 36268 5568
rect 36127 5528 36268 5556
rect 36127 5525 36139 5528
rect 36081 5519 36139 5525
rect 36262 5516 36268 5528
rect 36320 5516 36326 5568
rect 1104 5466 38824 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 34966 5466
rect 35018 5414 35030 5466
rect 35082 5414 35094 5466
rect 35146 5414 35158 5466
rect 35210 5414 38824 5466
rect 1104 5392 38824 5414
rect 27430 5352 27436 5364
rect 27391 5324 27436 5352
rect 27430 5312 27436 5324
rect 27488 5312 27494 5364
rect 27617 5355 27675 5361
rect 27617 5321 27629 5355
rect 27663 5352 27675 5355
rect 28902 5352 28908 5364
rect 27663 5324 28908 5352
rect 27663 5321 27675 5324
rect 27617 5315 27675 5321
rect 28902 5312 28908 5324
rect 28960 5312 28966 5364
rect 30374 5312 30380 5364
rect 30432 5352 30438 5364
rect 31205 5355 31263 5361
rect 31205 5352 31217 5355
rect 30432 5324 31217 5352
rect 30432 5312 30438 5324
rect 31205 5321 31217 5324
rect 31251 5321 31263 5355
rect 32398 5352 32404 5364
rect 32359 5324 32404 5352
rect 31205 5315 31263 5321
rect 28261 5219 28319 5225
rect 28261 5185 28273 5219
rect 28307 5216 28319 5219
rect 28718 5216 28724 5228
rect 28307 5188 28724 5216
rect 28307 5185 28319 5188
rect 28261 5179 28319 5185
rect 28718 5176 28724 5188
rect 28776 5176 28782 5228
rect 31220 5216 31248 5315
rect 32398 5312 32404 5324
rect 32456 5312 32462 5364
rect 33505 5355 33563 5361
rect 33505 5321 33517 5355
rect 33551 5352 33563 5355
rect 33594 5352 33600 5364
rect 33551 5324 33600 5352
rect 33551 5321 33563 5324
rect 33505 5315 33563 5321
rect 33594 5312 33600 5324
rect 33652 5312 33658 5364
rect 33870 5352 33876 5364
rect 33831 5324 33876 5352
rect 33870 5312 33876 5324
rect 33928 5312 33934 5364
rect 34238 5352 34244 5364
rect 34199 5324 34244 5352
rect 34238 5312 34244 5324
rect 34296 5312 34302 5364
rect 36170 5312 36176 5364
rect 36228 5352 36234 5364
rect 36817 5355 36875 5361
rect 36817 5352 36829 5355
rect 36228 5324 36829 5352
rect 36228 5312 36234 5324
rect 36817 5321 36829 5324
rect 36863 5321 36875 5355
rect 36817 5315 36875 5321
rect 31941 5219 31999 5225
rect 31941 5216 31953 5219
rect 31220 5188 31953 5216
rect 31941 5185 31953 5188
rect 31987 5216 31999 5219
rect 33042 5216 33048 5228
rect 31987 5188 33048 5216
rect 31987 5185 31999 5188
rect 31941 5179 31999 5185
rect 33042 5176 33048 5188
rect 33100 5176 33106 5228
rect 34422 5176 34428 5228
rect 34480 5216 34486 5228
rect 35158 5216 35164 5228
rect 34480 5188 35164 5216
rect 34480 5176 34486 5188
rect 34716 5160 34744 5188
rect 35158 5176 35164 5188
rect 35216 5216 35222 5228
rect 35437 5219 35495 5225
rect 35437 5216 35449 5219
rect 35216 5188 35449 5216
rect 35216 5176 35222 5188
rect 35437 5185 35449 5188
rect 35483 5185 35495 5219
rect 35437 5179 35495 5185
rect 29270 5148 29276 5160
rect 29231 5120 29276 5148
rect 29270 5108 29276 5120
rect 29328 5108 29334 5160
rect 34698 5108 34704 5160
rect 34756 5108 34762 5160
rect 28997 5083 29055 5089
rect 28997 5080 29009 5083
rect 28092 5052 29009 5080
rect 28092 5024 28120 5052
rect 28997 5049 29009 5052
rect 29043 5080 29055 5083
rect 29518 5083 29576 5089
rect 29518 5080 29530 5083
rect 29043 5052 29530 5080
rect 29043 5049 29055 5052
rect 28997 5043 29055 5049
rect 29518 5049 29530 5052
rect 29564 5049 29576 5083
rect 32861 5083 32919 5089
rect 32861 5080 32873 5083
rect 29518 5043 29576 5049
rect 32232 5052 32873 5080
rect 32232 5024 32260 5052
rect 32861 5049 32873 5052
rect 32907 5049 32919 5083
rect 32861 5043 32919 5049
rect 35704 5083 35762 5089
rect 35704 5049 35716 5083
rect 35750 5080 35762 5083
rect 36262 5080 36268 5092
rect 35750 5052 36268 5080
rect 35750 5049 35762 5052
rect 35704 5043 35762 5049
rect 36262 5040 36268 5052
rect 36320 5040 36326 5092
rect 26694 5012 26700 5024
rect 26655 4984 26700 5012
rect 26694 4972 26700 4984
rect 26752 4972 26758 5024
rect 27065 5015 27123 5021
rect 27065 4981 27077 5015
rect 27111 5012 27123 5015
rect 27890 5012 27896 5024
rect 27111 4984 27896 5012
rect 27111 4981 27123 4984
rect 27065 4975 27123 4981
rect 27890 4972 27896 4984
rect 27948 5012 27954 5024
rect 27985 5015 28043 5021
rect 27985 5012 27997 5015
rect 27948 4984 27997 5012
rect 27948 4972 27954 4984
rect 27985 4981 27997 4984
rect 28031 4981 28043 5015
rect 27985 4975 28043 4981
rect 28074 4972 28080 5024
rect 28132 5012 28138 5024
rect 28718 5012 28724 5024
rect 28132 4984 28177 5012
rect 28679 4984 28724 5012
rect 28132 4972 28138 4984
rect 28718 4972 28724 4984
rect 28776 4972 28782 5024
rect 30374 4972 30380 5024
rect 30432 5012 30438 5024
rect 30653 5015 30711 5021
rect 30653 5012 30665 5015
rect 30432 4984 30665 5012
rect 30432 4972 30438 4984
rect 30653 4981 30665 4984
rect 30699 4981 30711 5015
rect 32214 5012 32220 5024
rect 32175 4984 32220 5012
rect 30653 4975 30711 4981
rect 32214 4972 32220 4984
rect 32272 4972 32278 5024
rect 32766 5012 32772 5024
rect 32727 4984 32772 5012
rect 32766 4972 32772 4984
rect 32824 4972 32830 5024
rect 34701 5015 34759 5021
rect 34701 4981 34713 5015
rect 34747 5012 34759 5015
rect 34790 5012 34796 5024
rect 34747 4984 34796 5012
rect 34747 4981 34759 4984
rect 34701 4975 34759 4981
rect 34790 4972 34796 4984
rect 34848 4972 34854 5024
rect 35161 5015 35219 5021
rect 35161 4981 35173 5015
rect 35207 5012 35219 5015
rect 35250 5012 35256 5024
rect 35207 4984 35256 5012
rect 35207 4981 35219 4984
rect 35161 4975 35219 4981
rect 35250 4972 35256 4984
rect 35308 4972 35314 5024
rect 1104 4922 38824 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 38824 4922
rect 1104 4848 38824 4870
rect 27709 4811 27767 4817
rect 27709 4777 27721 4811
rect 27755 4808 27767 4811
rect 28074 4808 28080 4820
rect 27755 4780 28080 4808
rect 27755 4777 27767 4780
rect 27709 4771 27767 4777
rect 28074 4768 28080 4780
rect 28132 4808 28138 4820
rect 29273 4811 29331 4817
rect 29273 4808 29285 4811
rect 28132 4780 29285 4808
rect 28132 4768 28138 4780
rect 29273 4777 29285 4780
rect 29319 4777 29331 4811
rect 30190 4808 30196 4820
rect 30151 4780 30196 4808
rect 29273 4771 29331 4777
rect 30190 4768 30196 4780
rect 30248 4808 30254 4820
rect 30377 4811 30435 4817
rect 30377 4808 30389 4811
rect 30248 4780 30389 4808
rect 30248 4768 30254 4780
rect 30377 4777 30389 4780
rect 30423 4777 30435 4811
rect 30377 4771 30435 4777
rect 31754 4768 31760 4820
rect 31812 4808 31818 4820
rect 32309 4811 32367 4817
rect 32309 4808 32321 4811
rect 31812 4780 32321 4808
rect 31812 4768 31818 4780
rect 32309 4777 32321 4780
rect 32355 4777 32367 4811
rect 32309 4771 32367 4777
rect 33597 4811 33655 4817
rect 33597 4777 33609 4811
rect 33643 4777 33655 4811
rect 33597 4771 33655 4777
rect 27982 4700 27988 4752
rect 28040 4740 28046 4752
rect 28160 4743 28218 4749
rect 28160 4740 28172 4743
rect 28040 4712 28172 4740
rect 28040 4700 28046 4712
rect 28160 4709 28172 4712
rect 28206 4709 28218 4743
rect 33612 4740 33640 4771
rect 33778 4768 33784 4820
rect 33836 4808 33842 4820
rect 34057 4811 34115 4817
rect 34057 4808 34069 4811
rect 33836 4780 34069 4808
rect 33836 4768 33842 4780
rect 34057 4777 34069 4780
rect 34103 4808 34115 4811
rect 34422 4808 34428 4820
rect 34103 4780 34428 4808
rect 34103 4777 34115 4780
rect 34057 4771 34115 4777
rect 34422 4768 34428 4780
rect 34480 4768 34486 4820
rect 34698 4808 34704 4820
rect 34659 4780 34704 4808
rect 34698 4768 34704 4780
rect 34756 4768 34762 4820
rect 34606 4740 34612 4752
rect 33612 4712 34612 4740
rect 28160 4703 28218 4709
rect 34606 4700 34612 4712
rect 34664 4700 34670 4752
rect 26694 4632 26700 4684
rect 26752 4672 26758 4684
rect 27893 4675 27951 4681
rect 27893 4672 27905 4675
rect 26752 4644 27905 4672
rect 26752 4632 26758 4644
rect 27893 4641 27905 4644
rect 27939 4672 27951 4675
rect 28442 4672 28448 4684
rect 27939 4644 28448 4672
rect 27939 4641 27951 4644
rect 27893 4635 27951 4641
rect 28442 4632 28448 4644
rect 28500 4632 28506 4684
rect 30742 4672 30748 4684
rect 30703 4644 30748 4672
rect 30742 4632 30748 4644
rect 30800 4632 30806 4684
rect 30837 4675 30895 4681
rect 30837 4641 30849 4675
rect 30883 4672 30895 4675
rect 31202 4672 31208 4684
rect 30883 4644 31208 4672
rect 30883 4641 30895 4644
rect 30837 4635 30895 4641
rect 31202 4632 31208 4644
rect 31260 4632 31266 4684
rect 32122 4672 32128 4684
rect 32083 4644 32128 4672
rect 32122 4632 32128 4644
rect 32180 4672 32186 4684
rect 32677 4675 32735 4681
rect 32677 4672 32689 4675
rect 32180 4644 32689 4672
rect 32180 4632 32186 4644
rect 32677 4641 32689 4644
rect 32723 4641 32735 4675
rect 32677 4635 32735 4641
rect 33965 4675 34023 4681
rect 33965 4641 33977 4675
rect 34011 4672 34023 4675
rect 34054 4672 34060 4684
rect 34011 4644 34060 4672
rect 34011 4641 34023 4644
rect 33965 4635 34023 4641
rect 34054 4632 34060 4644
rect 34112 4632 34118 4684
rect 34698 4632 34704 4684
rect 34756 4672 34762 4684
rect 35417 4675 35475 4681
rect 35417 4672 35429 4675
rect 34756 4644 35429 4672
rect 34756 4632 34762 4644
rect 35417 4641 35429 4644
rect 35463 4641 35475 4675
rect 35417 4635 35475 4641
rect 31018 4604 31024 4616
rect 30979 4576 31024 4604
rect 31018 4564 31024 4576
rect 31076 4564 31082 4616
rect 33042 4564 33048 4616
rect 33100 4604 33106 4616
rect 33505 4607 33563 4613
rect 33505 4604 33517 4607
rect 33100 4576 33517 4604
rect 33100 4564 33106 4576
rect 33505 4573 33517 4576
rect 33551 4604 33563 4607
rect 34238 4604 34244 4616
rect 33551 4576 34244 4604
rect 33551 4573 33563 4576
rect 33505 4567 33563 4573
rect 34238 4564 34244 4576
rect 34296 4564 34302 4616
rect 34974 4604 34980 4616
rect 34935 4576 34980 4604
rect 34974 4564 34980 4576
rect 35032 4564 35038 4616
rect 35158 4604 35164 4616
rect 35119 4576 35164 4604
rect 35158 4564 35164 4576
rect 35216 4564 35222 4616
rect 28994 4428 29000 4480
rect 29052 4468 29058 4480
rect 29825 4471 29883 4477
rect 29825 4468 29837 4471
rect 29052 4440 29837 4468
rect 29052 4428 29058 4440
rect 29825 4437 29837 4440
rect 29871 4468 29883 4471
rect 30098 4468 30104 4480
rect 29871 4440 30104 4468
rect 29871 4437 29883 4440
rect 29825 4431 29883 4437
rect 30098 4428 30104 4440
rect 30156 4428 30162 4480
rect 35176 4468 35204 4564
rect 35526 4468 35532 4480
rect 35176 4440 35532 4468
rect 35526 4428 35532 4440
rect 35584 4428 35590 4480
rect 36262 4428 36268 4480
rect 36320 4468 36326 4480
rect 36541 4471 36599 4477
rect 36541 4468 36553 4471
rect 36320 4440 36553 4468
rect 36320 4428 36326 4440
rect 36541 4437 36553 4440
rect 36587 4437 36599 4471
rect 36541 4431 36599 4437
rect 1104 4378 38824 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 34966 4378
rect 35018 4326 35030 4378
rect 35082 4326 35094 4378
rect 35146 4326 35158 4378
rect 35210 4326 38824 4378
rect 1104 4304 38824 4326
rect 27982 4224 27988 4276
rect 28040 4264 28046 4276
rect 28629 4267 28687 4273
rect 28629 4264 28641 4267
rect 28040 4236 28641 4264
rect 28040 4224 28046 4236
rect 28629 4233 28641 4236
rect 28675 4233 28687 4267
rect 33778 4264 33784 4276
rect 33739 4236 33784 4264
rect 28629 4227 28687 4233
rect 33778 4224 33784 4236
rect 33836 4224 33842 4276
rect 34698 4264 34704 4276
rect 34659 4236 34704 4264
rect 34698 4224 34704 4236
rect 34756 4224 34762 4276
rect 27890 4156 27896 4208
rect 27948 4196 27954 4208
rect 27948 4168 28948 4196
rect 27948 4156 27954 4168
rect 27157 4131 27215 4137
rect 27157 4097 27169 4131
rect 27203 4128 27215 4131
rect 27982 4128 27988 4140
rect 27203 4100 27988 4128
rect 27203 4097 27215 4100
rect 27157 4091 27215 4097
rect 27982 4088 27988 4100
rect 28040 4088 28046 4140
rect 28166 4088 28172 4140
rect 28224 4128 28230 4140
rect 28261 4131 28319 4137
rect 28261 4128 28273 4131
rect 28224 4100 28273 4128
rect 28224 4088 28230 4100
rect 28261 4097 28273 4100
rect 28307 4128 28319 4131
rect 28718 4128 28724 4140
rect 28307 4100 28724 4128
rect 28307 4097 28319 4100
rect 28261 4091 28319 4097
rect 28718 4088 28724 4100
rect 28776 4088 28782 4140
rect 28920 4128 28948 4168
rect 29089 4131 29147 4137
rect 29089 4128 29101 4131
rect 28920 4100 29101 4128
rect 29089 4097 29101 4100
rect 29135 4128 29147 4131
rect 29135 4100 29408 4128
rect 29135 4097 29147 4100
rect 29089 4091 29147 4097
rect 27525 4063 27583 4069
rect 27525 4029 27537 4063
rect 27571 4060 27583 4063
rect 28077 4063 28135 4069
rect 28077 4060 28089 4063
rect 27571 4032 28089 4060
rect 27571 4029 27583 4032
rect 27525 4023 27583 4029
rect 28077 4029 28089 4032
rect 28123 4060 28135 4063
rect 28994 4060 29000 4072
rect 28123 4032 29000 4060
rect 28123 4029 28135 4032
rect 28077 4023 28135 4029
rect 28994 4020 29000 4032
rect 29052 4020 29058 4072
rect 29270 4060 29276 4072
rect 29231 4032 29276 4060
rect 29270 4020 29276 4032
rect 29328 4020 29334 4072
rect 29380 4060 29408 4100
rect 31110 4088 31116 4140
rect 31168 4128 31174 4140
rect 31168 4100 31800 4128
rect 31168 4088 31174 4100
rect 31772 4072 31800 4100
rect 29529 4063 29587 4069
rect 29529 4060 29541 4063
rect 29380 4032 29541 4060
rect 29529 4029 29541 4032
rect 29575 4060 29587 4063
rect 30282 4060 30288 4072
rect 29575 4032 30288 4060
rect 29575 4029 29587 4032
rect 29529 4023 29587 4029
rect 30282 4020 30288 4032
rect 30340 4020 30346 4072
rect 30742 4020 30748 4072
rect 30800 4060 30806 4072
rect 31573 4063 31631 4069
rect 31573 4060 31585 4063
rect 30800 4032 31585 4060
rect 30800 4020 30806 4032
rect 31573 4029 31585 4032
rect 31619 4029 31631 4063
rect 31754 4060 31760 4072
rect 31715 4032 31760 4060
rect 31573 4023 31631 4029
rect 28902 3992 28908 4004
rect 27632 3964 28908 3992
rect 26786 3924 26792 3936
rect 26747 3896 26792 3924
rect 26786 3884 26792 3896
rect 26844 3884 26850 3936
rect 27632 3933 27660 3964
rect 28902 3952 28908 3964
rect 28960 3952 28966 4004
rect 31202 3992 31208 4004
rect 31163 3964 31208 3992
rect 31202 3952 31208 3964
rect 31260 3952 31266 4004
rect 31588 3992 31616 4023
rect 31754 4020 31760 4032
rect 31812 4020 31818 4072
rect 35437 4063 35495 4069
rect 35437 4029 35449 4063
rect 35483 4060 35495 4063
rect 35526 4060 35532 4072
rect 35483 4032 35532 4060
rect 35483 4029 35495 4032
rect 35437 4023 35495 4029
rect 35526 4020 35532 4032
rect 35584 4020 35590 4072
rect 32002 3995 32060 4001
rect 32002 3992 32014 3995
rect 31588 3964 32014 3992
rect 32002 3961 32014 3964
rect 32048 3961 32060 3995
rect 32002 3955 32060 3961
rect 34790 3952 34796 4004
rect 34848 3992 34854 4004
rect 35345 3995 35403 4001
rect 35345 3992 35357 3995
rect 34848 3964 35357 3992
rect 34848 3952 34854 3964
rect 35345 3961 35357 3964
rect 35391 3992 35403 3995
rect 35704 3995 35762 4001
rect 35704 3992 35716 3995
rect 35391 3964 35716 3992
rect 35391 3961 35403 3964
rect 35345 3955 35403 3961
rect 35704 3961 35716 3964
rect 35750 3992 35762 3995
rect 35802 3992 35808 4004
rect 35750 3964 35808 3992
rect 35750 3961 35762 3964
rect 35704 3955 35762 3961
rect 35802 3952 35808 3964
rect 35860 3952 35866 4004
rect 27617 3927 27675 3933
rect 27617 3893 27629 3927
rect 27663 3893 27675 3927
rect 27982 3924 27988 3936
rect 27943 3896 27988 3924
rect 27617 3887 27675 3893
rect 27982 3884 27988 3896
rect 28040 3924 28046 3936
rect 29362 3924 29368 3936
rect 28040 3896 29368 3924
rect 28040 3884 28046 3896
rect 29362 3884 29368 3896
rect 29420 3884 29426 3936
rect 30650 3924 30656 3936
rect 30611 3896 30656 3924
rect 30650 3884 30656 3896
rect 30708 3884 30714 3936
rect 33134 3924 33140 3936
rect 33095 3896 33140 3924
rect 33134 3884 33140 3896
rect 33192 3884 33198 3936
rect 34146 3924 34152 3936
rect 34107 3896 34152 3924
rect 34146 3884 34152 3896
rect 34204 3884 34210 3936
rect 36814 3924 36820 3936
rect 36775 3896 36820 3924
rect 36814 3884 36820 3896
rect 36872 3884 36878 3936
rect 1104 3834 38824 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 38824 3834
rect 1104 3760 38824 3782
rect 27338 3720 27344 3732
rect 27299 3692 27344 3720
rect 27338 3680 27344 3692
rect 27396 3680 27402 3732
rect 28442 3720 28448 3732
rect 28403 3692 28448 3720
rect 28442 3680 28448 3692
rect 28500 3680 28506 3732
rect 28813 3723 28871 3729
rect 28813 3689 28825 3723
rect 28859 3720 28871 3723
rect 29270 3720 29276 3732
rect 28859 3692 29276 3720
rect 28859 3689 28871 3692
rect 28813 3683 28871 3689
rect 26786 3612 26792 3664
rect 26844 3652 26850 3664
rect 26844 3624 28028 3652
rect 26844 3612 26850 3624
rect 27706 3584 27712 3596
rect 27667 3556 27712 3584
rect 27706 3544 27712 3556
rect 27764 3544 27770 3596
rect 27798 3516 27804 3528
rect 27759 3488 27804 3516
rect 27798 3476 27804 3488
rect 27856 3476 27862 3528
rect 28000 3525 28028 3624
rect 28920 3593 28948 3692
rect 29270 3680 29276 3692
rect 29328 3680 29334 3732
rect 29362 3680 29368 3732
rect 29420 3720 29426 3732
rect 30285 3723 30343 3729
rect 30285 3720 30297 3723
rect 29420 3692 30297 3720
rect 29420 3680 29426 3692
rect 30285 3689 30297 3692
rect 30331 3689 30343 3723
rect 30285 3683 30343 3689
rect 31018 3680 31024 3732
rect 31076 3720 31082 3732
rect 31205 3723 31263 3729
rect 31205 3720 31217 3723
rect 31076 3692 31217 3720
rect 31076 3680 31082 3692
rect 31205 3689 31217 3692
rect 31251 3689 31263 3723
rect 31205 3683 31263 3689
rect 35437 3723 35495 3729
rect 35437 3689 35449 3723
rect 35483 3720 35495 3723
rect 35526 3720 35532 3732
rect 35483 3692 35532 3720
rect 35483 3689 35495 3692
rect 35437 3683 35495 3689
rect 35526 3680 35532 3692
rect 35584 3720 35590 3732
rect 35713 3723 35771 3729
rect 35713 3720 35725 3723
rect 35584 3692 35725 3720
rect 35584 3680 35590 3692
rect 35713 3689 35725 3692
rect 35759 3689 35771 3723
rect 35894 3720 35900 3732
rect 35855 3692 35900 3720
rect 35713 3683 35771 3689
rect 35894 3680 35900 3692
rect 35952 3680 35958 3732
rect 28994 3612 29000 3664
rect 29052 3652 29058 3664
rect 29172 3655 29230 3661
rect 29172 3652 29184 3655
rect 29052 3624 29184 3652
rect 29052 3612 29058 3624
rect 29172 3621 29184 3624
rect 29218 3652 29230 3655
rect 30650 3652 30656 3664
rect 29218 3624 30656 3652
rect 29218 3621 29230 3624
rect 29172 3615 29230 3621
rect 30650 3612 30656 3624
rect 30708 3612 30714 3664
rect 34698 3612 34704 3664
rect 34756 3652 34762 3664
rect 36357 3655 36415 3661
rect 36357 3652 36369 3655
rect 34756 3624 36369 3652
rect 34756 3612 34762 3624
rect 36357 3621 36369 3624
rect 36403 3652 36415 3655
rect 36814 3652 36820 3664
rect 36403 3624 36820 3652
rect 36403 3621 36415 3624
rect 36357 3615 36415 3621
rect 36814 3612 36820 3624
rect 36872 3612 36878 3664
rect 28905 3587 28963 3593
rect 28905 3553 28917 3587
rect 28951 3553 28963 3587
rect 28905 3547 28963 3553
rect 32309 3587 32367 3593
rect 32309 3553 32321 3587
rect 32355 3584 32367 3587
rect 32398 3584 32404 3596
rect 32355 3556 32404 3584
rect 32355 3553 32367 3556
rect 32309 3547 32367 3553
rect 32398 3544 32404 3556
rect 32456 3584 32462 3596
rect 33042 3584 33048 3596
rect 32456 3556 33048 3584
rect 32456 3544 32462 3556
rect 33042 3544 33048 3556
rect 33100 3544 33106 3596
rect 33686 3593 33692 3596
rect 33680 3584 33692 3593
rect 33647 3556 33692 3584
rect 33680 3547 33692 3556
rect 33686 3544 33692 3547
rect 33744 3544 33750 3596
rect 36262 3584 36268 3596
rect 36223 3556 36268 3584
rect 36262 3544 36268 3556
rect 36320 3544 36326 3596
rect 27985 3519 28043 3525
rect 27985 3485 27997 3519
rect 28031 3516 28043 3519
rect 28166 3516 28172 3528
rect 28031 3488 28172 3516
rect 28031 3485 28043 3488
rect 27985 3479 28043 3485
rect 28166 3476 28172 3488
rect 28224 3476 28230 3528
rect 31754 3476 31760 3528
rect 31812 3516 31818 3528
rect 31849 3519 31907 3525
rect 31849 3516 31861 3519
rect 31812 3488 31861 3516
rect 31812 3476 31818 3488
rect 31849 3485 31861 3488
rect 31895 3516 31907 3519
rect 32953 3519 33011 3525
rect 32953 3516 32965 3519
rect 31895 3488 32965 3516
rect 31895 3485 31907 3488
rect 31849 3479 31907 3485
rect 32953 3485 32965 3488
rect 32999 3516 33011 3519
rect 33410 3516 33416 3528
rect 32999 3488 33416 3516
rect 32999 3485 33011 3488
rect 32953 3479 33011 3485
rect 33410 3476 33416 3488
rect 33468 3476 33474 3528
rect 36446 3516 36452 3528
rect 36407 3488 36452 3516
rect 36446 3476 36452 3488
rect 36504 3476 36510 3528
rect 32490 3448 32496 3460
rect 32451 3420 32496 3448
rect 32490 3408 32496 3420
rect 32548 3408 32554 3460
rect 30742 3340 30748 3392
rect 30800 3380 30806 3392
rect 30837 3383 30895 3389
rect 30837 3380 30849 3383
rect 30800 3352 30849 3380
rect 30800 3340 30806 3352
rect 30837 3349 30849 3352
rect 30883 3349 30895 3383
rect 30837 3343 30895 3349
rect 34606 3340 34612 3392
rect 34664 3380 34670 3392
rect 34793 3383 34851 3389
rect 34793 3380 34805 3383
rect 34664 3352 34805 3380
rect 34664 3340 34670 3352
rect 34793 3349 34805 3352
rect 34839 3349 34851 3383
rect 34793 3343 34851 3349
rect 1104 3290 38824 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 34966 3290
rect 35018 3238 35030 3290
rect 35082 3238 35094 3290
rect 35146 3238 35158 3290
rect 35210 3238 38824 3290
rect 1104 3216 38824 3238
rect 27157 3179 27215 3185
rect 27157 3145 27169 3179
rect 27203 3176 27215 3179
rect 27798 3176 27804 3188
rect 27203 3148 27804 3176
rect 27203 3145 27215 3148
rect 27157 3139 27215 3145
rect 27798 3136 27804 3148
rect 27856 3136 27862 3188
rect 28994 3176 29000 3188
rect 28955 3148 29000 3176
rect 28994 3136 29000 3148
rect 29052 3136 29058 3188
rect 31570 3176 31576 3188
rect 31531 3148 31576 3176
rect 31570 3136 31576 3148
rect 31628 3176 31634 3188
rect 32030 3176 32036 3188
rect 31628 3148 32036 3176
rect 31628 3136 31634 3148
rect 32030 3136 32036 3148
rect 32088 3136 32094 3188
rect 36262 3136 36268 3188
rect 36320 3176 36326 3188
rect 37185 3179 37243 3185
rect 37185 3176 37197 3179
rect 36320 3148 37197 3176
rect 36320 3136 36326 3148
rect 37185 3145 37197 3148
rect 37231 3145 37243 3179
rect 37185 3139 37243 3145
rect 26789 3111 26847 3117
rect 26789 3077 26801 3111
rect 26835 3108 26847 3111
rect 27706 3108 27712 3120
rect 26835 3080 27712 3108
rect 26835 3077 26847 3080
rect 26789 3071 26847 3077
rect 27706 3068 27712 3080
rect 27764 3068 27770 3120
rect 36814 3108 36820 3120
rect 36775 3080 36820 3108
rect 36814 3068 36820 3080
rect 36872 3068 36878 3120
rect 27525 3043 27583 3049
rect 27525 3009 27537 3043
rect 27571 3040 27583 3043
rect 28074 3040 28080 3052
rect 27571 3012 28080 3040
rect 27571 3009 27583 3012
rect 27525 3003 27583 3009
rect 28074 3000 28080 3012
rect 28132 3000 28138 3052
rect 28166 3000 28172 3052
rect 28224 3040 28230 3052
rect 31294 3040 31300 3052
rect 28224 3012 28269 3040
rect 31207 3012 31300 3040
rect 28224 3000 28230 3012
rect 31294 3000 31300 3012
rect 31352 3040 31358 3052
rect 31754 3040 31760 3052
rect 31352 3012 31760 3040
rect 31352 3000 31358 3012
rect 31754 3000 31760 3012
rect 31812 3000 31818 3052
rect 33686 3040 33692 3052
rect 33647 3012 33692 3040
rect 33686 3000 33692 3012
rect 33744 3000 33750 3052
rect 36446 3000 36452 3052
rect 36504 3040 36510 3052
rect 37553 3043 37611 3049
rect 37553 3040 37565 3043
rect 36504 3012 37565 3040
rect 36504 3000 36510 3012
rect 37553 3009 37565 3012
rect 37599 3009 37611 3043
rect 37553 3003 37611 3009
rect 29270 2972 29276 2984
rect 29231 2944 29276 2972
rect 29270 2932 29276 2944
rect 29328 2932 29334 2984
rect 32030 2981 32036 2984
rect 32024 2972 32036 2981
rect 31943 2944 32036 2972
rect 32024 2935 32036 2944
rect 32088 2972 32094 2984
rect 33134 2972 33140 2984
rect 32088 2944 33140 2972
rect 32030 2932 32036 2935
rect 32088 2932 32094 2944
rect 33134 2932 33140 2944
rect 33192 2932 33198 2984
rect 33410 2932 33416 2984
rect 33468 2972 33474 2984
rect 34149 2975 34207 2981
rect 34149 2972 34161 2975
rect 33468 2944 34161 2972
rect 33468 2932 33474 2944
rect 34149 2941 34161 2944
rect 34195 2972 34207 2975
rect 34514 2972 34520 2984
rect 34195 2944 34520 2972
rect 34195 2941 34207 2944
rect 34149 2935 34207 2941
rect 34514 2932 34520 2944
rect 34572 2972 34578 2984
rect 34885 2975 34943 2981
rect 34885 2972 34897 2975
rect 34572 2944 34897 2972
rect 34572 2932 34578 2944
rect 34885 2941 34897 2944
rect 34931 2972 34943 2975
rect 35526 2972 35532 2984
rect 34931 2944 35532 2972
rect 34931 2941 34943 2944
rect 34885 2935 34943 2941
rect 35526 2932 35532 2944
rect 35584 2932 35590 2984
rect 29362 2864 29368 2916
rect 29420 2904 29426 2916
rect 29518 2907 29576 2913
rect 29518 2904 29530 2907
rect 29420 2876 29530 2904
rect 29420 2864 29426 2876
rect 29518 2873 29530 2876
rect 29564 2873 29576 2907
rect 35130 2907 35188 2913
rect 35130 2904 35142 2907
rect 29518 2867 29576 2873
rect 34624 2876 35142 2904
rect 34624 2848 34652 2876
rect 35130 2873 35142 2876
rect 35176 2873 35188 2907
rect 35130 2867 35188 2873
rect 27614 2836 27620 2848
rect 27575 2808 27620 2836
rect 27614 2796 27620 2808
rect 27672 2796 27678 2848
rect 27982 2836 27988 2848
rect 27943 2808 27988 2836
rect 27982 2796 27988 2808
rect 28040 2796 28046 2848
rect 30282 2796 30288 2848
rect 30340 2836 30346 2848
rect 30653 2839 30711 2845
rect 30653 2836 30665 2839
rect 30340 2808 30665 2836
rect 30340 2796 30346 2808
rect 30653 2805 30665 2808
rect 30699 2836 30711 2839
rect 31202 2836 31208 2848
rect 30699 2808 31208 2836
rect 30699 2805 30711 2808
rect 30653 2799 30711 2805
rect 31202 2796 31208 2808
rect 31260 2796 31266 2848
rect 33042 2796 33048 2848
rect 33100 2836 33106 2848
rect 33137 2839 33195 2845
rect 33137 2836 33149 2839
rect 33100 2808 33149 2836
rect 33100 2796 33106 2808
rect 33137 2805 33149 2808
rect 33183 2805 33195 2839
rect 34606 2836 34612 2848
rect 34567 2808 34612 2836
rect 33137 2799 33195 2805
rect 34606 2796 34612 2808
rect 34664 2796 34670 2848
rect 35802 2796 35808 2848
rect 35860 2836 35866 2848
rect 36265 2839 36323 2845
rect 36265 2836 36277 2839
rect 35860 2808 36277 2836
rect 35860 2796 35866 2808
rect 36265 2805 36277 2808
rect 36311 2805 36323 2839
rect 36265 2799 36323 2805
rect 1104 2746 38824 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 38824 2746
rect 1104 2672 38824 2694
rect 27709 2635 27767 2641
rect 27709 2601 27721 2635
rect 27755 2632 27767 2635
rect 27982 2632 27988 2644
rect 27755 2604 27988 2632
rect 27755 2601 27767 2604
rect 27709 2595 27767 2601
rect 27982 2592 27988 2604
rect 28040 2592 28046 2644
rect 28077 2635 28135 2641
rect 28077 2601 28089 2635
rect 28123 2632 28135 2635
rect 28166 2632 28172 2644
rect 28123 2604 28172 2632
rect 28123 2601 28135 2604
rect 28077 2595 28135 2601
rect 27341 2567 27399 2573
rect 27341 2533 27353 2567
rect 27387 2564 27399 2567
rect 28092 2564 28120 2595
rect 28166 2592 28172 2604
rect 28224 2592 28230 2644
rect 29362 2632 29368 2644
rect 29323 2604 29368 2632
rect 29362 2592 29368 2604
rect 29420 2592 29426 2644
rect 30742 2592 30748 2644
rect 30800 2632 30806 2644
rect 31113 2635 31171 2641
rect 31113 2632 31125 2635
rect 30800 2604 31125 2632
rect 30800 2592 30806 2604
rect 31113 2601 31125 2604
rect 31159 2601 31171 2635
rect 31938 2632 31944 2644
rect 31899 2604 31944 2632
rect 31113 2595 31171 2601
rect 31938 2592 31944 2604
rect 31996 2592 32002 2644
rect 32398 2632 32404 2644
rect 32359 2604 32404 2632
rect 32398 2592 32404 2604
rect 32456 2592 32462 2644
rect 33686 2592 33692 2644
rect 33744 2632 33750 2644
rect 33965 2635 34023 2641
rect 33965 2632 33977 2635
rect 33744 2604 33977 2632
rect 33744 2592 33750 2604
rect 33965 2601 33977 2604
rect 34011 2601 34023 2635
rect 34514 2632 34520 2644
rect 34475 2604 34520 2632
rect 33965 2595 34023 2601
rect 34514 2592 34520 2604
rect 34572 2592 34578 2644
rect 35250 2632 35256 2644
rect 35211 2604 35256 2632
rect 35250 2592 35256 2604
rect 35308 2592 35314 2644
rect 35986 2592 35992 2644
rect 36044 2632 36050 2644
rect 36817 2635 36875 2641
rect 36817 2632 36829 2635
rect 36044 2604 36829 2632
rect 36044 2592 36050 2604
rect 36817 2601 36829 2604
rect 36863 2601 36875 2635
rect 36817 2595 36875 2601
rect 27387 2536 28120 2564
rect 28997 2567 29055 2573
rect 27387 2533 27399 2536
rect 27341 2527 27399 2533
rect 28997 2533 29009 2567
rect 29043 2564 29055 2567
rect 29978 2567 30036 2573
rect 29978 2564 29990 2567
rect 29043 2536 29990 2564
rect 29043 2533 29055 2536
rect 28997 2527 29055 2533
rect 29978 2533 29990 2536
rect 30024 2564 30036 2567
rect 30282 2564 30288 2576
rect 30024 2536 30288 2564
rect 30024 2533 30036 2536
rect 29978 2527 30036 2533
rect 30282 2524 30288 2536
rect 30340 2524 30346 2576
rect 31956 2564 31984 2592
rect 32830 2567 32888 2573
rect 32830 2564 32842 2567
rect 31956 2536 32842 2564
rect 32830 2533 32842 2536
rect 32876 2564 32888 2567
rect 33042 2564 33048 2576
rect 32876 2536 33048 2564
rect 32876 2533 32888 2536
rect 32830 2527 32888 2533
rect 33042 2524 33048 2536
rect 33100 2524 33106 2576
rect 35268 2564 35296 2592
rect 35682 2567 35740 2573
rect 35682 2564 35694 2567
rect 35268 2536 35694 2564
rect 35682 2533 35694 2536
rect 35728 2564 35740 2567
rect 35802 2564 35808 2576
rect 35728 2536 35808 2564
rect 35728 2533 35740 2536
rect 35682 2527 35740 2533
rect 35802 2524 35808 2536
rect 35860 2524 35866 2576
rect 26697 2499 26755 2505
rect 26697 2465 26709 2499
rect 26743 2496 26755 2499
rect 28629 2499 28687 2505
rect 28629 2496 28641 2499
rect 26743 2468 28641 2496
rect 26743 2465 26755 2468
rect 26697 2459 26755 2465
rect 28629 2465 28641 2468
rect 28675 2496 28687 2499
rect 29270 2496 29276 2508
rect 28675 2468 29276 2496
rect 28675 2465 28687 2468
rect 28629 2459 28687 2465
rect 29270 2456 29276 2468
rect 29328 2496 29334 2508
rect 29733 2499 29791 2505
rect 29733 2496 29745 2499
rect 29328 2468 29745 2496
rect 29328 2456 29334 2468
rect 29733 2465 29745 2468
rect 29779 2496 29791 2499
rect 31294 2496 31300 2508
rect 29779 2468 31300 2496
rect 29779 2465 29791 2468
rect 29733 2459 29791 2465
rect 31294 2456 31300 2468
rect 31352 2456 31358 2508
rect 32585 2499 32643 2505
rect 32585 2465 32597 2499
rect 32631 2496 32643 2499
rect 33410 2496 33416 2508
rect 32631 2468 33416 2496
rect 32631 2465 32643 2468
rect 32585 2459 32643 2465
rect 33410 2456 33416 2468
rect 33468 2456 33474 2508
rect 35437 2499 35495 2505
rect 35437 2465 35449 2499
rect 35483 2496 35495 2499
rect 35526 2496 35532 2508
rect 35483 2468 35532 2496
rect 35483 2465 35495 2468
rect 35437 2459 35495 2465
rect 35526 2456 35532 2468
rect 35584 2496 35590 2508
rect 37369 2499 37427 2505
rect 37369 2496 37381 2499
rect 35584 2468 37381 2496
rect 35584 2456 35590 2468
rect 37369 2465 37381 2468
rect 37415 2465 37427 2499
rect 37369 2459 37427 2465
rect 8389 2295 8447 2301
rect 8389 2261 8401 2295
rect 8435 2292 8447 2295
rect 9950 2292 9956 2304
rect 8435 2264 9956 2292
rect 8435 2261 8447 2264
rect 8389 2255 8447 2261
rect 9950 2252 9956 2264
rect 10008 2252 10014 2304
rect 1104 2202 38824 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 34966 2202
rect 35018 2150 35030 2202
rect 35082 2150 35094 2202
rect 35146 2150 35158 2202
rect 35210 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 19606 37510 19658 37562
rect 19670 37510 19722 37562
rect 19734 37510 19786 37562
rect 19798 37510 19850 37562
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 34966 36966 35018 37018
rect 35030 36966 35082 37018
rect 35094 36966 35146 37018
rect 35158 36966 35210 37018
rect 19606 36422 19658 36474
rect 19670 36422 19722 36474
rect 19734 36422 19786 36474
rect 19798 36422 19850 36474
rect 6092 36320 6144 36372
rect 7196 36320 7248 36372
rect 5448 36227 5500 36236
rect 5448 36193 5457 36227
rect 5457 36193 5491 36227
rect 5491 36193 5500 36227
rect 5448 36184 5500 36193
rect 6644 36227 6696 36236
rect 6644 36193 6653 36227
rect 6653 36193 6687 36227
rect 6687 36193 6696 36227
rect 6644 36184 6696 36193
rect 22468 36184 22520 36236
rect 23848 36184 23900 36236
rect 14556 35980 14608 36032
rect 21456 36023 21508 36032
rect 21456 35989 21465 36023
rect 21465 35989 21499 36023
rect 21499 35989 21508 36023
rect 21456 35980 21508 35989
rect 22560 36023 22612 36032
rect 22560 35989 22569 36023
rect 22569 35989 22603 36023
rect 22603 35989 22612 36023
rect 22560 35980 22612 35989
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 34966 35878 35018 35930
rect 35030 35878 35082 35930
rect 35094 35878 35146 35930
rect 35158 35878 35210 35930
rect 4988 35776 5040 35828
rect 5264 35708 5316 35760
rect 6828 35776 6880 35828
rect 7472 35819 7524 35828
rect 7472 35785 7481 35819
rect 7481 35785 7515 35819
rect 7515 35785 7524 35819
rect 7472 35776 7524 35785
rect 8208 35776 8260 35828
rect 11888 35819 11940 35828
rect 11888 35785 11897 35819
rect 11897 35785 11931 35819
rect 11931 35785 11940 35819
rect 11888 35776 11940 35785
rect 22468 35819 22520 35828
rect 22468 35785 22477 35819
rect 22477 35785 22511 35819
rect 22511 35785 22520 35819
rect 22468 35776 22520 35785
rect 6644 35751 6696 35760
rect 6644 35717 6653 35751
rect 6653 35717 6687 35751
rect 6687 35717 6696 35751
rect 6644 35708 6696 35717
rect 15752 35708 15804 35760
rect 14924 35640 14976 35692
rect 22100 35640 22152 35692
rect 7472 35572 7524 35624
rect 11888 35572 11940 35624
rect 13544 35572 13596 35624
rect 14464 35615 14516 35624
rect 14464 35581 14473 35615
rect 14473 35581 14507 35615
rect 14507 35581 14516 35615
rect 14464 35572 14516 35581
rect 20996 35572 21048 35624
rect 21456 35572 21508 35624
rect 24768 35776 24820 35828
rect 35624 35819 35676 35828
rect 35624 35785 35633 35819
rect 35633 35785 35667 35819
rect 35667 35785 35676 35819
rect 35624 35776 35676 35785
rect 25688 35615 25740 35624
rect 25688 35581 25697 35615
rect 25697 35581 25731 35615
rect 25731 35581 25740 35615
rect 25688 35572 25740 35581
rect 35624 35572 35676 35624
rect 8576 35547 8628 35556
rect 8576 35513 8585 35547
rect 8585 35513 8619 35547
rect 8619 35513 8628 35547
rect 8576 35504 8628 35513
rect 25596 35547 25648 35556
rect 25596 35513 25605 35547
rect 25605 35513 25639 35547
rect 25639 35513 25648 35547
rect 25596 35504 25648 35513
rect 4988 35479 5040 35488
rect 4988 35445 4997 35479
rect 4997 35445 5031 35479
rect 5031 35445 5040 35479
rect 4988 35436 5040 35445
rect 5540 35479 5592 35488
rect 5540 35445 5549 35479
rect 5549 35445 5583 35479
rect 5583 35445 5592 35479
rect 5540 35436 5592 35445
rect 7472 35436 7524 35488
rect 11060 35436 11112 35488
rect 14556 35479 14608 35488
rect 14556 35445 14565 35479
rect 14565 35445 14599 35479
rect 14599 35445 14608 35479
rect 14556 35436 14608 35445
rect 16488 35436 16540 35488
rect 21180 35479 21232 35488
rect 21180 35445 21189 35479
rect 21189 35445 21223 35479
rect 21223 35445 21232 35479
rect 21180 35436 21232 35445
rect 21364 35479 21416 35488
rect 21364 35445 21373 35479
rect 21373 35445 21407 35479
rect 21407 35445 21416 35479
rect 21364 35436 21416 35445
rect 26976 35436 27028 35488
rect 19606 35334 19658 35386
rect 19670 35334 19722 35386
rect 19734 35334 19786 35386
rect 19798 35334 19850 35386
rect 1676 35232 1728 35284
rect 10876 35275 10928 35284
rect 10876 35241 10885 35275
rect 10885 35241 10919 35275
rect 10919 35241 10928 35275
rect 10876 35232 10928 35241
rect 15752 35275 15804 35284
rect 15752 35241 15761 35275
rect 15761 35241 15795 35275
rect 15795 35241 15804 35275
rect 15752 35232 15804 35241
rect 35532 35275 35584 35284
rect 35532 35241 35541 35275
rect 35541 35241 35575 35275
rect 35575 35241 35584 35275
rect 35532 35232 35584 35241
rect 8852 35164 8904 35216
rect 13728 35164 13780 35216
rect 21088 35164 21140 35216
rect 1400 35139 1452 35148
rect 1400 35105 1409 35139
rect 1409 35105 1443 35139
rect 1443 35105 1452 35139
rect 1400 35096 1452 35105
rect 4988 35139 5040 35148
rect 4988 35105 4997 35139
rect 4997 35105 5031 35139
rect 5031 35105 5040 35139
rect 4988 35096 5040 35105
rect 6828 35139 6880 35148
rect 6828 35105 6837 35139
rect 6837 35105 6871 35139
rect 6871 35105 6880 35139
rect 6828 35096 6880 35105
rect 8300 35139 8352 35148
rect 8300 35105 8309 35139
rect 8309 35105 8343 35139
rect 8343 35105 8352 35139
rect 8300 35096 8352 35105
rect 11244 35139 11296 35148
rect 11244 35105 11253 35139
rect 11253 35105 11287 35139
rect 11287 35105 11296 35139
rect 11244 35096 11296 35105
rect 13544 35139 13596 35148
rect 13544 35105 13553 35139
rect 13553 35105 13587 35139
rect 13587 35105 13596 35139
rect 13544 35096 13596 35105
rect 14832 35096 14884 35148
rect 16948 35096 17000 35148
rect 18328 35096 18380 35148
rect 21916 35096 21968 35148
rect 22928 35164 22980 35216
rect 22468 35096 22520 35148
rect 28080 35096 28132 35148
rect 35348 35139 35400 35148
rect 35348 35105 35357 35139
rect 35357 35105 35391 35139
rect 35391 35105 35400 35139
rect 35348 35096 35400 35105
rect 5080 35071 5132 35080
rect 5080 35037 5089 35071
rect 5089 35037 5123 35071
rect 5123 35037 5132 35071
rect 5080 35028 5132 35037
rect 5264 35071 5316 35080
rect 5264 35037 5273 35071
rect 5273 35037 5307 35071
rect 5307 35037 5316 35071
rect 5264 35028 5316 35037
rect 10048 35028 10100 35080
rect 11336 35071 11388 35080
rect 11336 35037 11345 35071
rect 11345 35037 11379 35071
rect 11379 35037 11388 35071
rect 11336 35028 11388 35037
rect 12532 35071 12584 35080
rect 12532 35037 12541 35071
rect 12541 35037 12575 35071
rect 12575 35037 12584 35071
rect 12532 35028 12584 35037
rect 14372 35028 14424 35080
rect 15200 35028 15252 35080
rect 15476 35028 15528 35080
rect 17868 35028 17920 35080
rect 4712 34960 4764 35012
rect 6920 34960 6972 35012
rect 13636 34960 13688 35012
rect 5448 34892 5500 34944
rect 7104 34892 7156 34944
rect 8484 34935 8536 34944
rect 8484 34901 8493 34935
rect 8493 34901 8527 34935
rect 8527 34901 8536 34935
rect 8484 34892 8536 34901
rect 9864 34892 9916 34944
rect 12072 34935 12124 34944
rect 12072 34901 12081 34935
rect 12081 34901 12115 34935
rect 12115 34901 12124 34935
rect 12072 34892 12124 34901
rect 14648 34935 14700 34944
rect 14648 34901 14657 34935
rect 14657 34901 14691 34935
rect 14691 34901 14700 34935
rect 14648 34892 14700 34901
rect 15752 34892 15804 34944
rect 17408 34892 17460 34944
rect 18512 34935 18564 34944
rect 18512 34901 18521 34935
rect 18521 34901 18555 34935
rect 18555 34901 18564 34935
rect 18512 34892 18564 34901
rect 21456 34935 21508 34944
rect 21456 34901 21465 34935
rect 21465 34901 21499 34935
rect 21499 34901 21508 34935
rect 21456 34892 21508 34901
rect 21916 34935 21968 34944
rect 21916 34901 21925 34935
rect 21925 34901 21959 34935
rect 21959 34901 21968 34935
rect 21916 34892 21968 34901
rect 24032 34892 24084 34944
rect 24216 34892 24268 34944
rect 25688 34892 25740 34944
rect 26700 34892 26752 34944
rect 28356 34892 28408 34944
rect 28816 34935 28868 34944
rect 28816 34901 28825 34935
rect 28825 34901 28859 34935
rect 28859 34901 28868 34935
rect 28816 34892 28868 34901
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 34966 34790 35018 34842
rect 35030 34790 35082 34842
rect 35094 34790 35146 34842
rect 35158 34790 35210 34842
rect 572 34688 624 34740
rect 2044 34731 2096 34740
rect 2044 34697 2053 34731
rect 2053 34697 2087 34731
rect 2087 34697 2096 34731
rect 2044 34688 2096 34697
rect 3148 34731 3200 34740
rect 3148 34697 3157 34731
rect 3157 34697 3191 34731
rect 3191 34697 3200 34731
rect 3148 34688 3200 34697
rect 5080 34688 5132 34740
rect 6828 34688 6880 34740
rect 8852 34731 8904 34740
rect 8852 34697 8861 34731
rect 8861 34697 8895 34731
rect 8895 34697 8904 34731
rect 8852 34688 8904 34697
rect 11244 34688 11296 34740
rect 13544 34688 13596 34740
rect 16948 34731 17000 34740
rect 16948 34697 16957 34731
rect 16957 34697 16991 34731
rect 16991 34697 17000 34731
rect 16948 34688 17000 34697
rect 17868 34731 17920 34740
rect 17868 34697 17877 34731
rect 17877 34697 17911 34731
rect 17911 34697 17920 34731
rect 17868 34688 17920 34697
rect 18052 34731 18104 34740
rect 18052 34697 18061 34731
rect 18061 34697 18095 34731
rect 18095 34697 18104 34731
rect 18052 34688 18104 34697
rect 20628 34731 20680 34740
rect 20628 34697 20637 34731
rect 20637 34697 20671 34731
rect 20671 34697 20680 34731
rect 20628 34688 20680 34697
rect 20996 34731 21048 34740
rect 20996 34697 21005 34731
rect 21005 34697 21039 34731
rect 21039 34697 21048 34731
rect 20996 34688 21048 34697
rect 22468 34731 22520 34740
rect 22468 34697 22477 34731
rect 22477 34697 22511 34731
rect 22511 34697 22520 34731
rect 22468 34688 22520 34697
rect 23388 34688 23440 34740
rect 25596 34731 25648 34740
rect 25596 34697 25605 34731
rect 25605 34697 25639 34731
rect 25639 34697 25648 34731
rect 25596 34688 25648 34697
rect 28080 34731 28132 34740
rect 28080 34697 28089 34731
rect 28089 34697 28123 34731
rect 28123 34697 28132 34731
rect 28080 34688 28132 34697
rect 35808 34688 35860 34740
rect 36728 34731 36780 34740
rect 36728 34697 36737 34731
rect 36737 34697 36771 34731
rect 36771 34697 36780 34731
rect 36728 34688 36780 34697
rect 2688 34663 2740 34672
rect 2688 34629 2697 34663
rect 2697 34629 2731 34663
rect 2731 34629 2740 34663
rect 2688 34620 2740 34629
rect 8300 34620 8352 34672
rect 5080 34552 5132 34604
rect 2044 34484 2096 34536
rect 3148 34484 3200 34536
rect 4620 34484 4672 34536
rect 5632 34484 5684 34536
rect 6920 34484 6972 34536
rect 8208 34484 8260 34536
rect 12072 34552 12124 34604
rect 14648 34552 14700 34604
rect 4712 34348 4764 34400
rect 6276 34391 6328 34400
rect 6276 34357 6285 34391
rect 6285 34357 6319 34391
rect 6319 34357 6328 34391
rect 6276 34348 6328 34357
rect 9864 34484 9916 34536
rect 14096 34484 14148 34536
rect 14832 34484 14884 34536
rect 17868 34552 17920 34604
rect 18512 34595 18564 34604
rect 18512 34561 18521 34595
rect 18521 34561 18555 34595
rect 18555 34561 18564 34595
rect 18512 34552 18564 34561
rect 19248 34552 19300 34604
rect 15200 34527 15252 34536
rect 10140 34416 10192 34468
rect 12532 34416 12584 34468
rect 13544 34416 13596 34468
rect 15200 34493 15234 34527
rect 15234 34493 15252 34527
rect 15200 34484 15252 34493
rect 17960 34484 18012 34536
rect 20628 34484 20680 34536
rect 21088 34527 21140 34536
rect 21088 34493 21097 34527
rect 21097 34493 21131 34527
rect 21131 34493 21140 34527
rect 21088 34484 21140 34493
rect 22928 34552 22980 34604
rect 24216 34595 24268 34604
rect 24216 34561 24225 34595
rect 24225 34561 24259 34595
rect 24259 34561 24268 34595
rect 24216 34552 24268 34561
rect 26700 34595 26752 34604
rect 26700 34561 26709 34595
rect 26709 34561 26743 34595
rect 26743 34561 26752 34595
rect 26700 34552 26752 34561
rect 26976 34527 27028 34536
rect 15292 34416 15344 34468
rect 22192 34416 22244 34468
rect 26608 34459 26660 34468
rect 26608 34425 26617 34459
rect 26617 34425 26651 34459
rect 26651 34425 26660 34459
rect 26976 34493 27010 34527
rect 27010 34493 27028 34527
rect 26976 34484 27028 34493
rect 35256 34527 35308 34536
rect 35256 34493 35265 34527
rect 35265 34493 35299 34527
rect 35299 34493 35308 34527
rect 35256 34484 35308 34493
rect 37096 34527 37148 34536
rect 37096 34493 37105 34527
rect 37105 34493 37139 34527
rect 37139 34493 37148 34527
rect 37096 34484 37148 34493
rect 26608 34416 26660 34425
rect 9772 34348 9824 34400
rect 11152 34391 11204 34400
rect 11152 34357 11161 34391
rect 11161 34357 11195 34391
rect 11195 34357 11204 34391
rect 11152 34348 11204 34357
rect 13268 34348 13320 34400
rect 14924 34348 14976 34400
rect 20168 34391 20220 34400
rect 20168 34357 20177 34391
rect 20177 34357 20211 34391
rect 20211 34357 20220 34391
rect 20168 34348 20220 34357
rect 24032 34391 24084 34400
rect 24032 34357 24041 34391
rect 24041 34357 24075 34391
rect 24075 34357 24084 34391
rect 24032 34348 24084 34357
rect 28356 34348 28408 34400
rect 30104 34348 30156 34400
rect 35348 34348 35400 34400
rect 19606 34246 19658 34298
rect 19670 34246 19722 34298
rect 19734 34246 19786 34298
rect 19798 34246 19850 34298
rect 1400 34144 1452 34196
rect 4160 34144 4212 34196
rect 6276 34144 6328 34196
rect 7196 34187 7248 34196
rect 7196 34153 7205 34187
rect 7205 34153 7239 34187
rect 7239 34153 7248 34187
rect 7196 34144 7248 34153
rect 4988 34076 5040 34128
rect 6828 34076 6880 34128
rect 4068 34051 4120 34060
rect 4068 34017 4077 34051
rect 4077 34017 4111 34051
rect 4111 34017 4120 34051
rect 4068 34008 4120 34017
rect 5540 34051 5592 34060
rect 5540 34017 5574 34051
rect 5574 34017 5592 34051
rect 5540 34008 5592 34017
rect 7932 34008 7984 34060
rect 8668 34008 8720 34060
rect 3976 33940 4028 33992
rect 9036 33940 9088 33992
rect 11336 34144 11388 34196
rect 13544 34187 13596 34196
rect 13544 34153 13553 34187
rect 13553 34153 13587 34187
rect 13587 34153 13596 34187
rect 13544 34144 13596 34153
rect 13820 34144 13872 34196
rect 16488 34144 16540 34196
rect 22192 34144 22244 34196
rect 22928 34187 22980 34196
rect 22928 34153 22937 34187
rect 22937 34153 22971 34187
rect 22971 34153 22980 34187
rect 22928 34144 22980 34153
rect 23480 34144 23532 34196
rect 28080 34144 28132 34196
rect 35624 34187 35676 34196
rect 35624 34153 35633 34187
rect 35633 34153 35667 34187
rect 35667 34153 35676 34187
rect 35624 34144 35676 34153
rect 9864 34076 9916 34128
rect 12164 34076 12216 34128
rect 9772 34008 9824 34060
rect 10692 34008 10744 34060
rect 14464 34008 14516 34060
rect 7472 33872 7524 33924
rect 5264 33804 5316 33856
rect 8024 33847 8076 33856
rect 8024 33813 8033 33847
rect 8033 33813 8067 33847
rect 8067 33813 8076 33847
rect 8024 33804 8076 33813
rect 8300 33804 8352 33856
rect 11796 33940 11848 33992
rect 15200 33940 15252 33992
rect 17776 34076 17828 34128
rect 18052 34008 18104 34060
rect 20720 34008 20772 34060
rect 21088 34076 21140 34128
rect 28816 34076 28868 34128
rect 21180 34051 21232 34060
rect 21180 34017 21214 34051
rect 21214 34017 21232 34051
rect 21180 34008 21232 34017
rect 23112 34008 23164 34060
rect 24032 34008 24084 34060
rect 25320 34051 25372 34060
rect 25320 34017 25329 34051
rect 25329 34017 25363 34051
rect 25363 34017 25372 34051
rect 25320 34008 25372 34017
rect 25964 34008 26016 34060
rect 28448 34008 28500 34060
rect 35900 34008 35952 34060
rect 22100 33940 22152 33992
rect 26424 33940 26476 33992
rect 15844 33915 15896 33924
rect 15844 33881 15853 33915
rect 15853 33881 15887 33915
rect 15887 33881 15896 33915
rect 15844 33872 15896 33881
rect 25780 33872 25832 33924
rect 14464 33847 14516 33856
rect 14464 33813 14473 33847
rect 14473 33813 14507 33847
rect 14507 33813 14516 33847
rect 14464 33804 14516 33813
rect 14832 33804 14884 33856
rect 15476 33847 15528 33856
rect 15476 33813 15485 33847
rect 15485 33813 15519 33847
rect 15519 33813 15528 33847
rect 15476 33804 15528 33813
rect 18788 33847 18840 33856
rect 18788 33813 18797 33847
rect 18797 33813 18831 33847
rect 18831 33813 18840 33847
rect 18788 33804 18840 33813
rect 23388 33847 23440 33856
rect 23388 33813 23397 33847
rect 23397 33813 23431 33847
rect 23431 33813 23440 33847
rect 23388 33804 23440 33813
rect 24400 33847 24452 33856
rect 24400 33813 24409 33847
rect 24409 33813 24443 33847
rect 24443 33813 24452 33847
rect 24400 33804 24452 33813
rect 25504 33847 25556 33856
rect 25504 33813 25513 33847
rect 25513 33813 25547 33847
rect 25547 33813 25556 33847
rect 25504 33804 25556 33813
rect 29092 33804 29144 33856
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 34966 33702 35018 33754
rect 35030 33702 35082 33754
rect 35094 33702 35146 33754
rect 35158 33702 35210 33754
rect 4068 33643 4120 33652
rect 4068 33609 4077 33643
rect 4077 33609 4111 33643
rect 4111 33609 4120 33643
rect 4068 33600 4120 33609
rect 5540 33600 5592 33652
rect 6828 33643 6880 33652
rect 4068 33464 4120 33516
rect 5540 33396 5592 33448
rect 4528 33371 4580 33380
rect 4528 33337 4562 33371
rect 4562 33337 4580 33371
rect 4528 33328 4580 33337
rect 4712 33328 4764 33380
rect 6828 33609 6837 33643
rect 6837 33609 6871 33643
rect 6871 33609 6880 33643
rect 6828 33600 6880 33609
rect 8300 33600 8352 33652
rect 10140 33643 10192 33652
rect 7472 33507 7524 33516
rect 7472 33473 7481 33507
rect 7481 33473 7515 33507
rect 7515 33473 7524 33507
rect 7472 33464 7524 33473
rect 10140 33609 10149 33643
rect 10149 33609 10183 33643
rect 10183 33609 10192 33643
rect 10140 33600 10192 33609
rect 10692 33643 10744 33652
rect 10692 33609 10701 33643
rect 10701 33609 10735 33643
rect 10735 33609 10744 33643
rect 10692 33600 10744 33609
rect 11152 33600 11204 33652
rect 12164 33643 12216 33652
rect 12164 33609 12173 33643
rect 12173 33609 12207 33643
rect 12207 33609 12216 33643
rect 12164 33600 12216 33609
rect 14372 33643 14424 33652
rect 14372 33609 14381 33643
rect 14381 33609 14415 33643
rect 14415 33609 14424 33643
rect 14372 33600 14424 33609
rect 14924 33643 14976 33652
rect 14924 33609 14933 33643
rect 14933 33609 14967 33643
rect 14967 33609 14976 33643
rect 14924 33600 14976 33609
rect 16488 33600 16540 33652
rect 19340 33600 19392 33652
rect 21364 33600 21416 33652
rect 23112 33643 23164 33652
rect 23112 33609 23121 33643
rect 23121 33609 23155 33643
rect 23155 33609 23164 33643
rect 23112 33600 23164 33609
rect 23480 33643 23532 33652
rect 23480 33609 23489 33643
rect 23489 33609 23523 33643
rect 23523 33609 23532 33643
rect 23480 33600 23532 33609
rect 23664 33643 23716 33652
rect 23664 33609 23673 33643
rect 23673 33609 23707 33643
rect 23707 33609 23716 33643
rect 23664 33600 23716 33609
rect 25596 33600 25648 33652
rect 9864 33532 9916 33584
rect 11796 33575 11848 33584
rect 11796 33541 11805 33575
rect 11805 33541 11839 33575
rect 11839 33541 11848 33575
rect 11796 33532 11848 33541
rect 8576 33464 8628 33516
rect 11244 33507 11296 33516
rect 11244 33473 11253 33507
rect 11253 33473 11287 33507
rect 11287 33473 11296 33507
rect 11244 33464 11296 33473
rect 21916 33532 21968 33584
rect 26240 33532 26292 33584
rect 7196 33439 7248 33448
rect 7196 33405 7205 33439
rect 7205 33405 7239 33439
rect 7239 33405 7248 33439
rect 7196 33396 7248 33405
rect 8852 33396 8904 33448
rect 9036 33439 9088 33448
rect 9036 33405 9070 33439
rect 9070 33405 9088 33439
rect 9036 33396 9088 33405
rect 12992 33439 13044 33448
rect 12992 33405 13001 33439
rect 13001 33405 13035 33439
rect 13035 33405 13044 33439
rect 12992 33396 13044 33405
rect 13268 33439 13320 33448
rect 13268 33405 13302 33439
rect 13302 33405 13320 33439
rect 13268 33396 13320 33405
rect 15292 33396 15344 33448
rect 20720 33507 20772 33516
rect 20720 33473 20729 33507
rect 20729 33473 20763 33507
rect 20763 33473 20772 33507
rect 20720 33464 20772 33473
rect 22100 33464 22152 33516
rect 24124 33507 24176 33516
rect 24124 33473 24133 33507
rect 24133 33473 24167 33507
rect 24167 33473 24176 33507
rect 24124 33464 24176 33473
rect 24400 33464 24452 33516
rect 26424 33507 26476 33516
rect 26424 33473 26433 33507
rect 26433 33473 26467 33507
rect 26467 33473 26476 33507
rect 26424 33464 26476 33473
rect 27620 33464 27672 33516
rect 18052 33439 18104 33448
rect 18052 33405 18061 33439
rect 18061 33405 18095 33439
rect 18095 33405 18104 33439
rect 18052 33396 18104 33405
rect 17960 33328 18012 33380
rect 18788 33396 18840 33448
rect 23388 33396 23440 33448
rect 24308 33396 24360 33448
rect 21732 33328 21784 33380
rect 23572 33328 23624 33380
rect 25872 33396 25924 33448
rect 26608 33396 26660 33448
rect 28080 33396 28132 33448
rect 24768 33328 24820 33380
rect 28816 33600 28868 33652
rect 35716 33600 35768 33652
rect 7932 33260 7984 33312
rect 15476 33260 15528 33312
rect 17776 33303 17828 33312
rect 17776 33269 17785 33303
rect 17785 33269 17819 33303
rect 17819 33269 17828 33303
rect 17776 33260 17828 33269
rect 25320 33260 25372 33312
rect 26240 33260 26292 33312
rect 26884 33260 26936 33312
rect 28356 33260 28408 33312
rect 35348 33303 35400 33312
rect 35348 33269 35357 33303
rect 35357 33269 35391 33303
rect 35391 33269 35400 33303
rect 35348 33260 35400 33269
rect 35900 33260 35952 33312
rect 19606 33158 19658 33210
rect 19670 33158 19722 33210
rect 19734 33158 19786 33210
rect 19798 33158 19850 33210
rect 4528 33056 4580 33108
rect 5540 33056 5592 33108
rect 8668 33099 8720 33108
rect 8668 33065 8677 33099
rect 8677 33065 8711 33099
rect 8711 33065 8720 33099
rect 8668 33056 8720 33065
rect 9036 33099 9088 33108
rect 9036 33065 9045 33099
rect 9045 33065 9079 33099
rect 9079 33065 9088 33099
rect 9036 33056 9088 33065
rect 10140 33099 10192 33108
rect 10140 33065 10149 33099
rect 10149 33065 10183 33099
rect 10183 33065 10192 33099
rect 10140 33056 10192 33065
rect 11336 33056 11388 33108
rect 11612 33099 11664 33108
rect 11612 33065 11621 33099
rect 11621 33065 11655 33099
rect 11655 33065 11664 33099
rect 11612 33056 11664 33065
rect 13268 33056 13320 33108
rect 13360 33099 13412 33108
rect 13360 33065 13369 33099
rect 13369 33065 13403 33099
rect 13403 33065 13412 33099
rect 15108 33099 15160 33108
rect 13360 33056 13412 33065
rect 15108 33065 15117 33099
rect 15117 33065 15151 33099
rect 15151 33065 15160 33099
rect 15108 33056 15160 33065
rect 17960 33056 18012 33108
rect 19340 33099 19392 33108
rect 19340 33065 19349 33099
rect 19349 33065 19383 33099
rect 19383 33065 19392 33099
rect 19340 33056 19392 33065
rect 20720 33099 20772 33108
rect 20720 33065 20729 33099
rect 20729 33065 20763 33099
rect 20763 33065 20772 33099
rect 20720 33056 20772 33065
rect 21180 33099 21232 33108
rect 21180 33065 21189 33099
rect 21189 33065 21223 33099
rect 21223 33065 21232 33099
rect 21180 33056 21232 33065
rect 23296 33099 23348 33108
rect 23296 33065 23305 33099
rect 23305 33065 23339 33099
rect 23339 33065 23348 33099
rect 23296 33056 23348 33065
rect 23940 33099 23992 33108
rect 23940 33065 23949 33099
rect 23949 33065 23983 33099
rect 23983 33065 23992 33099
rect 23940 33056 23992 33065
rect 24308 33099 24360 33108
rect 24308 33065 24317 33099
rect 24317 33065 24351 33099
rect 24351 33065 24360 33099
rect 24308 33056 24360 33065
rect 25504 33056 25556 33108
rect 25872 33099 25924 33108
rect 25872 33065 25881 33099
rect 25881 33065 25915 33099
rect 25915 33065 25924 33099
rect 25872 33056 25924 33065
rect 26240 33056 26292 33108
rect 26884 33099 26936 33108
rect 26884 33065 26893 33099
rect 26893 33065 26927 33099
rect 26927 33065 26936 33099
rect 26884 33056 26936 33065
rect 27620 33099 27672 33108
rect 27620 33065 27629 33099
rect 27629 33065 27663 33099
rect 27663 33065 27672 33099
rect 27620 33056 27672 33065
rect 28172 33056 28224 33108
rect 4620 32988 4672 33040
rect 8852 32988 8904 33040
rect 9220 32988 9272 33040
rect 10048 33031 10100 33040
rect 10048 32997 10057 33031
rect 10057 32997 10091 33031
rect 10091 32997 10100 33031
rect 10048 32988 10100 32997
rect 21732 33031 21784 33040
rect 4068 32963 4120 32972
rect 4068 32929 4077 32963
rect 4077 32929 4111 32963
rect 4111 32929 4120 32963
rect 4068 32920 4120 32929
rect 6920 32963 6972 32972
rect 6920 32929 6929 32963
rect 6929 32929 6963 32963
rect 6963 32929 6972 32963
rect 6920 32920 6972 32929
rect 8484 32920 8536 32972
rect 13268 32920 13320 32972
rect 13820 32963 13872 32972
rect 13820 32929 13829 32963
rect 13829 32929 13863 32963
rect 13863 32929 13872 32963
rect 13820 32920 13872 32929
rect 21732 32997 21741 33031
rect 21741 32997 21775 33031
rect 21775 32997 21784 33031
rect 21732 32988 21784 32997
rect 22560 32988 22612 33040
rect 23572 32988 23624 33040
rect 25228 33031 25280 33040
rect 25228 32997 25237 33031
rect 25237 32997 25271 33031
rect 25271 32997 25280 33031
rect 25228 32988 25280 32997
rect 25780 32988 25832 33040
rect 26332 32988 26384 33040
rect 27068 32988 27120 33040
rect 7012 32895 7064 32904
rect 7012 32861 7021 32895
rect 7021 32861 7055 32895
rect 7055 32861 7064 32895
rect 7012 32852 7064 32861
rect 7104 32895 7156 32904
rect 7104 32861 7113 32895
rect 7113 32861 7147 32895
rect 7147 32861 7156 32895
rect 7104 32852 7156 32861
rect 10232 32895 10284 32904
rect 10232 32861 10241 32895
rect 10241 32861 10275 32895
rect 10275 32861 10284 32895
rect 10232 32852 10284 32861
rect 11336 32852 11388 32904
rect 12164 32852 12216 32904
rect 13912 32895 13964 32904
rect 13912 32861 13921 32895
rect 13921 32861 13955 32895
rect 13955 32861 13964 32895
rect 13912 32852 13964 32861
rect 15844 32920 15896 32972
rect 17776 32920 17828 32972
rect 21824 32963 21876 32972
rect 21824 32929 21833 32963
rect 21833 32929 21867 32963
rect 21867 32929 21876 32963
rect 21824 32920 21876 32929
rect 14740 32852 14792 32904
rect 15752 32895 15804 32904
rect 15752 32861 15764 32895
rect 15764 32861 15798 32895
rect 15798 32861 15804 32895
rect 16028 32895 16080 32904
rect 15752 32852 15804 32861
rect 16028 32861 16037 32895
rect 16037 32861 16071 32895
rect 16071 32861 16080 32895
rect 16028 32852 16080 32861
rect 21916 32895 21968 32904
rect 3148 32759 3200 32768
rect 3148 32725 3157 32759
rect 3157 32725 3191 32759
rect 3191 32725 3200 32759
rect 3148 32716 3200 32725
rect 8116 32716 8168 32768
rect 8300 32759 8352 32768
rect 8300 32725 8309 32759
rect 8309 32725 8343 32759
rect 8343 32725 8352 32759
rect 8300 32716 8352 32725
rect 11612 32716 11664 32768
rect 12808 32759 12860 32768
rect 12808 32725 12817 32759
rect 12817 32725 12851 32759
rect 12851 32725 12860 32759
rect 12808 32716 12860 32725
rect 13728 32716 13780 32768
rect 13820 32716 13872 32768
rect 17132 32759 17184 32768
rect 17132 32725 17141 32759
rect 17141 32725 17175 32759
rect 17175 32725 17184 32759
rect 17132 32716 17184 32725
rect 17500 32759 17552 32768
rect 17500 32725 17509 32759
rect 17509 32725 17543 32759
rect 17543 32725 17552 32759
rect 21916 32861 21925 32895
rect 21925 32861 21959 32895
rect 21959 32861 21968 32895
rect 21916 32852 21968 32861
rect 23388 32895 23440 32904
rect 23388 32861 23397 32895
rect 23397 32861 23431 32895
rect 23431 32861 23440 32895
rect 23388 32852 23440 32861
rect 24676 32963 24728 32972
rect 24676 32929 24685 32963
rect 24685 32929 24719 32963
rect 24719 32929 24728 32963
rect 28632 32963 28684 32972
rect 24676 32920 24728 32929
rect 28632 32929 28666 32963
rect 28666 32929 28684 32963
rect 28632 32920 28684 32929
rect 26608 32852 26660 32904
rect 28356 32895 28408 32904
rect 28356 32861 28365 32895
rect 28365 32861 28399 32895
rect 28399 32861 28408 32895
rect 28356 32852 28408 32861
rect 17500 32716 17552 32725
rect 18144 32716 18196 32768
rect 23480 32716 23532 32768
rect 24860 32759 24912 32768
rect 24860 32725 24869 32759
rect 24869 32725 24903 32759
rect 24903 32725 24912 32759
rect 24860 32716 24912 32725
rect 26332 32759 26384 32768
rect 26332 32725 26341 32759
rect 26341 32725 26375 32759
rect 26375 32725 26384 32759
rect 26332 32716 26384 32725
rect 29000 32716 29052 32768
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 34966 32614 35018 32666
rect 35030 32614 35082 32666
rect 35094 32614 35146 32666
rect 35158 32614 35210 32666
rect 4620 32512 4672 32564
rect 5540 32555 5592 32564
rect 5540 32521 5549 32555
rect 5549 32521 5583 32555
rect 5583 32521 5592 32555
rect 5540 32512 5592 32521
rect 6460 32512 6512 32564
rect 7012 32512 7064 32564
rect 10048 32512 10100 32564
rect 10232 32555 10284 32564
rect 10232 32521 10241 32555
rect 10241 32521 10275 32555
rect 10275 32521 10284 32555
rect 10232 32512 10284 32521
rect 11612 32555 11664 32564
rect 11612 32521 11621 32555
rect 11621 32521 11655 32555
rect 11655 32521 11664 32555
rect 11612 32512 11664 32521
rect 12164 32512 12216 32564
rect 13176 32555 13228 32564
rect 13176 32521 13185 32555
rect 13185 32521 13219 32555
rect 13219 32521 13228 32555
rect 13176 32512 13228 32521
rect 13912 32512 13964 32564
rect 14648 32512 14700 32564
rect 6920 32444 6972 32496
rect 9496 32487 9548 32496
rect 9496 32453 9505 32487
rect 9505 32453 9539 32487
rect 9539 32453 9548 32487
rect 9496 32444 9548 32453
rect 13820 32487 13872 32496
rect 13820 32453 13829 32487
rect 13829 32453 13863 32487
rect 13863 32453 13872 32487
rect 13820 32444 13872 32453
rect 17500 32512 17552 32564
rect 18052 32512 18104 32564
rect 19064 32512 19116 32564
rect 20720 32512 20772 32564
rect 21732 32512 21784 32564
rect 3148 32419 3200 32428
rect 3148 32385 3157 32419
rect 3157 32385 3191 32419
rect 3191 32385 3200 32419
rect 3148 32376 3200 32385
rect 8300 32419 8352 32428
rect 8300 32385 8309 32419
rect 8309 32385 8343 32419
rect 8343 32385 8352 32419
rect 8300 32376 8352 32385
rect 15752 32376 15804 32428
rect 24216 32512 24268 32564
rect 25504 32512 25556 32564
rect 25964 32512 26016 32564
rect 27068 32555 27120 32564
rect 27068 32521 27077 32555
rect 27077 32521 27111 32555
rect 27111 32521 27120 32555
rect 27068 32512 27120 32521
rect 28632 32512 28684 32564
rect 25228 32487 25280 32496
rect 25228 32453 25237 32487
rect 25237 32453 25271 32487
rect 25271 32453 25280 32487
rect 25228 32444 25280 32453
rect 24124 32376 24176 32428
rect 24676 32376 24728 32428
rect 26148 32376 26200 32428
rect 29092 32487 29144 32496
rect 26608 32419 26660 32428
rect 26608 32385 26617 32419
rect 26617 32385 26651 32419
rect 26651 32385 26660 32419
rect 29092 32453 29101 32487
rect 29101 32453 29135 32487
rect 29135 32453 29144 32487
rect 29092 32444 29144 32453
rect 26608 32376 26660 32385
rect 28172 32419 28224 32428
rect 28172 32385 28181 32419
rect 28181 32385 28215 32419
rect 28215 32385 28224 32419
rect 28172 32376 28224 32385
rect 5540 32308 5592 32360
rect 8116 32351 8168 32360
rect 8116 32317 8125 32351
rect 8125 32317 8159 32351
rect 8159 32317 8168 32351
rect 8116 32308 8168 32317
rect 10876 32351 10928 32360
rect 10876 32317 10885 32351
rect 10885 32317 10919 32351
rect 10919 32317 10928 32351
rect 10876 32308 10928 32317
rect 11336 32351 11388 32360
rect 11336 32317 11345 32351
rect 11345 32317 11379 32351
rect 11379 32317 11388 32351
rect 11336 32308 11388 32317
rect 14740 32308 14792 32360
rect 15108 32351 15160 32360
rect 15108 32317 15117 32351
rect 15117 32317 15151 32351
rect 15151 32317 15160 32351
rect 15108 32308 15160 32317
rect 17040 32308 17092 32360
rect 18604 32308 18656 32360
rect 19248 32308 19300 32360
rect 21824 32308 21876 32360
rect 23940 32308 23992 32360
rect 26884 32308 26936 32360
rect 27712 32308 27764 32360
rect 28632 32308 28684 32360
rect 29276 32351 29328 32360
rect 29276 32317 29285 32351
rect 29285 32317 29319 32351
rect 29319 32317 29328 32351
rect 29276 32308 29328 32317
rect 3608 32240 3660 32292
rect 2044 32215 2096 32224
rect 2044 32181 2053 32215
rect 2053 32181 2087 32215
rect 2087 32181 2096 32215
rect 2044 32172 2096 32181
rect 2596 32172 2648 32224
rect 5816 32172 5868 32224
rect 8024 32240 8076 32292
rect 13268 32240 13320 32292
rect 16672 32240 16724 32292
rect 17776 32283 17828 32292
rect 17776 32249 17785 32283
rect 17785 32249 17819 32283
rect 17819 32249 17828 32283
rect 17776 32240 17828 32249
rect 23572 32240 23624 32292
rect 26332 32240 26384 32292
rect 27528 32240 27580 32292
rect 7748 32215 7800 32224
rect 7748 32181 7757 32215
rect 7757 32181 7791 32215
rect 7791 32181 7800 32215
rect 7748 32172 7800 32181
rect 9864 32172 9916 32224
rect 15844 32172 15896 32224
rect 16948 32215 17000 32224
rect 16948 32181 16957 32215
rect 16957 32181 16991 32215
rect 16991 32181 17000 32215
rect 16948 32172 17000 32181
rect 19340 32172 19392 32224
rect 19606 32070 19658 32122
rect 19670 32070 19722 32122
rect 19734 32070 19786 32122
rect 19798 32070 19850 32122
rect 2872 31968 2924 32020
rect 2780 31900 2832 31952
rect 3148 31968 3200 32020
rect 3608 31968 3660 32020
rect 4988 31968 5040 32020
rect 5172 31968 5224 32020
rect 5816 32011 5868 32020
rect 5816 31977 5825 32011
rect 5825 31977 5859 32011
rect 5859 31977 5868 32011
rect 5816 31968 5868 31977
rect 6552 31968 6604 32020
rect 7104 31968 7156 32020
rect 8484 32011 8536 32020
rect 4620 31900 4672 31952
rect 8484 31977 8493 32011
rect 8493 31977 8527 32011
rect 8527 31977 8536 32011
rect 8484 31968 8536 31977
rect 9588 31968 9640 32020
rect 10140 31968 10192 32020
rect 10876 31968 10928 32020
rect 14096 32011 14148 32020
rect 14096 31977 14105 32011
rect 14105 31977 14139 32011
rect 14139 31977 14148 32011
rect 14096 31968 14148 31977
rect 15108 31968 15160 32020
rect 16028 31968 16080 32020
rect 17500 32011 17552 32020
rect 17500 31977 17509 32011
rect 17509 31977 17543 32011
rect 17543 31977 17552 32011
rect 17500 31968 17552 31977
rect 17868 31968 17920 32020
rect 18604 32011 18656 32020
rect 18604 31977 18613 32011
rect 18613 31977 18647 32011
rect 18647 31977 18656 32011
rect 18604 31968 18656 31977
rect 19064 32011 19116 32020
rect 19064 31977 19073 32011
rect 19073 31977 19107 32011
rect 19107 31977 19116 32011
rect 19064 31968 19116 31977
rect 21824 31968 21876 32020
rect 8668 31900 8720 31952
rect 14740 31900 14792 31952
rect 16948 31900 17000 31952
rect 18052 31900 18104 31952
rect 21916 31900 21968 31952
rect 22008 31900 22060 31952
rect 23388 31968 23440 32020
rect 23572 31968 23624 32020
rect 24124 32011 24176 32020
rect 24124 31977 24133 32011
rect 24133 31977 24167 32011
rect 24167 31977 24176 32011
rect 24124 31968 24176 31977
rect 24860 31968 24912 32020
rect 26148 32011 26200 32020
rect 26148 31977 26157 32011
rect 26157 31977 26191 32011
rect 26191 31977 26200 32011
rect 26148 31968 26200 31977
rect 23296 31943 23348 31952
rect 23296 31909 23305 31943
rect 23305 31909 23339 31943
rect 23339 31909 23348 31943
rect 23296 31900 23348 31909
rect 24216 31900 24268 31952
rect 2044 31832 2096 31884
rect 6184 31875 6236 31884
rect 6184 31841 6193 31875
rect 6193 31841 6227 31875
rect 6227 31841 6236 31875
rect 6184 31832 6236 31841
rect 7748 31832 7800 31884
rect 8300 31832 8352 31884
rect 9220 31875 9272 31884
rect 9220 31841 9229 31875
rect 9229 31841 9263 31875
rect 9263 31841 9272 31875
rect 9220 31832 9272 31841
rect 9864 31832 9916 31884
rect 14832 31832 14884 31884
rect 17040 31875 17092 31884
rect 17040 31841 17049 31875
rect 17049 31841 17083 31875
rect 17083 31841 17092 31875
rect 17040 31832 17092 31841
rect 21548 31832 21600 31884
rect 23480 31875 23532 31884
rect 23480 31841 23489 31875
rect 23489 31841 23523 31875
rect 23523 31841 23532 31875
rect 23480 31832 23532 31841
rect 24768 31832 24820 31884
rect 26608 31900 26660 31952
rect 27068 31968 27120 32020
rect 35808 31968 35860 32020
rect 27712 31943 27764 31952
rect 27712 31909 27721 31943
rect 27721 31909 27755 31943
rect 27755 31909 27764 31943
rect 27712 31900 27764 31909
rect 26240 31832 26292 31884
rect 28724 31832 28776 31884
rect 35440 31875 35492 31884
rect 35440 31841 35449 31875
rect 35449 31841 35483 31875
rect 35483 31841 35492 31875
rect 35440 31832 35492 31841
rect 2596 31807 2648 31816
rect 1676 31628 1728 31680
rect 2596 31773 2605 31807
rect 2605 31773 2639 31807
rect 2639 31773 2648 31807
rect 2596 31764 2648 31773
rect 5816 31764 5868 31816
rect 6552 31764 6604 31816
rect 4988 31696 5040 31748
rect 17684 31696 17736 31748
rect 20996 31807 21048 31816
rect 17960 31696 18012 31748
rect 20996 31773 21005 31807
rect 21005 31773 21039 31807
rect 21039 31773 21048 31807
rect 20996 31764 21048 31773
rect 24124 31764 24176 31816
rect 26884 31807 26936 31816
rect 26884 31773 26893 31807
rect 26893 31773 26927 31807
rect 26927 31773 26936 31807
rect 26884 31764 26936 31773
rect 5080 31628 5132 31680
rect 5264 31628 5316 31680
rect 14740 31628 14792 31680
rect 15844 31671 15896 31680
rect 15844 31637 15853 31671
rect 15853 31637 15887 31671
rect 15887 31637 15896 31671
rect 15844 31628 15896 31637
rect 16212 31628 16264 31680
rect 24676 31671 24728 31680
rect 24676 31637 24685 31671
rect 24685 31637 24719 31671
rect 24719 31637 24728 31671
rect 24676 31628 24728 31637
rect 28356 31628 28408 31680
rect 28816 31628 28868 31680
rect 29276 31628 29328 31680
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 34966 31526 35018 31578
rect 35030 31526 35082 31578
rect 35094 31526 35146 31578
rect 35158 31526 35210 31578
rect 3608 31467 3660 31476
rect 3608 31433 3617 31467
rect 3617 31433 3651 31467
rect 3651 31433 3660 31467
rect 3608 31424 3660 31433
rect 6552 31467 6604 31476
rect 6552 31433 6561 31467
rect 6561 31433 6595 31467
rect 6595 31433 6604 31467
rect 6552 31424 6604 31433
rect 7932 31467 7984 31476
rect 7932 31433 7941 31467
rect 7941 31433 7975 31467
rect 7975 31433 7984 31467
rect 7932 31424 7984 31433
rect 8300 31424 8352 31476
rect 13176 31467 13228 31476
rect 13176 31433 13185 31467
rect 13185 31433 13219 31467
rect 13219 31433 13228 31467
rect 13176 31424 13228 31433
rect 14280 31467 14332 31476
rect 14280 31433 14289 31467
rect 14289 31433 14323 31467
rect 14323 31433 14332 31467
rect 14280 31424 14332 31433
rect 17960 31424 18012 31476
rect 22008 31424 22060 31476
rect 23480 31467 23532 31476
rect 23480 31433 23489 31467
rect 23489 31433 23523 31467
rect 23523 31433 23532 31467
rect 23480 31424 23532 31433
rect 24216 31467 24268 31476
rect 24216 31433 24225 31467
rect 24225 31433 24259 31467
rect 24259 31433 24268 31467
rect 24216 31424 24268 31433
rect 26240 31424 26292 31476
rect 27068 31467 27120 31476
rect 27068 31433 27077 31467
rect 27077 31433 27111 31467
rect 27111 31433 27120 31467
rect 27068 31424 27120 31433
rect 27620 31467 27672 31476
rect 27620 31433 27629 31467
rect 27629 31433 27663 31467
rect 27663 31433 27672 31467
rect 27620 31424 27672 31433
rect 1400 31220 1452 31272
rect 2780 31220 2832 31272
rect 2872 31152 2924 31204
rect 4620 31356 4672 31408
rect 17684 31399 17736 31408
rect 17684 31365 17693 31399
rect 17693 31365 17727 31399
rect 17727 31365 17736 31399
rect 17684 31356 17736 31365
rect 5172 31331 5224 31340
rect 5172 31297 5181 31331
rect 5181 31297 5215 31331
rect 5215 31297 5224 31331
rect 5172 31288 5224 31297
rect 5264 31331 5316 31340
rect 5264 31297 5273 31331
rect 5273 31297 5307 31331
rect 5307 31297 5316 31331
rect 5264 31288 5316 31297
rect 8852 31288 8904 31340
rect 10416 31288 10468 31340
rect 20996 31288 21048 31340
rect 21916 31356 21968 31408
rect 5080 31263 5132 31272
rect 5080 31229 5089 31263
rect 5089 31229 5123 31263
rect 5123 31229 5132 31263
rect 5080 31220 5132 31229
rect 8024 31220 8076 31272
rect 13176 31220 13228 31272
rect 14280 31220 14332 31272
rect 21548 31263 21600 31272
rect 9956 31152 10008 31204
rect 1676 31127 1728 31136
rect 1676 31093 1685 31127
rect 1685 31093 1719 31127
rect 1719 31093 1728 31127
rect 1676 31084 1728 31093
rect 4712 31127 4764 31136
rect 4712 31093 4721 31127
rect 4721 31093 4755 31127
rect 4755 31093 4764 31127
rect 4712 31084 4764 31093
rect 5816 31127 5868 31136
rect 5816 31093 5825 31127
rect 5825 31093 5859 31127
rect 5859 31093 5868 31127
rect 5816 31084 5868 31093
rect 6184 31084 6236 31136
rect 6828 31084 6880 31136
rect 8668 31084 8720 31136
rect 9680 31127 9732 31136
rect 9680 31093 9689 31127
rect 9689 31093 9723 31127
rect 9723 31093 9732 31127
rect 9680 31084 9732 31093
rect 10416 31127 10468 31136
rect 10416 31093 10425 31127
rect 10425 31093 10459 31127
rect 10459 31093 10468 31127
rect 10416 31084 10468 31093
rect 12256 31127 12308 31136
rect 12256 31093 12265 31127
rect 12265 31093 12299 31127
rect 12299 31093 12308 31127
rect 15476 31152 15528 31204
rect 16212 31152 16264 31204
rect 21548 31229 21557 31263
rect 21557 31229 21591 31263
rect 21591 31229 21600 31263
rect 21548 31220 21600 31229
rect 24032 31288 24084 31340
rect 28172 31331 28224 31340
rect 28172 31297 28181 31331
rect 28181 31297 28215 31331
rect 28215 31297 28224 31331
rect 28172 31288 28224 31297
rect 27068 31220 27120 31272
rect 21088 31195 21140 31204
rect 21088 31161 21097 31195
rect 21097 31161 21131 31195
rect 21131 31161 21140 31195
rect 21088 31152 21140 31161
rect 12256 31084 12308 31093
rect 12716 31084 12768 31136
rect 13820 31127 13872 31136
rect 13820 31093 13829 31127
rect 13829 31093 13863 31127
rect 13863 31093 13872 31127
rect 13820 31084 13872 31093
rect 16672 31127 16724 31136
rect 16672 31093 16681 31127
rect 16681 31093 16715 31127
rect 16715 31093 16724 31127
rect 16672 31084 16724 31093
rect 17592 31084 17644 31136
rect 18052 31084 18104 31136
rect 25320 31084 25372 31136
rect 28080 31127 28132 31136
rect 28080 31093 28089 31127
rect 28089 31093 28123 31127
rect 28123 31093 28132 31127
rect 28080 31084 28132 31093
rect 28724 31127 28776 31136
rect 28724 31093 28733 31127
rect 28733 31093 28767 31127
rect 28767 31093 28776 31127
rect 28724 31084 28776 31093
rect 28816 31084 28868 31136
rect 34704 31084 34756 31136
rect 35440 31127 35492 31136
rect 35440 31093 35449 31127
rect 35449 31093 35483 31127
rect 35483 31093 35492 31127
rect 35440 31084 35492 31093
rect 19606 30982 19658 31034
rect 19670 30982 19722 31034
rect 19734 30982 19786 31034
rect 19798 30982 19850 31034
rect 2872 30923 2924 30932
rect 2872 30889 2881 30923
rect 2881 30889 2915 30923
rect 2915 30889 2924 30923
rect 2872 30880 2924 30889
rect 4988 30880 5040 30932
rect 5080 30880 5132 30932
rect 6460 30880 6512 30932
rect 9864 30923 9916 30932
rect 9864 30889 9873 30923
rect 9873 30889 9907 30923
rect 9907 30889 9916 30923
rect 9864 30880 9916 30889
rect 14740 30923 14792 30932
rect 14740 30889 14749 30923
rect 14749 30889 14783 30923
rect 14783 30889 14792 30923
rect 14740 30880 14792 30889
rect 15200 30880 15252 30932
rect 17684 30880 17736 30932
rect 18972 30923 19024 30932
rect 18972 30889 18981 30923
rect 18981 30889 19015 30923
rect 19015 30889 19024 30923
rect 18972 30880 19024 30889
rect 21548 30880 21600 30932
rect 24032 30880 24084 30932
rect 4712 30812 4764 30864
rect 13636 30812 13688 30864
rect 21088 30812 21140 30864
rect 24676 30880 24728 30932
rect 28172 30880 28224 30932
rect 28724 30880 28776 30932
rect 35624 30923 35676 30932
rect 35624 30889 35633 30923
rect 35633 30889 35667 30923
rect 35667 30889 35676 30923
rect 35624 30880 35676 30889
rect 2044 30744 2096 30796
rect 4804 30787 4856 30796
rect 4804 30753 4813 30787
rect 4813 30753 4847 30787
rect 4847 30753 4856 30787
rect 4804 30744 4856 30753
rect 6000 30787 6052 30796
rect 6000 30753 6009 30787
rect 6009 30753 6043 30787
rect 6043 30753 6052 30787
rect 6000 30744 6052 30753
rect 8392 30787 8444 30796
rect 8392 30753 8401 30787
rect 8401 30753 8435 30787
rect 8435 30753 8444 30787
rect 8392 30744 8444 30753
rect 9680 30744 9732 30796
rect 10600 30744 10652 30796
rect 13728 30744 13780 30796
rect 15936 30787 15988 30796
rect 15936 30753 15945 30787
rect 15945 30753 15979 30787
rect 15979 30753 15988 30787
rect 15936 30744 15988 30753
rect 20168 30744 20220 30796
rect 20996 30744 21048 30796
rect 23480 30744 23532 30796
rect 24216 30744 24268 30796
rect 24584 30787 24636 30796
rect 24584 30753 24593 30787
rect 24593 30753 24627 30787
rect 24627 30753 24636 30787
rect 24584 30744 24636 30753
rect 24768 30744 24820 30796
rect 25044 30787 25096 30796
rect 25044 30753 25053 30787
rect 25053 30753 25087 30787
rect 25087 30753 25096 30787
rect 25044 30744 25096 30753
rect 26516 30787 26568 30796
rect 26516 30753 26525 30787
rect 26525 30753 26559 30787
rect 26559 30753 26568 30787
rect 26516 30744 26568 30753
rect 28080 30744 28132 30796
rect 28908 30744 28960 30796
rect 35532 30744 35584 30796
rect 1400 30676 1452 30728
rect 4896 30719 4948 30728
rect 4896 30685 4905 30719
rect 4905 30685 4939 30719
rect 4939 30685 4948 30719
rect 4896 30676 4948 30685
rect 3976 30608 4028 30660
rect 5264 30676 5316 30728
rect 8484 30719 8536 30728
rect 8484 30685 8493 30719
rect 8493 30685 8527 30719
rect 8527 30685 8536 30719
rect 8484 30676 8536 30685
rect 8116 30608 8168 30660
rect 8852 30676 8904 30728
rect 9588 30676 9640 30728
rect 10508 30719 10560 30728
rect 10508 30685 10517 30719
rect 10517 30685 10551 30719
rect 10551 30685 10560 30719
rect 10508 30676 10560 30685
rect 13544 30719 13596 30728
rect 13544 30685 13553 30719
rect 13553 30685 13587 30719
rect 13587 30685 13596 30719
rect 16028 30719 16080 30728
rect 13544 30676 13596 30685
rect 16028 30685 16037 30719
rect 16037 30685 16071 30719
rect 16071 30685 16080 30719
rect 16028 30676 16080 30685
rect 14924 30608 14976 30660
rect 16672 30676 16724 30728
rect 16948 30676 17000 30728
rect 5356 30540 5408 30592
rect 8024 30583 8076 30592
rect 8024 30549 8033 30583
rect 8033 30549 8067 30583
rect 8067 30549 8076 30583
rect 8024 30540 8076 30549
rect 12256 30540 12308 30592
rect 12624 30540 12676 30592
rect 12808 30583 12860 30592
rect 12808 30549 12817 30583
rect 12817 30549 12851 30583
rect 12851 30549 12860 30583
rect 12808 30540 12860 30549
rect 12992 30583 13044 30592
rect 12992 30549 13001 30583
rect 13001 30549 13035 30583
rect 13035 30549 13044 30583
rect 12992 30540 13044 30549
rect 14648 30540 14700 30592
rect 16120 30540 16172 30592
rect 17500 30676 17552 30728
rect 17592 30719 17644 30728
rect 17592 30685 17604 30719
rect 17604 30685 17638 30719
rect 17638 30685 17644 30719
rect 25320 30719 25372 30728
rect 17592 30676 17644 30685
rect 25320 30685 25329 30719
rect 25329 30685 25363 30719
rect 25363 30685 25372 30719
rect 25320 30676 25372 30685
rect 17776 30540 17828 30592
rect 23756 30583 23808 30592
rect 23756 30549 23765 30583
rect 23765 30549 23799 30583
rect 23799 30549 23808 30583
rect 23756 30540 23808 30549
rect 24768 30540 24820 30592
rect 28724 30540 28776 30592
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 34966 30438 35018 30490
rect 35030 30438 35082 30490
rect 35094 30438 35146 30490
rect 35158 30438 35210 30490
rect 4804 30336 4856 30388
rect 6000 30379 6052 30388
rect 6000 30345 6009 30379
rect 6009 30345 6043 30379
rect 6043 30345 6052 30379
rect 6000 30336 6052 30345
rect 6828 30336 6880 30388
rect 8208 30268 8260 30320
rect 8484 30336 8536 30388
rect 9956 30379 10008 30388
rect 9956 30345 9965 30379
rect 9965 30345 9999 30379
rect 9999 30345 10008 30379
rect 9956 30336 10008 30345
rect 14648 30336 14700 30388
rect 15660 30336 15712 30388
rect 15844 30336 15896 30388
rect 17500 30336 17552 30388
rect 21088 30336 21140 30388
rect 23480 30379 23532 30388
rect 23480 30345 23489 30379
rect 23489 30345 23523 30379
rect 23523 30345 23532 30379
rect 23480 30336 23532 30345
rect 23756 30336 23808 30388
rect 25044 30336 25096 30388
rect 26516 30336 26568 30388
rect 28080 30336 28132 30388
rect 24676 30268 24728 30320
rect 34612 30268 34664 30320
rect 35348 30268 35400 30320
rect 35716 30268 35768 30320
rect 4988 30200 5040 30252
rect 5356 30200 5408 30252
rect 8576 30243 8628 30252
rect 8576 30209 8585 30243
rect 8585 30209 8619 30243
rect 8619 30209 8628 30243
rect 8576 30200 8628 30209
rect 11888 30243 11940 30252
rect 1400 30175 1452 30184
rect 1400 30141 1409 30175
rect 1409 30141 1443 30175
rect 1443 30141 1452 30175
rect 1400 30132 1452 30141
rect 5540 30132 5592 30184
rect 11888 30209 11897 30243
rect 11897 30209 11931 30243
rect 11931 30209 11940 30243
rect 11888 30200 11940 30209
rect 12808 30200 12860 30252
rect 15752 30243 15804 30252
rect 15752 30209 15780 30243
rect 15780 30209 15804 30243
rect 15752 30200 15804 30209
rect 16120 30200 16172 30252
rect 18512 30243 18564 30252
rect 14188 30175 14240 30184
rect 1676 30107 1728 30116
rect 1676 30073 1710 30107
rect 1710 30073 1728 30107
rect 1676 30064 1728 30073
rect 5080 30107 5132 30116
rect 5080 30073 5089 30107
rect 5089 30073 5123 30107
rect 5123 30073 5132 30107
rect 5080 30064 5132 30073
rect 7932 30064 7984 30116
rect 8392 30064 8444 30116
rect 9312 30064 9364 30116
rect 10508 30064 10560 30116
rect 12072 30064 12124 30116
rect 2044 29996 2096 30048
rect 2964 29996 3016 30048
rect 3976 29996 4028 30048
rect 4160 30039 4212 30048
rect 4160 30005 4169 30039
rect 4169 30005 4203 30039
rect 4203 30005 4212 30039
rect 4160 29996 4212 30005
rect 5540 29996 5592 30048
rect 10600 30039 10652 30048
rect 10600 30005 10609 30039
rect 10609 30005 10643 30039
rect 10643 30005 10652 30039
rect 10600 29996 10652 30005
rect 11336 29996 11388 30048
rect 12348 29996 12400 30048
rect 12440 30039 12492 30048
rect 12440 30005 12449 30039
rect 12449 30005 12483 30039
rect 12483 30005 12492 30039
rect 12440 29996 12492 30005
rect 12624 29996 12676 30048
rect 14188 30141 14197 30175
rect 14197 30141 14231 30175
rect 14231 30141 14240 30175
rect 14188 30132 14240 30141
rect 15292 30175 15344 30184
rect 15292 30141 15301 30175
rect 15301 30141 15335 30175
rect 15335 30141 15344 30175
rect 15292 30132 15344 30141
rect 18512 30209 18521 30243
rect 18521 30209 18555 30243
rect 18555 30209 18564 30243
rect 18512 30200 18564 30209
rect 18696 30243 18748 30252
rect 18696 30209 18705 30243
rect 18705 30209 18739 30243
rect 18739 30209 18748 30243
rect 18696 30200 18748 30209
rect 19248 30200 19300 30252
rect 20168 30243 20220 30252
rect 20168 30209 20177 30243
rect 20177 30209 20211 30243
rect 20211 30209 20220 30243
rect 20168 30200 20220 30209
rect 24032 30132 24084 30184
rect 25320 30132 25372 30184
rect 35348 30132 35400 30184
rect 13636 30064 13688 30116
rect 17500 30107 17552 30116
rect 17500 30073 17509 30107
rect 17509 30073 17543 30107
rect 17543 30073 17552 30107
rect 17500 30064 17552 30073
rect 17960 30064 18012 30116
rect 13728 29996 13780 30048
rect 14372 30039 14424 30048
rect 14372 30005 14381 30039
rect 14381 30005 14415 30039
rect 14415 30005 14424 30039
rect 14372 29996 14424 30005
rect 15660 29996 15712 30048
rect 16028 29996 16080 30048
rect 17132 30039 17184 30048
rect 17132 30005 17141 30039
rect 17141 30005 17175 30039
rect 17175 30005 17184 30039
rect 17132 29996 17184 30005
rect 18052 30039 18104 30048
rect 18052 30005 18061 30039
rect 18061 30005 18095 30039
rect 18095 30005 18104 30039
rect 18052 29996 18104 30005
rect 19984 30039 20036 30048
rect 19984 30005 19993 30039
rect 19993 30005 20027 30039
rect 20027 30005 20036 30039
rect 19984 29996 20036 30005
rect 25780 29996 25832 30048
rect 28724 30039 28776 30048
rect 28724 30005 28733 30039
rect 28733 30005 28767 30039
rect 28767 30005 28776 30039
rect 28724 29996 28776 30005
rect 35532 29996 35584 30048
rect 19606 29894 19658 29946
rect 19670 29894 19722 29946
rect 19734 29894 19786 29946
rect 19798 29894 19850 29946
rect 1676 29792 1728 29844
rect 4896 29792 4948 29844
rect 5540 29792 5592 29844
rect 7932 29835 7984 29844
rect 7932 29801 7941 29835
rect 7941 29801 7975 29835
rect 7975 29801 7984 29835
rect 7932 29792 7984 29801
rect 8576 29792 8628 29844
rect 10600 29792 10652 29844
rect 13544 29835 13596 29844
rect 13544 29801 13553 29835
rect 13553 29801 13587 29835
rect 13587 29801 13596 29835
rect 13544 29792 13596 29801
rect 14188 29835 14240 29844
rect 14188 29801 14197 29835
rect 14197 29801 14231 29835
rect 14231 29801 14240 29835
rect 14188 29792 14240 29801
rect 14924 29792 14976 29844
rect 16028 29792 16080 29844
rect 17132 29792 17184 29844
rect 18696 29835 18748 29844
rect 18696 29801 18705 29835
rect 18705 29801 18739 29835
rect 18739 29801 18748 29835
rect 18696 29792 18748 29801
rect 21088 29835 21140 29844
rect 21088 29801 21097 29835
rect 21097 29801 21131 29835
rect 21131 29801 21140 29835
rect 21088 29792 21140 29801
rect 24124 29792 24176 29844
rect 25320 29792 25372 29844
rect 25780 29835 25832 29844
rect 25780 29801 25789 29835
rect 25789 29801 25823 29835
rect 25823 29801 25832 29835
rect 25780 29792 25832 29801
rect 35624 29835 35676 29844
rect 35624 29801 35633 29835
rect 35633 29801 35667 29835
rect 35667 29801 35676 29835
rect 35624 29792 35676 29801
rect 5080 29724 5132 29776
rect 7104 29724 7156 29776
rect 8668 29724 8720 29776
rect 9956 29767 10008 29776
rect 9956 29733 9990 29767
rect 9990 29733 10008 29767
rect 9956 29724 10008 29733
rect 14372 29724 14424 29776
rect 17592 29767 17644 29776
rect 17592 29733 17601 29767
rect 17601 29733 17635 29767
rect 17635 29733 17644 29767
rect 17592 29724 17644 29733
rect 20996 29724 21048 29776
rect 32680 29724 32732 29776
rect 1676 29699 1728 29708
rect 1676 29665 1710 29699
rect 1710 29665 1728 29699
rect 1676 29656 1728 29665
rect 5264 29656 5316 29708
rect 9680 29699 9732 29708
rect 9680 29665 9689 29699
rect 9689 29665 9723 29699
rect 9723 29665 9732 29699
rect 9680 29656 9732 29665
rect 10508 29656 10560 29708
rect 12256 29656 12308 29708
rect 15200 29656 15252 29708
rect 15752 29656 15804 29708
rect 17040 29656 17092 29708
rect 19524 29699 19576 29708
rect 19524 29665 19533 29699
rect 19533 29665 19567 29699
rect 19567 29665 19576 29699
rect 19524 29656 19576 29665
rect 23572 29699 23624 29708
rect 23572 29665 23581 29699
rect 23581 29665 23615 29699
rect 23615 29665 23624 29699
rect 23572 29656 23624 29665
rect 25044 29699 25096 29708
rect 25044 29665 25053 29699
rect 25053 29665 25087 29699
rect 25087 29665 25096 29699
rect 25044 29656 25096 29665
rect 27712 29699 27764 29708
rect 27712 29665 27721 29699
rect 27721 29665 27755 29699
rect 27755 29665 27764 29699
rect 27712 29656 27764 29665
rect 34520 29656 34572 29708
rect 1400 29631 1452 29640
rect 1400 29597 1409 29631
rect 1409 29597 1443 29631
rect 1443 29597 1452 29631
rect 1400 29588 1452 29597
rect 7472 29588 7524 29640
rect 8024 29588 8076 29640
rect 8668 29631 8720 29640
rect 8668 29597 8677 29631
rect 8677 29597 8711 29631
rect 8711 29597 8720 29631
rect 8668 29588 8720 29597
rect 12072 29588 12124 29640
rect 18144 29631 18196 29640
rect 7840 29452 7892 29504
rect 8024 29495 8076 29504
rect 8024 29461 8033 29495
rect 8033 29461 8067 29495
rect 8067 29461 8076 29495
rect 8024 29452 8076 29461
rect 15016 29452 15068 29504
rect 18144 29597 18153 29631
rect 18153 29597 18187 29631
rect 18187 29597 18196 29631
rect 18144 29588 18196 29597
rect 19248 29588 19300 29640
rect 18880 29520 18932 29572
rect 19984 29588 20036 29640
rect 24860 29588 24912 29640
rect 25320 29631 25372 29640
rect 25320 29597 25329 29631
rect 25329 29597 25363 29631
rect 25363 29597 25372 29631
rect 25320 29588 25372 29597
rect 25780 29588 25832 29640
rect 26148 29588 26200 29640
rect 31300 29631 31352 29640
rect 31300 29597 31309 29631
rect 31309 29597 31343 29631
rect 31343 29597 31352 29631
rect 31300 29588 31352 29597
rect 16028 29452 16080 29504
rect 16580 29452 16632 29504
rect 19064 29452 19116 29504
rect 19892 29452 19944 29504
rect 24492 29452 24544 29504
rect 26516 29452 26568 29504
rect 28724 29452 28776 29504
rect 33140 29452 33192 29504
rect 34796 29452 34848 29504
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 34966 29350 35018 29402
rect 35030 29350 35082 29402
rect 35094 29350 35146 29402
rect 35158 29350 35210 29402
rect 1676 29291 1728 29300
rect 1676 29257 1685 29291
rect 1685 29257 1719 29291
rect 1719 29257 1728 29291
rect 1676 29248 1728 29257
rect 2044 29291 2096 29300
rect 2044 29257 2053 29291
rect 2053 29257 2087 29291
rect 2087 29257 2096 29291
rect 2044 29248 2096 29257
rect 3332 29291 3384 29300
rect 3332 29257 3341 29291
rect 3341 29257 3375 29291
rect 3375 29257 3384 29291
rect 3332 29248 3384 29257
rect 5172 29248 5224 29300
rect 7104 29291 7156 29300
rect 7104 29257 7113 29291
rect 7113 29257 7147 29291
rect 7147 29257 7156 29291
rect 7104 29248 7156 29257
rect 7472 29291 7524 29300
rect 7472 29257 7481 29291
rect 7481 29257 7515 29291
rect 7515 29257 7524 29291
rect 7472 29248 7524 29257
rect 9312 29291 9364 29300
rect 9312 29257 9321 29291
rect 9321 29257 9355 29291
rect 9355 29257 9364 29291
rect 9312 29248 9364 29257
rect 9956 29291 10008 29300
rect 9956 29257 9965 29291
rect 9965 29257 9999 29291
rect 9999 29257 10008 29291
rect 9956 29248 10008 29257
rect 10416 29291 10468 29300
rect 10416 29257 10425 29291
rect 10425 29257 10459 29291
rect 10459 29257 10468 29291
rect 10416 29248 10468 29257
rect 12256 29291 12308 29300
rect 12256 29257 12265 29291
rect 12265 29257 12299 29291
rect 12299 29257 12308 29291
rect 12256 29248 12308 29257
rect 15476 29291 15528 29300
rect 15476 29257 15485 29291
rect 15485 29257 15519 29291
rect 15519 29257 15528 29291
rect 15476 29248 15528 29257
rect 12072 29180 12124 29232
rect 15936 29223 15988 29232
rect 15936 29189 15945 29223
rect 15945 29189 15979 29223
rect 15979 29189 15988 29223
rect 15936 29180 15988 29189
rect 1400 29112 1452 29164
rect 1952 29112 2004 29164
rect 10968 29155 11020 29164
rect 2688 29044 2740 29096
rect 4068 29044 4120 29096
rect 5264 29044 5316 29096
rect 7932 29087 7984 29096
rect 7932 29053 7941 29087
rect 7941 29053 7975 29087
rect 7975 29053 7984 29087
rect 7932 29044 7984 29053
rect 10968 29121 10977 29155
rect 10977 29121 11011 29155
rect 11011 29121 11020 29155
rect 10968 29112 11020 29121
rect 16396 29155 16448 29164
rect 16396 29121 16405 29155
rect 16405 29121 16439 29155
rect 16439 29121 16448 29155
rect 16396 29112 16448 29121
rect 18236 29248 18288 29300
rect 19524 29248 19576 29300
rect 19984 29248 20036 29300
rect 23572 29248 23624 29300
rect 27712 29248 27764 29300
rect 17040 29223 17092 29232
rect 17040 29189 17049 29223
rect 17049 29189 17083 29223
rect 17083 29189 17092 29223
rect 17040 29180 17092 29189
rect 18696 29180 18748 29232
rect 18880 29223 18932 29232
rect 18880 29189 18889 29223
rect 18889 29189 18923 29223
rect 18923 29189 18932 29223
rect 18880 29180 18932 29189
rect 25044 29180 25096 29232
rect 32680 29223 32732 29232
rect 32680 29189 32689 29223
rect 32689 29189 32723 29223
rect 32723 29189 32732 29223
rect 32680 29180 32732 29189
rect 31300 29155 31352 29164
rect 8208 29087 8260 29096
rect 8208 29053 8242 29087
rect 8242 29053 8260 29087
rect 8208 29044 8260 29053
rect 5448 28976 5500 29028
rect 13544 29044 13596 29096
rect 16212 29044 16264 29096
rect 17132 29044 17184 29096
rect 20168 29044 20220 29096
rect 24032 29044 24084 29096
rect 24584 29044 24636 29096
rect 25044 29087 25096 29096
rect 25044 29053 25053 29087
rect 25053 29053 25087 29087
rect 25087 29053 25096 29087
rect 25044 29044 25096 29053
rect 31300 29121 31309 29155
rect 31309 29121 31343 29155
rect 31343 29121 31352 29155
rect 31300 29112 31352 29121
rect 31944 29044 31996 29096
rect 9588 28908 9640 28960
rect 10508 28908 10560 28960
rect 17776 28976 17828 29028
rect 14372 28908 14424 28960
rect 15108 28908 15160 28960
rect 19248 28976 19300 29028
rect 19892 29019 19944 29028
rect 19892 28985 19926 29019
rect 19926 28985 19944 29019
rect 19892 28976 19944 28985
rect 24676 28976 24728 29028
rect 25320 29019 25372 29028
rect 25320 28985 25354 29019
rect 25354 28985 25372 29019
rect 25320 28976 25372 28985
rect 31576 29019 31628 29028
rect 31576 28985 31610 29019
rect 31610 28985 31628 29019
rect 31576 28976 31628 28985
rect 34520 28976 34572 29028
rect 34796 28976 34848 29028
rect 18880 28908 18932 28960
rect 24124 28951 24176 28960
rect 24124 28917 24133 28951
rect 24133 28917 24167 28951
rect 24167 28917 24176 28951
rect 24124 28908 24176 28917
rect 24860 28908 24912 28960
rect 26424 28951 26476 28960
rect 26424 28917 26433 28951
rect 26433 28917 26467 28951
rect 26467 28917 26476 28951
rect 26424 28908 26476 28917
rect 30840 28908 30892 28960
rect 34336 28951 34388 28960
rect 34336 28917 34345 28951
rect 34345 28917 34379 28951
rect 34379 28917 34388 28951
rect 34336 28908 34388 28917
rect 34888 28908 34940 28960
rect 19606 28806 19658 28858
rect 19670 28806 19722 28858
rect 19734 28806 19786 28858
rect 19798 28806 19850 28858
rect 1952 28747 2004 28756
rect 1952 28713 1961 28747
rect 1961 28713 1995 28747
rect 1995 28713 2004 28747
rect 1952 28704 2004 28713
rect 2688 28704 2740 28756
rect 5448 28747 5500 28756
rect 5448 28713 5457 28747
rect 5457 28713 5491 28747
rect 5491 28713 5500 28747
rect 5448 28704 5500 28713
rect 8300 28704 8352 28756
rect 10508 28747 10560 28756
rect 10508 28713 10517 28747
rect 10517 28713 10551 28747
rect 10551 28713 10560 28747
rect 10508 28704 10560 28713
rect 10968 28704 11020 28756
rect 12348 28704 12400 28756
rect 12808 28747 12860 28756
rect 7564 28636 7616 28688
rect 12808 28713 12817 28747
rect 12817 28713 12851 28747
rect 12851 28713 12860 28747
rect 12808 28704 12860 28713
rect 13544 28747 13596 28756
rect 13544 28713 13553 28747
rect 13553 28713 13587 28747
rect 13587 28713 13596 28747
rect 13544 28704 13596 28713
rect 13820 28704 13872 28756
rect 14372 28747 14424 28756
rect 14372 28713 14381 28747
rect 14381 28713 14415 28747
rect 14415 28713 14424 28747
rect 14372 28704 14424 28713
rect 15016 28704 15068 28756
rect 15200 28704 15252 28756
rect 15844 28747 15896 28756
rect 15844 28713 15853 28747
rect 15853 28713 15887 28747
rect 15887 28713 15896 28747
rect 15844 28704 15896 28713
rect 16396 28747 16448 28756
rect 16396 28713 16405 28747
rect 16405 28713 16439 28747
rect 16439 28713 16448 28747
rect 16396 28704 16448 28713
rect 18236 28747 18288 28756
rect 18236 28713 18245 28747
rect 18245 28713 18279 28747
rect 18279 28713 18288 28747
rect 18236 28704 18288 28713
rect 18972 28747 19024 28756
rect 18972 28713 18981 28747
rect 18981 28713 19015 28747
rect 19015 28713 19024 28747
rect 18972 28704 19024 28713
rect 19248 28747 19300 28756
rect 19248 28713 19257 28747
rect 19257 28713 19291 28747
rect 19291 28713 19300 28747
rect 19248 28704 19300 28713
rect 20168 28704 20220 28756
rect 24032 28747 24084 28756
rect 15752 28679 15804 28688
rect 2780 28611 2832 28620
rect 2780 28577 2789 28611
rect 2789 28577 2823 28611
rect 2823 28577 2832 28611
rect 3884 28611 3936 28620
rect 2780 28568 2832 28577
rect 3884 28577 3893 28611
rect 3893 28577 3927 28611
rect 3927 28577 3936 28611
rect 4068 28611 4120 28620
rect 3884 28568 3936 28577
rect 4068 28577 4077 28611
rect 4077 28577 4111 28611
rect 4111 28577 4120 28611
rect 4068 28568 4120 28577
rect 4620 28568 4672 28620
rect 5264 28568 5316 28620
rect 6644 28568 6696 28620
rect 7932 28568 7984 28620
rect 9680 28611 9732 28620
rect 9680 28577 9689 28611
rect 9689 28577 9723 28611
rect 9723 28577 9732 28611
rect 9680 28568 9732 28577
rect 11428 28611 11480 28620
rect 11428 28577 11437 28611
rect 11437 28577 11471 28611
rect 11471 28577 11480 28611
rect 11428 28568 11480 28577
rect 1860 28500 1912 28552
rect 2964 28543 3016 28552
rect 2964 28509 2973 28543
rect 2973 28509 3007 28543
rect 3007 28509 3016 28543
rect 11520 28543 11572 28552
rect 2964 28500 3016 28509
rect 11520 28509 11529 28543
rect 11529 28509 11563 28543
rect 11563 28509 11572 28543
rect 11520 28500 11572 28509
rect 15752 28645 15761 28679
rect 15761 28645 15795 28679
rect 15795 28645 15804 28679
rect 15752 28636 15804 28645
rect 19708 28636 19760 28688
rect 12716 28568 12768 28620
rect 13728 28611 13780 28620
rect 13728 28577 13737 28611
rect 13737 28577 13771 28611
rect 13771 28577 13780 28611
rect 13728 28568 13780 28577
rect 24032 28713 24041 28747
rect 24041 28713 24075 28747
rect 24075 28713 24084 28747
rect 24032 28704 24084 28713
rect 24768 28704 24820 28756
rect 25136 28704 25188 28756
rect 25688 28704 25740 28756
rect 26148 28704 26200 28756
rect 31576 28704 31628 28756
rect 33508 28747 33560 28756
rect 33508 28713 33517 28747
rect 33517 28713 33551 28747
rect 33551 28713 33560 28747
rect 33508 28704 33560 28713
rect 24676 28679 24728 28688
rect 24676 28645 24685 28679
rect 24685 28645 24719 28679
rect 24719 28645 24728 28679
rect 24676 28636 24728 28645
rect 26424 28636 26476 28688
rect 34888 28679 34940 28688
rect 34888 28645 34922 28679
rect 34922 28645 34940 28679
rect 34888 28636 34940 28645
rect 20720 28568 20772 28620
rect 21180 28611 21232 28620
rect 21180 28577 21214 28611
rect 21214 28577 21232 28611
rect 21180 28568 21232 28577
rect 32220 28568 32272 28620
rect 11796 28500 11848 28552
rect 16028 28543 16080 28552
rect 16028 28509 16037 28543
rect 16037 28509 16071 28543
rect 16071 28509 16080 28543
rect 16028 28500 16080 28509
rect 16488 28500 16540 28552
rect 19892 28543 19944 28552
rect 19892 28509 19901 28543
rect 19901 28509 19935 28543
rect 19935 28509 19944 28543
rect 19892 28500 19944 28509
rect 24584 28500 24636 28552
rect 25504 28543 25556 28552
rect 25504 28509 25513 28543
rect 25513 28509 25547 28543
rect 25547 28509 25556 28543
rect 25504 28500 25556 28509
rect 26516 28543 26568 28552
rect 19984 28432 20036 28484
rect 22284 28475 22336 28484
rect 22284 28441 22293 28475
rect 22293 28441 22327 28475
rect 22327 28441 22336 28475
rect 22284 28432 22336 28441
rect 25044 28364 25096 28416
rect 26148 28364 26200 28416
rect 26516 28509 26525 28543
rect 26525 28509 26559 28543
rect 26559 28509 26568 28543
rect 26516 28500 26568 28509
rect 30932 28543 30984 28552
rect 30932 28509 30941 28543
rect 30941 28509 30975 28543
rect 30975 28509 30984 28543
rect 30932 28500 30984 28509
rect 30840 28432 30892 28484
rect 27896 28407 27948 28416
rect 27896 28373 27905 28407
rect 27905 28373 27939 28407
rect 27939 28373 27948 28407
rect 27896 28364 27948 28373
rect 30012 28407 30064 28416
rect 30012 28373 30021 28407
rect 30021 28373 30055 28407
rect 30055 28373 30064 28407
rect 30012 28364 30064 28373
rect 30472 28407 30524 28416
rect 30472 28373 30481 28407
rect 30481 28373 30515 28407
rect 30515 28373 30524 28407
rect 30472 28364 30524 28373
rect 31944 28407 31996 28416
rect 31944 28373 31953 28407
rect 31953 28373 31987 28407
rect 31987 28373 31996 28407
rect 31944 28364 31996 28373
rect 34336 28364 34388 28416
rect 35992 28407 36044 28416
rect 35992 28373 36001 28407
rect 36001 28373 36035 28407
rect 36035 28373 36044 28407
rect 35992 28364 36044 28373
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 34966 28262 35018 28314
rect 35030 28262 35082 28314
rect 35094 28262 35146 28314
rect 35158 28262 35210 28314
rect 1860 28203 1912 28212
rect 1860 28169 1869 28203
rect 1869 28169 1903 28203
rect 1903 28169 1912 28203
rect 1860 28160 1912 28169
rect 4896 28160 4948 28212
rect 6644 28203 6696 28212
rect 6644 28169 6653 28203
rect 6653 28169 6687 28203
rect 6687 28169 6696 28203
rect 6644 28160 6696 28169
rect 9588 28160 9640 28212
rect 9680 28160 9732 28212
rect 11152 28203 11204 28212
rect 11152 28169 11161 28203
rect 11161 28169 11195 28203
rect 11195 28169 11204 28203
rect 11152 28160 11204 28169
rect 11520 28160 11572 28212
rect 11796 28203 11848 28212
rect 11796 28169 11805 28203
rect 11805 28169 11839 28203
rect 11839 28169 11848 28203
rect 11796 28160 11848 28169
rect 12716 28160 12768 28212
rect 13728 28203 13780 28212
rect 13728 28169 13737 28203
rect 13737 28169 13771 28203
rect 13771 28169 13780 28203
rect 13728 28160 13780 28169
rect 15752 28160 15804 28212
rect 16028 28160 16080 28212
rect 21640 28203 21692 28212
rect 21640 28169 21649 28203
rect 21649 28169 21683 28203
rect 21683 28169 21692 28203
rect 21640 28160 21692 28169
rect 24584 28203 24636 28212
rect 24584 28169 24593 28203
rect 24593 28169 24627 28203
rect 24627 28169 24636 28203
rect 24584 28160 24636 28169
rect 25688 28203 25740 28212
rect 25688 28169 25697 28203
rect 25697 28169 25731 28203
rect 25731 28169 25740 28203
rect 25688 28160 25740 28169
rect 26424 28160 26476 28212
rect 30932 28160 30984 28212
rect 32220 28203 32272 28212
rect 32220 28169 32229 28203
rect 32229 28169 32263 28203
rect 32263 28169 32272 28203
rect 32220 28160 32272 28169
rect 33968 28160 34020 28212
rect 34612 28160 34664 28212
rect 13636 28092 13688 28144
rect 34520 28092 34572 28144
rect 1952 28024 2004 28076
rect 5356 28067 5408 28076
rect 5356 28033 5365 28067
rect 5365 28033 5399 28067
rect 5399 28033 5408 28067
rect 5356 28024 5408 28033
rect 8116 28067 8168 28076
rect 8116 28033 8125 28067
rect 8125 28033 8159 28067
rect 8159 28033 8168 28067
rect 8116 28024 8168 28033
rect 15108 28024 15160 28076
rect 15844 28024 15896 28076
rect 19708 28067 19760 28076
rect 19708 28033 19717 28067
rect 19717 28033 19751 28067
rect 19751 28033 19760 28067
rect 19708 28024 19760 28033
rect 21180 28067 21232 28076
rect 21180 28033 21189 28067
rect 21189 28033 21223 28067
rect 21223 28033 21232 28067
rect 21180 28024 21232 28033
rect 22468 28024 22520 28076
rect 24860 28024 24912 28076
rect 25504 28024 25556 28076
rect 5448 27956 5500 28008
rect 8208 27956 8260 28008
rect 12440 27999 12492 28008
rect 12440 27965 12449 27999
rect 12449 27965 12483 27999
rect 12483 27965 12492 27999
rect 12440 27956 12492 27965
rect 18880 27956 18932 28008
rect 19064 27956 19116 28008
rect 19340 27956 19392 28008
rect 26148 27999 26200 28008
rect 26148 27965 26157 27999
rect 26157 27965 26191 27999
rect 26191 27965 26200 27999
rect 26148 27956 26200 27965
rect 30012 28024 30064 28076
rect 32956 28024 33008 28076
rect 27896 27956 27948 28008
rect 34796 28160 34848 28212
rect 34980 27999 35032 28008
rect 34980 27965 34989 27999
rect 34989 27965 35023 27999
rect 35023 27965 35032 27999
rect 34980 27956 35032 27965
rect 35072 27956 35124 28008
rect 35992 27956 36044 28008
rect 2688 27888 2740 27940
rect 4620 27888 4672 27940
rect 4160 27820 4212 27872
rect 5448 27820 5500 27872
rect 7288 27863 7340 27872
rect 7288 27829 7297 27863
rect 7297 27829 7331 27863
rect 7331 27829 7340 27863
rect 7288 27820 7340 27829
rect 7472 27863 7524 27872
rect 7472 27829 7481 27863
rect 7481 27829 7515 27863
rect 7515 27829 7524 27863
rect 7472 27820 7524 27829
rect 7564 27820 7616 27872
rect 11060 27820 11112 27872
rect 11428 27863 11480 27872
rect 11428 27829 11437 27863
rect 11437 27829 11471 27863
rect 11471 27829 11480 27863
rect 11428 27820 11480 27829
rect 17960 27820 18012 27872
rect 20628 27820 20680 27872
rect 20812 27863 20864 27872
rect 20812 27829 20821 27863
rect 20821 27829 20855 27863
rect 20855 27829 20864 27863
rect 20812 27820 20864 27829
rect 21456 27863 21508 27872
rect 21456 27829 21465 27863
rect 21465 27829 21499 27863
rect 21499 27829 21508 27863
rect 21456 27820 21508 27829
rect 21640 27820 21692 27872
rect 26332 27888 26384 27940
rect 30932 27888 30984 27940
rect 33324 27888 33376 27940
rect 24584 27820 24636 27872
rect 27252 27820 27304 27872
rect 32956 27820 33008 27872
rect 34336 27863 34388 27872
rect 34336 27829 34345 27863
rect 34345 27829 34379 27863
rect 34379 27829 34388 27863
rect 34336 27820 34388 27829
rect 34980 27820 35032 27872
rect 36360 27863 36412 27872
rect 36360 27829 36369 27863
rect 36369 27829 36403 27863
rect 36403 27829 36412 27863
rect 36360 27820 36412 27829
rect 19606 27718 19658 27770
rect 19670 27718 19722 27770
rect 19734 27718 19786 27770
rect 19798 27718 19850 27770
rect 1860 27616 1912 27668
rect 2780 27616 2832 27668
rect 4068 27616 4120 27668
rect 5448 27659 5500 27668
rect 5448 27625 5457 27659
rect 5457 27625 5491 27659
rect 5491 27625 5500 27659
rect 5448 27616 5500 27625
rect 7472 27616 7524 27668
rect 11152 27659 11204 27668
rect 2228 27548 2280 27600
rect 3884 27591 3936 27600
rect 2136 27480 2188 27532
rect 3884 27557 3893 27591
rect 3893 27557 3927 27591
rect 3927 27557 3936 27591
rect 3884 27548 3936 27557
rect 4160 27548 4212 27600
rect 4620 27548 4672 27600
rect 8116 27548 8168 27600
rect 11152 27625 11161 27659
rect 11161 27625 11195 27659
rect 11195 27625 11204 27659
rect 11152 27616 11204 27625
rect 9220 27548 9272 27600
rect 13452 27548 13504 27600
rect 14372 27616 14424 27668
rect 19340 27659 19392 27668
rect 19340 27625 19349 27659
rect 19349 27625 19383 27659
rect 19383 27625 19392 27659
rect 19340 27616 19392 27625
rect 16028 27548 16080 27600
rect 18972 27591 19024 27600
rect 18972 27557 18981 27591
rect 18981 27557 19015 27591
rect 19015 27557 19024 27591
rect 18972 27548 19024 27557
rect 21456 27616 21508 27668
rect 22468 27659 22520 27668
rect 22468 27625 22477 27659
rect 22477 27625 22511 27659
rect 22511 27625 22520 27659
rect 22468 27616 22520 27625
rect 26148 27616 26200 27668
rect 20720 27591 20772 27600
rect 20720 27557 20729 27591
rect 20729 27557 20763 27591
rect 20763 27557 20772 27591
rect 20720 27548 20772 27557
rect 20904 27548 20956 27600
rect 1768 27412 1820 27464
rect 5356 27480 5408 27532
rect 8852 27480 8904 27532
rect 11060 27480 11112 27532
rect 24768 27548 24820 27600
rect 21732 27480 21784 27532
rect 25136 27480 25188 27532
rect 25412 27480 25464 27532
rect 26148 27480 26200 27532
rect 8668 27455 8720 27464
rect 1952 27344 2004 27396
rect 3976 27344 4028 27396
rect 8668 27421 8677 27455
rect 8677 27421 8711 27455
rect 8711 27421 8720 27455
rect 8668 27412 8720 27421
rect 15568 27455 15620 27464
rect 15568 27421 15577 27455
rect 15577 27421 15611 27455
rect 15611 27421 15620 27455
rect 15568 27412 15620 27421
rect 25504 27455 25556 27464
rect 25504 27421 25513 27455
rect 25513 27421 25547 27455
rect 25547 27421 25556 27455
rect 25504 27412 25556 27421
rect 29828 27616 29880 27668
rect 30012 27616 30064 27668
rect 30472 27616 30524 27668
rect 33324 27659 33376 27668
rect 33324 27625 33333 27659
rect 33333 27625 33367 27659
rect 33367 27625 33376 27659
rect 33324 27616 33376 27625
rect 35072 27659 35124 27668
rect 35072 27625 35081 27659
rect 35081 27625 35115 27659
rect 35115 27625 35124 27659
rect 35072 27616 35124 27625
rect 32588 27591 32640 27600
rect 32588 27557 32597 27591
rect 32597 27557 32631 27591
rect 32631 27557 32640 27591
rect 32588 27548 32640 27557
rect 27252 27480 27304 27532
rect 29092 27480 29144 27532
rect 30748 27480 30800 27532
rect 32496 27523 32548 27532
rect 32496 27489 32505 27523
rect 32505 27489 32539 27523
rect 32539 27489 32548 27523
rect 32496 27480 32548 27489
rect 34152 27480 34204 27532
rect 34612 27480 34664 27532
rect 36360 27480 36412 27532
rect 26516 27455 26568 27464
rect 26516 27421 26525 27455
rect 26525 27421 26559 27455
rect 26559 27421 26568 27455
rect 26516 27412 26568 27421
rect 29552 27455 29604 27464
rect 29552 27421 29561 27455
rect 29561 27421 29595 27455
rect 29595 27421 29604 27455
rect 29552 27412 29604 27421
rect 8208 27344 8260 27396
rect 18880 27344 18932 27396
rect 20352 27344 20404 27396
rect 24952 27344 25004 27396
rect 27896 27387 27948 27396
rect 27896 27353 27905 27387
rect 27905 27353 27939 27387
rect 27939 27353 27948 27387
rect 27896 27344 27948 27353
rect 7564 27319 7616 27328
rect 7564 27285 7573 27319
rect 7573 27285 7607 27319
rect 7607 27285 7616 27319
rect 7564 27276 7616 27285
rect 16948 27319 17000 27328
rect 16948 27285 16957 27319
rect 16957 27285 16991 27319
rect 16991 27285 17000 27319
rect 16948 27276 17000 27285
rect 19984 27276 20036 27328
rect 24584 27319 24636 27328
rect 24584 27285 24593 27319
rect 24593 27285 24627 27319
rect 24627 27285 24636 27319
rect 24584 27276 24636 27285
rect 25228 27276 25280 27328
rect 30932 27319 30984 27328
rect 30932 27285 30941 27319
rect 30941 27285 30975 27319
rect 30975 27285 30984 27319
rect 30932 27276 30984 27285
rect 31576 27276 31628 27328
rect 34704 27455 34756 27464
rect 34704 27421 34713 27455
rect 34713 27421 34747 27455
rect 34747 27421 34756 27455
rect 34704 27412 34756 27421
rect 34980 27412 35032 27464
rect 32128 27319 32180 27328
rect 32128 27285 32137 27319
rect 32137 27285 32171 27319
rect 32171 27285 32180 27319
rect 32128 27276 32180 27285
rect 34244 27319 34296 27328
rect 34244 27285 34253 27319
rect 34253 27285 34287 27319
rect 34287 27285 34296 27319
rect 34244 27276 34296 27285
rect 35532 27276 35584 27328
rect 36820 27276 36872 27328
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 34966 27174 35018 27226
rect 35030 27174 35082 27226
rect 35094 27174 35146 27226
rect 35158 27174 35210 27226
rect 1768 27115 1820 27124
rect 1768 27081 1777 27115
rect 1777 27081 1811 27115
rect 1811 27081 1820 27115
rect 1768 27072 1820 27081
rect 2780 27072 2832 27124
rect 5356 27115 5408 27124
rect 4068 27004 4120 27056
rect 5356 27081 5365 27115
rect 5365 27081 5399 27115
rect 5399 27081 5408 27115
rect 5356 27072 5408 27081
rect 5724 27115 5776 27124
rect 5724 27081 5733 27115
rect 5733 27081 5767 27115
rect 5767 27081 5776 27115
rect 5724 27072 5776 27081
rect 7564 27072 7616 27124
rect 9220 27115 9272 27124
rect 9220 27081 9229 27115
rect 9229 27081 9263 27115
rect 9263 27081 9272 27115
rect 9220 27072 9272 27081
rect 10968 27072 11020 27124
rect 16028 27072 16080 27124
rect 18696 27115 18748 27124
rect 18696 27081 18705 27115
rect 18705 27081 18739 27115
rect 18739 27081 18748 27115
rect 18696 27072 18748 27081
rect 21640 27072 21692 27124
rect 25412 27072 25464 27124
rect 29092 27115 29144 27124
rect 29092 27081 29101 27115
rect 29101 27081 29135 27115
rect 29135 27081 29144 27115
rect 29092 27072 29144 27081
rect 32588 27072 32640 27124
rect 34152 27115 34204 27124
rect 34152 27081 34161 27115
rect 34161 27081 34195 27115
rect 34195 27081 34204 27115
rect 34152 27072 34204 27081
rect 34520 27072 34572 27124
rect 36360 27115 36412 27124
rect 8668 27004 8720 27056
rect 9864 27004 9916 27056
rect 11336 27004 11388 27056
rect 26516 27004 26568 27056
rect 29552 27004 29604 27056
rect 32496 27004 32548 27056
rect 6920 26979 6972 26988
rect 6920 26945 6929 26979
rect 6929 26945 6963 26979
rect 6963 26945 6972 26979
rect 6920 26936 6972 26945
rect 1492 26868 1544 26920
rect 1952 26868 2004 26920
rect 2136 26911 2188 26920
rect 2136 26877 2170 26911
rect 2170 26877 2188 26911
rect 2136 26868 2188 26877
rect 4620 26868 4672 26920
rect 9680 26868 9732 26920
rect 13452 26911 13504 26920
rect 13452 26877 13461 26911
rect 13461 26877 13495 26911
rect 13495 26877 13504 26911
rect 13452 26868 13504 26877
rect 15568 26936 15620 26988
rect 17132 26936 17184 26988
rect 21732 26979 21784 26988
rect 21732 26945 21741 26979
rect 21741 26945 21775 26979
rect 21775 26945 21784 26979
rect 21732 26936 21784 26945
rect 22284 26936 22336 26988
rect 25136 26936 25188 26988
rect 29828 26979 29880 26988
rect 13728 26911 13780 26920
rect 13728 26877 13762 26911
rect 13762 26877 13780 26911
rect 13728 26868 13780 26877
rect 18696 26868 18748 26920
rect 25228 26911 25280 26920
rect 25228 26877 25237 26911
rect 25237 26877 25271 26911
rect 25271 26877 25280 26911
rect 25228 26868 25280 26877
rect 29828 26945 29837 26979
rect 29837 26945 29871 26979
rect 29871 26945 29880 26979
rect 29828 26936 29880 26945
rect 32680 26936 32732 26988
rect 32956 26979 33008 26988
rect 32956 26945 32965 26979
rect 32965 26945 32999 26979
rect 32999 26945 33008 26979
rect 32956 26936 33008 26945
rect 36360 27081 36369 27115
rect 36369 27081 36403 27115
rect 36403 27081 36412 27115
rect 36360 27072 36412 27081
rect 34704 26936 34756 26988
rect 37004 26979 37056 26988
rect 37004 26945 37013 26979
rect 37013 26945 37047 26979
rect 37047 26945 37056 26979
rect 37004 26936 37056 26945
rect 36360 26868 36412 26920
rect 7288 26800 7340 26852
rect 8208 26800 8260 26852
rect 21916 26800 21968 26852
rect 25504 26843 25556 26852
rect 25504 26809 25538 26843
rect 25538 26809 25556 26843
rect 25504 26800 25556 26809
rect 29736 26843 29788 26852
rect 29736 26809 29745 26843
rect 29745 26809 29779 26843
rect 29779 26809 29788 26843
rect 29736 26800 29788 26809
rect 33048 26800 33100 26852
rect 34980 26800 35032 26852
rect 8852 26775 8904 26784
rect 8852 26741 8861 26775
rect 8861 26741 8895 26775
rect 8895 26741 8904 26775
rect 8852 26732 8904 26741
rect 11060 26775 11112 26784
rect 11060 26741 11069 26775
rect 11069 26741 11103 26775
rect 11103 26741 11112 26775
rect 11060 26732 11112 26741
rect 14832 26775 14884 26784
rect 14832 26741 14841 26775
rect 14841 26741 14875 26775
rect 14875 26741 14884 26775
rect 14832 26732 14884 26741
rect 17960 26732 18012 26784
rect 19340 26775 19392 26784
rect 19340 26741 19349 26775
rect 19349 26741 19383 26775
rect 19383 26741 19392 26775
rect 19340 26732 19392 26741
rect 20168 26775 20220 26784
rect 20168 26741 20177 26775
rect 20177 26741 20211 26775
rect 20211 26741 20220 26775
rect 20168 26732 20220 26741
rect 21272 26732 21324 26784
rect 22284 26775 22336 26784
rect 22284 26741 22293 26775
rect 22293 26741 22327 26775
rect 22327 26741 22336 26775
rect 22284 26732 22336 26741
rect 25320 26732 25372 26784
rect 27252 26775 27304 26784
rect 27252 26741 27261 26775
rect 27261 26741 27295 26775
rect 27295 26741 27304 26775
rect 27252 26732 27304 26741
rect 30748 26732 30800 26784
rect 31668 26732 31720 26784
rect 34428 26732 34480 26784
rect 36820 26775 36872 26784
rect 36820 26741 36829 26775
rect 36829 26741 36863 26775
rect 36863 26741 36872 26775
rect 36820 26732 36872 26741
rect 37832 26775 37884 26784
rect 37832 26741 37841 26775
rect 37841 26741 37875 26775
rect 37875 26741 37884 26775
rect 37832 26732 37884 26741
rect 19606 26630 19658 26682
rect 19670 26630 19722 26682
rect 19734 26630 19786 26682
rect 19798 26630 19850 26682
rect 2136 26528 2188 26580
rect 4620 26571 4672 26580
rect 4620 26537 4629 26571
rect 4629 26537 4663 26571
rect 4663 26537 4672 26571
rect 4620 26528 4672 26537
rect 6460 26571 6512 26580
rect 6460 26537 6469 26571
rect 6469 26537 6503 26571
rect 6503 26537 6512 26571
rect 6460 26528 6512 26537
rect 6644 26528 6696 26580
rect 6920 26528 6972 26580
rect 11060 26528 11112 26580
rect 11336 26528 11388 26580
rect 13544 26528 13596 26580
rect 14832 26528 14884 26580
rect 19156 26528 19208 26580
rect 19340 26528 19392 26580
rect 22284 26571 22336 26580
rect 22284 26537 22293 26571
rect 22293 26537 22327 26571
rect 22327 26537 22336 26571
rect 22284 26528 22336 26537
rect 25504 26528 25556 26580
rect 29368 26571 29420 26580
rect 29368 26537 29377 26571
rect 29377 26537 29411 26571
rect 29411 26537 29420 26571
rect 29368 26528 29420 26537
rect 29552 26528 29604 26580
rect 30748 26571 30800 26580
rect 30748 26537 30757 26571
rect 30757 26537 30791 26571
rect 30791 26537 30800 26571
rect 30748 26528 30800 26537
rect 30840 26528 30892 26580
rect 32680 26528 32732 26580
rect 32956 26528 33008 26580
rect 34244 26528 34296 26580
rect 34980 26571 35032 26580
rect 34980 26537 34989 26571
rect 34989 26537 35023 26571
rect 35023 26537 35032 26571
rect 34980 26528 35032 26537
rect 37004 26528 37056 26580
rect 1768 26503 1820 26512
rect 1768 26469 1802 26503
rect 1802 26469 1820 26503
rect 1768 26460 1820 26469
rect 16120 26460 16172 26512
rect 16948 26460 17000 26512
rect 19432 26460 19484 26512
rect 20168 26460 20220 26512
rect 25320 26460 25372 26512
rect 31944 26503 31996 26512
rect 31944 26469 31953 26503
rect 31953 26469 31987 26503
rect 31987 26469 31996 26503
rect 31944 26460 31996 26469
rect 1492 26435 1544 26444
rect 1492 26401 1501 26435
rect 1501 26401 1535 26435
rect 1535 26401 1544 26435
rect 1492 26392 1544 26401
rect 6736 26392 6788 26444
rect 9036 26392 9088 26444
rect 11612 26435 11664 26444
rect 11612 26401 11621 26435
rect 11621 26401 11655 26435
rect 11655 26401 11664 26435
rect 11612 26392 11664 26401
rect 13176 26435 13228 26444
rect 13176 26401 13185 26435
rect 13185 26401 13219 26435
rect 13219 26401 13228 26435
rect 13176 26392 13228 26401
rect 15568 26435 15620 26444
rect 15568 26401 15577 26435
rect 15577 26401 15611 26435
rect 15611 26401 15620 26435
rect 15568 26392 15620 26401
rect 18328 26392 18380 26444
rect 19248 26392 19300 26444
rect 6828 26256 6880 26308
rect 8116 26324 8168 26376
rect 8484 26367 8536 26376
rect 8484 26333 8493 26367
rect 8493 26333 8527 26367
rect 8527 26333 8536 26367
rect 8484 26324 8536 26333
rect 8576 26367 8628 26376
rect 8576 26333 8585 26367
rect 8585 26333 8619 26367
rect 8619 26333 8628 26367
rect 8576 26324 8628 26333
rect 11428 26324 11480 26376
rect 20076 26392 20128 26444
rect 22008 26392 22060 26444
rect 24952 26392 25004 26444
rect 26424 26392 26476 26444
rect 28908 26392 28960 26444
rect 29184 26435 29236 26444
rect 29184 26401 29193 26435
rect 29193 26401 29227 26435
rect 29227 26401 29236 26435
rect 29184 26392 29236 26401
rect 30932 26392 30984 26444
rect 31484 26392 31536 26444
rect 34060 26435 34112 26444
rect 20904 26367 20956 26376
rect 5816 26188 5868 26240
rect 9680 26256 9732 26308
rect 8576 26188 8628 26240
rect 10600 26188 10652 26240
rect 20904 26333 20913 26367
rect 20913 26333 20947 26367
rect 20947 26333 20956 26367
rect 20904 26324 20956 26333
rect 24124 26324 24176 26376
rect 24584 26324 24636 26376
rect 25320 26367 25372 26376
rect 25320 26333 25329 26367
rect 25329 26333 25363 26367
rect 25363 26333 25372 26367
rect 25320 26324 25372 26333
rect 20352 26299 20404 26308
rect 12440 26188 12492 26240
rect 16488 26188 16540 26240
rect 17960 26188 18012 26240
rect 20352 26265 20361 26299
rect 20361 26265 20395 26299
rect 20395 26265 20404 26299
rect 20352 26256 20404 26265
rect 20536 26256 20588 26308
rect 19800 26188 19852 26240
rect 26240 26299 26292 26308
rect 22928 26188 22980 26240
rect 24584 26188 24636 26240
rect 26240 26265 26249 26299
rect 26249 26265 26283 26299
rect 26283 26265 26292 26299
rect 26700 26324 26752 26376
rect 26976 26367 27028 26376
rect 26976 26333 26988 26367
rect 26988 26333 27022 26367
rect 27022 26333 27028 26367
rect 26976 26324 27028 26333
rect 30840 26367 30892 26376
rect 30840 26333 30849 26367
rect 30849 26333 30883 26367
rect 30883 26333 30892 26367
rect 30840 26324 30892 26333
rect 26240 26256 26292 26265
rect 28264 26256 28316 26308
rect 31668 26324 31720 26376
rect 34060 26401 34069 26435
rect 34069 26401 34103 26435
rect 34103 26401 34112 26435
rect 34060 26392 34112 26401
rect 34612 26392 34664 26444
rect 35532 26460 35584 26512
rect 35256 26392 35308 26444
rect 36820 26392 36872 26444
rect 25044 26188 25096 26240
rect 32312 26256 32364 26308
rect 31576 26231 31628 26240
rect 31576 26197 31585 26231
rect 31585 26197 31619 26231
rect 31619 26197 31628 26231
rect 33048 26324 33100 26376
rect 31576 26188 31628 26197
rect 35532 26188 35584 26240
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 34966 26086 35018 26138
rect 35030 26086 35082 26138
rect 35094 26086 35146 26138
rect 35158 26086 35210 26138
rect 2228 26027 2280 26036
rect 2228 25993 2237 26027
rect 2237 25993 2271 26027
rect 2271 25993 2280 26027
rect 2228 25984 2280 25993
rect 5816 26027 5868 26036
rect 5816 25993 5825 26027
rect 5825 25993 5859 26027
rect 5859 25993 5868 26027
rect 5816 25984 5868 25993
rect 8208 26027 8260 26036
rect 8208 25993 8217 26027
rect 8217 25993 8251 26027
rect 8251 25993 8260 26027
rect 8208 25984 8260 25993
rect 8484 25984 8536 26036
rect 9588 25984 9640 26036
rect 11336 26027 11388 26036
rect 11336 25993 11345 26027
rect 11345 25993 11379 26027
rect 11379 25993 11388 26027
rect 11336 25984 11388 25993
rect 6644 25848 6696 25900
rect 9864 25891 9916 25900
rect 9864 25857 9873 25891
rect 9873 25857 9907 25891
rect 9907 25857 9916 25891
rect 9864 25848 9916 25857
rect 16120 25891 16172 25900
rect 16120 25857 16129 25891
rect 16129 25857 16163 25891
rect 16163 25857 16172 25891
rect 16120 25848 16172 25857
rect 16304 25891 16356 25900
rect 16304 25857 16313 25891
rect 16313 25857 16347 25891
rect 16347 25857 16356 25891
rect 17868 25984 17920 26036
rect 18328 26027 18380 26036
rect 18328 25993 18337 26027
rect 18337 25993 18371 26027
rect 18371 25993 18380 26027
rect 18328 25984 18380 25993
rect 19156 25984 19208 26036
rect 21916 25984 21968 26036
rect 22928 26027 22980 26036
rect 17132 25959 17184 25968
rect 17132 25925 17141 25959
rect 17141 25925 17175 25959
rect 17175 25925 17184 25959
rect 17132 25916 17184 25925
rect 22928 25993 22937 26027
rect 22937 25993 22971 26027
rect 22971 25993 22980 26027
rect 22928 25984 22980 25993
rect 26332 25984 26384 26036
rect 28908 25984 28960 26036
rect 31760 26027 31812 26036
rect 31760 25993 31769 26027
rect 31769 25993 31803 26027
rect 31803 25993 31812 26027
rect 31760 25984 31812 25993
rect 34060 26027 34112 26036
rect 24308 25916 24360 25968
rect 26424 25916 26476 25968
rect 33324 25916 33376 25968
rect 34060 25993 34069 26027
rect 34069 25993 34103 26027
rect 34103 25993 34112 26027
rect 34060 25984 34112 25993
rect 34612 26027 34664 26036
rect 34612 25993 34621 26027
rect 34621 25993 34655 26027
rect 34655 25993 34664 26027
rect 34612 25984 34664 25993
rect 35716 25984 35768 26036
rect 16304 25848 16356 25857
rect 19248 25848 19300 25900
rect 19800 25891 19852 25900
rect 19800 25857 19809 25891
rect 19809 25857 19843 25891
rect 19843 25857 19852 25891
rect 19800 25848 19852 25857
rect 20536 25848 20588 25900
rect 20996 25848 21048 25900
rect 21272 25891 21324 25900
rect 21272 25857 21284 25891
rect 21284 25857 21318 25891
rect 21318 25857 21324 25891
rect 21272 25848 21324 25857
rect 9680 25823 9732 25832
rect 9680 25789 9689 25823
rect 9689 25789 9723 25823
rect 9723 25789 9732 25823
rect 9680 25780 9732 25789
rect 12440 25823 12492 25832
rect 12440 25789 12449 25823
rect 12449 25789 12483 25823
rect 12483 25789 12492 25823
rect 12440 25780 12492 25789
rect 1768 25712 1820 25764
rect 2688 25712 2740 25764
rect 6736 25712 6788 25764
rect 7104 25755 7156 25764
rect 7104 25721 7138 25755
rect 7138 25721 7156 25755
rect 7104 25712 7156 25721
rect 13544 25780 13596 25832
rect 15108 25780 15160 25832
rect 16028 25823 16080 25832
rect 16028 25789 16037 25823
rect 16037 25789 16071 25823
rect 16071 25789 16080 25823
rect 16028 25780 16080 25789
rect 16488 25780 16540 25832
rect 19984 25780 20036 25832
rect 20628 25780 20680 25832
rect 20904 25780 20956 25832
rect 23480 25823 23532 25832
rect 23480 25789 23489 25823
rect 23489 25789 23523 25823
rect 23523 25789 23532 25823
rect 24400 25823 24452 25832
rect 23480 25780 23532 25789
rect 24400 25789 24409 25823
rect 24409 25789 24443 25823
rect 24443 25789 24452 25823
rect 24400 25780 24452 25789
rect 24584 25848 24636 25900
rect 27252 25848 27304 25900
rect 27712 25891 27764 25900
rect 27712 25857 27721 25891
rect 27721 25857 27755 25891
rect 27755 25857 27764 25891
rect 27712 25848 27764 25857
rect 31484 25848 31536 25900
rect 33692 25891 33744 25900
rect 33692 25857 33701 25891
rect 33701 25857 33735 25891
rect 33735 25857 33744 25891
rect 33692 25848 33744 25857
rect 24952 25780 25004 25832
rect 27068 25780 27120 25832
rect 29184 25780 29236 25832
rect 29828 25780 29880 25832
rect 31760 25780 31812 25832
rect 33048 25780 33100 25832
rect 35532 25780 35584 25832
rect 19340 25712 19392 25764
rect 28264 25712 28316 25764
rect 30012 25755 30064 25764
rect 30012 25721 30046 25755
rect 30046 25721 30064 25755
rect 30012 25712 30064 25721
rect 35716 25712 35768 25764
rect 1952 25644 2004 25696
rect 6828 25644 6880 25696
rect 9036 25644 9088 25696
rect 9680 25644 9732 25696
rect 11612 25687 11664 25696
rect 11612 25653 11621 25687
rect 11621 25653 11655 25687
rect 11655 25653 11664 25687
rect 11612 25644 11664 25653
rect 13820 25687 13872 25696
rect 13820 25653 13829 25687
rect 13829 25653 13863 25687
rect 13863 25653 13872 25687
rect 13820 25644 13872 25653
rect 15660 25687 15712 25696
rect 15660 25653 15669 25687
rect 15669 25653 15703 25687
rect 15703 25653 15712 25687
rect 15660 25644 15712 25653
rect 20260 25687 20312 25696
rect 20260 25653 20269 25687
rect 20269 25653 20303 25687
rect 20303 25653 20312 25687
rect 20260 25644 20312 25653
rect 20720 25687 20772 25696
rect 20720 25653 20729 25687
rect 20729 25653 20763 25687
rect 20763 25653 20772 25687
rect 20720 25644 20772 25653
rect 26608 25687 26660 25696
rect 26608 25653 26617 25687
rect 26617 25653 26651 25687
rect 26651 25653 26660 25687
rect 26608 25644 26660 25653
rect 28908 25687 28960 25696
rect 28908 25653 28917 25687
rect 28917 25653 28951 25687
rect 28951 25653 28960 25687
rect 28908 25644 28960 25653
rect 31116 25687 31168 25696
rect 31116 25653 31125 25687
rect 31125 25653 31159 25687
rect 31159 25653 31168 25687
rect 31116 25644 31168 25653
rect 32864 25687 32916 25696
rect 32864 25653 32873 25687
rect 32873 25653 32907 25687
rect 32907 25653 32916 25687
rect 32864 25644 32916 25653
rect 33140 25644 33192 25696
rect 36820 25687 36872 25696
rect 36820 25653 36829 25687
rect 36829 25653 36863 25687
rect 36863 25653 36872 25687
rect 36820 25644 36872 25653
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 7104 25440 7156 25492
rect 8576 25440 8628 25492
rect 11612 25440 11664 25492
rect 13544 25483 13596 25492
rect 13544 25449 13553 25483
rect 13553 25449 13587 25483
rect 13587 25449 13596 25483
rect 13544 25440 13596 25449
rect 14556 25483 14608 25492
rect 14556 25449 14565 25483
rect 14565 25449 14599 25483
rect 14599 25449 14608 25483
rect 14556 25440 14608 25449
rect 18420 25483 18472 25492
rect 18420 25449 18429 25483
rect 18429 25449 18463 25483
rect 18463 25449 18472 25483
rect 18420 25440 18472 25449
rect 19340 25483 19392 25492
rect 19340 25449 19349 25483
rect 19349 25449 19383 25483
rect 19383 25449 19392 25483
rect 19340 25440 19392 25449
rect 20076 25483 20128 25492
rect 20076 25449 20085 25483
rect 20085 25449 20119 25483
rect 20119 25449 20128 25483
rect 20076 25440 20128 25449
rect 20812 25440 20864 25492
rect 22100 25440 22152 25492
rect 24124 25483 24176 25492
rect 24124 25449 24133 25483
rect 24133 25449 24167 25483
rect 24167 25449 24176 25483
rect 24124 25440 24176 25449
rect 24308 25440 24360 25492
rect 24584 25483 24636 25492
rect 24584 25449 24593 25483
rect 24593 25449 24627 25483
rect 24627 25449 24636 25483
rect 24584 25440 24636 25449
rect 25228 25440 25280 25492
rect 26976 25440 27028 25492
rect 6644 25304 6696 25356
rect 6828 25304 6880 25356
rect 10140 25304 10192 25356
rect 12440 25372 12492 25424
rect 16028 25372 16080 25424
rect 19892 25372 19944 25424
rect 21456 25372 21508 25424
rect 11888 25347 11940 25356
rect 11888 25313 11922 25347
rect 11922 25313 11940 25347
rect 11888 25304 11940 25313
rect 14464 25304 14516 25356
rect 18604 25304 18656 25356
rect 24768 25304 24820 25356
rect 26240 25304 26292 25356
rect 27528 25440 27580 25492
rect 27712 25483 27764 25492
rect 27712 25449 27721 25483
rect 27721 25449 27755 25483
rect 27755 25449 27764 25483
rect 27712 25440 27764 25449
rect 29736 25483 29788 25492
rect 29736 25449 29745 25483
rect 29745 25449 29779 25483
rect 29779 25449 29788 25483
rect 29736 25440 29788 25449
rect 30196 25483 30248 25492
rect 30196 25449 30205 25483
rect 30205 25449 30239 25483
rect 30239 25449 30248 25483
rect 30196 25440 30248 25449
rect 31668 25483 31720 25492
rect 31668 25449 31677 25483
rect 31677 25449 31711 25483
rect 31711 25449 31720 25483
rect 31668 25440 31720 25449
rect 31760 25483 31812 25492
rect 31760 25449 31769 25483
rect 31769 25449 31803 25483
rect 31803 25449 31812 25483
rect 31760 25440 31812 25449
rect 34244 25483 34296 25492
rect 31116 25372 31168 25424
rect 31576 25372 31628 25424
rect 34244 25449 34253 25483
rect 34253 25449 34287 25483
rect 34287 25449 34296 25483
rect 34244 25440 34296 25449
rect 34612 25440 34664 25492
rect 35256 25483 35308 25492
rect 35256 25449 35265 25483
rect 35265 25449 35299 25483
rect 35299 25449 35308 25483
rect 35256 25440 35308 25449
rect 33876 25372 33928 25424
rect 27344 25304 27396 25356
rect 28908 25304 28960 25356
rect 29828 25304 29880 25356
rect 30012 25304 30064 25356
rect 30656 25347 30708 25356
rect 30656 25313 30665 25347
rect 30665 25313 30699 25347
rect 30699 25313 30708 25347
rect 30656 25304 30708 25313
rect 31944 25347 31996 25356
rect 31944 25313 31945 25347
rect 31945 25313 31979 25347
rect 31979 25313 31996 25347
rect 31944 25304 31996 25313
rect 32496 25347 32548 25356
rect 32496 25313 32505 25347
rect 32505 25313 32539 25347
rect 32539 25313 32548 25347
rect 32496 25304 32548 25313
rect 34060 25304 34112 25356
rect 35900 25304 35952 25356
rect 10508 25279 10560 25288
rect 10508 25245 10517 25279
rect 10517 25245 10551 25279
rect 10551 25245 10560 25279
rect 10508 25236 10560 25245
rect 10600 25279 10652 25288
rect 10600 25245 10609 25279
rect 10609 25245 10643 25279
rect 10643 25245 10652 25279
rect 10600 25236 10652 25245
rect 15384 25236 15436 25288
rect 17960 25236 18012 25288
rect 20720 25236 20772 25288
rect 20904 25279 20956 25288
rect 20904 25245 20913 25279
rect 20913 25245 20947 25279
rect 20947 25245 20956 25279
rect 20904 25236 20956 25245
rect 25044 25279 25096 25288
rect 25044 25245 25053 25279
rect 25053 25245 25087 25279
rect 25087 25245 25096 25279
rect 25044 25236 25096 25245
rect 24860 25168 24912 25220
rect 26148 25236 26200 25288
rect 30840 25279 30892 25288
rect 30840 25245 30849 25279
rect 30849 25245 30883 25279
rect 30883 25245 30892 25279
rect 30840 25236 30892 25245
rect 32128 25236 32180 25288
rect 31576 25168 31628 25220
rect 34336 25279 34388 25288
rect 34336 25245 34345 25279
rect 34345 25245 34379 25279
rect 34379 25245 34388 25279
rect 34336 25236 34388 25245
rect 33692 25168 33744 25220
rect 34520 25168 34572 25220
rect 35716 25168 35768 25220
rect 36820 25236 36872 25288
rect 1952 25100 2004 25152
rect 9680 25100 9732 25152
rect 10140 25100 10192 25152
rect 12992 25143 13044 25152
rect 12992 25109 13001 25143
rect 13001 25109 13035 25143
rect 13035 25109 13044 25143
rect 12992 25100 13044 25109
rect 16580 25100 16632 25152
rect 17868 25100 17920 25152
rect 29184 25100 29236 25152
rect 32220 25100 32272 25152
rect 33140 25143 33192 25152
rect 33140 25109 33149 25143
rect 33149 25109 33183 25143
rect 33183 25109 33192 25143
rect 33140 25100 33192 25109
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 34966 24998 35018 25050
rect 35030 24998 35082 25050
rect 35094 24998 35146 25050
rect 35158 24998 35210 25050
rect 6644 24896 6696 24948
rect 6828 24896 6880 24948
rect 8576 24896 8628 24948
rect 10508 24896 10560 24948
rect 11888 24939 11940 24948
rect 11888 24905 11897 24939
rect 11897 24905 11931 24939
rect 11931 24905 11940 24939
rect 11888 24896 11940 24905
rect 6920 24735 6972 24744
rect 6920 24701 6929 24735
rect 6929 24701 6963 24735
rect 6963 24701 6972 24735
rect 6920 24692 6972 24701
rect 9036 24692 9088 24744
rect 9864 24735 9916 24744
rect 9864 24701 9873 24735
rect 9873 24701 9907 24735
rect 9907 24701 9916 24735
rect 9864 24692 9916 24701
rect 10140 24735 10192 24744
rect 10140 24701 10174 24735
rect 10174 24701 10192 24735
rect 10140 24692 10192 24701
rect 10508 24692 10560 24744
rect 12716 24896 12768 24948
rect 15108 24939 15160 24948
rect 15108 24905 15117 24939
rect 15117 24905 15151 24939
rect 15151 24905 15160 24939
rect 15108 24896 15160 24905
rect 18420 24896 18472 24948
rect 20260 24896 20312 24948
rect 21272 24896 21324 24948
rect 21456 24939 21508 24948
rect 21456 24905 21465 24939
rect 21465 24905 21499 24939
rect 21499 24905 21508 24939
rect 21456 24896 21508 24905
rect 27344 24939 27396 24948
rect 27344 24905 27353 24939
rect 27353 24905 27387 24939
rect 27387 24905 27396 24939
rect 27344 24896 27396 24905
rect 30656 24896 30708 24948
rect 31944 24896 31996 24948
rect 32496 24896 32548 24948
rect 34060 24896 34112 24948
rect 34244 24939 34296 24948
rect 34244 24905 34253 24939
rect 34253 24905 34287 24939
rect 34287 24905 34296 24939
rect 34244 24896 34296 24905
rect 36820 24896 36872 24948
rect 25044 24828 25096 24880
rect 24768 24760 24820 24812
rect 32680 24803 32732 24812
rect 32680 24769 32689 24803
rect 32689 24769 32723 24803
rect 32723 24769 32732 24803
rect 32680 24760 32732 24769
rect 34612 24760 34664 24812
rect 12716 24735 12768 24744
rect 12716 24701 12750 24735
rect 12750 24701 12768 24735
rect 12716 24692 12768 24701
rect 12992 24692 13044 24744
rect 15384 24692 15436 24744
rect 18972 24735 19024 24744
rect 11244 24599 11296 24608
rect 11244 24565 11253 24599
rect 11253 24565 11287 24599
rect 11287 24565 11296 24599
rect 11244 24556 11296 24565
rect 12440 24556 12492 24608
rect 15936 24624 15988 24676
rect 18972 24701 18981 24735
rect 18981 24701 19015 24735
rect 19015 24701 19024 24735
rect 18972 24692 19024 24701
rect 19892 24692 19944 24744
rect 20904 24692 20956 24744
rect 24860 24692 24912 24744
rect 25136 24692 25188 24744
rect 25320 24735 25372 24744
rect 25320 24701 25354 24735
rect 25354 24701 25372 24735
rect 25320 24692 25372 24701
rect 29736 24692 29788 24744
rect 20260 24624 20312 24676
rect 30932 24624 30984 24676
rect 33784 24692 33836 24744
rect 34428 24692 34480 24744
rect 13820 24599 13872 24608
rect 13820 24565 13829 24599
rect 13829 24565 13863 24599
rect 13863 24565 13872 24599
rect 13820 24556 13872 24565
rect 14464 24599 14516 24608
rect 14464 24565 14473 24599
rect 14473 24565 14507 24599
rect 14507 24565 14516 24599
rect 14464 24556 14516 24565
rect 16672 24599 16724 24608
rect 16672 24565 16681 24599
rect 16681 24565 16715 24599
rect 16715 24565 16724 24599
rect 16672 24556 16724 24565
rect 17776 24599 17828 24608
rect 17776 24565 17785 24599
rect 17785 24565 17819 24599
rect 17819 24565 17828 24599
rect 17776 24556 17828 24565
rect 18604 24599 18656 24608
rect 18604 24565 18613 24599
rect 18613 24565 18647 24599
rect 18647 24565 18656 24599
rect 18604 24556 18656 24565
rect 22376 24599 22428 24608
rect 22376 24565 22385 24599
rect 22385 24565 22419 24599
rect 22419 24565 22428 24599
rect 22376 24556 22428 24565
rect 26148 24556 26200 24608
rect 26424 24599 26476 24608
rect 26424 24565 26433 24599
rect 26433 24565 26467 24599
rect 26467 24565 26476 24599
rect 26424 24556 26476 24565
rect 30840 24556 30892 24608
rect 31116 24556 31168 24608
rect 35532 24624 35584 24676
rect 32128 24556 32180 24608
rect 35164 24556 35216 24608
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 6828 24395 6880 24404
rect 6828 24361 6837 24395
rect 6837 24361 6871 24395
rect 6871 24361 6880 24395
rect 6828 24352 6880 24361
rect 8484 24395 8536 24404
rect 8484 24361 8493 24395
rect 8493 24361 8527 24395
rect 8527 24361 8536 24395
rect 8484 24352 8536 24361
rect 15476 24395 15528 24404
rect 15476 24361 15485 24395
rect 15485 24361 15519 24395
rect 15519 24361 15528 24395
rect 15476 24352 15528 24361
rect 15936 24395 15988 24404
rect 15936 24361 15945 24395
rect 15945 24361 15979 24395
rect 15979 24361 15988 24395
rect 15936 24352 15988 24361
rect 16488 24352 16540 24404
rect 20812 24352 20864 24404
rect 24768 24352 24820 24404
rect 25136 24352 25188 24404
rect 26240 24395 26292 24404
rect 26240 24361 26249 24395
rect 26249 24361 26283 24395
rect 26283 24361 26292 24395
rect 26240 24352 26292 24361
rect 30932 24395 30984 24404
rect 30932 24361 30941 24395
rect 30941 24361 30975 24395
rect 30975 24361 30984 24395
rect 30932 24352 30984 24361
rect 31944 24395 31996 24404
rect 31944 24361 31953 24395
rect 31953 24361 31987 24395
rect 31987 24361 31996 24395
rect 31944 24352 31996 24361
rect 32128 24395 32180 24404
rect 32128 24361 32137 24395
rect 32137 24361 32171 24395
rect 32171 24361 32180 24395
rect 32128 24352 32180 24361
rect 33784 24395 33836 24404
rect 33784 24361 33793 24395
rect 33793 24361 33827 24395
rect 33827 24361 33836 24395
rect 33784 24352 33836 24361
rect 34336 24352 34388 24404
rect 10600 24284 10652 24336
rect 11244 24284 11296 24336
rect 12440 24284 12492 24336
rect 14556 24284 14608 24336
rect 15384 24284 15436 24336
rect 20720 24284 20772 24336
rect 25320 24284 25372 24336
rect 32036 24284 32088 24336
rect 35900 24327 35952 24336
rect 35900 24293 35909 24327
rect 35909 24293 35943 24327
rect 35943 24293 35952 24327
rect 35900 24284 35952 24293
rect 7196 24216 7248 24268
rect 7748 24216 7800 24268
rect 9864 24216 9916 24268
rect 10416 24216 10468 24268
rect 16672 24216 16724 24268
rect 17132 24216 17184 24268
rect 17868 24216 17920 24268
rect 18512 24216 18564 24268
rect 18972 24259 19024 24268
rect 18972 24225 18981 24259
rect 18981 24225 19015 24259
rect 19015 24225 19024 24259
rect 18972 24216 19024 24225
rect 20904 24216 20956 24268
rect 22376 24216 22428 24268
rect 29092 24216 29144 24268
rect 31116 24216 31168 24268
rect 32128 24216 32180 24268
rect 34612 24216 34664 24268
rect 36912 24216 36964 24268
rect 16304 24148 16356 24200
rect 18788 24148 18840 24200
rect 12992 24080 13044 24132
rect 18236 24080 18288 24132
rect 21088 24148 21140 24200
rect 32588 24191 32640 24200
rect 19340 24080 19392 24132
rect 20260 24080 20312 24132
rect 11152 24055 11204 24064
rect 11152 24021 11161 24055
rect 11161 24021 11195 24055
rect 11195 24021 11204 24055
rect 11152 24012 11204 24021
rect 17224 24055 17276 24064
rect 17224 24021 17233 24055
rect 17233 24021 17267 24055
rect 17267 24021 17276 24055
rect 17224 24012 17276 24021
rect 18420 24055 18472 24064
rect 18420 24021 18429 24055
rect 18429 24021 18463 24055
rect 18463 24021 18472 24055
rect 18420 24012 18472 24021
rect 18604 24055 18656 24064
rect 18604 24021 18613 24055
rect 18613 24021 18647 24055
rect 18647 24021 18656 24055
rect 18604 24012 18656 24021
rect 19524 24012 19576 24064
rect 19800 24012 19852 24064
rect 32588 24157 32597 24191
rect 32597 24157 32631 24191
rect 32631 24157 32640 24191
rect 32588 24148 32640 24157
rect 32680 24191 32732 24200
rect 32680 24157 32689 24191
rect 32689 24157 32723 24191
rect 32723 24157 32732 24191
rect 32680 24148 32732 24157
rect 34428 24148 34480 24200
rect 35164 24191 35216 24200
rect 35164 24157 35173 24191
rect 35173 24157 35207 24191
rect 35207 24157 35216 24191
rect 35164 24148 35216 24157
rect 33324 24080 33376 24132
rect 35716 24080 35768 24132
rect 29736 24012 29788 24064
rect 34520 24055 34572 24064
rect 34520 24021 34529 24055
rect 34529 24021 34563 24055
rect 34563 24021 34572 24055
rect 34520 24012 34572 24021
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 34966 23910 35018 23962
rect 35030 23910 35082 23962
rect 35094 23910 35146 23962
rect 35158 23910 35210 23962
rect 7196 23851 7248 23860
rect 7196 23817 7205 23851
rect 7205 23817 7239 23851
rect 7239 23817 7248 23851
rect 7196 23808 7248 23817
rect 9036 23851 9088 23860
rect 9036 23817 9045 23851
rect 9045 23817 9079 23851
rect 9079 23817 9088 23851
rect 9036 23808 9088 23817
rect 9680 23808 9732 23860
rect 10232 23672 10284 23724
rect 10600 23715 10652 23724
rect 10600 23681 10609 23715
rect 10609 23681 10643 23715
rect 10643 23681 10652 23715
rect 10600 23672 10652 23681
rect 10692 23715 10744 23724
rect 10692 23681 10701 23715
rect 10701 23681 10735 23715
rect 10735 23681 10744 23715
rect 16672 23808 16724 23860
rect 17132 23851 17184 23860
rect 17132 23817 17141 23851
rect 17141 23817 17175 23851
rect 17175 23817 17184 23851
rect 17132 23808 17184 23817
rect 19064 23851 19116 23860
rect 19064 23817 19073 23851
rect 19073 23817 19107 23851
rect 19107 23817 19116 23851
rect 19064 23808 19116 23817
rect 20260 23851 20312 23860
rect 20260 23817 20269 23851
rect 20269 23817 20303 23851
rect 20303 23817 20312 23851
rect 20260 23808 20312 23817
rect 20720 23851 20772 23860
rect 20720 23817 20729 23851
rect 20729 23817 20763 23851
rect 20763 23817 20772 23851
rect 20720 23808 20772 23817
rect 22008 23808 22060 23860
rect 29092 23851 29144 23860
rect 29092 23817 29101 23851
rect 29101 23817 29135 23851
rect 29135 23817 29144 23851
rect 29092 23808 29144 23817
rect 31116 23851 31168 23860
rect 31116 23817 31125 23851
rect 31125 23817 31159 23851
rect 31159 23817 31168 23851
rect 31116 23808 31168 23817
rect 32128 23851 32180 23860
rect 32128 23817 32137 23851
rect 32137 23817 32171 23851
rect 32171 23817 32180 23851
rect 32128 23808 32180 23817
rect 33048 23808 33100 23860
rect 34244 23808 34296 23860
rect 34612 23851 34664 23860
rect 34612 23817 34621 23851
rect 34621 23817 34655 23851
rect 34655 23817 34664 23851
rect 34612 23808 34664 23817
rect 36912 23851 36964 23860
rect 36912 23817 36921 23851
rect 36921 23817 36955 23851
rect 36955 23817 36964 23851
rect 36912 23808 36964 23817
rect 32680 23740 32732 23792
rect 10692 23672 10744 23681
rect 8484 23604 8536 23656
rect 10508 23647 10560 23656
rect 10508 23613 10517 23647
rect 10517 23613 10551 23647
rect 10551 23613 10560 23647
rect 11152 23647 11204 23656
rect 10508 23604 10560 23613
rect 11152 23613 11161 23647
rect 11161 23613 11195 23647
rect 11195 23613 11204 23647
rect 11152 23604 11204 23613
rect 12992 23604 13044 23656
rect 14556 23647 14608 23656
rect 14556 23613 14565 23647
rect 14565 23613 14599 23647
rect 14599 23613 14608 23647
rect 14556 23604 14608 23613
rect 19432 23672 19484 23724
rect 19800 23715 19852 23724
rect 19800 23681 19809 23715
rect 19809 23681 19843 23715
rect 19843 23681 19852 23715
rect 19800 23672 19852 23681
rect 18420 23604 18472 23656
rect 19064 23604 19116 23656
rect 19524 23647 19576 23656
rect 19524 23613 19533 23647
rect 19533 23613 19567 23647
rect 19567 23613 19576 23647
rect 19524 23604 19576 23613
rect 29736 23647 29788 23656
rect 29736 23613 29745 23647
rect 29745 23613 29779 23647
rect 29779 23613 29788 23647
rect 29736 23604 29788 23613
rect 32312 23604 32364 23656
rect 34336 23740 34388 23792
rect 36544 23604 36596 23656
rect 7748 23536 7800 23588
rect 21548 23536 21600 23588
rect 30932 23536 30984 23588
rect 32588 23536 32640 23588
rect 34336 23536 34388 23588
rect 35256 23536 35308 23588
rect 35900 23536 35952 23588
rect 10416 23468 10468 23520
rect 12348 23468 12400 23520
rect 15200 23468 15252 23520
rect 16580 23468 16632 23520
rect 18512 23468 18564 23520
rect 18696 23511 18748 23520
rect 18696 23477 18705 23511
rect 18705 23477 18739 23511
rect 18739 23477 18748 23511
rect 18696 23468 18748 23477
rect 19156 23511 19208 23520
rect 19156 23477 19165 23511
rect 19165 23477 19199 23511
rect 19199 23477 19208 23511
rect 19156 23468 19208 23477
rect 19340 23468 19392 23520
rect 28724 23511 28776 23520
rect 28724 23477 28733 23511
rect 28733 23477 28767 23511
rect 28767 23477 28776 23511
rect 28724 23468 28776 23477
rect 31760 23468 31812 23520
rect 34428 23468 34480 23520
rect 36268 23511 36320 23520
rect 36268 23477 36277 23511
rect 36277 23477 36311 23511
rect 36311 23477 36320 23511
rect 36268 23468 36320 23477
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 7748 23307 7800 23316
rect 7748 23273 7757 23307
rect 7757 23273 7791 23307
rect 7791 23273 7800 23307
rect 7748 23264 7800 23273
rect 10232 23307 10284 23316
rect 10232 23273 10241 23307
rect 10241 23273 10275 23307
rect 10275 23273 10284 23307
rect 10232 23264 10284 23273
rect 10416 23307 10468 23316
rect 10416 23273 10425 23307
rect 10425 23273 10459 23307
rect 10459 23273 10468 23307
rect 10416 23264 10468 23273
rect 10692 23264 10744 23316
rect 14096 23307 14148 23316
rect 14096 23273 14105 23307
rect 14105 23273 14139 23307
rect 14139 23273 14148 23307
rect 14096 23264 14148 23273
rect 15108 23264 15160 23316
rect 16396 23264 16448 23316
rect 17224 23264 17276 23316
rect 18236 23307 18288 23316
rect 18236 23273 18245 23307
rect 18245 23273 18279 23307
rect 18279 23273 18288 23307
rect 18236 23264 18288 23273
rect 18788 23264 18840 23316
rect 20260 23264 20312 23316
rect 21088 23307 21140 23316
rect 21088 23273 21097 23307
rect 21097 23273 21131 23307
rect 21131 23273 21140 23307
rect 21088 23264 21140 23273
rect 25136 23307 25188 23316
rect 25136 23273 25145 23307
rect 25145 23273 25179 23307
rect 25179 23273 25188 23307
rect 25136 23264 25188 23273
rect 30932 23307 30984 23316
rect 30932 23273 30941 23307
rect 30941 23273 30975 23307
rect 30975 23273 30984 23307
rect 30932 23264 30984 23273
rect 32128 23264 32180 23316
rect 32864 23264 32916 23316
rect 34244 23264 34296 23316
rect 34428 23307 34480 23316
rect 34428 23273 34437 23307
rect 34437 23273 34471 23307
rect 34471 23273 34480 23307
rect 34428 23264 34480 23273
rect 34520 23264 34572 23316
rect 35900 23307 35952 23316
rect 35900 23273 35909 23307
rect 35909 23273 35943 23307
rect 35943 23273 35952 23307
rect 35900 23264 35952 23273
rect 15936 23239 15988 23248
rect 15936 23205 15945 23239
rect 15945 23205 15979 23239
rect 15979 23205 15988 23239
rect 15936 23196 15988 23205
rect 16304 23239 16356 23248
rect 16304 23205 16313 23239
rect 16313 23205 16347 23239
rect 16347 23205 16356 23239
rect 16304 23196 16356 23205
rect 19432 23196 19484 23248
rect 27160 23196 27212 23248
rect 10600 23171 10652 23180
rect 10600 23137 10609 23171
rect 10609 23137 10643 23171
rect 10643 23137 10652 23171
rect 10600 23128 10652 23137
rect 14004 23171 14056 23180
rect 14004 23137 14013 23171
rect 14013 23137 14047 23171
rect 14047 23137 14056 23171
rect 14004 23128 14056 23137
rect 15292 23171 15344 23180
rect 15292 23137 15301 23171
rect 15301 23137 15335 23171
rect 15335 23137 15344 23171
rect 15292 23128 15344 23137
rect 13544 23103 13596 23112
rect 13544 23069 13553 23103
rect 13553 23069 13587 23103
rect 13587 23069 13596 23103
rect 13544 23060 13596 23069
rect 18144 23128 18196 23180
rect 18696 23128 18748 23180
rect 19156 23128 19208 23180
rect 19892 23128 19944 23180
rect 26792 23128 26844 23180
rect 29736 23196 29788 23248
rect 34336 23196 34388 23248
rect 29644 23128 29696 23180
rect 31024 23128 31076 23180
rect 32220 23128 32272 23180
rect 33324 23128 33376 23180
rect 34704 23128 34756 23180
rect 17040 23103 17092 23112
rect 17040 23069 17049 23103
rect 17049 23069 17083 23103
rect 17083 23069 17092 23103
rect 17040 23060 17092 23069
rect 17408 23060 17460 23112
rect 35256 23060 35308 23112
rect 36268 23060 36320 23112
rect 18788 22992 18840 23044
rect 13636 22967 13688 22976
rect 13636 22933 13645 22967
rect 13645 22933 13679 22967
rect 13679 22933 13688 22967
rect 13636 22924 13688 22933
rect 21548 22967 21600 22976
rect 21548 22933 21557 22967
rect 21557 22933 21591 22967
rect 21591 22933 21600 22967
rect 21548 22924 21600 22933
rect 26148 22924 26200 22976
rect 34520 22967 34572 22976
rect 34520 22933 34529 22967
rect 34529 22933 34563 22967
rect 34563 22933 34572 22967
rect 34520 22924 34572 22933
rect 35532 22967 35584 22976
rect 35532 22933 35541 22967
rect 35541 22933 35575 22967
rect 35575 22933 35584 22967
rect 35532 22924 35584 22933
rect 36544 22967 36596 22976
rect 36544 22933 36553 22967
rect 36553 22933 36587 22967
rect 36587 22933 36596 22967
rect 36544 22924 36596 22933
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 34966 22822 35018 22874
rect 35030 22822 35082 22874
rect 35094 22822 35146 22874
rect 35158 22822 35210 22874
rect 6920 22720 6972 22772
rect 8576 22720 8628 22772
rect 10600 22720 10652 22772
rect 13176 22720 13228 22772
rect 14004 22720 14056 22772
rect 17224 22720 17276 22772
rect 19064 22720 19116 22772
rect 19432 22720 19484 22772
rect 27160 22763 27212 22772
rect 27160 22729 27169 22763
rect 27169 22729 27203 22763
rect 27203 22729 27212 22763
rect 27160 22720 27212 22729
rect 31024 22763 31076 22772
rect 31024 22729 31033 22763
rect 31033 22729 31067 22763
rect 31067 22729 31076 22763
rect 31024 22720 31076 22729
rect 31668 22720 31720 22772
rect 32220 22720 32272 22772
rect 32956 22763 33008 22772
rect 32956 22729 32965 22763
rect 32965 22729 32999 22763
rect 32999 22729 33008 22763
rect 32956 22720 33008 22729
rect 33324 22720 33376 22772
rect 34704 22720 34756 22772
rect 35440 22720 35492 22772
rect 36268 22720 36320 22772
rect 16488 22652 16540 22704
rect 18420 22652 18472 22704
rect 17040 22627 17092 22636
rect 17040 22593 17049 22627
rect 17049 22593 17083 22627
rect 17083 22593 17092 22627
rect 17040 22584 17092 22593
rect 17408 22584 17460 22636
rect 13912 22516 13964 22568
rect 14648 22516 14700 22568
rect 18788 22584 18840 22636
rect 26792 22652 26844 22704
rect 25136 22627 25188 22636
rect 19156 22559 19208 22568
rect 19156 22525 19165 22559
rect 19165 22525 19199 22559
rect 19199 22525 19208 22559
rect 19156 22516 19208 22525
rect 25136 22593 25145 22627
rect 25145 22593 25179 22627
rect 25179 22593 25188 22627
rect 25136 22584 25188 22593
rect 36084 22584 36136 22636
rect 19984 22516 20036 22568
rect 28724 22559 28776 22568
rect 28724 22525 28733 22559
rect 28733 22525 28767 22559
rect 28767 22525 28776 22559
rect 28724 22516 28776 22525
rect 29736 22516 29788 22568
rect 32956 22516 33008 22568
rect 33876 22516 33928 22568
rect 35532 22516 35584 22568
rect 35900 22516 35952 22568
rect 14096 22491 14148 22500
rect 14096 22457 14130 22491
rect 14130 22457 14148 22491
rect 14096 22448 14148 22457
rect 17040 22448 17092 22500
rect 25320 22448 25372 22500
rect 29552 22491 29604 22500
rect 29552 22457 29561 22491
rect 29561 22457 29595 22491
rect 29595 22457 29604 22491
rect 29552 22448 29604 22457
rect 16856 22423 16908 22432
rect 16856 22389 16865 22423
rect 16865 22389 16899 22423
rect 16899 22389 16908 22423
rect 16856 22380 16908 22389
rect 22376 22423 22428 22432
rect 22376 22389 22385 22423
rect 22385 22389 22419 22423
rect 22419 22389 22428 22423
rect 22376 22380 22428 22389
rect 32128 22423 32180 22432
rect 32128 22389 32137 22423
rect 32137 22389 32171 22423
rect 32171 22389 32180 22423
rect 32128 22380 32180 22389
rect 34428 22380 34480 22432
rect 35164 22380 35216 22432
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 13544 22219 13596 22228
rect 13544 22185 13553 22219
rect 13553 22185 13587 22219
rect 13587 22185 13596 22219
rect 13544 22176 13596 22185
rect 14096 22176 14148 22228
rect 14648 22219 14700 22228
rect 14648 22185 14657 22219
rect 14657 22185 14691 22219
rect 14691 22185 14700 22219
rect 14648 22176 14700 22185
rect 15292 22219 15344 22228
rect 15292 22185 15301 22219
rect 15301 22185 15335 22219
rect 15335 22185 15344 22219
rect 15292 22176 15344 22185
rect 16396 22219 16448 22228
rect 16396 22185 16405 22219
rect 16405 22185 16439 22219
rect 16439 22185 16448 22219
rect 16396 22176 16448 22185
rect 17040 22219 17092 22228
rect 17040 22185 17049 22219
rect 17049 22185 17083 22219
rect 17083 22185 17092 22219
rect 17040 22176 17092 22185
rect 17408 22219 17460 22228
rect 17408 22185 17417 22219
rect 17417 22185 17451 22219
rect 17451 22185 17460 22219
rect 17408 22176 17460 22185
rect 18144 22219 18196 22228
rect 18144 22185 18153 22219
rect 18153 22185 18187 22219
rect 18187 22185 18196 22219
rect 18144 22176 18196 22185
rect 29644 22219 29696 22228
rect 29644 22185 29653 22219
rect 29653 22185 29687 22219
rect 29687 22185 29696 22219
rect 29644 22176 29696 22185
rect 33876 22176 33928 22228
rect 34612 22176 34664 22228
rect 12256 22040 12308 22092
rect 14648 22040 14700 22092
rect 16856 22083 16908 22092
rect 12440 21972 12492 22024
rect 13544 21972 13596 22024
rect 15016 21972 15068 22024
rect 12992 21947 13044 21956
rect 12992 21913 13001 21947
rect 13001 21913 13035 21947
rect 13035 21913 13044 21947
rect 12992 21904 13044 21913
rect 16856 22049 16865 22083
rect 16865 22049 16899 22083
rect 16899 22049 16908 22083
rect 16856 22040 16908 22049
rect 18604 22083 18656 22092
rect 18604 22049 18613 22083
rect 18613 22049 18647 22083
rect 18647 22049 18656 22083
rect 18604 22040 18656 22049
rect 19432 22108 19484 22160
rect 26792 22151 26844 22160
rect 26792 22117 26826 22151
rect 26826 22117 26844 22151
rect 26792 22108 26844 22117
rect 34336 22108 34388 22160
rect 35164 22176 35216 22228
rect 35256 22108 35308 22160
rect 35624 22108 35676 22160
rect 35808 22108 35860 22160
rect 36176 22108 36228 22160
rect 22284 22040 22336 22092
rect 23112 22040 23164 22092
rect 24032 22040 24084 22092
rect 35716 22040 35768 22092
rect 15752 22015 15804 22024
rect 15752 21981 15761 22015
rect 15761 21981 15795 22015
rect 15795 21981 15804 22015
rect 15752 21972 15804 21981
rect 16028 21972 16080 22024
rect 22376 21972 22428 22024
rect 23020 22015 23072 22024
rect 23020 21981 23029 22015
rect 23029 21981 23063 22015
rect 23063 21981 23072 22015
rect 23020 21972 23072 21981
rect 26516 22015 26568 22024
rect 15844 21904 15896 21956
rect 19248 21904 19300 21956
rect 19156 21836 19208 21888
rect 21088 21836 21140 21888
rect 22284 21879 22336 21888
rect 22284 21845 22293 21879
rect 22293 21845 22327 21879
rect 22327 21845 22336 21879
rect 22284 21836 22336 21845
rect 23480 21836 23532 21888
rect 23664 21836 23716 21888
rect 26516 21981 26525 22015
rect 26525 21981 26559 22015
rect 26559 21981 26568 22015
rect 26516 21972 26568 21981
rect 32128 21972 32180 22024
rect 34612 22015 34664 22024
rect 34612 21981 34621 22015
rect 34621 21981 34655 22015
rect 34655 21981 34664 22015
rect 34612 21972 34664 21981
rect 25136 21836 25188 21888
rect 25320 21879 25372 21888
rect 25320 21845 25329 21879
rect 25329 21845 25363 21879
rect 25363 21845 25372 21879
rect 25320 21836 25372 21845
rect 27160 21836 27212 21888
rect 29736 21836 29788 21888
rect 30564 21836 30616 21888
rect 35348 21836 35400 21888
rect 36176 21904 36228 21956
rect 35992 21879 36044 21888
rect 35992 21845 36001 21879
rect 36001 21845 36035 21879
rect 36035 21845 36044 21879
rect 35992 21836 36044 21845
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 34966 21734 35018 21786
rect 35030 21734 35082 21786
rect 35094 21734 35146 21786
rect 35158 21734 35210 21786
rect 8576 21675 8628 21684
rect 8576 21641 8585 21675
rect 8585 21641 8619 21675
rect 8619 21641 8628 21675
rect 8576 21632 8628 21641
rect 13176 21675 13228 21684
rect 13176 21641 13185 21675
rect 13185 21641 13219 21675
rect 13219 21641 13228 21675
rect 13176 21632 13228 21641
rect 14648 21675 14700 21684
rect 14648 21641 14657 21675
rect 14657 21641 14691 21675
rect 14691 21641 14700 21675
rect 14648 21632 14700 21641
rect 15752 21632 15804 21684
rect 15844 21632 15896 21684
rect 16856 21632 16908 21684
rect 19984 21675 20036 21684
rect 19984 21641 19993 21675
rect 19993 21641 20027 21675
rect 20027 21641 20036 21675
rect 19984 21632 20036 21641
rect 22284 21632 22336 21684
rect 12440 21428 12492 21480
rect 17132 21496 17184 21548
rect 17776 21496 17828 21548
rect 26148 21632 26200 21684
rect 26792 21675 26844 21684
rect 26792 21641 26801 21675
rect 26801 21641 26835 21675
rect 26835 21641 26844 21675
rect 26792 21632 26844 21641
rect 27896 21675 27948 21684
rect 27896 21641 27905 21675
rect 27905 21641 27939 21675
rect 27939 21641 27948 21675
rect 27896 21632 27948 21641
rect 29552 21632 29604 21684
rect 35256 21632 35308 21684
rect 35808 21632 35860 21684
rect 36084 21632 36136 21684
rect 26332 21564 26384 21616
rect 19156 21428 19208 21480
rect 21088 21471 21140 21480
rect 21088 21437 21097 21471
rect 21097 21437 21131 21471
rect 21131 21437 21140 21471
rect 21088 21428 21140 21437
rect 23664 21471 23716 21480
rect 23664 21437 23673 21471
rect 23673 21437 23707 21471
rect 23707 21437 23716 21471
rect 23664 21428 23716 21437
rect 26148 21471 26200 21480
rect 26148 21437 26157 21471
rect 26157 21437 26191 21471
rect 26191 21437 26200 21471
rect 26148 21428 26200 21437
rect 27896 21428 27948 21480
rect 30564 21428 30616 21480
rect 34612 21428 34664 21480
rect 34888 21471 34940 21480
rect 34888 21437 34897 21471
rect 34897 21437 34931 21471
rect 34931 21437 34940 21471
rect 34888 21428 34940 21437
rect 12992 21360 13044 21412
rect 14648 21360 14700 21412
rect 9128 21335 9180 21344
rect 9128 21301 9137 21335
rect 9137 21301 9171 21335
rect 9171 21301 9180 21335
rect 9128 21292 9180 21301
rect 12256 21335 12308 21344
rect 12256 21301 12265 21335
rect 12265 21301 12299 21335
rect 12299 21301 12308 21335
rect 12256 21292 12308 21301
rect 14096 21292 14148 21344
rect 16764 21335 16816 21344
rect 16764 21301 16773 21335
rect 16773 21301 16807 21335
rect 16807 21301 16816 21335
rect 16764 21292 16816 21301
rect 16856 21335 16908 21344
rect 16856 21301 16865 21335
rect 16865 21301 16899 21335
rect 16899 21301 16908 21335
rect 16856 21292 16908 21301
rect 17960 21292 18012 21344
rect 19248 21360 19300 21412
rect 25136 21360 25188 21412
rect 26516 21360 26568 21412
rect 27620 21360 27672 21412
rect 30196 21360 30248 21412
rect 33324 21360 33376 21412
rect 35992 21428 36044 21480
rect 23112 21335 23164 21344
rect 23112 21301 23121 21335
rect 23121 21301 23155 21335
rect 23155 21301 23164 21335
rect 23112 21292 23164 21301
rect 24032 21292 24084 21344
rect 24952 21292 25004 21344
rect 26240 21292 26292 21344
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 13728 21088 13780 21140
rect 14096 21131 14148 21140
rect 14096 21097 14105 21131
rect 14105 21097 14139 21131
rect 14139 21097 14148 21131
rect 14096 21088 14148 21097
rect 15292 21131 15344 21140
rect 15292 21097 15301 21131
rect 15301 21097 15335 21131
rect 15335 21097 15344 21131
rect 15292 21088 15344 21097
rect 16764 21131 16816 21140
rect 16764 21097 16773 21131
rect 16773 21097 16807 21131
rect 16807 21097 16816 21131
rect 16764 21088 16816 21097
rect 18604 21088 18656 21140
rect 19340 21088 19392 21140
rect 21088 21131 21140 21140
rect 21088 21097 21097 21131
rect 21097 21097 21131 21131
rect 21131 21097 21140 21131
rect 21088 21088 21140 21097
rect 23112 21131 23164 21140
rect 23112 21097 23121 21131
rect 23121 21097 23155 21131
rect 23155 21097 23164 21131
rect 23112 21088 23164 21097
rect 24032 21131 24084 21140
rect 24032 21097 24041 21131
rect 24041 21097 24075 21131
rect 24075 21097 24084 21131
rect 24032 21088 24084 21097
rect 25504 21131 25556 21140
rect 25504 21097 25513 21131
rect 25513 21097 25547 21131
rect 25547 21097 25556 21131
rect 25504 21088 25556 21097
rect 26608 21088 26660 21140
rect 30564 21088 30616 21140
rect 32128 21088 32180 21140
rect 33324 21131 33376 21140
rect 33324 21097 33333 21131
rect 33333 21097 33367 21131
rect 33367 21097 33376 21131
rect 33324 21088 33376 21097
rect 35900 21088 35952 21140
rect 12992 21063 13044 21072
rect 12992 21029 13026 21063
rect 13026 21029 13044 21063
rect 12992 21020 13044 21029
rect 17132 21063 17184 21072
rect 17132 21029 17141 21063
rect 17141 21029 17175 21063
rect 17175 21029 17184 21063
rect 17132 21020 17184 21029
rect 12440 20952 12492 21004
rect 16488 20952 16540 21004
rect 15752 20927 15804 20936
rect 15752 20893 15761 20927
rect 15761 20893 15795 20927
rect 15795 20893 15804 20927
rect 15752 20884 15804 20893
rect 16028 20884 16080 20936
rect 17960 20952 18012 21004
rect 18328 20952 18380 21004
rect 19156 20952 19208 21004
rect 19524 20952 19576 21004
rect 21732 20995 21784 21004
rect 21732 20961 21741 20995
rect 21741 20961 21775 20995
rect 21775 20961 21784 20995
rect 21732 20952 21784 20961
rect 22008 20995 22060 21004
rect 22008 20961 22042 20995
rect 22042 20961 22060 20995
rect 22008 20952 22060 20961
rect 24216 20995 24268 21004
rect 24216 20961 24225 20995
rect 24225 20961 24259 20995
rect 24259 20961 24268 20995
rect 24216 20952 24268 20961
rect 28080 20995 28132 21004
rect 28080 20961 28089 20995
rect 28089 20961 28123 20995
rect 28123 20961 28132 20995
rect 28080 20952 28132 20961
rect 29828 20995 29880 21004
rect 29828 20961 29837 20995
rect 29837 20961 29871 20995
rect 29871 20961 29880 20995
rect 29828 20952 29880 20961
rect 18236 20927 18288 20936
rect 18236 20893 18245 20927
rect 18245 20893 18279 20927
rect 18279 20893 18288 20927
rect 18236 20884 18288 20893
rect 26976 20927 27028 20936
rect 26976 20893 26985 20927
rect 26985 20893 27019 20927
rect 27019 20893 27028 20927
rect 26976 20884 27028 20893
rect 27160 20927 27212 20936
rect 27160 20893 27169 20927
rect 27169 20893 27203 20927
rect 27203 20893 27212 20927
rect 27160 20884 27212 20893
rect 30288 20952 30340 21004
rect 16856 20816 16908 20868
rect 17868 20816 17920 20868
rect 29092 20816 29144 20868
rect 29552 20816 29604 20868
rect 33692 20884 33744 20936
rect 34152 20884 34204 20936
rect 34428 20927 34480 20936
rect 34428 20893 34440 20927
rect 34440 20893 34474 20927
rect 34474 20893 34480 20927
rect 34428 20884 34480 20893
rect 34612 20884 34664 20936
rect 34888 20884 34940 20936
rect 16672 20748 16724 20800
rect 20536 20748 20588 20800
rect 23020 20748 23072 20800
rect 26516 20791 26568 20800
rect 26516 20757 26525 20791
rect 26525 20757 26559 20791
rect 26559 20757 26568 20791
rect 26516 20748 26568 20757
rect 27620 20791 27672 20800
rect 27620 20757 27629 20791
rect 27629 20757 27663 20791
rect 27663 20757 27672 20791
rect 27620 20748 27672 20757
rect 29460 20791 29512 20800
rect 29460 20757 29469 20791
rect 29469 20757 29503 20791
rect 29503 20757 29512 20791
rect 29460 20748 29512 20757
rect 35348 20748 35400 20800
rect 35900 20748 35952 20800
rect 36544 20748 36596 20800
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 34966 20646 35018 20698
rect 35030 20646 35082 20698
rect 35094 20646 35146 20698
rect 35158 20646 35210 20698
rect 10048 20587 10100 20596
rect 10048 20553 10057 20587
rect 10057 20553 10091 20587
rect 10091 20553 10100 20587
rect 10048 20544 10100 20553
rect 12992 20544 13044 20596
rect 15752 20544 15804 20596
rect 16580 20544 16632 20596
rect 17960 20544 18012 20596
rect 19340 20544 19392 20596
rect 19524 20544 19576 20596
rect 26608 20587 26660 20596
rect 26608 20553 26617 20587
rect 26617 20553 26651 20587
rect 26651 20553 26660 20587
rect 26608 20544 26660 20553
rect 28080 20544 28132 20596
rect 29092 20587 29144 20596
rect 29092 20553 29101 20587
rect 29101 20553 29135 20587
rect 29135 20553 29144 20587
rect 29092 20544 29144 20553
rect 29828 20544 29880 20596
rect 34336 20544 34388 20596
rect 34428 20544 34480 20596
rect 9128 20476 9180 20528
rect 10048 20340 10100 20392
rect 23388 20476 23440 20528
rect 15016 20408 15068 20460
rect 16396 20408 16448 20460
rect 23020 20408 23072 20460
rect 23480 20408 23532 20460
rect 24492 20476 24544 20528
rect 24952 20451 25004 20460
rect 24952 20417 24961 20451
rect 24961 20417 24995 20451
rect 24995 20417 25004 20451
rect 24952 20408 25004 20417
rect 25136 20451 25188 20460
rect 25136 20417 25145 20451
rect 25145 20417 25179 20451
rect 25179 20417 25188 20451
rect 26148 20451 26200 20460
rect 25136 20408 25188 20417
rect 13268 20340 13320 20392
rect 13728 20340 13780 20392
rect 18052 20383 18104 20392
rect 18052 20349 18061 20383
rect 18061 20349 18095 20383
rect 18095 20349 18104 20383
rect 18052 20340 18104 20349
rect 22100 20340 22152 20392
rect 25320 20340 25372 20392
rect 14004 20272 14056 20324
rect 12256 20204 12308 20256
rect 12624 20204 12676 20256
rect 13728 20204 13780 20256
rect 18328 20315 18380 20324
rect 18328 20281 18362 20315
rect 18362 20281 18380 20315
rect 18328 20272 18380 20281
rect 15752 20204 15804 20256
rect 21456 20204 21508 20256
rect 26148 20417 26157 20451
rect 26157 20417 26191 20451
rect 26191 20417 26200 20451
rect 26148 20408 26200 20417
rect 33876 20476 33928 20528
rect 34152 20476 34204 20528
rect 30564 20451 30616 20460
rect 30564 20417 30573 20451
rect 30573 20417 30607 20451
rect 30607 20417 30616 20451
rect 30564 20408 30616 20417
rect 33324 20408 33376 20460
rect 33416 20340 33468 20392
rect 34244 20340 34296 20392
rect 21916 20204 21968 20256
rect 22100 20247 22152 20256
rect 22100 20213 22109 20247
rect 22109 20213 22143 20247
rect 22143 20213 22152 20247
rect 23664 20247 23716 20256
rect 22100 20204 22152 20213
rect 23664 20213 23673 20247
rect 23673 20213 23707 20247
rect 23707 20213 23716 20247
rect 23664 20204 23716 20213
rect 25872 20272 25924 20324
rect 26332 20272 26384 20324
rect 27160 20272 27212 20324
rect 27620 20272 27672 20324
rect 30932 20272 30984 20324
rect 34612 20272 34664 20324
rect 28080 20247 28132 20256
rect 28080 20213 28089 20247
rect 28089 20213 28123 20247
rect 28123 20213 28132 20247
rect 28080 20204 28132 20213
rect 31944 20247 31996 20256
rect 31944 20213 31953 20247
rect 31953 20213 31987 20247
rect 31987 20213 31996 20247
rect 31944 20204 31996 20213
rect 35072 20340 35124 20392
rect 35808 20340 35860 20392
rect 35808 20204 35860 20256
rect 36176 20204 36228 20256
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 2780 20043 2832 20052
rect 2780 20009 2789 20043
rect 2789 20009 2823 20043
rect 2823 20009 2832 20043
rect 2780 20000 2832 20009
rect 12440 20000 12492 20052
rect 13268 20043 13320 20052
rect 13268 20009 13277 20043
rect 13277 20009 13311 20043
rect 13311 20009 13320 20043
rect 13268 20000 13320 20009
rect 13452 20000 13504 20052
rect 14004 20043 14056 20052
rect 14004 20009 14013 20043
rect 14013 20009 14047 20043
rect 14047 20009 14056 20043
rect 14004 20000 14056 20009
rect 15016 20043 15068 20052
rect 15016 20009 15025 20043
rect 15025 20009 15059 20043
rect 15059 20009 15068 20043
rect 15016 20000 15068 20009
rect 15752 20043 15804 20052
rect 15752 20009 15761 20043
rect 15761 20009 15795 20043
rect 15795 20009 15804 20043
rect 15752 20000 15804 20009
rect 17960 20000 18012 20052
rect 1584 19932 1636 19984
rect 1952 19864 2004 19916
rect 12624 19864 12676 19916
rect 13544 19864 13596 19916
rect 16672 19932 16724 19984
rect 16212 19907 16264 19916
rect 16212 19873 16246 19907
rect 16246 19873 16264 19907
rect 16212 19864 16264 19873
rect 18788 19907 18840 19916
rect 18788 19873 18797 19907
rect 18797 19873 18831 19907
rect 18831 19873 18840 19907
rect 18788 19864 18840 19873
rect 21732 20000 21784 20052
rect 22100 20000 22152 20052
rect 23388 20043 23440 20052
rect 23388 20009 23397 20043
rect 23397 20009 23431 20043
rect 23431 20009 23440 20043
rect 23388 20000 23440 20009
rect 23480 20000 23532 20052
rect 24952 20000 25004 20052
rect 25412 20000 25464 20052
rect 26976 20000 27028 20052
rect 27252 20000 27304 20052
rect 29460 20000 29512 20052
rect 30380 20043 30432 20052
rect 30380 20009 30389 20043
rect 30389 20009 30423 20043
rect 30423 20009 30432 20043
rect 30380 20000 30432 20009
rect 33416 20000 33468 20052
rect 28080 19932 28132 19984
rect 30196 19932 30248 19984
rect 21456 19864 21508 19916
rect 25320 19864 25372 19916
rect 26608 19864 26660 19916
rect 27620 19864 27672 19916
rect 28724 19864 28776 19916
rect 30748 19907 30800 19916
rect 30748 19873 30757 19907
rect 30757 19873 30791 19907
rect 30791 19873 30800 19907
rect 30748 19864 30800 19873
rect 17868 19796 17920 19848
rect 23848 19839 23900 19848
rect 23848 19805 23857 19839
rect 23857 19805 23891 19839
rect 23891 19805 23900 19839
rect 23848 19796 23900 19805
rect 24768 19728 24820 19780
rect 26148 19796 26200 19848
rect 29092 19796 29144 19848
rect 34060 19932 34112 19984
rect 34428 19932 34480 19984
rect 35072 19975 35124 19984
rect 35072 19941 35081 19975
rect 35081 19941 35115 19975
rect 35115 19941 35124 19975
rect 35072 19932 35124 19941
rect 35532 19907 35584 19916
rect 35532 19873 35541 19907
rect 35541 19873 35575 19907
rect 35575 19873 35584 19907
rect 35532 19864 35584 19873
rect 31944 19796 31996 19848
rect 33784 19796 33836 19848
rect 34244 19839 34296 19848
rect 34244 19805 34253 19839
rect 34253 19805 34287 19839
rect 34287 19805 34296 19839
rect 34244 19796 34296 19805
rect 35716 19839 35768 19848
rect 35716 19805 35725 19839
rect 35725 19805 35759 19839
rect 35759 19805 35768 19839
rect 35716 19796 35768 19805
rect 34612 19728 34664 19780
rect 35256 19728 35308 19780
rect 17960 19703 18012 19712
rect 17960 19669 17969 19703
rect 17969 19669 18003 19703
rect 18003 19669 18012 19703
rect 18236 19703 18288 19712
rect 17960 19660 18012 19669
rect 18236 19669 18245 19703
rect 18245 19669 18279 19703
rect 18279 19669 18288 19703
rect 18236 19660 18288 19669
rect 24216 19660 24268 19712
rect 25780 19660 25832 19712
rect 25872 19703 25924 19712
rect 25872 19669 25881 19703
rect 25881 19669 25915 19703
rect 25915 19669 25924 19703
rect 25872 19660 25924 19669
rect 26056 19660 26108 19712
rect 29000 19660 29052 19712
rect 30932 19660 30984 19712
rect 32404 19703 32456 19712
rect 32404 19669 32413 19703
rect 32413 19669 32447 19703
rect 32447 19669 32456 19703
rect 32404 19660 32456 19669
rect 35348 19660 35400 19712
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 34966 19558 35018 19610
rect 35030 19558 35082 19610
rect 35094 19558 35146 19610
rect 35158 19558 35210 19610
rect 1584 19499 1636 19508
rect 1584 19465 1593 19499
rect 1593 19465 1627 19499
rect 1627 19465 1636 19499
rect 1584 19456 1636 19465
rect 1952 19499 2004 19508
rect 1952 19465 1961 19499
rect 1961 19465 1995 19499
rect 1995 19465 2004 19499
rect 1952 19456 2004 19465
rect 14832 19499 14884 19508
rect 14832 19465 14841 19499
rect 14841 19465 14875 19499
rect 14875 19465 14884 19499
rect 14832 19456 14884 19465
rect 15752 19456 15804 19508
rect 17868 19499 17920 19508
rect 17868 19465 17877 19499
rect 17877 19465 17911 19499
rect 17911 19465 17920 19499
rect 17868 19456 17920 19465
rect 18328 19456 18380 19508
rect 24860 19456 24912 19508
rect 25412 19456 25464 19508
rect 26056 19499 26108 19508
rect 26056 19465 26065 19499
rect 26065 19465 26099 19499
rect 26099 19465 26108 19499
rect 26056 19456 26108 19465
rect 26608 19499 26660 19508
rect 26608 19465 26617 19499
rect 26617 19465 26651 19499
rect 26651 19465 26660 19499
rect 26608 19456 26660 19465
rect 28080 19499 28132 19508
rect 28080 19465 28089 19499
rect 28089 19465 28123 19499
rect 28123 19465 28132 19499
rect 28080 19456 28132 19465
rect 34060 19499 34112 19508
rect 34060 19465 34069 19499
rect 34069 19465 34103 19499
rect 34103 19465 34112 19499
rect 34060 19456 34112 19465
rect 13452 19363 13504 19372
rect 13452 19329 13461 19363
rect 13461 19329 13495 19363
rect 13495 19329 13504 19363
rect 13452 19320 13504 19329
rect 16396 19320 16448 19372
rect 13728 19295 13780 19304
rect 13728 19261 13762 19295
rect 13762 19261 13780 19295
rect 13728 19252 13780 19261
rect 16212 19252 16264 19304
rect 17960 19320 18012 19372
rect 25412 19320 25464 19372
rect 29460 19320 29512 19372
rect 30196 19320 30248 19372
rect 30564 19320 30616 19372
rect 32404 19320 32456 19372
rect 35808 19456 35860 19508
rect 18052 19295 18104 19304
rect 18052 19261 18061 19295
rect 18061 19261 18095 19295
rect 18095 19261 18104 19295
rect 18052 19252 18104 19261
rect 20628 19252 20680 19304
rect 21732 19252 21784 19304
rect 24768 19252 24820 19304
rect 26516 19252 26568 19304
rect 27804 19252 27856 19304
rect 15844 19227 15896 19236
rect 15844 19193 15853 19227
rect 15853 19193 15887 19227
rect 15887 19193 15896 19227
rect 15844 19184 15896 19193
rect 18144 19184 18196 19236
rect 18788 19184 18840 19236
rect 20168 19184 20220 19236
rect 16488 19116 16540 19168
rect 19984 19159 20036 19168
rect 19984 19125 19993 19159
rect 19993 19125 20027 19159
rect 20027 19125 20036 19159
rect 19984 19116 20036 19125
rect 21456 19116 21508 19168
rect 24124 19159 24176 19168
rect 24124 19125 24133 19159
rect 24133 19125 24167 19159
rect 24167 19125 24176 19159
rect 24124 19116 24176 19125
rect 24308 19116 24360 19168
rect 26884 19227 26936 19236
rect 26884 19193 26893 19227
rect 26893 19193 26927 19227
rect 26927 19193 26936 19227
rect 26884 19184 26936 19193
rect 30748 19252 30800 19304
rect 33048 19252 33100 19304
rect 32128 19184 32180 19236
rect 34244 19184 34296 19236
rect 36176 19252 36228 19304
rect 35808 19184 35860 19236
rect 24584 19159 24636 19168
rect 24584 19125 24593 19159
rect 24593 19125 24627 19159
rect 24627 19125 24636 19159
rect 24584 19116 24636 19125
rect 24676 19116 24728 19168
rect 28356 19116 28408 19168
rect 28632 19159 28684 19168
rect 28632 19125 28641 19159
rect 28641 19125 28675 19159
rect 28675 19125 28684 19159
rect 28632 19116 28684 19125
rect 29368 19116 29420 19168
rect 30380 19116 30432 19168
rect 31300 19116 31352 19168
rect 32312 19159 32364 19168
rect 32312 19125 32321 19159
rect 32321 19125 32355 19159
rect 32355 19125 32364 19159
rect 32312 19116 32364 19125
rect 32772 19159 32824 19168
rect 32772 19125 32781 19159
rect 32781 19125 32815 19159
rect 32815 19125 32824 19159
rect 32772 19116 32824 19125
rect 33784 19116 33836 19168
rect 33968 19116 34020 19168
rect 35532 19116 35584 19168
rect 35716 19116 35768 19168
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 13544 18955 13596 18964
rect 13544 18921 13553 18955
rect 13553 18921 13587 18955
rect 13587 18921 13596 18955
rect 13544 18912 13596 18921
rect 16212 18912 16264 18964
rect 18144 18955 18196 18964
rect 18144 18921 18153 18955
rect 18153 18921 18187 18955
rect 18187 18921 18196 18955
rect 18144 18912 18196 18921
rect 20536 18955 20588 18964
rect 20536 18921 20545 18955
rect 20545 18921 20579 18955
rect 20579 18921 20588 18955
rect 20536 18912 20588 18921
rect 21456 18955 21508 18964
rect 21456 18921 21465 18955
rect 21465 18921 21499 18955
rect 21499 18921 21508 18955
rect 21456 18912 21508 18921
rect 24676 18955 24728 18964
rect 24676 18921 24685 18955
rect 24685 18921 24719 18955
rect 24719 18921 24728 18955
rect 24676 18912 24728 18921
rect 24860 18955 24912 18964
rect 24860 18921 24869 18955
rect 24869 18921 24903 18955
rect 24903 18921 24912 18955
rect 24860 18912 24912 18921
rect 25504 18912 25556 18964
rect 27804 18955 27856 18964
rect 27804 18921 27813 18955
rect 27813 18921 27847 18955
rect 27847 18921 27856 18955
rect 27804 18912 27856 18921
rect 28356 18955 28408 18964
rect 28356 18921 28365 18955
rect 28365 18921 28399 18955
rect 28399 18921 28408 18955
rect 28356 18912 28408 18921
rect 28724 18912 28776 18964
rect 29092 18912 29144 18964
rect 30932 18955 30984 18964
rect 30932 18921 30941 18955
rect 30941 18921 30975 18955
rect 30975 18921 30984 18955
rect 30932 18912 30984 18921
rect 32128 18955 32180 18964
rect 32128 18921 32137 18955
rect 32137 18921 32171 18955
rect 32171 18921 32180 18955
rect 32128 18912 32180 18921
rect 34244 18912 34296 18964
rect 35256 18912 35308 18964
rect 35532 18912 35584 18964
rect 15844 18844 15896 18896
rect 22100 18844 22152 18896
rect 18420 18819 18472 18828
rect 18420 18785 18429 18819
rect 18429 18785 18463 18819
rect 18463 18785 18472 18819
rect 18420 18776 18472 18785
rect 25596 18844 25648 18896
rect 25964 18887 26016 18896
rect 25964 18853 25973 18887
rect 25973 18853 26007 18887
rect 26007 18853 26016 18887
rect 25964 18844 26016 18853
rect 28816 18844 28868 18896
rect 30288 18844 30340 18896
rect 36176 18887 36228 18896
rect 36176 18853 36185 18887
rect 36185 18853 36219 18887
rect 36219 18853 36228 18887
rect 36176 18844 36228 18853
rect 14004 18708 14056 18760
rect 20076 18708 20128 18760
rect 20260 18708 20312 18760
rect 22928 18776 22980 18828
rect 23664 18776 23716 18828
rect 25228 18819 25280 18828
rect 25228 18785 25237 18819
rect 25237 18785 25271 18819
rect 25271 18785 25280 18819
rect 25228 18776 25280 18785
rect 25780 18776 25832 18828
rect 26884 18819 26936 18828
rect 26884 18785 26893 18819
rect 26893 18785 26927 18819
rect 26927 18785 26936 18819
rect 26884 18776 26936 18785
rect 22376 18751 22428 18760
rect 22376 18717 22385 18751
rect 22385 18717 22419 18751
rect 22419 18717 22428 18751
rect 22376 18708 22428 18717
rect 24492 18708 24544 18760
rect 25412 18751 25464 18760
rect 25412 18717 25421 18751
rect 25421 18717 25455 18751
rect 25455 18717 25464 18751
rect 25412 18708 25464 18717
rect 28448 18751 28500 18760
rect 28448 18717 28457 18751
rect 28457 18717 28491 18751
rect 28491 18717 28500 18751
rect 28448 18708 28500 18717
rect 28908 18708 28960 18760
rect 29092 18708 29144 18760
rect 30196 18776 30248 18828
rect 33692 18776 33744 18828
rect 33876 18776 33928 18828
rect 34060 18751 34112 18760
rect 26976 18640 27028 18692
rect 30564 18640 30616 18692
rect 34060 18717 34072 18751
rect 34072 18717 34106 18751
rect 34106 18717 34112 18751
rect 34060 18708 34112 18717
rect 34336 18751 34388 18760
rect 34336 18717 34345 18751
rect 34345 18717 34379 18751
rect 34379 18717 34388 18751
rect 34336 18708 34388 18717
rect 16304 18572 16356 18624
rect 18052 18572 18104 18624
rect 23388 18572 23440 18624
rect 28816 18572 28868 18624
rect 32128 18572 32180 18624
rect 32772 18572 32824 18624
rect 35716 18615 35768 18624
rect 35716 18581 35725 18615
rect 35725 18581 35759 18615
rect 35759 18581 35768 18615
rect 35716 18572 35768 18581
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 34966 18470 35018 18522
rect 35030 18470 35082 18522
rect 35094 18470 35146 18522
rect 35158 18470 35210 18522
rect 15844 18368 15896 18420
rect 17868 18411 17920 18420
rect 17868 18377 17877 18411
rect 17877 18377 17911 18411
rect 17911 18377 17920 18411
rect 17868 18368 17920 18377
rect 22376 18368 22428 18420
rect 22928 18411 22980 18420
rect 22928 18377 22937 18411
rect 22937 18377 22971 18411
rect 22971 18377 22980 18411
rect 22928 18368 22980 18377
rect 23664 18368 23716 18420
rect 24400 18411 24452 18420
rect 24400 18377 24409 18411
rect 24409 18377 24443 18411
rect 24443 18377 24452 18411
rect 24400 18368 24452 18377
rect 25504 18411 25556 18420
rect 25504 18377 25513 18411
rect 25513 18377 25547 18411
rect 25547 18377 25556 18411
rect 25504 18368 25556 18377
rect 25780 18411 25832 18420
rect 25780 18377 25789 18411
rect 25789 18377 25823 18411
rect 25823 18377 25832 18411
rect 25780 18368 25832 18377
rect 28448 18411 28500 18420
rect 28448 18377 28457 18411
rect 28457 18377 28491 18411
rect 28491 18377 28500 18411
rect 28448 18368 28500 18377
rect 28724 18411 28776 18420
rect 28724 18377 28733 18411
rect 28733 18377 28767 18411
rect 28767 18377 28776 18411
rect 28724 18368 28776 18377
rect 30380 18411 30432 18420
rect 30380 18377 30389 18411
rect 30389 18377 30423 18411
rect 30423 18377 30432 18411
rect 30380 18368 30432 18377
rect 19984 18300 20036 18352
rect 20536 18300 20588 18352
rect 23848 18300 23900 18352
rect 25228 18300 25280 18352
rect 13452 18164 13504 18216
rect 14004 18207 14056 18216
rect 14004 18173 14013 18207
rect 14013 18173 14047 18207
rect 14047 18173 14056 18207
rect 14004 18164 14056 18173
rect 14832 18164 14884 18216
rect 18052 18207 18104 18216
rect 18052 18173 18061 18207
rect 18061 18173 18095 18207
rect 18095 18173 18104 18207
rect 18052 18164 18104 18173
rect 20628 18275 20680 18284
rect 20628 18241 20637 18275
rect 20637 18241 20671 18275
rect 20671 18241 20680 18275
rect 20628 18232 20680 18241
rect 24492 18232 24544 18284
rect 28632 18232 28684 18284
rect 35808 18368 35860 18420
rect 33876 18300 33928 18352
rect 25964 18207 26016 18216
rect 25964 18173 25973 18207
rect 25973 18173 26007 18207
rect 26007 18173 26016 18207
rect 25964 18164 26016 18173
rect 27804 18207 27856 18216
rect 27804 18173 27813 18207
rect 27813 18173 27847 18207
rect 27847 18173 27856 18207
rect 27804 18164 27856 18173
rect 30564 18207 30616 18216
rect 30564 18173 30573 18207
rect 30573 18173 30607 18207
rect 30607 18173 30616 18207
rect 30564 18164 30616 18173
rect 20720 18096 20772 18148
rect 24860 18139 24912 18148
rect 24860 18105 24869 18139
rect 24869 18105 24903 18139
rect 24903 18105 24912 18139
rect 24860 18096 24912 18105
rect 30380 18096 30432 18148
rect 31300 18207 31352 18216
rect 31300 18173 31309 18207
rect 31309 18173 31343 18207
rect 31343 18173 31352 18207
rect 31300 18164 31352 18173
rect 31760 18164 31812 18216
rect 33600 18207 33652 18216
rect 33600 18173 33609 18207
rect 33609 18173 33643 18207
rect 33643 18173 33652 18207
rect 33600 18164 33652 18173
rect 34336 18164 34388 18216
rect 35900 18164 35952 18216
rect 33416 18096 33468 18148
rect 35716 18096 35768 18148
rect 16304 18071 16356 18080
rect 16304 18037 16313 18071
rect 16313 18037 16347 18071
rect 16347 18037 16356 18071
rect 16304 18028 16356 18037
rect 20168 18071 20220 18080
rect 20168 18037 20177 18071
rect 20177 18037 20211 18071
rect 20211 18037 20220 18071
rect 20168 18028 20220 18037
rect 24768 18071 24820 18080
rect 24768 18037 24777 18071
rect 24777 18037 24811 18071
rect 24811 18037 24820 18071
rect 24768 18028 24820 18037
rect 29552 18071 29604 18080
rect 29552 18037 29561 18071
rect 29561 18037 29595 18071
rect 29595 18037 29604 18071
rect 29552 18028 29604 18037
rect 32588 18028 32640 18080
rect 33232 18071 33284 18080
rect 33232 18037 33241 18071
rect 33241 18037 33275 18071
rect 33275 18037 33284 18071
rect 33232 18028 33284 18037
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 14004 17867 14056 17876
rect 14004 17833 14013 17867
rect 14013 17833 14047 17867
rect 14047 17833 14056 17867
rect 14004 17824 14056 17833
rect 16304 17824 16356 17876
rect 18052 17867 18104 17876
rect 18052 17833 18061 17867
rect 18061 17833 18095 17867
rect 18095 17833 18104 17867
rect 18052 17824 18104 17833
rect 20168 17867 20220 17876
rect 20168 17833 20177 17867
rect 20177 17833 20211 17867
rect 20211 17833 20220 17867
rect 20168 17824 20220 17833
rect 20812 17824 20864 17876
rect 24308 17824 24360 17876
rect 24860 17867 24912 17876
rect 24860 17833 24869 17867
rect 24869 17833 24903 17867
rect 24903 17833 24912 17867
rect 24860 17824 24912 17833
rect 25412 17824 25464 17876
rect 26516 17867 26568 17876
rect 26516 17833 26525 17867
rect 26525 17833 26559 17867
rect 26559 17833 26568 17867
rect 26516 17824 26568 17833
rect 27804 17867 27856 17876
rect 27804 17833 27813 17867
rect 27813 17833 27847 17867
rect 27847 17833 27856 17867
rect 27804 17824 27856 17833
rect 31300 17867 31352 17876
rect 31300 17833 31309 17867
rect 31309 17833 31343 17867
rect 31343 17833 31352 17867
rect 31300 17824 31352 17833
rect 31760 17824 31812 17876
rect 32496 17867 32548 17876
rect 32496 17833 32505 17867
rect 32505 17833 32539 17867
rect 32539 17833 32548 17867
rect 32496 17824 32548 17833
rect 32588 17867 32640 17876
rect 32588 17833 32597 17867
rect 32597 17833 32631 17867
rect 32631 17833 32640 17867
rect 33600 17867 33652 17876
rect 32588 17824 32640 17833
rect 33600 17833 33609 17867
rect 33609 17833 33643 17867
rect 33643 17833 33652 17867
rect 33600 17824 33652 17833
rect 34060 17867 34112 17876
rect 34060 17833 34069 17867
rect 34069 17833 34103 17867
rect 34103 17833 34112 17867
rect 34060 17824 34112 17833
rect 35900 17867 35952 17876
rect 35900 17833 35909 17867
rect 35909 17833 35943 17867
rect 35943 17833 35952 17867
rect 35900 17824 35952 17833
rect 19616 17756 19668 17808
rect 20536 17756 20588 17808
rect 24768 17756 24820 17808
rect 28908 17756 28960 17808
rect 29460 17756 29512 17808
rect 33416 17756 33468 17808
rect 35348 17756 35400 17808
rect 36268 17756 36320 17808
rect 22192 17731 22244 17740
rect 22192 17697 22201 17731
rect 22201 17697 22235 17731
rect 22235 17697 22244 17731
rect 22192 17688 22244 17697
rect 22468 17688 22520 17740
rect 23388 17731 23440 17740
rect 23388 17697 23397 17731
rect 23397 17697 23431 17731
rect 23431 17697 23440 17731
rect 23388 17688 23440 17697
rect 24492 17688 24544 17740
rect 25228 17731 25280 17740
rect 25228 17697 25237 17731
rect 25237 17697 25271 17731
rect 25271 17697 25280 17731
rect 25228 17688 25280 17697
rect 26884 17731 26936 17740
rect 26884 17697 26893 17731
rect 26893 17697 26927 17731
rect 26927 17697 26936 17731
rect 26884 17688 26936 17697
rect 35256 17688 35308 17740
rect 25320 17663 25372 17672
rect 25320 17629 25329 17663
rect 25329 17629 25363 17663
rect 25363 17629 25372 17663
rect 25320 17620 25372 17629
rect 26976 17663 27028 17672
rect 25136 17552 25188 17604
rect 26976 17629 26985 17663
rect 26985 17629 27019 17663
rect 27019 17629 27028 17663
rect 26976 17620 27028 17629
rect 18420 17527 18472 17536
rect 18420 17493 18429 17527
rect 18429 17493 18463 17527
rect 18463 17493 18472 17527
rect 18420 17484 18472 17493
rect 20720 17527 20772 17536
rect 20720 17493 20729 17527
rect 20729 17493 20763 17527
rect 20763 17493 20772 17527
rect 20720 17484 20772 17493
rect 21824 17527 21876 17536
rect 21824 17493 21833 17527
rect 21833 17493 21867 17527
rect 21867 17493 21876 17527
rect 21824 17484 21876 17493
rect 24952 17484 25004 17536
rect 25872 17484 25924 17536
rect 32772 17663 32824 17672
rect 32772 17629 32781 17663
rect 32781 17629 32815 17663
rect 32815 17629 32824 17663
rect 32772 17620 32824 17629
rect 34060 17620 34112 17672
rect 35348 17620 35400 17672
rect 32128 17595 32180 17604
rect 32128 17561 32137 17595
rect 32137 17561 32171 17595
rect 32171 17561 32180 17595
rect 32128 17552 32180 17561
rect 34244 17552 34296 17604
rect 34520 17552 34572 17604
rect 35624 17552 35676 17604
rect 35900 17552 35952 17604
rect 27896 17484 27948 17536
rect 29092 17527 29144 17536
rect 29092 17493 29101 17527
rect 29101 17493 29135 17527
rect 29135 17493 29144 17527
rect 29092 17484 29144 17493
rect 30472 17484 30524 17536
rect 35716 17484 35768 17536
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 34966 17382 35018 17434
rect 35030 17382 35082 17434
rect 35094 17382 35146 17434
rect 35158 17382 35210 17434
rect 18972 17323 19024 17332
rect 18972 17289 18981 17323
rect 18981 17289 19015 17323
rect 19015 17289 19024 17323
rect 18972 17280 19024 17289
rect 20720 17280 20772 17332
rect 22192 17280 22244 17332
rect 23388 17323 23440 17332
rect 23388 17289 23397 17323
rect 23397 17289 23431 17323
rect 23431 17289 23440 17323
rect 23388 17280 23440 17289
rect 23848 17323 23900 17332
rect 23848 17289 23857 17323
rect 23857 17289 23891 17323
rect 23891 17289 23900 17323
rect 23848 17280 23900 17289
rect 27436 17323 27488 17332
rect 27436 17289 27445 17323
rect 27445 17289 27479 17323
rect 27479 17289 27488 17323
rect 27436 17280 27488 17289
rect 27896 17323 27948 17332
rect 27896 17289 27905 17323
rect 27905 17289 27939 17323
rect 27939 17289 27948 17323
rect 27896 17280 27948 17289
rect 29092 17323 29144 17332
rect 29092 17289 29101 17323
rect 29101 17289 29135 17323
rect 29135 17289 29144 17323
rect 29092 17280 29144 17289
rect 29460 17323 29512 17332
rect 29460 17289 29469 17323
rect 29469 17289 29503 17323
rect 29503 17289 29512 17323
rect 29460 17280 29512 17289
rect 30380 17280 30432 17332
rect 32772 17280 32824 17332
rect 33232 17280 33284 17332
rect 34060 17323 34112 17332
rect 34060 17289 34069 17323
rect 34069 17289 34103 17323
rect 34103 17289 34112 17323
rect 34060 17280 34112 17289
rect 35256 17280 35308 17332
rect 32496 17255 32548 17264
rect 32496 17221 32505 17255
rect 32505 17221 32539 17255
rect 32539 17221 32548 17255
rect 32496 17212 32548 17221
rect 33692 17255 33744 17264
rect 33692 17221 33701 17255
rect 33701 17221 33735 17255
rect 33735 17221 33744 17255
rect 33692 17212 33744 17221
rect 19616 17187 19668 17196
rect 19616 17153 19625 17187
rect 19625 17153 19659 17187
rect 19659 17153 19668 17187
rect 19616 17144 19668 17153
rect 19892 17144 19944 17196
rect 32588 17144 32640 17196
rect 35716 17280 35768 17332
rect 20628 17076 20680 17128
rect 22468 17119 22520 17128
rect 22468 17085 22477 17119
rect 22477 17085 22511 17119
rect 22511 17085 22520 17119
rect 22468 17076 22520 17085
rect 23664 17119 23716 17128
rect 23664 17085 23673 17119
rect 23673 17085 23707 17119
rect 23707 17085 23716 17119
rect 23664 17076 23716 17085
rect 24860 17119 24912 17128
rect 24860 17085 24869 17119
rect 24869 17085 24903 17119
rect 24903 17085 24912 17119
rect 24860 17076 24912 17085
rect 24952 17076 25004 17128
rect 26976 17076 27028 17128
rect 27620 17119 27672 17128
rect 27620 17085 27629 17119
rect 27629 17085 27663 17119
rect 27663 17085 27672 17119
rect 27620 17076 27672 17085
rect 30288 17076 30340 17128
rect 30472 17119 30524 17128
rect 19064 17008 19116 17060
rect 22284 17008 22336 17060
rect 24124 17008 24176 17060
rect 25320 17008 25372 17060
rect 30472 17085 30506 17119
rect 30506 17085 30524 17119
rect 30472 17076 30524 17085
rect 35808 17008 35860 17060
rect 20168 16940 20220 16992
rect 25228 16940 25280 16992
rect 26240 16983 26292 16992
rect 26240 16949 26249 16983
rect 26249 16949 26283 16983
rect 26283 16949 26292 16983
rect 26240 16940 26292 16949
rect 26884 16940 26936 16992
rect 35348 16940 35400 16992
rect 36912 16940 36964 16992
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 19064 16779 19116 16788
rect 19064 16745 19073 16779
rect 19073 16745 19107 16779
rect 19107 16745 19116 16779
rect 19064 16736 19116 16745
rect 19248 16779 19300 16788
rect 19248 16745 19257 16779
rect 19257 16745 19291 16779
rect 19291 16745 19300 16779
rect 19248 16736 19300 16745
rect 22284 16779 22336 16788
rect 22284 16745 22293 16779
rect 22293 16745 22327 16779
rect 22327 16745 22336 16779
rect 22284 16736 22336 16745
rect 23664 16779 23716 16788
rect 23664 16745 23673 16779
rect 23673 16745 23707 16779
rect 23707 16745 23716 16779
rect 23664 16736 23716 16745
rect 25228 16736 25280 16788
rect 20168 16668 20220 16720
rect 22100 16668 22152 16720
rect 24124 16668 24176 16720
rect 24860 16668 24912 16720
rect 19616 16643 19668 16652
rect 19616 16609 19625 16643
rect 19625 16609 19659 16643
rect 19659 16609 19668 16643
rect 19616 16600 19668 16609
rect 20720 16600 20772 16652
rect 26976 16736 27028 16788
rect 29920 16779 29972 16788
rect 29920 16745 29929 16779
rect 29929 16745 29963 16779
rect 29963 16745 29972 16779
rect 29920 16736 29972 16745
rect 30380 16736 30432 16788
rect 35808 16736 35860 16788
rect 29552 16668 29604 16720
rect 30196 16668 30248 16720
rect 27068 16600 27120 16652
rect 29000 16600 29052 16652
rect 19708 16575 19760 16584
rect 19708 16541 19717 16575
rect 19717 16541 19751 16575
rect 19751 16541 19760 16575
rect 19708 16532 19760 16541
rect 19892 16575 19944 16584
rect 19892 16541 19901 16575
rect 19901 16541 19935 16575
rect 19935 16541 19944 16575
rect 19892 16532 19944 16541
rect 26516 16575 26568 16584
rect 26516 16541 26525 16575
rect 26525 16541 26559 16575
rect 26559 16541 26568 16575
rect 26516 16532 26568 16541
rect 30380 16575 30432 16584
rect 30380 16541 30389 16575
rect 30389 16541 30423 16575
rect 30423 16541 30432 16575
rect 30380 16532 30432 16541
rect 30472 16575 30524 16584
rect 30472 16541 30481 16575
rect 30481 16541 30515 16575
rect 30515 16541 30524 16575
rect 30472 16532 30524 16541
rect 35440 16532 35492 16584
rect 36636 16532 36688 16584
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 34966 16294 35018 16346
rect 35030 16294 35082 16346
rect 35094 16294 35146 16346
rect 35158 16294 35210 16346
rect 19892 16192 19944 16244
rect 20168 16235 20220 16244
rect 20168 16201 20177 16235
rect 20177 16201 20211 16235
rect 20211 16201 20220 16235
rect 20168 16192 20220 16201
rect 22100 16235 22152 16244
rect 22100 16201 22109 16235
rect 22109 16201 22143 16235
rect 22143 16201 22152 16235
rect 22100 16192 22152 16201
rect 24124 16192 24176 16244
rect 27068 16192 27120 16244
rect 29920 16235 29972 16244
rect 29920 16201 29929 16235
rect 29929 16201 29963 16235
rect 29963 16201 29972 16235
rect 29920 16192 29972 16201
rect 30196 16235 30248 16244
rect 30196 16201 30205 16235
rect 30205 16201 30239 16235
rect 30239 16201 30248 16235
rect 30196 16192 30248 16201
rect 30472 16192 30524 16244
rect 25136 16124 25188 16176
rect 33048 16124 33100 16176
rect 34612 16124 34664 16176
rect 19708 16056 19760 16108
rect 20628 16056 20680 16108
rect 28632 16099 28684 16108
rect 20720 16031 20772 16040
rect 20720 15997 20729 16031
rect 20729 15997 20763 16031
rect 20763 15997 20772 16031
rect 20720 15988 20772 15997
rect 24584 15988 24636 16040
rect 24860 15988 24912 16040
rect 26516 15988 26568 16040
rect 28632 16065 28641 16099
rect 28641 16065 28675 16099
rect 28675 16065 28684 16099
rect 28632 16056 28684 16065
rect 29920 15988 29972 16040
rect 19616 15920 19668 15972
rect 22284 15920 22336 15972
rect 25780 15963 25832 15972
rect 25780 15929 25814 15963
rect 25814 15929 25832 15963
rect 25780 15920 25832 15929
rect 27160 15852 27212 15904
rect 29460 15895 29512 15904
rect 29460 15861 29469 15895
rect 29469 15861 29503 15895
rect 29503 15861 29512 15895
rect 29460 15852 29512 15861
rect 33048 15852 33100 15904
rect 35808 15852 35860 15904
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 22284 15691 22336 15700
rect 22284 15657 22293 15691
rect 22293 15657 22327 15691
rect 22327 15657 22336 15691
rect 22284 15648 22336 15657
rect 30380 15691 30432 15700
rect 30380 15657 30389 15691
rect 30389 15657 30423 15691
rect 30423 15657 30432 15691
rect 30380 15648 30432 15657
rect 35716 15648 35768 15700
rect 35992 15691 36044 15700
rect 35992 15657 36001 15691
rect 36001 15657 36035 15691
rect 36035 15657 36044 15691
rect 35992 15648 36044 15657
rect 20628 15512 20680 15564
rect 22008 15512 22060 15564
rect 27988 15512 28040 15564
rect 29736 15555 29788 15564
rect 29736 15521 29745 15555
rect 29745 15521 29779 15555
rect 29779 15521 29788 15555
rect 29736 15512 29788 15521
rect 32220 15512 32272 15564
rect 33048 15512 33100 15564
rect 35440 15555 35492 15564
rect 35440 15521 35449 15555
rect 35449 15521 35483 15555
rect 35483 15521 35492 15555
rect 35440 15512 35492 15521
rect 20720 15487 20772 15496
rect 20720 15453 20729 15487
rect 20729 15453 20763 15487
rect 20763 15453 20772 15487
rect 20904 15487 20956 15496
rect 20720 15444 20772 15453
rect 20904 15453 20913 15487
rect 20913 15453 20947 15487
rect 20947 15453 20956 15487
rect 20904 15444 20956 15453
rect 27804 15487 27856 15496
rect 27804 15453 27813 15487
rect 27813 15453 27847 15487
rect 27847 15453 27856 15487
rect 27804 15444 27856 15453
rect 27896 15487 27948 15496
rect 27896 15453 27905 15487
rect 27905 15453 27939 15487
rect 27939 15453 27948 15487
rect 27896 15444 27948 15453
rect 29460 15444 29512 15496
rect 31760 15444 31812 15496
rect 32956 15487 33008 15496
rect 32956 15453 32965 15487
rect 32965 15453 32999 15487
rect 32999 15453 33008 15487
rect 32956 15444 33008 15453
rect 27160 15376 27212 15428
rect 26516 15308 26568 15360
rect 27068 15351 27120 15360
rect 27068 15317 27077 15351
rect 27077 15317 27111 15351
rect 27111 15317 27120 15351
rect 27068 15308 27120 15317
rect 27344 15351 27396 15360
rect 27344 15317 27353 15351
rect 27353 15317 27387 15351
rect 27387 15317 27396 15351
rect 27344 15308 27396 15317
rect 30196 15308 30248 15360
rect 32404 15351 32456 15360
rect 32404 15317 32413 15351
rect 32413 15317 32447 15351
rect 32447 15317 32456 15351
rect 32404 15308 32456 15317
rect 34520 15308 34572 15360
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 34966 15206 35018 15258
rect 35030 15206 35082 15258
rect 35094 15206 35146 15258
rect 35158 15206 35210 15258
rect 20628 15147 20680 15156
rect 20628 15113 20637 15147
rect 20637 15113 20671 15147
rect 20671 15113 20680 15147
rect 20628 15104 20680 15113
rect 22100 15104 22152 15156
rect 27804 15104 27856 15156
rect 27988 15147 28040 15156
rect 27988 15113 27997 15147
rect 27997 15113 28031 15147
rect 28031 15113 28040 15147
rect 27988 15104 28040 15113
rect 29736 15104 29788 15156
rect 31760 15147 31812 15156
rect 31760 15113 31769 15147
rect 31769 15113 31803 15147
rect 31803 15113 31812 15147
rect 32220 15147 32272 15156
rect 31760 15104 31812 15113
rect 32220 15113 32229 15147
rect 32229 15113 32263 15147
rect 32263 15113 32272 15147
rect 32220 15104 32272 15113
rect 32956 15104 33008 15156
rect 35440 15104 35492 15156
rect 27068 15036 27120 15088
rect 28080 15036 28132 15088
rect 27160 15011 27212 15020
rect 20904 14900 20956 14952
rect 27160 14977 27169 15011
rect 27169 14977 27203 15011
rect 27203 14977 27212 15011
rect 27160 14968 27212 14977
rect 30564 15011 30616 15020
rect 30564 14977 30573 15011
rect 30573 14977 30607 15011
rect 30607 14977 30616 15011
rect 30564 14968 30616 14977
rect 21364 14943 21416 14952
rect 21364 14909 21398 14943
rect 21398 14909 21416 14943
rect 21364 14900 21416 14909
rect 27344 14900 27396 14952
rect 30012 14943 30064 14952
rect 30012 14909 30021 14943
rect 30021 14909 30055 14943
rect 30055 14909 30064 14943
rect 30012 14900 30064 14909
rect 21180 14832 21232 14884
rect 26516 14875 26568 14884
rect 26516 14841 26525 14875
rect 26525 14841 26559 14875
rect 26559 14841 26568 14875
rect 26516 14832 26568 14841
rect 30748 14900 30800 14952
rect 32312 14943 32364 14952
rect 32312 14909 32321 14943
rect 32321 14909 32355 14943
rect 32355 14909 32364 14943
rect 32312 14900 32364 14909
rect 35256 14900 35308 14952
rect 35992 14900 36044 14952
rect 32772 14832 32824 14884
rect 36452 14832 36504 14884
rect 26608 14807 26660 14816
rect 26608 14773 26617 14807
rect 26617 14773 26651 14807
rect 26651 14773 26660 14807
rect 26608 14764 26660 14773
rect 33784 14764 33836 14816
rect 35532 14764 35584 14816
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 24584 14603 24636 14612
rect 24584 14569 24593 14603
rect 24593 14569 24627 14603
rect 24627 14569 24636 14603
rect 24584 14560 24636 14569
rect 26516 14603 26568 14612
rect 26516 14569 26525 14603
rect 26525 14569 26559 14603
rect 26559 14569 26568 14603
rect 26516 14560 26568 14569
rect 27068 14492 27120 14544
rect 23848 14467 23900 14476
rect 23848 14433 23857 14467
rect 23857 14433 23891 14467
rect 23891 14433 23900 14467
rect 23848 14424 23900 14433
rect 23940 14399 23992 14408
rect 23940 14365 23949 14399
rect 23949 14365 23983 14399
rect 23983 14365 23992 14399
rect 23940 14356 23992 14365
rect 26976 14399 27028 14408
rect 23112 14288 23164 14340
rect 26976 14365 26985 14399
rect 26985 14365 27019 14399
rect 27019 14365 27028 14399
rect 26976 14356 27028 14365
rect 27344 14356 27396 14408
rect 27896 14560 27948 14612
rect 30012 14560 30064 14612
rect 32220 14603 32272 14612
rect 32220 14569 32229 14603
rect 32229 14569 32263 14603
rect 32263 14569 32272 14603
rect 32220 14560 32272 14569
rect 33876 14560 33928 14612
rect 34612 14560 34664 14612
rect 35532 14603 35584 14612
rect 27988 14492 28040 14544
rect 28724 14492 28776 14544
rect 35532 14569 35541 14603
rect 35541 14569 35575 14603
rect 35575 14569 35584 14603
rect 35532 14560 35584 14569
rect 36176 14560 36228 14612
rect 36084 14492 36136 14544
rect 28080 14356 28132 14408
rect 30288 14424 30340 14476
rect 21180 14263 21232 14272
rect 21180 14229 21189 14263
rect 21189 14229 21223 14263
rect 21223 14229 21232 14263
rect 21180 14220 21232 14229
rect 24032 14220 24084 14272
rect 32312 14220 32364 14272
rect 32772 14263 32824 14272
rect 32772 14229 32781 14263
rect 32781 14229 32815 14263
rect 32815 14229 32824 14263
rect 32772 14220 32824 14229
rect 34428 14424 34480 14476
rect 33600 14356 33652 14408
rect 33784 14356 33836 14408
rect 36176 14356 36228 14408
rect 36452 14399 36504 14408
rect 36452 14365 36461 14399
rect 36461 14365 36495 14399
rect 36495 14365 36504 14399
rect 36452 14356 36504 14365
rect 33232 14220 33284 14272
rect 35900 14263 35952 14272
rect 35900 14229 35909 14263
rect 35909 14229 35943 14263
rect 35943 14229 35952 14263
rect 35900 14220 35952 14229
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 34966 14118 35018 14170
rect 35030 14118 35082 14170
rect 35094 14118 35146 14170
rect 35158 14118 35210 14170
rect 23112 14016 23164 14068
rect 23848 14016 23900 14068
rect 26148 14016 26200 14068
rect 26976 14016 27028 14068
rect 27804 14016 27856 14068
rect 28724 14059 28776 14068
rect 28724 14025 28733 14059
rect 28733 14025 28767 14059
rect 28767 14025 28776 14059
rect 28724 14016 28776 14025
rect 29000 14016 29052 14068
rect 30012 14016 30064 14068
rect 32680 14016 32732 14068
rect 33600 14016 33652 14068
rect 33876 14016 33928 14068
rect 36084 14016 36136 14068
rect 36452 14016 36504 14068
rect 36820 13991 36872 14000
rect 36820 13957 36829 13991
rect 36829 13957 36863 13991
rect 36863 13957 36872 13991
rect 36820 13948 36872 13957
rect 33784 13880 33836 13932
rect 23664 13855 23716 13864
rect 23664 13821 23673 13855
rect 23673 13821 23707 13855
rect 23707 13821 23716 13855
rect 23664 13812 23716 13821
rect 23940 13855 23992 13864
rect 23940 13821 23963 13855
rect 23963 13821 23992 13855
rect 23940 13812 23992 13821
rect 26700 13855 26752 13864
rect 26700 13821 26709 13855
rect 26709 13821 26743 13855
rect 26743 13821 26752 13855
rect 26700 13812 26752 13821
rect 28080 13812 28132 13864
rect 30012 13855 30064 13864
rect 30012 13821 30046 13855
rect 30046 13821 30064 13855
rect 23020 13719 23072 13728
rect 23020 13685 23029 13719
rect 23029 13685 23063 13719
rect 23063 13685 23072 13719
rect 27068 13744 27120 13796
rect 30012 13812 30064 13821
rect 32312 13855 32364 13864
rect 32312 13821 32321 13855
rect 32321 13821 32355 13855
rect 32355 13821 32364 13855
rect 32312 13812 32364 13821
rect 35256 13812 35308 13864
rect 35532 13812 35584 13864
rect 30288 13744 30340 13796
rect 23020 13676 23072 13685
rect 30932 13676 30984 13728
rect 32128 13719 32180 13728
rect 32128 13685 32137 13719
rect 32137 13685 32171 13719
rect 32171 13685 32180 13719
rect 32128 13676 32180 13685
rect 33692 13719 33744 13728
rect 33692 13685 33701 13719
rect 33701 13685 33735 13719
rect 33735 13685 33744 13719
rect 33692 13676 33744 13685
rect 34796 13676 34848 13728
rect 35348 13676 35400 13728
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 23848 13472 23900 13524
rect 25596 13472 25648 13524
rect 26148 13472 26200 13524
rect 27344 13472 27396 13524
rect 29000 13515 29052 13524
rect 29000 13481 29009 13515
rect 29009 13481 29043 13515
rect 29043 13481 29052 13515
rect 29000 13472 29052 13481
rect 30288 13472 30340 13524
rect 30472 13515 30524 13524
rect 30472 13481 30481 13515
rect 30481 13481 30515 13515
rect 30515 13481 30524 13515
rect 30472 13472 30524 13481
rect 30748 13472 30800 13524
rect 24676 13404 24728 13456
rect 27804 13404 27856 13456
rect 28080 13404 28132 13456
rect 30656 13404 30708 13456
rect 32312 13472 32364 13524
rect 32404 13472 32456 13524
rect 23664 13336 23716 13388
rect 23756 13336 23808 13388
rect 24584 13336 24636 13388
rect 26608 13336 26660 13388
rect 30380 13336 30432 13388
rect 32772 13472 32824 13524
rect 33876 13472 33928 13524
rect 34428 13472 34480 13524
rect 34796 13472 34848 13524
rect 35256 13472 35308 13524
rect 35808 13515 35860 13524
rect 35808 13481 35817 13515
rect 35817 13481 35851 13515
rect 35851 13481 35860 13515
rect 35808 13472 35860 13481
rect 36176 13472 36228 13524
rect 22836 13311 22888 13320
rect 22836 13277 22845 13311
rect 22845 13277 22879 13311
rect 22879 13277 22888 13311
rect 22836 13268 22888 13277
rect 23112 13268 23164 13320
rect 30564 13311 30616 13320
rect 30564 13277 30573 13311
rect 30573 13277 30607 13311
rect 30607 13277 30616 13311
rect 30564 13268 30616 13277
rect 32680 13311 32732 13320
rect 32680 13277 32689 13311
rect 32689 13277 32723 13311
rect 32723 13277 32732 13311
rect 32680 13268 32732 13277
rect 35532 13336 35584 13388
rect 33416 13311 33468 13320
rect 33416 13277 33425 13311
rect 33425 13277 33459 13311
rect 33459 13277 33468 13311
rect 33416 13268 33468 13277
rect 35900 13311 35952 13320
rect 35900 13277 35909 13311
rect 35909 13277 35943 13311
rect 35943 13277 35952 13311
rect 35900 13268 35952 13277
rect 36084 13268 36136 13320
rect 34244 13200 34296 13252
rect 35532 13200 35584 13252
rect 22376 13175 22428 13184
rect 22376 13141 22385 13175
rect 22385 13141 22419 13175
rect 22419 13141 22428 13175
rect 22376 13132 22428 13141
rect 27620 13132 27672 13184
rect 30012 13132 30064 13184
rect 35256 13175 35308 13184
rect 35256 13141 35265 13175
rect 35265 13141 35299 13175
rect 35299 13141 35308 13175
rect 35256 13132 35308 13141
rect 35992 13132 36044 13184
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 34966 13030 35018 13082
rect 35030 13030 35082 13082
rect 35094 13030 35146 13082
rect 35158 13030 35210 13082
rect 23020 12928 23072 12980
rect 24676 12971 24728 12980
rect 24676 12937 24685 12971
rect 24685 12937 24719 12971
rect 24719 12937 24728 12971
rect 24676 12928 24728 12937
rect 25596 12971 25648 12980
rect 25596 12937 25605 12971
rect 25605 12937 25639 12971
rect 25639 12937 25648 12971
rect 25596 12928 25648 12937
rect 27068 12971 27120 12980
rect 27068 12937 27077 12971
rect 27077 12937 27111 12971
rect 27111 12937 27120 12971
rect 27068 12928 27120 12937
rect 27804 12928 27856 12980
rect 28080 12971 28132 12980
rect 28080 12937 28089 12971
rect 28089 12937 28123 12971
rect 28123 12937 28132 12971
rect 28080 12928 28132 12937
rect 30196 12971 30248 12980
rect 30196 12937 30205 12971
rect 30205 12937 30239 12971
rect 30239 12937 30248 12971
rect 30196 12928 30248 12937
rect 30564 12928 30616 12980
rect 32772 12971 32824 12980
rect 32772 12937 32781 12971
rect 32781 12937 32815 12971
rect 32815 12937 32824 12971
rect 32772 12928 32824 12937
rect 33048 12928 33100 12980
rect 35808 12928 35860 12980
rect 35900 12928 35952 12980
rect 24860 12860 24912 12912
rect 22376 12792 22428 12844
rect 24124 12835 24176 12844
rect 24124 12801 24133 12835
rect 24133 12801 24167 12835
rect 24167 12801 24176 12835
rect 24124 12792 24176 12801
rect 24584 12792 24636 12844
rect 30380 12860 30432 12912
rect 30472 12903 30524 12912
rect 30472 12869 30481 12903
rect 30481 12869 30515 12903
rect 30515 12869 30524 12903
rect 30472 12860 30524 12869
rect 33876 12860 33928 12912
rect 36452 12860 36504 12912
rect 30656 12835 30708 12844
rect 21180 12724 21232 12776
rect 24032 12767 24084 12776
rect 24032 12733 24041 12767
rect 24041 12733 24075 12767
rect 24075 12733 24084 12767
rect 24032 12724 24084 12733
rect 25688 12767 25740 12776
rect 25688 12733 25697 12767
rect 25697 12733 25731 12767
rect 25731 12733 25740 12767
rect 25688 12724 25740 12733
rect 30656 12801 30665 12835
rect 30665 12801 30699 12835
rect 30699 12801 30708 12835
rect 30656 12792 30708 12801
rect 33784 12835 33836 12844
rect 33784 12801 33793 12835
rect 33793 12801 33827 12835
rect 33827 12801 33836 12835
rect 33784 12792 33836 12801
rect 34336 12792 34388 12844
rect 29644 12724 29696 12776
rect 30012 12724 30064 12776
rect 30932 12767 30984 12776
rect 30932 12733 30966 12767
rect 30966 12733 30984 12767
rect 30932 12724 30984 12733
rect 22376 12656 22428 12708
rect 22836 12656 22888 12708
rect 33140 12656 33192 12708
rect 33416 12656 33468 12708
rect 23664 12588 23716 12640
rect 31760 12588 31812 12640
rect 32128 12588 32180 12640
rect 33600 12631 33652 12640
rect 33600 12597 33609 12631
rect 33609 12597 33643 12631
rect 33643 12597 33652 12631
rect 33600 12588 33652 12597
rect 33784 12588 33836 12640
rect 34152 12588 34204 12640
rect 34796 12792 34848 12844
rect 35256 12724 35308 12776
rect 35716 12724 35768 12776
rect 34428 12588 34480 12640
rect 34520 12588 34572 12640
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 23664 12427 23716 12436
rect 23664 12393 23673 12427
rect 23673 12393 23707 12427
rect 23707 12393 23716 12427
rect 23664 12384 23716 12393
rect 24124 12384 24176 12436
rect 26608 12384 26660 12436
rect 27436 12427 27488 12436
rect 27436 12393 27445 12427
rect 27445 12393 27479 12427
rect 27479 12393 27488 12427
rect 27436 12384 27488 12393
rect 29644 12427 29696 12436
rect 29644 12393 29653 12427
rect 29653 12393 29687 12427
rect 29687 12393 29696 12427
rect 29644 12384 29696 12393
rect 30288 12384 30340 12436
rect 30380 12384 30432 12436
rect 33140 12384 33192 12436
rect 33324 12384 33376 12436
rect 34244 12427 34296 12436
rect 22376 12316 22428 12368
rect 30196 12316 30248 12368
rect 34244 12393 34253 12427
rect 34253 12393 34287 12427
rect 34287 12393 34296 12427
rect 34244 12384 34296 12393
rect 34336 12384 34388 12436
rect 36084 12384 36136 12436
rect 24860 12248 24912 12300
rect 27620 12248 27672 12300
rect 27804 12291 27856 12300
rect 27804 12257 27813 12291
rect 27813 12257 27847 12291
rect 27847 12257 27856 12291
rect 27804 12248 27856 12257
rect 29000 12291 29052 12300
rect 29000 12257 29009 12291
rect 29009 12257 29043 12291
rect 29043 12257 29052 12291
rect 29000 12248 29052 12257
rect 30104 12248 30156 12300
rect 33140 12291 33192 12300
rect 33140 12257 33149 12291
rect 33149 12257 33183 12291
rect 33183 12257 33192 12291
rect 33140 12248 33192 12257
rect 33600 12248 33652 12300
rect 33876 12248 33928 12300
rect 34612 12291 34664 12300
rect 34612 12257 34646 12291
rect 34646 12257 34664 12291
rect 34612 12248 34664 12257
rect 21180 12223 21232 12232
rect 21180 12189 21189 12223
rect 21189 12189 21223 12223
rect 21223 12189 21232 12223
rect 22284 12223 22336 12232
rect 21180 12180 21232 12189
rect 22284 12189 22293 12223
rect 22293 12189 22327 12223
rect 22327 12189 22336 12223
rect 22284 12180 22336 12189
rect 26608 12180 26660 12232
rect 28080 12223 28132 12232
rect 28080 12189 28089 12223
rect 28089 12189 28123 12223
rect 28123 12189 28132 12223
rect 28080 12180 28132 12189
rect 30656 12223 30708 12232
rect 30656 12189 30665 12223
rect 30665 12189 30699 12223
rect 30699 12189 30708 12223
rect 30656 12180 30708 12189
rect 30932 12180 30984 12232
rect 33232 12223 33284 12232
rect 33232 12189 33241 12223
rect 33241 12189 33275 12223
rect 33275 12189 33284 12223
rect 33232 12180 33284 12189
rect 33692 12180 33744 12232
rect 31484 12155 31536 12164
rect 31484 12121 31493 12155
rect 31493 12121 31527 12155
rect 31527 12121 31536 12155
rect 31484 12112 31536 12121
rect 32680 12112 32732 12164
rect 24584 12087 24636 12096
rect 24584 12053 24593 12087
rect 24593 12053 24627 12087
rect 24627 12053 24636 12087
rect 24584 12044 24636 12053
rect 25504 12044 25556 12096
rect 25688 12087 25740 12096
rect 25688 12053 25697 12087
rect 25697 12053 25731 12087
rect 25731 12053 25740 12087
rect 25688 12044 25740 12053
rect 29184 12087 29236 12096
rect 29184 12053 29193 12087
rect 29193 12053 29227 12087
rect 29227 12053 29236 12087
rect 29184 12044 29236 12053
rect 31944 12087 31996 12096
rect 31944 12053 31953 12087
rect 31953 12053 31987 12087
rect 31987 12053 31996 12087
rect 31944 12044 31996 12053
rect 32772 12087 32824 12096
rect 32772 12053 32781 12087
rect 32781 12053 32815 12087
rect 32815 12053 32824 12087
rect 32772 12044 32824 12053
rect 33692 12044 33744 12096
rect 34336 12044 34388 12096
rect 34612 12044 34664 12096
rect 35440 12044 35492 12096
rect 35716 12087 35768 12096
rect 35716 12053 35725 12087
rect 35725 12053 35759 12087
rect 35759 12053 35768 12087
rect 35716 12044 35768 12053
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 34966 11942 35018 11994
rect 35030 11942 35082 11994
rect 35094 11942 35146 11994
rect 35158 11942 35210 11994
rect 24860 11840 24912 11892
rect 25504 11840 25556 11892
rect 26700 11883 26752 11892
rect 26700 11849 26709 11883
rect 26709 11849 26743 11883
rect 26743 11849 26752 11883
rect 26700 11840 26752 11849
rect 27804 11840 27856 11892
rect 29000 11883 29052 11892
rect 29000 11849 29009 11883
rect 29009 11849 29043 11883
rect 29043 11849 29052 11883
rect 29000 11840 29052 11849
rect 29184 11840 29236 11892
rect 30104 11883 30156 11892
rect 30104 11849 30113 11883
rect 30113 11849 30147 11883
rect 30147 11849 30156 11883
rect 30104 11840 30156 11849
rect 30380 11840 30432 11892
rect 22284 11772 22336 11824
rect 23388 11772 23440 11824
rect 26608 11815 26660 11824
rect 26608 11781 26617 11815
rect 26617 11781 26651 11815
rect 26651 11781 26660 11815
rect 26608 11772 26660 11781
rect 30656 11772 30708 11824
rect 23664 11704 23716 11756
rect 22560 11636 22612 11688
rect 27436 11704 27488 11756
rect 28080 11747 28132 11756
rect 28080 11713 28089 11747
rect 28089 11713 28123 11747
rect 28123 11713 28132 11747
rect 28080 11704 28132 11713
rect 31484 11704 31536 11756
rect 33232 11840 33284 11892
rect 33692 11840 33744 11892
rect 33876 11883 33928 11892
rect 33876 11849 33885 11883
rect 33885 11849 33919 11883
rect 33919 11849 33928 11883
rect 33876 11840 33928 11849
rect 34336 11883 34388 11892
rect 34336 11849 34345 11883
rect 34345 11849 34379 11883
rect 34379 11849 34388 11883
rect 34336 11840 34388 11849
rect 34612 11840 34664 11892
rect 35348 11840 35400 11892
rect 35716 11840 35768 11892
rect 36268 11840 36320 11892
rect 35256 11772 35308 11824
rect 36084 11772 36136 11824
rect 33140 11747 33192 11756
rect 23480 11568 23532 11620
rect 27344 11636 27396 11688
rect 31392 11636 31444 11688
rect 31576 11636 31628 11688
rect 33140 11713 33149 11747
rect 33149 11713 33183 11747
rect 33183 11713 33192 11747
rect 33140 11704 33192 11713
rect 35440 11747 35492 11756
rect 35440 11713 35449 11747
rect 35449 11713 35483 11747
rect 35483 11713 35492 11747
rect 35440 11704 35492 11713
rect 35348 11679 35400 11688
rect 35348 11645 35357 11679
rect 35357 11645 35391 11679
rect 35391 11645 35400 11679
rect 35348 11636 35400 11645
rect 28724 11568 28776 11620
rect 32128 11568 32180 11620
rect 35072 11568 35124 11620
rect 22376 11543 22428 11552
rect 22376 11509 22385 11543
rect 22385 11509 22419 11543
rect 22419 11509 22428 11543
rect 22376 11500 22428 11509
rect 23756 11543 23808 11552
rect 23756 11509 23765 11543
rect 23765 11509 23799 11543
rect 23799 11509 23808 11543
rect 23756 11500 23808 11509
rect 26240 11543 26292 11552
rect 26240 11509 26249 11543
rect 26249 11509 26283 11543
rect 26283 11509 26292 11543
rect 26240 11500 26292 11509
rect 27896 11543 27948 11552
rect 27896 11509 27905 11543
rect 27905 11509 27939 11543
rect 27939 11509 27948 11543
rect 27896 11500 27948 11509
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 22376 11296 22428 11348
rect 27160 11296 27212 11348
rect 28080 11296 28132 11348
rect 28724 11339 28776 11348
rect 28724 11305 28733 11339
rect 28733 11305 28767 11339
rect 28767 11305 28776 11339
rect 28724 11296 28776 11305
rect 31392 11339 31444 11348
rect 31392 11305 31401 11339
rect 31401 11305 31435 11339
rect 31435 11305 31444 11339
rect 31392 11296 31444 11305
rect 32128 11339 32180 11348
rect 32128 11305 32137 11339
rect 32137 11305 32171 11339
rect 32171 11305 32180 11339
rect 32128 11296 32180 11305
rect 35072 11339 35124 11348
rect 35072 11305 35081 11339
rect 35081 11305 35115 11339
rect 35115 11305 35124 11339
rect 35072 11296 35124 11305
rect 27528 11228 27580 11280
rect 35440 11228 35492 11280
rect 22468 11160 22520 11212
rect 22652 11203 22704 11212
rect 22652 11169 22686 11203
rect 22686 11169 22704 11203
rect 22652 11160 22704 11169
rect 25320 11203 25372 11212
rect 25320 11169 25329 11203
rect 25329 11169 25363 11203
rect 25363 11169 25372 11203
rect 25320 11160 25372 11169
rect 26424 11160 26476 11212
rect 28540 11203 28592 11212
rect 28540 11169 28549 11203
rect 28549 11169 28583 11203
rect 28583 11169 28592 11203
rect 28540 11160 28592 11169
rect 33876 11160 33928 11212
rect 27436 11092 27488 11144
rect 35440 11092 35492 11144
rect 27896 11024 27948 11076
rect 29184 11067 29236 11076
rect 29184 11033 29193 11067
rect 29193 11033 29227 11067
rect 29227 11033 29236 11067
rect 29184 11024 29236 11033
rect 22560 10956 22612 11008
rect 24308 10999 24360 11008
rect 24308 10965 24317 10999
rect 24317 10965 24351 10999
rect 24351 10965 24360 10999
rect 24308 10956 24360 10965
rect 26976 10999 27028 11008
rect 26976 10965 26985 10999
rect 26985 10965 27019 10999
rect 27019 10965 27028 10999
rect 26976 10956 27028 10965
rect 30288 10956 30340 11008
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 34966 10854 35018 10906
rect 35030 10854 35082 10906
rect 35094 10854 35146 10906
rect 35158 10854 35210 10906
rect 23756 10752 23808 10804
rect 27344 10752 27396 10804
rect 28264 10752 28316 10804
rect 30104 10752 30156 10804
rect 22560 10659 22612 10668
rect 22560 10625 22569 10659
rect 22569 10625 22603 10659
rect 22603 10625 22612 10659
rect 22560 10616 22612 10625
rect 25320 10727 25372 10736
rect 25320 10693 25329 10727
rect 25329 10693 25363 10727
rect 25363 10693 25372 10727
rect 25320 10684 25372 10693
rect 28540 10727 28592 10736
rect 28540 10693 28549 10727
rect 28549 10693 28583 10727
rect 28583 10693 28592 10727
rect 28540 10684 28592 10693
rect 24584 10659 24636 10668
rect 24584 10625 24593 10659
rect 24593 10625 24627 10659
rect 24627 10625 24636 10659
rect 24584 10616 24636 10625
rect 26976 10659 27028 10668
rect 26976 10625 26985 10659
rect 26985 10625 27019 10659
rect 27019 10625 27028 10659
rect 26976 10616 27028 10625
rect 27160 10659 27212 10668
rect 27160 10625 27169 10659
rect 27169 10625 27203 10659
rect 27203 10625 27212 10659
rect 27160 10616 27212 10625
rect 30196 10616 30248 10668
rect 35440 10659 35492 10668
rect 35440 10625 35449 10659
rect 35449 10625 35483 10659
rect 35483 10625 35492 10659
rect 35440 10616 35492 10625
rect 22284 10548 22336 10600
rect 22652 10548 22704 10600
rect 23112 10548 23164 10600
rect 28908 10548 28960 10600
rect 24308 10523 24360 10532
rect 24308 10489 24317 10523
rect 24317 10489 24351 10523
rect 24351 10489 24360 10523
rect 24308 10480 24360 10489
rect 27160 10480 27212 10532
rect 27436 10480 27488 10532
rect 30104 10480 30156 10532
rect 35808 10480 35860 10532
rect 22284 10412 22336 10464
rect 22928 10412 22980 10464
rect 23112 10455 23164 10464
rect 23112 10421 23121 10455
rect 23121 10421 23155 10455
rect 23155 10421 23164 10455
rect 23112 10412 23164 10421
rect 26424 10455 26476 10464
rect 26424 10421 26433 10455
rect 26433 10421 26467 10455
rect 26467 10421 26476 10455
rect 26424 10412 26476 10421
rect 26608 10412 26660 10464
rect 27620 10455 27672 10464
rect 27620 10421 27629 10455
rect 27629 10421 27663 10455
rect 27663 10421 27672 10455
rect 27620 10412 27672 10421
rect 29920 10412 29972 10464
rect 30288 10455 30340 10464
rect 30288 10421 30297 10455
rect 30297 10421 30331 10455
rect 30331 10421 30340 10455
rect 30288 10412 30340 10421
rect 34520 10412 34572 10464
rect 36820 10455 36872 10464
rect 36820 10421 36829 10455
rect 36829 10421 36863 10455
rect 36863 10421 36872 10455
rect 36820 10412 36872 10421
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 23112 10208 23164 10260
rect 26424 10208 26476 10260
rect 30104 10208 30156 10260
rect 30564 10208 30616 10260
rect 32496 10251 32548 10260
rect 32496 10217 32505 10251
rect 32505 10217 32539 10251
rect 32539 10217 32548 10251
rect 32496 10208 32548 10217
rect 35440 10251 35492 10260
rect 35440 10217 35449 10251
rect 35449 10217 35483 10251
rect 35483 10217 35492 10251
rect 35440 10208 35492 10217
rect 35532 10208 35584 10260
rect 33140 10140 33192 10192
rect 23020 10115 23072 10124
rect 23020 10081 23054 10115
rect 23054 10081 23072 10115
rect 23020 10072 23072 10081
rect 27620 10072 27672 10124
rect 29092 10072 29144 10124
rect 33048 10115 33100 10124
rect 33048 10081 33057 10115
rect 33057 10081 33091 10115
rect 33091 10081 33100 10115
rect 33048 10072 33100 10081
rect 33876 10140 33928 10192
rect 33508 10072 33560 10124
rect 36268 10115 36320 10124
rect 36268 10081 36277 10115
rect 36277 10081 36311 10115
rect 36311 10081 36320 10115
rect 36268 10072 36320 10081
rect 29920 10047 29972 10056
rect 29920 10013 29929 10047
rect 29929 10013 29963 10047
rect 29963 10013 29972 10047
rect 29920 10004 29972 10013
rect 30104 10047 30156 10056
rect 30104 10013 30113 10047
rect 30113 10013 30147 10047
rect 30147 10013 30156 10047
rect 30104 10004 30156 10013
rect 36360 10047 36412 10056
rect 36360 10013 36369 10047
rect 36369 10013 36403 10047
rect 36403 10013 36412 10047
rect 36360 10004 36412 10013
rect 36820 10004 36872 10056
rect 29828 9936 29880 9988
rect 22468 9911 22520 9920
rect 22468 9877 22477 9911
rect 22477 9877 22511 9911
rect 22511 9877 22520 9911
rect 22468 9868 22520 9877
rect 26332 9911 26384 9920
rect 26332 9877 26341 9911
rect 26341 9877 26375 9911
rect 26375 9877 26384 9911
rect 26332 9868 26384 9877
rect 26608 9868 26660 9920
rect 29460 9911 29512 9920
rect 29460 9877 29469 9911
rect 29469 9877 29503 9911
rect 29503 9877 29512 9911
rect 29460 9868 29512 9877
rect 34796 9911 34848 9920
rect 34796 9877 34805 9911
rect 34805 9877 34839 9911
rect 34839 9877 34848 9911
rect 34796 9868 34848 9877
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 34966 9766 35018 9818
rect 35030 9766 35082 9818
rect 35094 9766 35146 9818
rect 35158 9766 35210 9818
rect 23020 9664 23072 9716
rect 29092 9707 29144 9716
rect 23480 9639 23532 9648
rect 23480 9605 23489 9639
rect 23489 9605 23523 9639
rect 23523 9605 23532 9639
rect 23480 9596 23532 9605
rect 29092 9673 29101 9707
rect 29101 9673 29135 9707
rect 29135 9673 29144 9707
rect 29092 9664 29144 9673
rect 28724 9639 28776 9648
rect 28724 9605 28733 9639
rect 28733 9605 28767 9639
rect 28767 9605 28776 9639
rect 30104 9664 30156 9716
rect 30288 9664 30340 9716
rect 33048 9664 33100 9716
rect 35808 9664 35860 9716
rect 28724 9596 28776 9605
rect 31852 9596 31904 9648
rect 29460 9528 29512 9580
rect 30564 9571 30616 9580
rect 30564 9537 30573 9571
rect 30573 9537 30607 9571
rect 30607 9537 30616 9571
rect 30564 9528 30616 9537
rect 33508 9571 33560 9580
rect 33508 9537 33517 9571
rect 33517 9537 33551 9571
rect 33551 9537 33560 9571
rect 33508 9528 33560 9537
rect 22468 9435 22520 9444
rect 22468 9401 22477 9435
rect 22477 9401 22511 9435
rect 22511 9401 22520 9435
rect 22468 9392 22520 9401
rect 23480 9392 23532 9444
rect 24860 9460 24912 9512
rect 25688 9503 25740 9512
rect 25688 9469 25697 9503
rect 25697 9469 25731 9503
rect 25731 9469 25740 9503
rect 25688 9460 25740 9469
rect 26240 9460 26292 9512
rect 29828 9503 29880 9512
rect 29828 9469 29837 9503
rect 29837 9469 29871 9503
rect 29871 9469 29880 9503
rect 29828 9460 29880 9469
rect 32496 9460 32548 9512
rect 24492 9392 24544 9444
rect 26056 9435 26108 9444
rect 26056 9401 26065 9435
rect 26065 9401 26099 9435
rect 26099 9401 26108 9435
rect 26056 9392 26108 9401
rect 27528 9367 27580 9376
rect 27528 9333 27537 9367
rect 27537 9333 27571 9367
rect 27571 9333 27580 9367
rect 27528 9324 27580 9333
rect 27620 9324 27672 9376
rect 28908 9324 28960 9376
rect 29644 9367 29696 9376
rect 29644 9333 29653 9367
rect 29653 9333 29687 9367
rect 29687 9333 29696 9367
rect 29644 9324 29696 9333
rect 32496 9367 32548 9376
rect 32496 9333 32505 9367
rect 32505 9333 32539 9367
rect 32539 9333 32548 9367
rect 32496 9324 32548 9333
rect 33140 9392 33192 9444
rect 36268 9460 36320 9512
rect 34796 9392 34848 9444
rect 35440 9392 35492 9444
rect 33324 9324 33376 9376
rect 34888 9324 34940 9376
rect 35992 9324 36044 9376
rect 36820 9367 36872 9376
rect 36820 9333 36829 9367
rect 36829 9333 36863 9367
rect 36863 9333 36872 9367
rect 36820 9324 36872 9333
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 24860 9163 24912 9172
rect 24860 9129 24869 9163
rect 24869 9129 24903 9163
rect 24903 9129 24912 9163
rect 24860 9120 24912 9129
rect 29920 9120 29972 9172
rect 30196 9120 30248 9172
rect 32956 9120 33008 9172
rect 34244 9120 34296 9172
rect 36268 9163 36320 9172
rect 29828 9095 29880 9104
rect 29828 9061 29862 9095
rect 29862 9061 29880 9095
rect 29828 9052 29880 9061
rect 36268 9129 36277 9163
rect 36277 9129 36311 9163
rect 36311 9129 36320 9163
rect 36268 9120 36320 9129
rect 36360 9120 36412 9172
rect 23480 9027 23532 9036
rect 23480 8993 23489 9027
rect 23489 8993 23523 9027
rect 23523 8993 23532 9027
rect 23480 8984 23532 8993
rect 23756 9027 23808 9036
rect 23756 8993 23790 9027
rect 23790 8993 23808 9027
rect 23756 8984 23808 8993
rect 26148 9027 26200 9036
rect 26148 8993 26157 9027
rect 26157 8993 26191 9027
rect 26191 8993 26200 9027
rect 26148 8984 26200 8993
rect 26424 8984 26476 9036
rect 27712 8984 27764 9036
rect 35348 8984 35400 9036
rect 24492 8848 24544 8900
rect 26240 8916 26292 8968
rect 26516 8959 26568 8968
rect 26516 8925 26525 8959
rect 26525 8925 26559 8959
rect 26559 8925 26568 8959
rect 26516 8916 26568 8925
rect 29368 8916 29420 8968
rect 31944 8916 31996 8968
rect 33048 8959 33100 8968
rect 33048 8925 33060 8959
rect 33060 8925 33094 8959
rect 33094 8925 33100 8959
rect 33324 8959 33376 8968
rect 33048 8916 33100 8925
rect 33324 8925 33333 8959
rect 33333 8925 33367 8959
rect 33367 8925 33376 8959
rect 33324 8916 33376 8925
rect 35440 8848 35492 8900
rect 35808 8959 35860 8968
rect 35808 8925 35817 8959
rect 35817 8925 35851 8959
rect 35851 8925 35860 8959
rect 35808 8916 35860 8925
rect 35900 8848 35952 8900
rect 27896 8823 27948 8832
rect 27896 8789 27905 8823
rect 27905 8789 27939 8823
rect 27939 8789 27948 8823
rect 27896 8780 27948 8789
rect 29184 8780 29236 8832
rect 32036 8780 32088 8832
rect 32864 8780 32916 8832
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 34966 8678 35018 8730
rect 35030 8678 35082 8730
rect 35094 8678 35146 8730
rect 35158 8678 35210 8730
rect 23756 8576 23808 8628
rect 26056 8619 26108 8628
rect 26056 8585 26065 8619
rect 26065 8585 26099 8619
rect 26099 8585 26108 8619
rect 26056 8576 26108 8585
rect 26424 8619 26476 8628
rect 26424 8585 26433 8619
rect 26433 8585 26467 8619
rect 26467 8585 26476 8619
rect 26424 8576 26476 8585
rect 26608 8619 26660 8628
rect 26608 8585 26617 8619
rect 26617 8585 26651 8619
rect 26651 8585 26660 8619
rect 26608 8576 26660 8585
rect 27712 8576 27764 8628
rect 29736 8576 29788 8628
rect 30380 8576 30432 8628
rect 31852 8619 31904 8628
rect 31852 8585 31861 8619
rect 31861 8585 31895 8619
rect 31895 8585 31904 8619
rect 31852 8576 31904 8585
rect 32496 8576 32548 8628
rect 27896 8508 27948 8560
rect 33508 8508 33560 8560
rect 27160 8483 27212 8492
rect 27160 8449 27169 8483
rect 27169 8449 27203 8483
rect 27203 8449 27212 8483
rect 29368 8483 29420 8492
rect 27160 8440 27212 8449
rect 29368 8449 29377 8483
rect 29377 8449 29411 8483
rect 29411 8449 29420 8483
rect 29368 8440 29420 8449
rect 24124 8415 24176 8424
rect 24124 8381 24133 8415
rect 24133 8381 24167 8415
rect 24167 8381 24176 8415
rect 24124 8372 24176 8381
rect 26884 8372 26936 8424
rect 27528 8372 27580 8424
rect 30196 8304 30248 8356
rect 30380 8304 30432 8356
rect 32036 8415 32088 8424
rect 32036 8381 32045 8415
rect 32045 8381 32079 8415
rect 32079 8381 32088 8415
rect 32036 8372 32088 8381
rect 33140 8372 33192 8424
rect 32864 8304 32916 8356
rect 34520 8576 34572 8628
rect 34704 8508 34756 8560
rect 35164 8508 35216 8560
rect 35808 8576 35860 8628
rect 37096 8619 37148 8628
rect 37096 8585 37105 8619
rect 37105 8585 37139 8619
rect 37139 8585 37148 8619
rect 37096 8576 37148 8585
rect 35900 8551 35952 8560
rect 35900 8517 35909 8551
rect 35909 8517 35943 8551
rect 35943 8517 35952 8551
rect 35900 8508 35952 8517
rect 35440 8483 35492 8492
rect 35440 8449 35449 8483
rect 35449 8449 35483 8483
rect 35483 8449 35492 8483
rect 35440 8440 35492 8449
rect 37096 8372 37148 8424
rect 35808 8304 35860 8356
rect 36084 8304 36136 8356
rect 28356 8236 28408 8288
rect 31760 8279 31812 8288
rect 31760 8245 31769 8279
rect 31769 8245 31803 8279
rect 31803 8245 31812 8279
rect 36636 8279 36688 8288
rect 31760 8236 31812 8245
rect 36636 8245 36645 8279
rect 36645 8245 36679 8279
rect 36679 8245 36688 8279
rect 36636 8236 36688 8245
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 24124 8032 24176 8084
rect 24492 8032 24544 8084
rect 26148 8032 26200 8084
rect 26884 8032 26936 8084
rect 27160 8075 27212 8084
rect 27160 8041 27169 8075
rect 27169 8041 27203 8075
rect 27203 8041 27212 8075
rect 27160 8032 27212 8041
rect 29000 8032 29052 8084
rect 30380 8075 30432 8084
rect 30380 8041 30389 8075
rect 30389 8041 30423 8075
rect 30423 8041 30432 8075
rect 30380 8032 30432 8041
rect 31760 8032 31812 8084
rect 33048 8032 33100 8084
rect 33324 8032 33376 8084
rect 35348 8075 35400 8084
rect 35348 8041 35357 8075
rect 35357 8041 35391 8075
rect 35391 8041 35400 8075
rect 35348 8032 35400 8041
rect 28724 7964 28776 8016
rect 31944 8007 31996 8016
rect 31944 7973 31953 8007
rect 31953 7973 31987 8007
rect 31987 7973 31996 8007
rect 31944 7964 31996 7973
rect 32956 7964 33008 8016
rect 35624 7964 35676 8016
rect 32128 7939 32180 7948
rect 32128 7905 32137 7939
rect 32137 7905 32171 7939
rect 32171 7905 32180 7939
rect 32128 7896 32180 7905
rect 33140 7896 33192 7948
rect 33324 7896 33376 7948
rect 36176 7896 36228 7948
rect 28356 7871 28408 7880
rect 28356 7837 28365 7871
rect 28365 7837 28399 7871
rect 28399 7837 28408 7871
rect 28356 7828 28408 7837
rect 32036 7828 32088 7880
rect 35532 7760 35584 7812
rect 36360 7760 36412 7812
rect 34612 7735 34664 7744
rect 34612 7701 34621 7735
rect 34621 7701 34655 7735
rect 34655 7701 34664 7735
rect 34612 7692 34664 7701
rect 34796 7692 34848 7744
rect 35716 7692 35768 7744
rect 36084 7735 36136 7744
rect 36084 7701 36093 7735
rect 36093 7701 36127 7735
rect 36127 7701 36136 7735
rect 36084 7692 36136 7701
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 34966 7590 35018 7642
rect 35030 7590 35082 7642
rect 35094 7590 35146 7642
rect 35158 7590 35210 7642
rect 28724 7488 28776 7540
rect 32036 7531 32088 7540
rect 32036 7497 32045 7531
rect 32045 7497 32079 7531
rect 32079 7497 32088 7531
rect 32036 7488 32088 7497
rect 32404 7488 32456 7540
rect 33140 7488 33192 7540
rect 35624 7488 35676 7540
rect 29092 7352 29144 7404
rect 32864 7395 32916 7404
rect 32864 7361 32873 7395
rect 32873 7361 32907 7395
rect 32907 7361 32916 7395
rect 32864 7352 32916 7361
rect 32036 7284 32088 7336
rect 33324 7327 33376 7336
rect 33324 7293 33333 7327
rect 33333 7293 33367 7327
rect 33367 7293 33376 7327
rect 35440 7327 35492 7336
rect 33324 7284 33376 7293
rect 31208 7216 31260 7268
rect 32680 7259 32732 7268
rect 32680 7225 32689 7259
rect 32689 7225 32723 7259
rect 32723 7225 32732 7259
rect 32680 7216 32732 7225
rect 27620 7148 27672 7200
rect 28356 7148 28408 7200
rect 31300 7191 31352 7200
rect 31300 7157 31309 7191
rect 31309 7157 31343 7191
rect 31343 7157 31352 7191
rect 31300 7148 31352 7157
rect 35440 7293 35449 7327
rect 35449 7293 35483 7327
rect 35483 7293 35492 7327
rect 35440 7284 35492 7293
rect 36176 7216 36228 7268
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 32128 6944 32180 6996
rect 32680 6987 32732 6996
rect 32680 6953 32689 6987
rect 32689 6953 32723 6987
rect 32723 6953 32732 6987
rect 32680 6944 32732 6953
rect 34796 6944 34848 6996
rect 35440 6944 35492 6996
rect 31300 6876 31352 6928
rect 32772 6876 32824 6928
rect 33324 6876 33376 6928
rect 26792 6851 26844 6860
rect 26792 6817 26826 6851
rect 26826 6817 26844 6851
rect 26792 6808 26844 6817
rect 30288 6851 30340 6860
rect 30288 6817 30297 6851
rect 30297 6817 30331 6851
rect 30331 6817 30340 6851
rect 30288 6808 30340 6817
rect 31852 6808 31904 6860
rect 31944 6808 31996 6860
rect 34244 6851 34296 6860
rect 26516 6783 26568 6792
rect 26516 6749 26525 6783
rect 26525 6749 26559 6783
rect 26559 6749 26568 6783
rect 26516 6740 26568 6749
rect 34244 6817 34253 6851
rect 34253 6817 34287 6851
rect 34287 6817 34296 6851
rect 34244 6808 34296 6817
rect 35440 6808 35492 6860
rect 37004 6808 37056 6860
rect 32404 6672 32456 6724
rect 26516 6604 26568 6656
rect 27528 6604 27580 6656
rect 27896 6647 27948 6656
rect 27896 6613 27905 6647
rect 27905 6613 27939 6647
rect 27939 6613 27948 6647
rect 27896 6604 27948 6613
rect 29828 6604 29880 6656
rect 30840 6604 30892 6656
rect 31392 6647 31444 6656
rect 31392 6613 31401 6647
rect 31401 6613 31435 6647
rect 31435 6613 31444 6647
rect 31392 6604 31444 6613
rect 33784 6647 33836 6656
rect 33784 6613 33793 6647
rect 33793 6613 33827 6647
rect 33827 6613 33836 6647
rect 33784 6604 33836 6613
rect 35532 6647 35584 6656
rect 35532 6613 35541 6647
rect 35541 6613 35575 6647
rect 35575 6613 35584 6647
rect 35532 6604 35584 6613
rect 36176 6604 36228 6656
rect 36452 6604 36504 6656
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 34966 6502 35018 6554
rect 35030 6502 35082 6554
rect 35094 6502 35146 6554
rect 35158 6502 35210 6554
rect 26792 6400 26844 6452
rect 30840 6443 30892 6452
rect 30840 6409 30849 6443
rect 30849 6409 30883 6443
rect 30883 6409 30892 6443
rect 30840 6400 30892 6409
rect 32404 6443 32456 6452
rect 32404 6409 32413 6443
rect 32413 6409 32447 6443
rect 32447 6409 32456 6443
rect 32404 6400 32456 6409
rect 32772 6443 32824 6452
rect 32772 6409 32781 6443
rect 32781 6409 32815 6443
rect 32815 6409 32824 6443
rect 32772 6400 32824 6409
rect 36544 6443 36596 6452
rect 36544 6409 36553 6443
rect 36553 6409 36587 6443
rect 36587 6409 36596 6443
rect 36544 6400 36596 6409
rect 37004 6443 37056 6452
rect 37004 6409 37013 6443
rect 37013 6409 37047 6443
rect 37047 6409 37056 6443
rect 37004 6400 37056 6409
rect 30288 6375 30340 6384
rect 27896 6264 27948 6316
rect 28724 6264 28776 6316
rect 30288 6341 30297 6375
rect 30297 6341 30331 6375
rect 30331 6341 30340 6375
rect 30288 6332 30340 6341
rect 29828 6307 29880 6316
rect 29828 6273 29837 6307
rect 29837 6273 29871 6307
rect 29871 6273 29880 6307
rect 29828 6264 29880 6273
rect 34244 6375 34296 6384
rect 34244 6341 34253 6375
rect 34253 6341 34287 6375
rect 34287 6341 34296 6375
rect 34244 6332 34296 6341
rect 31392 6264 31444 6316
rect 33416 6264 33468 6316
rect 33784 6264 33836 6316
rect 37280 6375 37332 6384
rect 37280 6341 37289 6375
rect 37289 6341 37323 6375
rect 37323 6341 37332 6375
rect 37280 6332 37332 6341
rect 32128 6196 32180 6248
rect 33140 6196 33192 6248
rect 31852 6128 31904 6180
rect 36084 6196 36136 6248
rect 26516 6060 26568 6112
rect 26700 6060 26752 6112
rect 27988 6103 28040 6112
rect 27988 6069 27997 6103
rect 27997 6069 28031 6103
rect 28031 6069 28040 6103
rect 27988 6060 28040 6069
rect 28724 6103 28776 6112
rect 28724 6069 28733 6103
rect 28733 6069 28767 6103
rect 28767 6069 28776 6103
rect 28724 6060 28776 6069
rect 29000 6060 29052 6112
rect 31116 6060 31168 6112
rect 31300 6103 31352 6112
rect 31300 6069 31309 6103
rect 31309 6069 31343 6103
rect 31343 6069 31352 6103
rect 31300 6060 31352 6069
rect 31668 6103 31720 6112
rect 31668 6069 31677 6103
rect 31677 6069 31711 6103
rect 31711 6069 31720 6103
rect 31668 6060 31720 6069
rect 32956 6060 33008 6112
rect 34612 6103 34664 6112
rect 34612 6069 34621 6103
rect 34621 6069 34655 6103
rect 34655 6069 34664 6103
rect 34612 6060 34664 6069
rect 35072 6103 35124 6112
rect 35072 6069 35081 6103
rect 35081 6069 35115 6103
rect 35115 6069 35124 6103
rect 35072 6060 35124 6069
rect 35440 6103 35492 6112
rect 35440 6069 35449 6103
rect 35449 6069 35483 6103
rect 35483 6069 35492 6103
rect 35440 6060 35492 6069
rect 35900 6060 35952 6112
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 27988 5856 28040 5908
rect 31668 5856 31720 5908
rect 33876 5856 33928 5908
rect 35072 5856 35124 5908
rect 27436 5788 27488 5840
rect 27896 5788 27948 5840
rect 29828 5788 29880 5840
rect 30288 5788 30340 5840
rect 31300 5788 31352 5840
rect 31944 5831 31996 5840
rect 30196 5763 30248 5772
rect 30196 5729 30205 5763
rect 30205 5729 30239 5763
rect 30239 5729 30248 5763
rect 30196 5720 30248 5729
rect 31944 5797 31953 5831
rect 31953 5797 31987 5831
rect 31987 5797 31996 5831
rect 31944 5788 31996 5797
rect 32956 5831 33008 5840
rect 32956 5797 32965 5831
rect 32965 5797 32999 5831
rect 32999 5797 33008 5831
rect 32956 5788 33008 5797
rect 33600 5831 33652 5840
rect 33600 5797 33609 5831
rect 33609 5797 33643 5831
rect 33643 5797 33652 5831
rect 33600 5788 33652 5797
rect 35532 5788 35584 5840
rect 26700 5652 26752 5704
rect 30104 5652 30156 5704
rect 34796 5720 34848 5772
rect 33416 5652 33468 5704
rect 34244 5652 34296 5704
rect 34428 5652 34480 5704
rect 34888 5695 34940 5704
rect 34888 5661 34897 5695
rect 34897 5661 34931 5695
rect 34931 5661 34940 5695
rect 34888 5652 34940 5661
rect 35256 5652 35308 5704
rect 35532 5695 35584 5704
rect 35532 5661 35541 5695
rect 35541 5661 35575 5695
rect 35575 5661 35584 5695
rect 35532 5652 35584 5661
rect 31116 5584 31168 5636
rect 33140 5627 33192 5636
rect 33140 5593 33149 5627
rect 33149 5593 33183 5627
rect 33183 5593 33192 5627
rect 33140 5584 33192 5593
rect 34520 5584 34572 5636
rect 29000 5516 29052 5568
rect 29828 5559 29880 5568
rect 29828 5525 29837 5559
rect 29837 5525 29871 5559
rect 29871 5525 29880 5559
rect 29828 5516 29880 5525
rect 32772 5516 32824 5568
rect 36268 5516 36320 5568
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 34966 5414 35018 5466
rect 35030 5414 35082 5466
rect 35094 5414 35146 5466
rect 35158 5414 35210 5466
rect 27436 5355 27488 5364
rect 27436 5321 27445 5355
rect 27445 5321 27479 5355
rect 27479 5321 27488 5355
rect 27436 5312 27488 5321
rect 28908 5312 28960 5364
rect 30380 5312 30432 5364
rect 32404 5355 32456 5364
rect 28724 5176 28776 5228
rect 32404 5321 32413 5355
rect 32413 5321 32447 5355
rect 32447 5321 32456 5355
rect 32404 5312 32456 5321
rect 33600 5312 33652 5364
rect 33876 5355 33928 5364
rect 33876 5321 33885 5355
rect 33885 5321 33919 5355
rect 33919 5321 33928 5355
rect 33876 5312 33928 5321
rect 34244 5355 34296 5364
rect 34244 5321 34253 5355
rect 34253 5321 34287 5355
rect 34287 5321 34296 5355
rect 34244 5312 34296 5321
rect 36176 5312 36228 5364
rect 33048 5219 33100 5228
rect 33048 5185 33057 5219
rect 33057 5185 33091 5219
rect 33091 5185 33100 5219
rect 33048 5176 33100 5185
rect 34428 5176 34480 5228
rect 35164 5176 35216 5228
rect 29276 5151 29328 5160
rect 29276 5117 29285 5151
rect 29285 5117 29319 5151
rect 29319 5117 29328 5151
rect 29276 5108 29328 5117
rect 34704 5108 34756 5160
rect 36268 5040 36320 5092
rect 26700 5015 26752 5024
rect 26700 4981 26709 5015
rect 26709 4981 26743 5015
rect 26743 4981 26752 5015
rect 26700 4972 26752 4981
rect 27896 4972 27948 5024
rect 28080 5015 28132 5024
rect 28080 4981 28089 5015
rect 28089 4981 28123 5015
rect 28123 4981 28132 5015
rect 28724 5015 28776 5024
rect 28080 4972 28132 4981
rect 28724 4981 28733 5015
rect 28733 4981 28767 5015
rect 28767 4981 28776 5015
rect 28724 4972 28776 4981
rect 30380 4972 30432 5024
rect 32220 5015 32272 5024
rect 32220 4981 32229 5015
rect 32229 4981 32263 5015
rect 32263 4981 32272 5015
rect 32220 4972 32272 4981
rect 32772 5015 32824 5024
rect 32772 4981 32781 5015
rect 32781 4981 32815 5015
rect 32815 4981 32824 5015
rect 32772 4972 32824 4981
rect 34796 4972 34848 5024
rect 35256 4972 35308 5024
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 28080 4768 28132 4820
rect 30196 4811 30248 4820
rect 30196 4777 30205 4811
rect 30205 4777 30239 4811
rect 30239 4777 30248 4811
rect 30196 4768 30248 4777
rect 31760 4768 31812 4820
rect 27988 4700 28040 4752
rect 33784 4768 33836 4820
rect 34428 4768 34480 4820
rect 34704 4811 34756 4820
rect 34704 4777 34713 4811
rect 34713 4777 34747 4811
rect 34747 4777 34756 4811
rect 34704 4768 34756 4777
rect 34612 4700 34664 4752
rect 26700 4632 26752 4684
rect 28448 4632 28500 4684
rect 30748 4675 30800 4684
rect 30748 4641 30757 4675
rect 30757 4641 30791 4675
rect 30791 4641 30800 4675
rect 30748 4632 30800 4641
rect 31208 4632 31260 4684
rect 32128 4675 32180 4684
rect 32128 4641 32137 4675
rect 32137 4641 32171 4675
rect 32171 4641 32180 4675
rect 32128 4632 32180 4641
rect 34060 4632 34112 4684
rect 34704 4632 34756 4684
rect 31024 4607 31076 4616
rect 31024 4573 31033 4607
rect 31033 4573 31067 4607
rect 31067 4573 31076 4607
rect 31024 4564 31076 4573
rect 33048 4564 33100 4616
rect 34244 4607 34296 4616
rect 34244 4573 34253 4607
rect 34253 4573 34287 4607
rect 34287 4573 34296 4607
rect 34244 4564 34296 4573
rect 34980 4607 35032 4616
rect 34980 4573 34989 4607
rect 34989 4573 35023 4607
rect 35023 4573 35032 4607
rect 34980 4564 35032 4573
rect 35164 4607 35216 4616
rect 35164 4573 35173 4607
rect 35173 4573 35207 4607
rect 35207 4573 35216 4607
rect 35164 4564 35216 4573
rect 29000 4428 29052 4480
rect 30104 4428 30156 4480
rect 35532 4428 35584 4480
rect 36268 4428 36320 4480
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 34966 4326 35018 4378
rect 35030 4326 35082 4378
rect 35094 4326 35146 4378
rect 35158 4326 35210 4378
rect 27988 4224 28040 4276
rect 33784 4267 33836 4276
rect 33784 4233 33793 4267
rect 33793 4233 33827 4267
rect 33827 4233 33836 4267
rect 33784 4224 33836 4233
rect 34704 4267 34756 4276
rect 34704 4233 34713 4267
rect 34713 4233 34747 4267
rect 34747 4233 34756 4267
rect 34704 4224 34756 4233
rect 27896 4156 27948 4208
rect 27988 4088 28040 4140
rect 28172 4088 28224 4140
rect 28724 4088 28776 4140
rect 29000 4020 29052 4072
rect 29276 4063 29328 4072
rect 29276 4029 29285 4063
rect 29285 4029 29319 4063
rect 29319 4029 29328 4063
rect 29276 4020 29328 4029
rect 31116 4088 31168 4140
rect 30288 4020 30340 4072
rect 30748 4020 30800 4072
rect 31760 4063 31812 4072
rect 26792 3927 26844 3936
rect 26792 3893 26801 3927
rect 26801 3893 26835 3927
rect 26835 3893 26844 3927
rect 26792 3884 26844 3893
rect 28908 3952 28960 4004
rect 31208 3995 31260 4004
rect 31208 3961 31217 3995
rect 31217 3961 31251 3995
rect 31251 3961 31260 3995
rect 31208 3952 31260 3961
rect 31760 4029 31769 4063
rect 31769 4029 31803 4063
rect 31803 4029 31812 4063
rect 31760 4020 31812 4029
rect 35532 4020 35584 4072
rect 34796 3952 34848 4004
rect 35808 3952 35860 4004
rect 27988 3927 28040 3936
rect 27988 3893 27997 3927
rect 27997 3893 28031 3927
rect 28031 3893 28040 3927
rect 27988 3884 28040 3893
rect 29368 3884 29420 3936
rect 30656 3927 30708 3936
rect 30656 3893 30665 3927
rect 30665 3893 30699 3927
rect 30699 3893 30708 3927
rect 30656 3884 30708 3893
rect 33140 3927 33192 3936
rect 33140 3893 33149 3927
rect 33149 3893 33183 3927
rect 33183 3893 33192 3927
rect 33140 3884 33192 3893
rect 34152 3927 34204 3936
rect 34152 3893 34161 3927
rect 34161 3893 34195 3927
rect 34195 3893 34204 3927
rect 34152 3884 34204 3893
rect 36820 3927 36872 3936
rect 36820 3893 36829 3927
rect 36829 3893 36863 3927
rect 36863 3893 36872 3927
rect 36820 3884 36872 3893
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 27344 3723 27396 3732
rect 27344 3689 27353 3723
rect 27353 3689 27387 3723
rect 27387 3689 27396 3723
rect 27344 3680 27396 3689
rect 28448 3723 28500 3732
rect 28448 3689 28457 3723
rect 28457 3689 28491 3723
rect 28491 3689 28500 3723
rect 28448 3680 28500 3689
rect 26792 3612 26844 3664
rect 27712 3587 27764 3596
rect 27712 3553 27721 3587
rect 27721 3553 27755 3587
rect 27755 3553 27764 3587
rect 27712 3544 27764 3553
rect 27804 3519 27856 3528
rect 27804 3485 27813 3519
rect 27813 3485 27847 3519
rect 27847 3485 27856 3519
rect 27804 3476 27856 3485
rect 29276 3680 29328 3732
rect 29368 3680 29420 3732
rect 31024 3680 31076 3732
rect 35532 3680 35584 3732
rect 35900 3723 35952 3732
rect 35900 3689 35909 3723
rect 35909 3689 35943 3723
rect 35943 3689 35952 3723
rect 35900 3680 35952 3689
rect 29000 3612 29052 3664
rect 30656 3612 30708 3664
rect 34704 3612 34756 3664
rect 36820 3612 36872 3664
rect 32404 3544 32456 3596
rect 33048 3544 33100 3596
rect 33692 3587 33744 3596
rect 33692 3553 33726 3587
rect 33726 3553 33744 3587
rect 33692 3544 33744 3553
rect 36268 3587 36320 3596
rect 36268 3553 36277 3587
rect 36277 3553 36311 3587
rect 36311 3553 36320 3587
rect 36268 3544 36320 3553
rect 28172 3476 28224 3528
rect 31760 3476 31812 3528
rect 33416 3519 33468 3528
rect 33416 3485 33425 3519
rect 33425 3485 33459 3519
rect 33459 3485 33468 3519
rect 33416 3476 33468 3485
rect 36452 3519 36504 3528
rect 36452 3485 36461 3519
rect 36461 3485 36495 3519
rect 36495 3485 36504 3519
rect 36452 3476 36504 3485
rect 32496 3451 32548 3460
rect 32496 3417 32505 3451
rect 32505 3417 32539 3451
rect 32539 3417 32548 3451
rect 32496 3408 32548 3417
rect 30748 3340 30800 3392
rect 34612 3340 34664 3392
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 34966 3238 35018 3290
rect 35030 3238 35082 3290
rect 35094 3238 35146 3290
rect 35158 3238 35210 3290
rect 27804 3136 27856 3188
rect 29000 3179 29052 3188
rect 29000 3145 29009 3179
rect 29009 3145 29043 3179
rect 29043 3145 29052 3179
rect 29000 3136 29052 3145
rect 31576 3179 31628 3188
rect 31576 3145 31585 3179
rect 31585 3145 31619 3179
rect 31619 3145 31628 3179
rect 31576 3136 31628 3145
rect 32036 3136 32088 3188
rect 36268 3136 36320 3188
rect 27712 3068 27764 3120
rect 36820 3111 36872 3120
rect 36820 3077 36829 3111
rect 36829 3077 36863 3111
rect 36863 3077 36872 3111
rect 36820 3068 36872 3077
rect 28080 3043 28132 3052
rect 28080 3009 28089 3043
rect 28089 3009 28123 3043
rect 28123 3009 28132 3043
rect 28080 3000 28132 3009
rect 28172 3043 28224 3052
rect 28172 3009 28181 3043
rect 28181 3009 28215 3043
rect 28215 3009 28224 3043
rect 31300 3043 31352 3052
rect 28172 3000 28224 3009
rect 31300 3009 31309 3043
rect 31309 3009 31343 3043
rect 31343 3009 31352 3043
rect 31760 3043 31812 3052
rect 31300 3000 31352 3009
rect 31760 3009 31769 3043
rect 31769 3009 31803 3043
rect 31803 3009 31812 3043
rect 31760 3000 31812 3009
rect 33692 3043 33744 3052
rect 33692 3009 33701 3043
rect 33701 3009 33735 3043
rect 33735 3009 33744 3043
rect 33692 3000 33744 3009
rect 36452 3000 36504 3052
rect 29276 2975 29328 2984
rect 29276 2941 29285 2975
rect 29285 2941 29319 2975
rect 29319 2941 29328 2975
rect 29276 2932 29328 2941
rect 32036 2975 32088 2984
rect 32036 2941 32070 2975
rect 32070 2941 32088 2975
rect 32036 2932 32088 2941
rect 33140 2932 33192 2984
rect 33416 2932 33468 2984
rect 34520 2932 34572 2984
rect 35532 2932 35584 2984
rect 29368 2864 29420 2916
rect 27620 2839 27672 2848
rect 27620 2805 27629 2839
rect 27629 2805 27663 2839
rect 27663 2805 27672 2839
rect 27620 2796 27672 2805
rect 27988 2839 28040 2848
rect 27988 2805 27997 2839
rect 27997 2805 28031 2839
rect 28031 2805 28040 2839
rect 27988 2796 28040 2805
rect 30288 2796 30340 2848
rect 31208 2796 31260 2848
rect 33048 2796 33100 2848
rect 34612 2839 34664 2848
rect 34612 2805 34621 2839
rect 34621 2805 34655 2839
rect 34655 2805 34664 2839
rect 34612 2796 34664 2805
rect 35808 2796 35860 2848
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 27988 2592 28040 2644
rect 28172 2592 28224 2644
rect 29368 2635 29420 2644
rect 29368 2601 29377 2635
rect 29377 2601 29411 2635
rect 29411 2601 29420 2635
rect 29368 2592 29420 2601
rect 30748 2592 30800 2644
rect 31944 2635 31996 2644
rect 31944 2601 31953 2635
rect 31953 2601 31987 2635
rect 31987 2601 31996 2635
rect 31944 2592 31996 2601
rect 32404 2635 32456 2644
rect 32404 2601 32413 2635
rect 32413 2601 32447 2635
rect 32447 2601 32456 2635
rect 32404 2592 32456 2601
rect 33692 2592 33744 2644
rect 34520 2635 34572 2644
rect 34520 2601 34529 2635
rect 34529 2601 34563 2635
rect 34563 2601 34572 2635
rect 34520 2592 34572 2601
rect 35256 2635 35308 2644
rect 35256 2601 35265 2635
rect 35265 2601 35299 2635
rect 35299 2601 35308 2635
rect 35256 2592 35308 2601
rect 35992 2592 36044 2644
rect 30288 2524 30340 2576
rect 33048 2524 33100 2576
rect 35808 2524 35860 2576
rect 29276 2456 29328 2508
rect 31300 2456 31352 2508
rect 33416 2456 33468 2508
rect 35532 2456 35584 2508
rect 9956 2252 10008 2304
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 34966 2150 35018 2202
rect 35030 2150 35082 2202
rect 35094 2150 35146 2202
rect 35158 2150 35210 2202
<< metal2 >>
rect 570 39520 626 40000
rect 1674 39520 1730 40000
rect 2778 39520 2834 40000
rect 3882 39520 3938 40000
rect 4986 39520 5042 40000
rect 6090 39520 6146 40000
rect 7194 39520 7250 40000
rect 8298 39520 8354 40000
rect 9402 39520 9458 40000
rect 10506 39520 10562 40000
rect 11610 39520 11666 40000
rect 12714 39520 12770 40000
rect 13910 39520 13966 40000
rect 15014 39520 15070 40000
rect 16118 39520 16174 40000
rect 17222 39520 17278 40000
rect 18326 39520 18382 40000
rect 19430 39520 19486 40000
rect 20534 39520 20590 40000
rect 21638 39520 21694 40000
rect 22742 39520 22798 40000
rect 23846 39520 23902 40000
rect 24950 39520 25006 40000
rect 26054 39522 26110 40000
rect 26054 39520 26188 39522
rect 27250 39520 27306 40000
rect 28354 39520 28410 40000
rect 29458 39520 29514 40000
rect 30562 39520 30618 40000
rect 31666 39520 31722 40000
rect 32770 39520 32826 40000
rect 33874 39520 33930 40000
rect 34978 39520 35034 40000
rect 36082 39520 36138 40000
rect 37186 39520 37242 40000
rect 38290 39520 38346 40000
rect 39394 39520 39450 40000
rect 584 34746 612 39520
rect 1398 35320 1454 35329
rect 1688 35290 1716 39520
rect 1398 35255 1454 35264
rect 1676 35284 1728 35290
rect 1412 35154 1440 35255
rect 1676 35226 1728 35232
rect 1400 35148 1452 35154
rect 1400 35090 1452 35096
rect 572 34740 624 34746
rect 572 34682 624 34688
rect 1412 34202 1440 35090
rect 2042 35048 2098 35057
rect 2042 34983 2098 34992
rect 2056 34746 2084 34983
rect 2044 34740 2096 34746
rect 2044 34682 2096 34688
rect 2056 34542 2084 34682
rect 2688 34672 2740 34678
rect 2792 34626 2820 39520
rect 3146 36136 3202 36145
rect 3146 36071 3202 36080
rect 3160 34746 3188 36071
rect 3896 34898 3924 39520
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4220 36944 4516 36964
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4220 35856 4516 35876
rect 5000 35834 5028 39520
rect 6104 36378 6132 39520
rect 7208 36378 7236 39520
rect 6092 36372 6144 36378
rect 6092 36314 6144 36320
rect 7196 36372 7248 36378
rect 7196 36314 7248 36320
rect 5448 36236 5500 36242
rect 5448 36178 5500 36184
rect 6644 36236 6696 36242
rect 6644 36178 6696 36184
rect 5460 35986 5488 36178
rect 5460 35958 5580 35986
rect 4988 35828 5040 35834
rect 4988 35770 5040 35776
rect 5264 35760 5316 35766
rect 5264 35702 5316 35708
rect 4988 35488 5040 35494
rect 4986 35456 4988 35465
rect 5040 35456 5042 35465
rect 4986 35391 5042 35400
rect 4988 35148 5040 35154
rect 4988 35090 5040 35096
rect 4712 35012 4764 35018
rect 4712 34954 4764 34960
rect 3896 34870 4108 34898
rect 3148 34740 3200 34746
rect 3148 34682 3200 34688
rect 2740 34620 2820 34626
rect 2688 34614 2820 34620
rect 2700 34598 2820 34614
rect 3160 34542 3188 34682
rect 4080 34626 4108 34870
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4220 34768 4516 34788
rect 4080 34598 4200 34626
rect 2044 34536 2096 34542
rect 2044 34478 2096 34484
rect 3148 34536 3200 34542
rect 3148 34478 3200 34484
rect 4172 34202 4200 34598
rect 4620 34536 4672 34542
rect 4620 34478 4672 34484
rect 1400 34196 1452 34202
rect 1400 34138 1452 34144
rect 4160 34196 4212 34202
rect 4160 34138 4212 34144
rect 4068 34060 4120 34066
rect 4068 34002 4120 34008
rect 3976 33992 4028 33998
rect 4080 33969 4108 34002
rect 3976 33934 4028 33940
rect 4066 33960 4122 33969
rect 3988 33538 4016 33934
rect 4066 33895 4122 33904
rect 4080 33658 4108 33895
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4220 33680 4516 33700
rect 4068 33652 4120 33658
rect 4068 33594 4120 33600
rect 3988 33522 4108 33538
rect 3988 33516 4120 33522
rect 3988 33510 4068 33516
rect 4068 33458 4120 33464
rect 4080 32978 4108 33458
rect 4528 33380 4580 33386
rect 4528 33322 4580 33328
rect 4540 33114 4568 33322
rect 4528 33108 4580 33114
rect 4528 33050 4580 33056
rect 4632 33046 4660 34478
rect 4724 34406 4752 34954
rect 4712 34400 4764 34406
rect 4712 34342 4764 34348
rect 4724 33386 4752 34342
rect 5000 34134 5028 35090
rect 5276 35086 5304 35702
rect 5552 35494 5580 35958
rect 6656 35766 6684 36178
rect 7470 35864 7526 35873
rect 6828 35828 6880 35834
rect 8312 35850 8340 39520
rect 8220 35834 8340 35850
rect 7470 35799 7472 35808
rect 6828 35770 6880 35776
rect 7524 35799 7526 35808
rect 8208 35828 8340 35834
rect 7472 35770 7524 35776
rect 8260 35822 8340 35828
rect 8208 35770 8260 35776
rect 6644 35760 6696 35766
rect 6642 35728 6644 35737
rect 6840 35737 6868 35770
rect 6696 35728 6698 35737
rect 6642 35663 6698 35672
rect 6826 35728 6882 35737
rect 6826 35663 6882 35672
rect 7484 35630 7512 35770
rect 7472 35624 7524 35630
rect 7472 35566 7524 35572
rect 8574 35592 8630 35601
rect 8574 35527 8576 35536
rect 8628 35527 8630 35536
rect 8576 35498 8628 35504
rect 5540 35488 5592 35494
rect 5538 35456 5540 35465
rect 7472 35488 7524 35494
rect 5592 35456 5594 35465
rect 7472 35430 7524 35436
rect 5538 35391 5594 35400
rect 6826 35184 6882 35193
rect 6826 35119 6828 35128
rect 6880 35119 6882 35128
rect 6828 35090 6880 35096
rect 5080 35080 5132 35086
rect 5080 35022 5132 35028
rect 5264 35080 5316 35086
rect 5264 35022 5316 35028
rect 5092 34746 5120 35022
rect 5080 34740 5132 34746
rect 5080 34682 5132 34688
rect 5078 34640 5134 34649
rect 5078 34575 5080 34584
rect 5132 34575 5134 34584
rect 5080 34546 5132 34552
rect 4988 34128 5040 34134
rect 4988 34070 5040 34076
rect 4712 33380 4764 33386
rect 4712 33322 4764 33328
rect 4620 33040 4672 33046
rect 4620 32982 4672 32988
rect 4068 32972 4120 32978
rect 4068 32914 4120 32920
rect 3148 32768 3200 32774
rect 3148 32710 3200 32716
rect 3160 32434 3188 32710
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 4632 32570 4660 32982
rect 4620 32564 4672 32570
rect 4620 32506 4672 32512
rect 3148 32428 3200 32434
rect 3148 32370 3200 32376
rect 2044 32224 2096 32230
rect 2044 32166 2096 32172
rect 2596 32224 2648 32230
rect 2596 32166 2648 32172
rect 2056 31890 2084 32166
rect 2044 31884 2096 31890
rect 2044 31826 2096 31832
rect 1676 31680 1728 31686
rect 1676 31622 1728 31628
rect 1400 31272 1452 31278
rect 1400 31214 1452 31220
rect 1412 30734 1440 31214
rect 1688 31142 1716 31622
rect 1676 31136 1728 31142
rect 1676 31078 1728 31084
rect 1400 30728 1452 30734
rect 1400 30670 1452 30676
rect 1412 30190 1440 30670
rect 1400 30184 1452 30190
rect 1400 30126 1452 30132
rect 1412 29646 1440 30126
rect 1688 30122 1716 31078
rect 2056 30802 2084 31826
rect 2608 31822 2636 32166
rect 2870 32056 2926 32065
rect 3160 32026 3188 32370
rect 3608 32292 3660 32298
rect 3608 32234 3660 32240
rect 3620 32026 3648 32234
rect 4986 32056 5042 32065
rect 2870 31991 2872 32000
rect 2924 31991 2926 32000
rect 3148 32020 3200 32026
rect 2872 31962 2924 31968
rect 3148 31962 3200 31968
rect 3608 32020 3660 32026
rect 4986 31991 4988 32000
rect 3608 31962 3660 31968
rect 5040 31991 5042 32000
rect 4988 31962 5040 31968
rect 2780 31952 2832 31958
rect 2780 31894 2832 31900
rect 2596 31816 2648 31822
rect 2596 31758 2648 31764
rect 2792 31278 2820 31894
rect 3620 31482 3648 31962
rect 4620 31952 4672 31958
rect 5092 31906 5120 34546
rect 5276 33862 5304 35022
rect 5448 34944 5500 34950
rect 5448 34886 5500 34892
rect 5264 33856 5316 33862
rect 5264 33798 5316 33804
rect 5172 32020 5224 32026
rect 5172 31962 5224 31968
rect 4620 31894 4672 31900
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4220 31504 4516 31524
rect 3608 31476 3660 31482
rect 3608 31418 3660 31424
rect 4632 31414 4660 31894
rect 5000 31878 5120 31906
rect 5000 31754 5028 31878
rect 4988 31748 5040 31754
rect 4988 31690 5040 31696
rect 4620 31408 4672 31414
rect 4620 31350 4672 31356
rect 2780 31272 2832 31278
rect 2780 31214 2832 31220
rect 2872 31204 2924 31210
rect 2872 31146 2924 31152
rect 2884 30938 2912 31146
rect 4712 31136 4764 31142
rect 3330 31104 3386 31113
rect 4712 31078 4764 31084
rect 3330 31039 3386 31048
rect 2872 30932 2924 30938
rect 2872 30874 2924 30880
rect 2044 30796 2096 30802
rect 2044 30738 2096 30744
rect 1676 30116 1728 30122
rect 1676 30058 1728 30064
rect 1688 29850 1716 30058
rect 2056 30054 2084 30738
rect 2044 30048 2096 30054
rect 2044 29990 2096 29996
rect 2964 30048 3016 30054
rect 2964 29990 3016 29996
rect 1676 29844 1728 29850
rect 1676 29786 1728 29792
rect 1674 29744 1730 29753
rect 1674 29679 1676 29688
rect 1728 29679 1730 29688
rect 1676 29650 1728 29656
rect 1400 29640 1452 29646
rect 1400 29582 1452 29588
rect 1412 29170 1440 29582
rect 1688 29306 1716 29650
rect 2056 29306 2084 29990
rect 1676 29300 1728 29306
rect 1676 29242 1728 29248
rect 2044 29300 2096 29306
rect 2044 29242 2096 29248
rect 1400 29164 1452 29170
rect 1400 29106 1452 29112
rect 1952 29164 2004 29170
rect 1952 29106 2004 29112
rect 1964 28762 1992 29106
rect 2688 29096 2740 29102
rect 2688 29038 2740 29044
rect 2700 28762 2728 29038
rect 1952 28756 2004 28762
rect 1952 28698 2004 28704
rect 2688 28756 2740 28762
rect 2688 28698 2740 28704
rect 1860 28552 1912 28558
rect 1860 28494 1912 28500
rect 1872 28218 1900 28494
rect 1860 28212 1912 28218
rect 1860 28154 1912 28160
rect 1872 27674 1900 28154
rect 1964 28082 1992 28698
rect 2780 28620 2832 28626
rect 2780 28562 2832 28568
rect 1952 28076 2004 28082
rect 1952 28018 2004 28024
rect 2688 27940 2740 27946
rect 2688 27882 2740 27888
rect 1860 27668 1912 27674
rect 1860 27610 1912 27616
rect 2228 27600 2280 27606
rect 2228 27542 2280 27548
rect 2136 27532 2188 27538
rect 2136 27474 2188 27480
rect 1768 27464 1820 27470
rect 1768 27406 1820 27412
rect 1780 27130 1808 27406
rect 1952 27396 2004 27402
rect 1952 27338 2004 27344
rect 1768 27124 1820 27130
rect 1768 27066 1820 27072
rect 1492 26920 1544 26926
rect 1492 26862 1544 26868
rect 1504 26450 1532 26862
rect 1780 26518 1808 27066
rect 1964 26926 1992 27338
rect 2148 26926 2176 27474
rect 1952 26920 2004 26926
rect 1952 26862 2004 26868
rect 2136 26920 2188 26926
rect 2136 26862 2188 26868
rect 1768 26512 1820 26518
rect 1768 26454 1820 26460
rect 1492 26444 1544 26450
rect 1492 26386 1544 26392
rect 1780 25770 1808 26454
rect 1768 25764 1820 25770
rect 1768 25706 1820 25712
rect 1964 25702 1992 26862
rect 2148 26586 2176 26862
rect 2136 26580 2188 26586
rect 2136 26522 2188 26528
rect 2240 26042 2268 27542
rect 2700 27010 2728 27882
rect 2792 27674 2820 28562
rect 2976 28558 3004 29990
rect 3344 29306 3372 31039
rect 4724 30870 4752 31078
rect 5000 30938 5028 31690
rect 5080 31680 5132 31686
rect 5080 31622 5132 31628
rect 5092 31278 5120 31622
rect 5184 31346 5212 31962
rect 5276 31686 5304 33798
rect 5460 32450 5488 34886
rect 6840 34746 6868 35090
rect 6920 35012 6972 35018
rect 6920 34954 6972 34960
rect 6828 34740 6880 34746
rect 6828 34682 6880 34688
rect 6932 34542 6960 34954
rect 7104 34944 7156 34950
rect 7104 34886 7156 34892
rect 5632 34536 5684 34542
rect 5632 34478 5684 34484
rect 6920 34536 6972 34542
rect 6920 34478 6972 34484
rect 5540 34060 5592 34066
rect 5540 34002 5592 34008
rect 5552 33658 5580 34002
rect 5540 33652 5592 33658
rect 5540 33594 5592 33600
rect 5644 33538 5672 34478
rect 6276 34400 6328 34406
rect 6276 34342 6328 34348
rect 6288 34202 6316 34342
rect 6276 34196 6328 34202
rect 6276 34138 6328 34144
rect 6828 34128 6880 34134
rect 6828 34070 6880 34076
rect 6840 33658 6868 34070
rect 6828 33652 6880 33658
rect 6828 33594 6880 33600
rect 5552 33510 5672 33538
rect 5552 33454 5580 33510
rect 5540 33448 5592 33454
rect 5540 33390 5592 33396
rect 5552 33114 5580 33390
rect 5540 33108 5592 33114
rect 5540 33050 5592 33056
rect 5552 32570 5580 33050
rect 6920 32972 6972 32978
rect 6920 32914 6972 32920
rect 5540 32564 5592 32570
rect 5540 32506 5592 32512
rect 6460 32564 6512 32570
rect 6460 32506 6512 32512
rect 5460 32422 5580 32450
rect 5552 32366 5580 32422
rect 5540 32360 5592 32366
rect 5540 32302 5592 32308
rect 5816 32224 5868 32230
rect 5816 32166 5868 32172
rect 5828 32026 5856 32166
rect 5816 32020 5868 32026
rect 5816 31962 5868 31968
rect 6184 31884 6236 31890
rect 6184 31826 6236 31832
rect 5816 31816 5868 31822
rect 5816 31758 5868 31764
rect 5264 31680 5316 31686
rect 5264 31622 5316 31628
rect 5276 31346 5304 31622
rect 5172 31340 5224 31346
rect 5172 31282 5224 31288
rect 5264 31340 5316 31346
rect 5264 31282 5316 31288
rect 5080 31272 5132 31278
rect 5080 31214 5132 31220
rect 5092 30938 5120 31214
rect 4988 30932 5040 30938
rect 4988 30874 5040 30880
rect 5080 30932 5132 30938
rect 5080 30874 5132 30880
rect 4712 30864 4764 30870
rect 4712 30806 4764 30812
rect 4804 30796 4856 30802
rect 4804 30738 4856 30744
rect 3976 30660 4028 30666
rect 3976 30602 4028 30608
rect 3988 30054 4016 30602
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 4816 30394 4844 30738
rect 4896 30728 4948 30734
rect 4896 30670 4948 30676
rect 4804 30388 4856 30394
rect 4804 30330 4856 30336
rect 3976 30048 4028 30054
rect 3976 29990 4028 29996
rect 4160 30048 4212 30054
rect 4160 29990 4212 29996
rect 4172 29753 4200 29990
rect 4908 29850 4936 30670
rect 5000 30258 5028 30874
rect 5276 30734 5304 31282
rect 5828 31142 5856 31758
rect 6196 31142 6224 31826
rect 5816 31136 5868 31142
rect 5814 31104 5816 31113
rect 6184 31136 6236 31142
rect 5868 31104 5870 31113
rect 6184 31078 6236 31084
rect 5814 31039 5870 31048
rect 6472 30938 6500 32506
rect 6932 32502 6960 32914
rect 7116 32910 7144 34886
rect 7484 34649 7512 35430
rect 8852 35216 8904 35222
rect 9416 35193 9444 39520
rect 10520 35737 10548 39520
rect 11624 35873 11652 39520
rect 11610 35864 11666 35873
rect 11610 35799 11666 35808
rect 11886 35864 11942 35873
rect 11886 35799 11888 35808
rect 11940 35799 11942 35808
rect 11888 35770 11940 35776
rect 10506 35728 10562 35737
rect 10506 35663 10562 35672
rect 11900 35630 11928 35770
rect 11888 35624 11940 35630
rect 11888 35566 11940 35572
rect 11060 35488 11112 35494
rect 11060 35430 11112 35436
rect 10874 35320 10930 35329
rect 10874 35255 10876 35264
rect 10928 35255 10930 35264
rect 10876 35226 10928 35232
rect 8852 35158 8904 35164
rect 9402 35184 9458 35193
rect 8300 35148 8352 35154
rect 8300 35090 8352 35096
rect 8312 34678 8340 35090
rect 8484 34944 8536 34950
rect 8484 34886 8536 34892
rect 8300 34672 8352 34678
rect 7470 34640 7526 34649
rect 8300 34614 8352 34620
rect 7470 34575 7526 34584
rect 7196 34196 7248 34202
rect 7196 34138 7248 34144
rect 7208 33454 7236 34138
rect 7484 33930 7512 34575
rect 8208 34536 8260 34542
rect 8208 34478 8260 34484
rect 7932 34060 7984 34066
rect 7932 34002 7984 34008
rect 7472 33924 7524 33930
rect 7472 33866 7524 33872
rect 7484 33522 7512 33866
rect 7472 33516 7524 33522
rect 7472 33458 7524 33464
rect 7196 33448 7248 33454
rect 7196 33390 7248 33396
rect 7944 33318 7972 34002
rect 8024 33856 8076 33862
rect 8024 33798 8076 33804
rect 7932 33312 7984 33318
rect 7932 33254 7984 33260
rect 7012 32904 7064 32910
rect 7012 32846 7064 32852
rect 7104 32904 7156 32910
rect 7104 32846 7156 32852
rect 7024 32570 7052 32846
rect 7012 32564 7064 32570
rect 7012 32506 7064 32512
rect 6920 32496 6972 32502
rect 6920 32438 6972 32444
rect 7116 32026 7144 32846
rect 7748 32224 7800 32230
rect 7748 32166 7800 32172
rect 6552 32020 6604 32026
rect 6552 31962 6604 31968
rect 7104 32020 7156 32026
rect 7104 31962 7156 31968
rect 6564 31822 6592 31962
rect 7760 31890 7788 32166
rect 7748 31884 7800 31890
rect 7748 31826 7800 31832
rect 6552 31816 6604 31822
rect 6552 31758 6604 31764
rect 6564 31482 6592 31758
rect 7944 31482 7972 33254
rect 8036 33153 8064 33798
rect 8220 33674 8248 34478
rect 8300 33856 8352 33862
rect 8300 33798 8352 33804
rect 8312 33674 8340 33798
rect 8220 33658 8340 33674
rect 8220 33652 8352 33658
rect 8220 33646 8300 33652
rect 8300 33594 8352 33600
rect 8022 33144 8078 33153
rect 8022 33079 8078 33088
rect 8496 32978 8524 34886
rect 8864 34785 8892 35158
rect 9402 35119 9458 35128
rect 10048 35080 10100 35086
rect 10888 35057 10916 35226
rect 10048 35022 10100 35028
rect 10874 35048 10930 35057
rect 9864 34944 9916 34950
rect 9864 34886 9916 34892
rect 8850 34776 8906 34785
rect 8850 34711 8852 34720
rect 8904 34711 8906 34720
rect 8852 34682 8904 34688
rect 9876 34542 9904 34886
rect 9864 34536 9916 34542
rect 9864 34478 9916 34484
rect 9772 34400 9824 34406
rect 9772 34342 9824 34348
rect 9784 34066 9812 34342
rect 9876 34134 9904 34478
rect 9864 34128 9916 34134
rect 9864 34070 9916 34076
rect 8668 34060 8720 34066
rect 8668 34002 8720 34008
rect 9772 34060 9824 34066
rect 9772 34002 9824 34008
rect 8576 33516 8628 33522
rect 8576 33458 8628 33464
rect 8484 32972 8536 32978
rect 8484 32914 8536 32920
rect 8116 32768 8168 32774
rect 8116 32710 8168 32716
rect 8300 32768 8352 32774
rect 8300 32710 8352 32716
rect 8128 32366 8156 32710
rect 8312 32434 8340 32710
rect 8300 32428 8352 32434
rect 8300 32370 8352 32376
rect 8116 32360 8168 32366
rect 8116 32302 8168 32308
rect 8024 32292 8076 32298
rect 8024 32234 8076 32240
rect 6552 31476 6604 31482
rect 6552 31418 6604 31424
rect 7932 31476 7984 31482
rect 7932 31418 7984 31424
rect 8036 31278 8064 32234
rect 8496 32026 8524 32914
rect 8484 32020 8536 32026
rect 8484 31962 8536 31968
rect 8300 31884 8352 31890
rect 8300 31826 8352 31832
rect 8312 31482 8340 31826
rect 8300 31476 8352 31482
rect 8300 31418 8352 31424
rect 8024 31272 8076 31278
rect 8024 31214 8076 31220
rect 6828 31136 6880 31142
rect 6828 31078 6880 31084
rect 6460 30932 6512 30938
rect 6460 30874 6512 30880
rect 6000 30796 6052 30802
rect 6000 30738 6052 30744
rect 5264 30728 5316 30734
rect 5264 30670 5316 30676
rect 5356 30592 5408 30598
rect 5408 30552 5488 30580
rect 5356 30534 5408 30540
rect 5460 30274 5488 30552
rect 6012 30394 6040 30738
rect 6840 30394 6868 31078
rect 8392 30796 8444 30802
rect 8392 30738 8444 30744
rect 8116 30660 8168 30666
rect 8116 30602 8168 30608
rect 8024 30592 8076 30598
rect 8024 30534 8076 30540
rect 6000 30388 6052 30394
rect 6000 30330 6052 30336
rect 6828 30388 6880 30394
rect 6828 30330 6880 30336
rect 4988 30252 5040 30258
rect 4988 30194 5040 30200
rect 5356 30252 5408 30258
rect 5460 30246 5580 30274
rect 5356 30194 5408 30200
rect 5080 30116 5132 30122
rect 5080 30058 5132 30064
rect 4896 29844 4948 29850
rect 4896 29786 4948 29792
rect 4158 29744 4214 29753
rect 4158 29679 4214 29688
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4220 29328 4516 29348
rect 3332 29300 3384 29306
rect 3332 29242 3384 29248
rect 4068 29096 4120 29102
rect 4068 29038 4120 29044
rect 4080 28626 4108 29038
rect 3884 28620 3936 28626
rect 3884 28562 3936 28568
rect 4068 28620 4120 28626
rect 4068 28562 4120 28568
rect 4620 28620 4672 28626
rect 4620 28562 4672 28568
rect 2964 28552 3016 28558
rect 2964 28494 3016 28500
rect 2780 27668 2832 27674
rect 2780 27610 2832 27616
rect 3896 27606 3924 28562
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 4632 27946 4660 28562
rect 4908 28218 4936 29786
rect 5092 29782 5120 30058
rect 5080 29776 5132 29782
rect 5080 29718 5132 29724
rect 5092 29322 5120 29718
rect 5264 29708 5316 29714
rect 5264 29650 5316 29656
rect 5092 29306 5212 29322
rect 5092 29300 5224 29306
rect 5092 29294 5172 29300
rect 5172 29242 5224 29248
rect 5276 29102 5304 29650
rect 5264 29096 5316 29102
rect 5264 29038 5316 29044
rect 5276 28626 5304 29038
rect 5264 28620 5316 28626
rect 5264 28562 5316 28568
rect 4896 28212 4948 28218
rect 4896 28154 4948 28160
rect 5368 28082 5396 30194
rect 5552 30190 5580 30246
rect 5540 30184 5592 30190
rect 5540 30126 5592 30132
rect 7932 30116 7984 30122
rect 7932 30058 7984 30064
rect 5540 30048 5592 30054
rect 5540 29990 5592 29996
rect 5552 29850 5580 29990
rect 7944 29850 7972 30058
rect 5540 29844 5592 29850
rect 5540 29786 5592 29792
rect 7932 29844 7984 29850
rect 7932 29786 7984 29792
rect 7104 29776 7156 29782
rect 7104 29718 7156 29724
rect 7116 29306 7144 29718
rect 8036 29646 8064 30534
rect 7472 29640 7524 29646
rect 7472 29582 7524 29588
rect 8024 29640 8076 29646
rect 8024 29582 8076 29588
rect 7484 29306 7512 29582
rect 7840 29504 7892 29510
rect 7840 29446 7892 29452
rect 8024 29504 8076 29510
rect 8024 29446 8076 29452
rect 7104 29300 7156 29306
rect 7104 29242 7156 29248
rect 7472 29300 7524 29306
rect 7472 29242 7524 29248
rect 7852 29186 7880 29446
rect 7930 29200 7986 29209
rect 7852 29158 7930 29186
rect 7930 29135 7986 29144
rect 7944 29102 7972 29135
rect 7932 29096 7984 29102
rect 7932 29038 7984 29044
rect 5448 29028 5500 29034
rect 5448 28970 5500 28976
rect 5460 28762 5488 28970
rect 5448 28756 5500 28762
rect 5448 28698 5500 28704
rect 5356 28076 5408 28082
rect 5356 28018 5408 28024
rect 4620 27940 4672 27946
rect 4620 27882 4672 27888
rect 4160 27872 4212 27878
rect 4160 27814 4212 27820
rect 4068 27668 4120 27674
rect 4068 27610 4120 27616
rect 3884 27600 3936 27606
rect 3884 27542 3936 27548
rect 3974 27432 4030 27441
rect 3974 27367 3976 27376
rect 4028 27367 4030 27376
rect 3976 27338 4028 27344
rect 2780 27124 2832 27130
rect 2780 27066 2832 27072
rect 2792 27010 2820 27066
rect 4080 27062 4108 27610
rect 4172 27606 4200 27814
rect 4160 27600 4212 27606
rect 4160 27542 4212 27548
rect 4620 27600 4672 27606
rect 4620 27542 4672 27548
rect 4220 27228 4516 27248
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 2700 26982 2820 27010
rect 4068 27056 4120 27062
rect 4068 26998 4120 27004
rect 4632 26926 4660 27542
rect 5368 27538 5396 28018
rect 5460 28014 5488 28698
rect 7564 28688 7616 28694
rect 7564 28630 7616 28636
rect 6644 28620 6696 28626
rect 6644 28562 6696 28568
rect 6656 28218 6684 28562
rect 6644 28212 6696 28218
rect 6644 28154 6696 28160
rect 5448 28008 5500 28014
rect 5448 27950 5500 27956
rect 7576 27878 7604 28630
rect 7944 28626 7972 29038
rect 8036 28665 8064 29446
rect 8022 28656 8078 28665
rect 7932 28620 7984 28626
rect 8022 28591 8078 28600
rect 7932 28562 7984 28568
rect 8128 28082 8156 30602
rect 8208 30320 8260 30326
rect 8208 30262 8260 30268
rect 8220 29102 8248 30262
rect 8404 30122 8432 30738
rect 8484 30728 8536 30734
rect 8484 30670 8536 30676
rect 8496 30394 8524 30670
rect 8484 30388 8536 30394
rect 8484 30330 8536 30336
rect 8588 30258 8616 33458
rect 8680 33114 8708 34002
rect 9036 33992 9088 33998
rect 9036 33934 9088 33940
rect 9048 33454 9076 33934
rect 9876 33590 9904 34070
rect 9864 33584 9916 33590
rect 9864 33526 9916 33532
rect 8852 33448 8904 33454
rect 8852 33390 8904 33396
rect 9036 33448 9088 33454
rect 9036 33390 9088 33396
rect 8668 33108 8720 33114
rect 8668 33050 8720 33056
rect 8680 31958 8708 33050
rect 8864 33046 8892 33390
rect 9048 33114 9076 33390
rect 9036 33108 9088 33114
rect 9036 33050 9088 33056
rect 10060 33046 10088 35022
rect 10874 34983 10930 34992
rect 10140 34468 10192 34474
rect 10140 34410 10192 34416
rect 10152 33658 10180 34410
rect 10692 34060 10744 34066
rect 10692 34002 10744 34008
rect 10704 33658 10732 34002
rect 10140 33652 10192 33658
rect 10140 33594 10192 33600
rect 10692 33652 10744 33658
rect 10692 33594 10744 33600
rect 10152 33402 10180 33594
rect 10152 33374 10272 33402
rect 10138 33144 10194 33153
rect 10138 33079 10140 33088
rect 10192 33079 10194 33088
rect 10140 33050 10192 33056
rect 8852 33040 8904 33046
rect 8852 32982 8904 32988
rect 9220 33040 9272 33046
rect 9220 32982 9272 32988
rect 10048 33040 10100 33046
rect 10048 32982 10100 32988
rect 8668 31952 8720 31958
rect 8668 31894 8720 31900
rect 9232 31890 9260 32982
rect 10060 32570 10088 32982
rect 10048 32564 10100 32570
rect 10048 32506 10100 32512
rect 9496 32496 9548 32502
rect 9494 32464 9496 32473
rect 9548 32464 9550 32473
rect 9494 32399 9550 32408
rect 9864 32224 9916 32230
rect 9864 32166 9916 32172
rect 9588 32020 9640 32026
rect 9588 31962 9640 31968
rect 9220 31884 9272 31890
rect 9220 31826 9272 31832
rect 8852 31340 8904 31346
rect 8852 31282 8904 31288
rect 8668 31136 8720 31142
rect 8668 31078 8720 31084
rect 8576 30252 8628 30258
rect 8576 30194 8628 30200
rect 8392 30116 8444 30122
rect 8392 30058 8444 30064
rect 8588 29850 8616 30194
rect 8576 29844 8628 29850
rect 8576 29786 8628 29792
rect 8680 29782 8708 31078
rect 8864 30734 8892 31282
rect 9600 30734 9628 31962
rect 9876 31890 9904 32166
rect 10152 32026 10180 33050
rect 10244 32910 10272 33374
rect 10232 32904 10284 32910
rect 10232 32846 10284 32852
rect 10244 32570 10272 32846
rect 10874 32736 10930 32745
rect 10874 32671 10930 32680
rect 10232 32564 10284 32570
rect 10232 32506 10284 32512
rect 10888 32366 10916 32671
rect 10876 32360 10928 32366
rect 10876 32302 10928 32308
rect 10888 32026 10916 32302
rect 10140 32020 10192 32026
rect 10140 31962 10192 31968
rect 10876 32020 10928 32026
rect 10876 31962 10928 31968
rect 9864 31884 9916 31890
rect 9864 31826 9916 31832
rect 9680 31136 9732 31142
rect 9680 31078 9732 31084
rect 9692 30802 9720 31078
rect 9876 30938 9904 31826
rect 10416 31340 10468 31346
rect 10416 31282 10468 31288
rect 9956 31204 10008 31210
rect 9956 31146 10008 31152
rect 9864 30932 9916 30938
rect 9864 30874 9916 30880
rect 9680 30796 9732 30802
rect 9680 30738 9732 30744
rect 8852 30728 8904 30734
rect 8852 30670 8904 30676
rect 9588 30728 9640 30734
rect 9588 30670 9640 30676
rect 9968 30394 9996 31146
rect 10428 31142 10456 31282
rect 10416 31136 10468 31142
rect 10414 31104 10416 31113
rect 10468 31104 10470 31113
rect 10414 31039 10470 31048
rect 10600 30796 10652 30802
rect 10600 30738 10652 30744
rect 10508 30728 10560 30734
rect 10508 30670 10560 30676
rect 9956 30388 10008 30394
rect 9956 30330 10008 30336
rect 9312 30116 9364 30122
rect 9312 30058 9364 30064
rect 8668 29776 8720 29782
rect 8668 29718 8720 29724
rect 8668 29640 8720 29646
rect 8668 29582 8720 29588
rect 8208 29096 8260 29102
rect 8260 29056 8340 29084
rect 8208 29038 8260 29044
rect 8312 28762 8340 29056
rect 8300 28756 8352 28762
rect 8300 28698 8352 28704
rect 8116 28076 8168 28082
rect 8116 28018 8168 28024
rect 5448 27872 5500 27878
rect 5448 27814 5500 27820
rect 7288 27872 7340 27878
rect 7288 27814 7340 27820
rect 7472 27872 7524 27878
rect 7472 27814 7524 27820
rect 7564 27872 7616 27878
rect 7564 27814 7616 27820
rect 5460 27674 5488 27814
rect 5448 27668 5500 27674
rect 5448 27610 5500 27616
rect 5356 27532 5408 27538
rect 5356 27474 5408 27480
rect 5368 27130 5396 27474
rect 5722 27432 5778 27441
rect 5722 27367 5778 27376
rect 5736 27130 5764 27367
rect 5356 27124 5408 27130
rect 5356 27066 5408 27072
rect 5724 27124 5776 27130
rect 5724 27066 5776 27072
rect 6920 26988 6972 26994
rect 6920 26930 6972 26936
rect 4620 26920 4672 26926
rect 4620 26862 4672 26868
rect 4632 26586 4660 26862
rect 6458 26752 6514 26761
rect 6458 26687 6514 26696
rect 6472 26586 6500 26687
rect 6932 26586 6960 26930
rect 7300 26858 7328 27814
rect 7484 27674 7512 27814
rect 7472 27668 7524 27674
rect 7472 27610 7524 27616
rect 7576 27334 7604 27814
rect 8128 27606 8156 28018
rect 8208 28008 8260 28014
rect 8208 27950 8260 27956
rect 8116 27600 8168 27606
rect 8116 27542 8168 27548
rect 7564 27328 7616 27334
rect 7564 27270 7616 27276
rect 7576 27130 7604 27270
rect 7564 27124 7616 27130
rect 7564 27066 7616 27072
rect 8128 27010 8156 27542
rect 8220 27402 8248 27950
rect 8680 27470 8708 29582
rect 9324 29306 9352 30058
rect 9968 29782 9996 30330
rect 10520 30122 10548 30670
rect 10508 30116 10560 30122
rect 10508 30058 10560 30064
rect 10414 30016 10470 30025
rect 10414 29951 10470 29960
rect 9956 29776 10008 29782
rect 9956 29718 10008 29724
rect 9680 29708 9732 29714
rect 9680 29650 9732 29656
rect 9312 29300 9364 29306
rect 9312 29242 9364 29248
rect 9692 29209 9720 29650
rect 9968 29306 9996 29718
rect 10428 29306 10456 29951
rect 10520 29714 10548 30058
rect 10612 30054 10640 30738
rect 10600 30048 10652 30054
rect 10600 29990 10652 29996
rect 10612 29850 10640 29990
rect 10600 29844 10652 29850
rect 10600 29786 10652 29792
rect 10508 29708 10560 29714
rect 10508 29650 10560 29656
rect 9956 29300 10008 29306
rect 9956 29242 10008 29248
rect 10416 29300 10468 29306
rect 10416 29242 10468 29248
rect 9678 29200 9734 29209
rect 11072 29186 11100 35430
rect 11244 35148 11296 35154
rect 11244 35090 11296 35096
rect 11256 34746 11284 35090
rect 11336 35080 11388 35086
rect 11336 35022 11388 35028
rect 12532 35080 12584 35086
rect 12532 35022 12584 35028
rect 11244 34740 11296 34746
rect 11244 34682 11296 34688
rect 11152 34400 11204 34406
rect 11152 34342 11204 34348
rect 11164 33658 11192 34342
rect 11152 33652 11204 33658
rect 11152 33594 11204 33600
rect 11256 33522 11284 34682
rect 11348 34202 11376 35022
rect 12072 34944 12124 34950
rect 12072 34886 12124 34892
rect 12084 34610 12112 34886
rect 12072 34604 12124 34610
rect 12072 34546 12124 34552
rect 12544 34474 12572 35022
rect 12728 34785 12756 39520
rect 13924 35873 13952 39520
rect 14556 36032 14608 36038
rect 14556 35974 14608 35980
rect 13910 35864 13966 35873
rect 13910 35799 13966 35808
rect 14462 35728 14518 35737
rect 14462 35663 14518 35672
rect 14476 35630 14504 35663
rect 13544 35624 13596 35630
rect 13544 35566 13596 35572
rect 14464 35624 14516 35630
rect 14464 35566 14516 35572
rect 13556 35154 13584 35566
rect 14568 35494 14596 35974
rect 14924 35692 14976 35698
rect 14924 35634 14976 35640
rect 14556 35488 14608 35494
rect 14556 35430 14608 35436
rect 13728 35216 13780 35222
rect 13634 35184 13690 35193
rect 13544 35148 13596 35154
rect 13728 35158 13780 35164
rect 13634 35119 13690 35128
rect 13544 35090 13596 35096
rect 12714 34776 12770 34785
rect 13556 34746 13584 35090
rect 13648 35018 13676 35119
rect 13636 35012 13688 35018
rect 13636 34954 13688 34960
rect 13648 34921 13676 34954
rect 13634 34912 13690 34921
rect 13634 34847 13690 34856
rect 12714 34711 12770 34720
rect 13544 34740 13596 34746
rect 13544 34682 13596 34688
rect 12532 34468 12584 34474
rect 12532 34410 12584 34416
rect 13544 34468 13596 34474
rect 13544 34410 13596 34416
rect 13268 34400 13320 34406
rect 13268 34342 13320 34348
rect 11336 34196 11388 34202
rect 11336 34138 11388 34144
rect 11244 33516 11296 33522
rect 11244 33458 11296 33464
rect 11348 33114 11376 34138
rect 12164 34128 12216 34134
rect 12164 34070 12216 34076
rect 11796 33992 11848 33998
rect 11796 33934 11848 33940
rect 11808 33590 11836 33934
rect 12176 33658 12204 34070
rect 12164 33652 12216 33658
rect 12164 33594 12216 33600
rect 11796 33584 11848 33590
rect 11796 33526 11848 33532
rect 11610 33144 11666 33153
rect 11336 33108 11388 33114
rect 11610 33079 11612 33088
rect 11336 33050 11388 33056
rect 11664 33079 11666 33088
rect 11612 33050 11664 33056
rect 11336 32904 11388 32910
rect 11336 32846 11388 32852
rect 11348 32366 11376 32846
rect 11624 32774 11652 33050
rect 12176 32910 12204 33594
rect 13280 33454 13308 34342
rect 13556 34202 13584 34410
rect 13544 34196 13596 34202
rect 13544 34138 13596 34144
rect 13740 34184 13768 35158
rect 14372 35080 14424 35086
rect 14372 35022 14424 35028
rect 14096 34536 14148 34542
rect 14096 34478 14148 34484
rect 13820 34196 13872 34202
rect 13740 34156 13820 34184
rect 12992 33448 13044 33454
rect 12992 33390 13044 33396
rect 13268 33448 13320 33454
rect 13268 33390 13320 33396
rect 13004 33289 13032 33390
rect 12990 33280 13046 33289
rect 12990 33215 13046 33224
rect 13280 33130 13308 33390
rect 13358 33280 13414 33289
rect 13358 33215 13414 33224
rect 13188 33114 13308 33130
rect 13372 33114 13400 33215
rect 13188 33108 13320 33114
rect 13188 33102 13268 33108
rect 12164 32904 12216 32910
rect 12164 32846 12216 32852
rect 11612 32768 11664 32774
rect 11612 32710 11664 32716
rect 11624 32570 11652 32710
rect 12176 32570 12204 32846
rect 12808 32768 12860 32774
rect 12806 32736 12808 32745
rect 12860 32736 12862 32745
rect 12806 32671 12862 32680
rect 13188 32570 13216 33102
rect 13268 33050 13320 33056
rect 13360 33108 13412 33114
rect 13360 33050 13412 33056
rect 13268 32972 13320 32978
rect 13268 32914 13320 32920
rect 11612 32564 11664 32570
rect 11612 32506 11664 32512
rect 12164 32564 12216 32570
rect 12164 32506 12216 32512
rect 13176 32564 13228 32570
rect 13176 32506 13228 32512
rect 11336 32360 11388 32366
rect 11334 32328 11336 32337
rect 11388 32328 11390 32337
rect 13280 32298 13308 32914
rect 13740 32774 13768 34156
rect 13820 34138 13872 34144
rect 13820 32972 13872 32978
rect 13820 32914 13872 32920
rect 13832 32774 13860 32914
rect 13912 32904 13964 32910
rect 13912 32846 13964 32852
rect 13728 32768 13780 32774
rect 13728 32710 13780 32716
rect 13820 32768 13872 32774
rect 13820 32710 13872 32716
rect 13832 32502 13860 32710
rect 13924 32570 13952 32846
rect 13912 32564 13964 32570
rect 13912 32506 13964 32512
rect 13820 32496 13872 32502
rect 13818 32464 13820 32473
rect 13872 32464 13874 32473
rect 13818 32399 13874 32408
rect 11334 32263 11390 32272
rect 13268 32292 13320 32298
rect 13268 32234 13320 32240
rect 13174 31648 13230 31657
rect 13174 31583 13230 31592
rect 13188 31482 13216 31583
rect 13176 31476 13228 31482
rect 13176 31418 13228 31424
rect 13188 31278 13216 31418
rect 13176 31272 13228 31278
rect 13176 31214 13228 31220
rect 12256 31136 12308 31142
rect 12256 31078 12308 31084
rect 12716 31136 12768 31142
rect 12716 31078 12768 31084
rect 12268 30598 12296 31078
rect 12256 30592 12308 30598
rect 12256 30534 12308 30540
rect 12624 30592 12676 30598
rect 12624 30534 12676 30540
rect 11886 30288 11942 30297
rect 11886 30223 11888 30232
rect 11940 30223 11942 30232
rect 11888 30194 11940 30200
rect 12072 30116 12124 30122
rect 12072 30058 12124 30064
rect 11336 30048 11388 30054
rect 11336 29990 11388 29996
rect 10980 29170 11100 29186
rect 9678 29135 9734 29144
rect 10968 29164 11100 29170
rect 11020 29158 11100 29164
rect 10968 29106 11020 29112
rect 9588 28960 9640 28966
rect 9588 28902 9640 28908
rect 10508 28960 10560 28966
rect 10508 28902 10560 28908
rect 9600 28218 9628 28902
rect 10520 28762 10548 28902
rect 10980 28762 11008 29106
rect 10508 28756 10560 28762
rect 10508 28698 10560 28704
rect 10968 28756 11020 28762
rect 10968 28698 11020 28704
rect 9678 28656 9734 28665
rect 9678 28591 9680 28600
rect 9732 28591 9734 28600
rect 9680 28562 9732 28568
rect 9692 28218 9720 28562
rect 9588 28212 9640 28218
rect 9588 28154 9640 28160
rect 9680 28212 9732 28218
rect 9680 28154 9732 28160
rect 11152 28212 11204 28218
rect 11152 28154 11204 28160
rect 11060 27872 11112 27878
rect 10980 27820 11060 27826
rect 10980 27814 11112 27820
rect 10980 27798 11100 27814
rect 9220 27600 9272 27606
rect 9220 27542 9272 27548
rect 8852 27532 8904 27538
rect 8852 27474 8904 27480
rect 8668 27464 8720 27470
rect 8668 27406 8720 27412
rect 8208 27396 8260 27402
rect 8208 27338 8260 27344
rect 8680 27062 8708 27406
rect 8668 27056 8720 27062
rect 8128 26982 8524 27010
rect 8668 26998 8720 27004
rect 7288 26852 7340 26858
rect 7288 26794 7340 26800
rect 4620 26580 4672 26586
rect 4620 26522 4672 26528
rect 6460 26580 6512 26586
rect 6460 26522 6512 26528
rect 6644 26580 6696 26586
rect 6644 26522 6696 26528
rect 6920 26580 6972 26586
rect 6920 26522 6972 26528
rect 5816 26240 5868 26246
rect 5816 26182 5868 26188
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 5828 26042 5856 26182
rect 2228 26036 2280 26042
rect 2228 25978 2280 25984
rect 5816 26036 5868 26042
rect 5816 25978 5868 25984
rect 6656 25906 6684 26522
rect 6736 26444 6788 26450
rect 6736 26386 6788 26392
rect 6644 25900 6696 25906
rect 6644 25842 6696 25848
rect 2688 25764 2740 25770
rect 2740 25724 2820 25752
rect 2688 25706 2740 25712
rect 1952 25696 2004 25702
rect 1952 25638 2004 25644
rect 1964 25158 1992 25638
rect 1952 25152 2004 25158
rect 1952 25094 2004 25100
rect 1582 20088 1638 20097
rect 1582 20023 1638 20032
rect 1596 19990 1624 20023
rect 1584 19984 1636 19990
rect 1584 19926 1636 19932
rect 1596 19514 1624 19926
rect 1964 19922 1992 25094
rect 2792 20058 2820 25724
rect 6656 25362 6684 25842
rect 6748 25770 6776 26386
rect 8128 26382 8156 26982
rect 8496 26874 8524 26982
rect 8208 26852 8260 26858
rect 8496 26846 8616 26874
rect 8208 26794 8260 26800
rect 8116 26376 8168 26382
rect 8116 26318 8168 26324
rect 6828 26308 6880 26314
rect 6828 26250 6880 26256
rect 6736 25764 6788 25770
rect 6736 25706 6788 25712
rect 6840 25702 6868 26250
rect 8220 26042 8248 26794
rect 8588 26382 8616 26846
rect 8864 26790 8892 27474
rect 9232 27130 9260 27542
rect 10980 27130 11008 27798
rect 11164 27674 11192 28154
rect 11152 27668 11204 27674
rect 11152 27610 11204 27616
rect 11060 27532 11112 27538
rect 11060 27474 11112 27480
rect 9220 27124 9272 27130
rect 9220 27066 9272 27072
rect 10968 27124 11020 27130
rect 10968 27066 11020 27072
rect 9864 27056 9916 27062
rect 9864 26998 9916 27004
rect 9680 26920 9732 26926
rect 9600 26868 9680 26874
rect 9600 26862 9732 26868
rect 9600 26846 9720 26862
rect 8852 26784 8904 26790
rect 8850 26752 8852 26761
rect 8904 26752 8906 26761
rect 8850 26687 8906 26696
rect 9036 26444 9088 26450
rect 9036 26386 9088 26392
rect 8484 26376 8536 26382
rect 8484 26318 8536 26324
rect 8576 26376 8628 26382
rect 8576 26318 8628 26324
rect 8496 26042 8524 26318
rect 8588 26246 8616 26318
rect 8576 26240 8628 26246
rect 8576 26182 8628 26188
rect 8208 26036 8260 26042
rect 8208 25978 8260 25984
rect 8484 26036 8536 26042
rect 8484 25978 8536 25984
rect 7104 25764 7156 25770
rect 7104 25706 7156 25712
rect 6828 25696 6880 25702
rect 6828 25638 6880 25644
rect 6840 25362 6868 25638
rect 7116 25498 7144 25706
rect 7104 25492 7156 25498
rect 7104 25434 7156 25440
rect 6644 25356 6696 25362
rect 6644 25298 6696 25304
rect 6828 25356 6880 25362
rect 6828 25298 6880 25304
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 6656 24954 6684 25298
rect 6840 24954 6868 25298
rect 6644 24948 6696 24954
rect 6644 24890 6696 24896
rect 6828 24948 6880 24954
rect 6828 24890 6880 24896
rect 6840 24410 6868 24890
rect 6920 24744 6972 24750
rect 6920 24686 6972 24692
rect 6828 24404 6880 24410
rect 6828 24346 6880 24352
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 6932 22778 6960 24686
rect 8496 24410 8524 25978
rect 8588 25498 8616 26182
rect 9048 25702 9076 26386
rect 9600 26042 9628 26846
rect 9680 26308 9732 26314
rect 9680 26250 9732 26256
rect 9588 26036 9640 26042
rect 9588 25978 9640 25984
rect 9692 25838 9720 26250
rect 9876 25906 9904 26998
rect 11072 26790 11100 27474
rect 11348 27062 11376 29990
rect 12084 29646 12112 30058
rect 12268 29714 12296 30534
rect 12636 30054 12664 30534
rect 12348 30048 12400 30054
rect 12348 29990 12400 29996
rect 12440 30048 12492 30054
rect 12624 30048 12676 30054
rect 12440 29990 12492 29996
rect 12622 30016 12624 30025
rect 12676 30016 12678 30025
rect 12256 29708 12308 29714
rect 12256 29650 12308 29656
rect 12072 29640 12124 29646
rect 12072 29582 12124 29588
rect 12084 29238 12112 29582
rect 12268 29306 12296 29650
rect 12256 29300 12308 29306
rect 12256 29242 12308 29248
rect 12072 29232 12124 29238
rect 12072 29174 12124 29180
rect 12360 28762 12388 29990
rect 12348 28756 12400 28762
rect 12348 28698 12400 28704
rect 11428 28620 11480 28626
rect 11428 28562 11480 28568
rect 11440 27878 11468 28562
rect 11520 28552 11572 28558
rect 11520 28494 11572 28500
rect 11796 28552 11848 28558
rect 11796 28494 11848 28500
rect 11532 28218 11560 28494
rect 11808 28218 11836 28494
rect 11520 28212 11572 28218
rect 11520 28154 11572 28160
rect 11796 28212 11848 28218
rect 11796 28154 11848 28160
rect 12452 28014 12480 29990
rect 12622 29951 12678 29960
rect 12728 28626 12756 31078
rect 12808 30592 12860 30598
rect 12808 30534 12860 30540
rect 12992 30592 13044 30598
rect 12992 30534 13044 30540
rect 12820 30258 12848 30534
rect 12808 30252 12860 30258
rect 12808 30194 12860 30200
rect 12820 28762 12848 30194
rect 13004 29345 13032 30534
rect 12990 29336 13046 29345
rect 12990 29271 13046 29280
rect 12808 28756 12860 28762
rect 12808 28698 12860 28704
rect 12716 28620 12768 28626
rect 12716 28562 12768 28568
rect 12728 28218 12756 28562
rect 12716 28212 12768 28218
rect 12716 28154 12768 28160
rect 12440 28008 12492 28014
rect 12440 27950 12492 27956
rect 11428 27872 11480 27878
rect 11428 27814 11480 27820
rect 11336 27056 11388 27062
rect 11336 26998 11388 27004
rect 11060 26784 11112 26790
rect 11060 26726 11112 26732
rect 11348 26738 11376 26998
rect 11072 26586 11100 26726
rect 11348 26710 11468 26738
rect 11060 26580 11112 26586
rect 11060 26522 11112 26528
rect 11336 26580 11388 26586
rect 11336 26522 11388 26528
rect 10600 26240 10652 26246
rect 10600 26182 10652 26188
rect 9864 25900 9916 25906
rect 9864 25842 9916 25848
rect 9680 25832 9732 25838
rect 9680 25774 9732 25780
rect 9036 25696 9088 25702
rect 9036 25638 9088 25644
rect 9680 25696 9732 25702
rect 9680 25638 9732 25644
rect 8576 25492 8628 25498
rect 8576 25434 8628 25440
rect 8588 24954 8616 25434
rect 8576 24948 8628 24954
rect 8576 24890 8628 24896
rect 9048 24750 9076 25638
rect 9692 25158 9720 25638
rect 10140 25356 10192 25362
rect 10140 25298 10192 25304
rect 10152 25158 10180 25298
rect 10612 25294 10640 26182
rect 11348 26042 11376 26522
rect 11440 26382 11468 26710
rect 11612 26444 11664 26450
rect 11612 26386 11664 26392
rect 13176 26444 13228 26450
rect 13176 26386 13228 26392
rect 11428 26376 11480 26382
rect 11428 26318 11480 26324
rect 11336 26036 11388 26042
rect 11336 25978 11388 25984
rect 11624 25702 11652 26386
rect 12440 26240 12492 26246
rect 12440 26182 12492 26188
rect 12452 25838 12480 26182
rect 12440 25832 12492 25838
rect 12440 25774 12492 25780
rect 11612 25696 11664 25702
rect 11612 25638 11664 25644
rect 11624 25498 11652 25638
rect 11886 25528 11942 25537
rect 11612 25492 11664 25498
rect 11886 25463 11942 25472
rect 11612 25434 11664 25440
rect 11900 25362 11928 25463
rect 12452 25430 12480 25774
rect 13188 25537 13216 26386
rect 13280 25673 13308 32234
rect 14108 32026 14136 34478
rect 14384 33658 14412 35022
rect 14464 34060 14516 34066
rect 14464 34002 14516 34008
rect 14476 33862 14504 34002
rect 14464 33856 14516 33862
rect 14464 33798 14516 33804
rect 14372 33652 14424 33658
rect 14372 33594 14424 33600
rect 14476 32745 14504 33798
rect 14568 33153 14596 35430
rect 14832 35148 14884 35154
rect 14832 35090 14884 35096
rect 14648 34944 14700 34950
rect 14648 34886 14700 34892
rect 14660 34610 14688 34886
rect 14648 34604 14700 34610
rect 14648 34546 14700 34552
rect 14844 34542 14872 35090
rect 14832 34536 14884 34542
rect 14832 34478 14884 34484
rect 14936 34406 14964 35634
rect 14924 34400 14976 34406
rect 14924 34342 14976 34348
rect 14832 33856 14884 33862
rect 14832 33798 14884 33804
rect 14554 33144 14610 33153
rect 14554 33079 14610 33088
rect 14740 32904 14792 32910
rect 14740 32846 14792 32852
rect 14462 32736 14518 32745
rect 14462 32671 14518 32680
rect 14648 32564 14700 32570
rect 14648 32506 14700 32512
rect 14096 32020 14148 32026
rect 14096 31962 14148 31968
rect 14278 31512 14334 31521
rect 14278 31447 14280 31456
rect 14332 31447 14334 31456
rect 14280 31418 14332 31424
rect 14292 31278 14320 31418
rect 14280 31272 14332 31278
rect 14280 31214 14332 31220
rect 13820 31136 13872 31142
rect 13818 31104 13820 31113
rect 13872 31104 13874 31113
rect 13818 31039 13874 31048
rect 13636 30864 13688 30870
rect 13636 30806 13688 30812
rect 13544 30728 13596 30734
rect 13544 30670 13596 30676
rect 13556 29850 13584 30670
rect 13648 30122 13676 30806
rect 13728 30796 13780 30802
rect 13728 30738 13780 30744
rect 13636 30116 13688 30122
rect 13636 30058 13688 30064
rect 13544 29844 13596 29850
rect 13544 29786 13596 29792
rect 13556 29102 13584 29786
rect 13544 29096 13596 29102
rect 13544 29038 13596 29044
rect 13556 28762 13584 29038
rect 13544 28756 13596 28762
rect 13544 28698 13596 28704
rect 13648 28150 13676 30058
rect 13740 30054 13768 30738
rect 14660 30598 14688 32506
rect 14752 32366 14780 32846
rect 14740 32360 14792 32366
rect 14740 32302 14792 32308
rect 14752 31958 14780 32302
rect 14740 31952 14792 31958
rect 14740 31894 14792 31900
rect 14752 31686 14780 31894
rect 14844 31890 14872 33798
rect 14936 33658 14964 34342
rect 14924 33652 14976 33658
rect 14924 33594 14976 33600
rect 14832 31884 14884 31890
rect 14832 31826 14884 31832
rect 14740 31680 14792 31686
rect 14740 31622 14792 31628
rect 14752 30938 14780 31622
rect 14740 30932 14792 30938
rect 14740 30874 14792 30880
rect 14924 30660 14976 30666
rect 14924 30602 14976 30608
rect 14648 30592 14700 30598
rect 14648 30534 14700 30540
rect 14660 30394 14688 30534
rect 14648 30388 14700 30394
rect 14648 30330 14700 30336
rect 14188 30184 14240 30190
rect 14188 30126 14240 30132
rect 13728 30048 13780 30054
rect 13780 30008 13860 30036
rect 13728 29990 13780 29996
rect 13832 28762 13860 30008
rect 14200 29850 14228 30126
rect 14372 30048 14424 30054
rect 14372 29990 14424 29996
rect 14188 29844 14240 29850
rect 14188 29786 14240 29792
rect 14384 29782 14412 29990
rect 14936 29850 14964 30602
rect 15028 30297 15056 39520
rect 15752 35760 15804 35766
rect 15752 35702 15804 35708
rect 15764 35290 15792 35702
rect 15752 35284 15804 35290
rect 15752 35226 15804 35232
rect 15200 35080 15252 35086
rect 15200 35022 15252 35028
rect 15476 35080 15528 35086
rect 15476 35022 15528 35028
rect 15212 34542 15240 35022
rect 15200 34536 15252 34542
rect 15200 34478 15252 34484
rect 15292 34468 15344 34474
rect 15292 34410 15344 34416
rect 15200 33992 15252 33998
rect 15200 33934 15252 33940
rect 15212 33130 15240 33934
rect 15304 33454 15332 34410
rect 15488 33862 15516 35022
rect 15752 34944 15804 34950
rect 15752 34886 15804 34892
rect 15476 33856 15528 33862
rect 15476 33798 15528 33804
rect 15292 33448 15344 33454
rect 15292 33390 15344 33396
rect 15304 33289 15332 33390
rect 15488 33318 15516 33798
rect 15476 33312 15528 33318
rect 15290 33280 15346 33289
rect 15476 33254 15528 33260
rect 15290 33215 15346 33224
rect 15120 33114 15240 33130
rect 15108 33108 15240 33114
rect 15160 33102 15240 33108
rect 15108 33050 15160 33056
rect 15106 32464 15162 32473
rect 15106 32399 15162 32408
rect 15120 32366 15148 32399
rect 15108 32360 15160 32366
rect 15108 32302 15160 32308
rect 15120 32026 15148 32302
rect 15108 32020 15160 32026
rect 15108 31962 15160 31968
rect 15212 30938 15240 33102
rect 15488 31362 15516 33254
rect 15764 32910 15792 34886
rect 15842 33960 15898 33969
rect 15842 33895 15844 33904
rect 15896 33895 15898 33904
rect 15844 33866 15896 33872
rect 15844 32972 15896 32978
rect 15844 32914 15896 32920
rect 15752 32904 15804 32910
rect 15752 32846 15804 32852
rect 15764 32434 15792 32846
rect 15752 32428 15804 32434
rect 15752 32370 15804 32376
rect 15856 32230 15884 32914
rect 16028 32904 16080 32910
rect 16028 32846 16080 32852
rect 16040 32609 16068 32846
rect 16026 32600 16082 32609
rect 16026 32535 16082 32544
rect 15844 32224 15896 32230
rect 15844 32166 15896 32172
rect 15856 31686 15884 32166
rect 16040 32026 16068 32535
rect 16028 32020 16080 32026
rect 16028 31962 16080 31968
rect 15844 31680 15896 31686
rect 15844 31622 15896 31628
rect 15396 31334 15516 31362
rect 15200 30932 15252 30938
rect 15200 30874 15252 30880
rect 15014 30288 15070 30297
rect 15014 30223 15070 30232
rect 15290 30288 15346 30297
rect 15290 30223 15346 30232
rect 15304 30190 15332 30223
rect 15292 30184 15344 30190
rect 15292 30126 15344 30132
rect 14924 29844 14976 29850
rect 14924 29786 14976 29792
rect 14372 29776 14424 29782
rect 14372 29718 14424 29724
rect 15200 29708 15252 29714
rect 15200 29650 15252 29656
rect 15016 29504 15068 29510
rect 15016 29446 15068 29452
rect 14372 28960 14424 28966
rect 14372 28902 14424 28908
rect 14384 28762 14412 28902
rect 15028 28762 15056 29446
rect 15108 28960 15160 28966
rect 15108 28902 15160 28908
rect 13820 28756 13872 28762
rect 13820 28698 13872 28704
rect 14372 28756 14424 28762
rect 14372 28698 14424 28704
rect 15016 28756 15068 28762
rect 15016 28698 15068 28704
rect 13728 28620 13780 28626
rect 13728 28562 13780 28568
rect 13740 28218 13768 28562
rect 13728 28212 13780 28218
rect 13728 28154 13780 28160
rect 13636 28144 13688 28150
rect 13636 28086 13688 28092
rect 14384 27674 14412 28698
rect 15120 28082 15148 28902
rect 15212 28762 15240 29650
rect 15200 28756 15252 28762
rect 15200 28698 15252 28704
rect 15108 28076 15160 28082
rect 15108 28018 15160 28024
rect 14372 27668 14424 27674
rect 14372 27610 14424 27616
rect 13452 27600 13504 27606
rect 13452 27542 13504 27548
rect 13464 26926 13492 27542
rect 15396 27033 15424 31334
rect 15476 31204 15528 31210
rect 15476 31146 15528 31152
rect 15488 29306 15516 31146
rect 15856 30394 15884 31622
rect 16132 31521 16160 39520
rect 16488 35488 16540 35494
rect 16488 35430 16540 35436
rect 16500 34202 16528 35430
rect 16948 35148 17000 35154
rect 16948 35090 17000 35096
rect 16960 34746 16988 35090
rect 16948 34740 17000 34746
rect 16948 34682 17000 34688
rect 16488 34196 16540 34202
rect 16488 34138 16540 34144
rect 16500 33658 16528 34138
rect 16488 33652 16540 33658
rect 16488 33594 16540 33600
rect 17132 32768 17184 32774
rect 17132 32710 17184 32716
rect 17144 32473 17172 32710
rect 17130 32464 17186 32473
rect 17130 32399 17186 32408
rect 17040 32360 17092 32366
rect 17040 32302 17092 32308
rect 16672 32292 16724 32298
rect 16672 32234 16724 32240
rect 16212 31680 16264 31686
rect 16212 31622 16264 31628
rect 16118 31512 16174 31521
rect 16118 31447 16174 31456
rect 16224 31210 16252 31622
rect 16212 31204 16264 31210
rect 16212 31146 16264 31152
rect 15936 30796 15988 30802
rect 15936 30738 15988 30744
rect 15948 30433 15976 30738
rect 16028 30728 16080 30734
rect 16028 30670 16080 30676
rect 15934 30424 15990 30433
rect 15660 30388 15712 30394
rect 15660 30330 15712 30336
rect 15844 30388 15896 30394
rect 15934 30359 15990 30368
rect 15844 30330 15896 30336
rect 15672 30054 15700 30330
rect 15752 30252 15804 30258
rect 15752 30194 15804 30200
rect 15660 30048 15712 30054
rect 15660 29990 15712 29996
rect 15764 29714 15792 30194
rect 15752 29708 15804 29714
rect 15752 29650 15804 29656
rect 15476 29300 15528 29306
rect 15476 29242 15528 29248
rect 15948 29238 15976 30359
rect 16040 30054 16068 30670
rect 16120 30592 16172 30598
rect 16120 30534 16172 30540
rect 16132 30258 16160 30534
rect 16120 30252 16172 30258
rect 16120 30194 16172 30200
rect 16028 30048 16080 30054
rect 16028 29990 16080 29996
rect 16040 29850 16068 29990
rect 16028 29844 16080 29850
rect 16028 29786 16080 29792
rect 16028 29504 16080 29510
rect 16224 29458 16252 31146
rect 16684 31142 16712 32234
rect 16948 32224 17000 32230
rect 16948 32166 17000 32172
rect 16960 31958 16988 32166
rect 16948 31952 17000 31958
rect 16948 31894 17000 31900
rect 16672 31136 16724 31142
rect 16672 31078 16724 31084
rect 16684 30734 16712 31078
rect 16960 30734 16988 31894
rect 17052 31890 17080 32302
rect 17236 31906 17264 39520
rect 18050 36136 18106 36145
rect 18050 36071 18106 36080
rect 17868 35080 17920 35086
rect 17868 35022 17920 35028
rect 17408 34944 17460 34950
rect 17408 34886 17460 34892
rect 17040 31884 17092 31890
rect 17040 31826 17092 31832
rect 17144 31878 17264 31906
rect 17144 31770 17172 31878
rect 17052 31742 17172 31770
rect 17052 31657 17080 31742
rect 17038 31648 17094 31657
rect 17038 31583 17094 31592
rect 16672 30728 16724 30734
rect 16672 30670 16724 30676
rect 16948 30728 17000 30734
rect 16948 30670 17000 30676
rect 16960 30297 16988 30670
rect 16946 30288 17002 30297
rect 16946 30223 17002 30232
rect 17132 30048 17184 30054
rect 17132 29990 17184 29996
rect 17144 29850 17172 29990
rect 17132 29844 17184 29850
rect 17132 29786 17184 29792
rect 17040 29708 17092 29714
rect 17040 29650 17092 29656
rect 16080 29452 16252 29458
rect 16028 29446 16252 29452
rect 16580 29504 16632 29510
rect 16580 29446 16632 29452
rect 16040 29430 16252 29446
rect 15936 29232 15988 29238
rect 15750 29200 15806 29209
rect 15936 29174 15988 29180
rect 15750 29135 15806 29144
rect 15764 28694 15792 29135
rect 16224 29102 16252 29430
rect 16394 29336 16450 29345
rect 16394 29271 16450 29280
rect 16408 29170 16436 29271
rect 16396 29164 16448 29170
rect 16396 29106 16448 29112
rect 16212 29096 16264 29102
rect 15842 29064 15898 29073
rect 16212 29038 16264 29044
rect 15842 28999 15898 29008
rect 15856 28762 15884 28999
rect 16408 28762 16436 29106
rect 15844 28756 15896 28762
rect 15844 28698 15896 28704
rect 16396 28756 16448 28762
rect 16396 28698 16448 28704
rect 15752 28688 15804 28694
rect 15752 28630 15804 28636
rect 15764 28218 15792 28630
rect 15752 28212 15804 28218
rect 15752 28154 15804 28160
rect 15856 28082 15884 28698
rect 16592 28642 16620 29446
rect 17052 29238 17080 29650
rect 17040 29232 17092 29238
rect 17040 29174 17092 29180
rect 17132 29096 17184 29102
rect 17132 29038 17184 29044
rect 16500 28614 16620 28642
rect 16500 28558 16528 28614
rect 16028 28552 16080 28558
rect 16028 28494 16080 28500
rect 16488 28552 16540 28558
rect 16488 28494 16540 28500
rect 16040 28218 16068 28494
rect 16028 28212 16080 28218
rect 16028 28154 16080 28160
rect 15844 28076 15896 28082
rect 15844 28018 15896 28024
rect 16040 27606 16068 28154
rect 16028 27600 16080 27606
rect 16028 27542 16080 27548
rect 15568 27464 15620 27470
rect 15568 27406 15620 27412
rect 13726 27024 13782 27033
rect 13726 26959 13782 26968
rect 15382 27024 15438 27033
rect 15580 26994 15608 27406
rect 16040 27130 16068 27542
rect 16948 27328 17000 27334
rect 16948 27270 17000 27276
rect 16028 27124 16080 27130
rect 16028 27066 16080 27072
rect 15382 26959 15438 26968
rect 15568 26988 15620 26994
rect 13740 26926 13768 26959
rect 15568 26930 15620 26936
rect 13452 26920 13504 26926
rect 13452 26862 13504 26868
rect 13728 26920 13780 26926
rect 13728 26862 13780 26868
rect 14832 26784 14884 26790
rect 14832 26726 14884 26732
rect 14844 26586 14872 26726
rect 13544 26580 13596 26586
rect 13544 26522 13596 26528
rect 14832 26580 14884 26586
rect 14832 26522 14884 26528
rect 13556 25838 13584 26522
rect 15580 26450 15608 26930
rect 16960 26518 16988 27270
rect 17144 26994 17172 29038
rect 17132 26988 17184 26994
rect 17132 26930 17184 26936
rect 16120 26512 16172 26518
rect 16120 26454 16172 26460
rect 16948 26512 17000 26518
rect 16948 26454 17000 26460
rect 15568 26444 15620 26450
rect 15568 26386 15620 26392
rect 16132 25906 16160 26454
rect 16488 26240 16540 26246
rect 16488 26182 16540 26188
rect 16120 25900 16172 25906
rect 16120 25842 16172 25848
rect 16304 25900 16356 25906
rect 16304 25842 16356 25848
rect 13544 25832 13596 25838
rect 13544 25774 13596 25780
rect 15108 25832 15160 25838
rect 15108 25774 15160 25780
rect 16028 25832 16080 25838
rect 16028 25774 16080 25780
rect 13266 25664 13322 25673
rect 13266 25599 13322 25608
rect 13174 25528 13230 25537
rect 13174 25463 13230 25472
rect 12440 25424 12492 25430
rect 12440 25366 12492 25372
rect 11888 25356 11940 25362
rect 11888 25298 11940 25304
rect 10508 25288 10560 25294
rect 10508 25230 10560 25236
rect 10600 25288 10652 25294
rect 10652 25236 10732 25242
rect 10600 25230 10732 25236
rect 9680 25152 9732 25158
rect 9680 25094 9732 25100
rect 10140 25152 10192 25158
rect 10140 25094 10192 25100
rect 9036 24744 9088 24750
rect 9036 24686 9088 24692
rect 8484 24404 8536 24410
rect 8484 24346 8536 24352
rect 7196 24268 7248 24274
rect 7196 24210 7248 24216
rect 7748 24268 7800 24274
rect 7748 24210 7800 24216
rect 7208 23866 7236 24210
rect 7196 23860 7248 23866
rect 7196 23802 7248 23808
rect 7208 23769 7236 23802
rect 7194 23760 7250 23769
rect 7194 23695 7250 23704
rect 7760 23594 7788 24210
rect 8496 23662 8524 24346
rect 9048 23866 9076 24686
rect 9692 23866 9720 25094
rect 10152 24750 10180 25094
rect 10520 24954 10548 25230
rect 10612 25214 10732 25230
rect 10508 24948 10560 24954
rect 10508 24890 10560 24896
rect 10520 24750 10548 24890
rect 9864 24744 9916 24750
rect 10140 24744 10192 24750
rect 9864 24686 9916 24692
rect 10138 24712 10140 24721
rect 10508 24744 10560 24750
rect 10192 24712 10194 24721
rect 9876 24274 9904 24686
rect 10508 24686 10560 24692
rect 10138 24647 10194 24656
rect 10600 24336 10652 24342
rect 10600 24278 10652 24284
rect 9864 24268 9916 24274
rect 9864 24210 9916 24216
rect 10416 24268 10468 24274
rect 10416 24210 10468 24216
rect 9036 23860 9088 23866
rect 9036 23802 9088 23808
rect 9680 23860 9732 23866
rect 9680 23802 9732 23808
rect 10232 23724 10284 23730
rect 10232 23666 10284 23672
rect 8484 23656 8536 23662
rect 8484 23598 8536 23604
rect 7748 23588 7800 23594
rect 7748 23530 7800 23536
rect 7760 23322 7788 23530
rect 10244 23322 10272 23666
rect 10428 23526 10456 24210
rect 10506 23760 10562 23769
rect 10612 23730 10640 24278
rect 10704 23730 10732 25214
rect 11900 24954 11928 25298
rect 11888 24948 11940 24954
rect 11888 24890 11940 24896
rect 12452 24614 12480 25366
rect 12992 25152 13044 25158
rect 12992 25094 13044 25100
rect 12716 24948 12768 24954
rect 12716 24890 12768 24896
rect 12728 24750 12756 24890
rect 13004 24750 13032 25094
rect 12716 24744 12768 24750
rect 12716 24686 12768 24692
rect 12992 24744 13044 24750
rect 12992 24686 13044 24692
rect 11244 24608 11296 24614
rect 11244 24550 11296 24556
rect 12440 24608 12492 24614
rect 12440 24550 12492 24556
rect 11256 24342 11284 24550
rect 12452 24342 12480 24550
rect 11244 24336 11296 24342
rect 11244 24278 11296 24284
rect 12440 24336 12492 24342
rect 12440 24278 12492 24284
rect 12992 24132 13044 24138
rect 12992 24074 13044 24080
rect 11152 24064 11204 24070
rect 11152 24006 11204 24012
rect 10506 23695 10562 23704
rect 10600 23724 10652 23730
rect 10520 23662 10548 23695
rect 10600 23666 10652 23672
rect 10692 23724 10744 23730
rect 10692 23666 10744 23672
rect 10508 23656 10560 23662
rect 10508 23598 10560 23604
rect 10416 23520 10468 23526
rect 10416 23462 10468 23468
rect 10428 23322 10456 23462
rect 10704 23322 10732 23666
rect 11164 23662 11192 24006
rect 13004 23662 13032 24074
rect 11152 23656 11204 23662
rect 11152 23598 11204 23604
rect 12992 23656 13044 23662
rect 12992 23598 13044 23604
rect 12348 23520 12400 23526
rect 12400 23480 12480 23508
rect 12348 23462 12400 23468
rect 7748 23316 7800 23322
rect 7748 23258 7800 23264
rect 10232 23316 10284 23322
rect 10232 23258 10284 23264
rect 10416 23316 10468 23322
rect 10416 23258 10468 23264
rect 10692 23316 10744 23322
rect 10692 23258 10744 23264
rect 10600 23180 10652 23186
rect 10600 23122 10652 23128
rect 10612 22778 10640 23122
rect 6920 22772 6972 22778
rect 6920 22714 6972 22720
rect 8576 22772 8628 22778
rect 8576 22714 8628 22720
rect 10600 22772 10652 22778
rect 10600 22714 10652 22720
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 8588 21690 8616 22714
rect 12256 22092 12308 22098
rect 12256 22034 12308 22040
rect 8576 21684 8628 21690
rect 8576 21626 8628 21632
rect 12268 21350 12296 22034
rect 12452 22030 12480 23480
rect 12440 22024 12492 22030
rect 12440 21966 12492 21972
rect 12452 21486 12480 21966
rect 13004 21962 13032 23598
rect 13176 22772 13228 22778
rect 13176 22714 13228 22720
rect 12992 21956 13044 21962
rect 12992 21898 13044 21904
rect 13188 21690 13216 22714
rect 13176 21684 13228 21690
rect 13176 21626 13228 21632
rect 12440 21480 12492 21486
rect 12440 21422 12492 21428
rect 9128 21344 9180 21350
rect 9128 21286 9180 21292
rect 12256 21344 12308 21350
rect 12256 21286 12308 21292
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 9140 20534 9168 21286
rect 10046 20632 10102 20641
rect 10046 20567 10048 20576
rect 10100 20567 10102 20576
rect 10048 20538 10100 20544
rect 9128 20528 9180 20534
rect 9128 20470 9180 20476
rect 10060 20398 10088 20538
rect 10048 20392 10100 20398
rect 10048 20334 10100 20340
rect 12268 20262 12296 21286
rect 12452 21010 12480 21422
rect 12992 21412 13044 21418
rect 12992 21354 13044 21360
rect 13004 21078 13032 21354
rect 12992 21072 13044 21078
rect 12992 21014 13044 21020
rect 12440 21004 12492 21010
rect 12440 20946 12492 20952
rect 12256 20256 12308 20262
rect 12256 20198 12308 20204
rect 12452 20058 12480 20946
rect 13004 20602 13032 21014
rect 13280 20641 13308 25599
rect 13556 25498 13584 25774
rect 13820 25696 13872 25702
rect 13820 25638 13872 25644
rect 14554 25664 14610 25673
rect 13832 25537 13860 25638
rect 14554 25599 14610 25608
rect 13818 25528 13874 25537
rect 13544 25492 13596 25498
rect 14568 25498 14596 25599
rect 13818 25463 13874 25472
rect 14556 25492 14608 25498
rect 13544 25434 13596 25440
rect 14556 25434 14608 25440
rect 14464 25356 14516 25362
rect 14464 25298 14516 25304
rect 13818 24712 13874 24721
rect 13818 24647 13874 24656
rect 13832 24614 13860 24647
rect 14476 24614 14504 25298
rect 15120 24954 15148 25774
rect 15660 25696 15712 25702
rect 15660 25638 15712 25644
rect 15672 25537 15700 25638
rect 15658 25528 15714 25537
rect 15658 25463 15714 25472
rect 16040 25430 16068 25774
rect 16028 25424 16080 25430
rect 16028 25366 16080 25372
rect 15384 25288 15436 25294
rect 15384 25230 15436 25236
rect 15108 24948 15160 24954
rect 15108 24890 15160 24896
rect 15396 24750 15424 25230
rect 15384 24744 15436 24750
rect 15384 24686 15436 24692
rect 13820 24608 13872 24614
rect 13820 24550 13872 24556
rect 14464 24608 14516 24614
rect 14464 24550 14516 24556
rect 14476 24313 14504 24550
rect 15396 24342 15424 24686
rect 15936 24676 15988 24682
rect 15936 24618 15988 24624
rect 15474 24576 15530 24585
rect 15474 24511 15530 24520
rect 15488 24410 15516 24511
rect 15948 24410 15976 24618
rect 15476 24404 15528 24410
rect 15476 24346 15528 24352
rect 15936 24404 15988 24410
rect 15936 24346 15988 24352
rect 14556 24336 14608 24342
rect 14462 24304 14518 24313
rect 14556 24278 14608 24284
rect 15384 24336 15436 24342
rect 15384 24278 15436 24284
rect 14462 24239 14518 24248
rect 14568 23662 14596 24278
rect 14556 23656 14608 23662
rect 14556 23598 14608 23604
rect 15200 23520 15252 23526
rect 15200 23462 15252 23468
rect 15212 23338 15240 23462
rect 15120 23322 15240 23338
rect 14096 23316 14148 23322
rect 14096 23258 14148 23264
rect 15108 23316 15240 23322
rect 15160 23310 15240 23316
rect 15108 23258 15160 23264
rect 14004 23180 14056 23186
rect 14004 23122 14056 23128
rect 13544 23112 13596 23118
rect 13544 23054 13596 23060
rect 13556 22234 13584 23054
rect 13636 22976 13688 22982
rect 13636 22918 13688 22924
rect 13544 22228 13596 22234
rect 13544 22170 13596 22176
rect 13556 22030 13584 22170
rect 13544 22024 13596 22030
rect 13648 22001 13676 22918
rect 14016 22778 14044 23122
rect 14004 22772 14056 22778
rect 14004 22714 14056 22720
rect 13912 22568 13964 22574
rect 13912 22510 13964 22516
rect 13924 22250 13952 22510
rect 14108 22506 14136 23258
rect 15948 23254 15976 24346
rect 16316 24206 16344 25842
rect 16500 25838 16528 26182
rect 17144 25974 17172 26930
rect 17132 25968 17184 25974
rect 17132 25910 17184 25916
rect 16488 25832 16540 25838
rect 16488 25774 16540 25780
rect 16580 25152 16632 25158
rect 16580 25094 16632 25100
rect 16592 24426 16620 25094
rect 16672 24608 16724 24614
rect 16672 24550 16724 24556
rect 16500 24410 16620 24426
rect 16488 24404 16620 24410
rect 16540 24398 16620 24404
rect 16488 24346 16540 24352
rect 16684 24274 16712 24550
rect 16672 24268 16724 24274
rect 16672 24210 16724 24216
rect 17132 24268 17184 24274
rect 17132 24210 17184 24216
rect 16304 24200 16356 24206
rect 16304 24142 16356 24148
rect 16316 23254 16344 24142
rect 16684 23866 16712 24210
rect 17144 23866 17172 24210
rect 17224 24064 17276 24070
rect 17224 24006 17276 24012
rect 16672 23860 16724 23866
rect 16672 23802 16724 23808
rect 17132 23860 17184 23866
rect 17132 23802 17184 23808
rect 16580 23520 16632 23526
rect 16580 23462 16632 23468
rect 16396 23316 16448 23322
rect 16396 23258 16448 23264
rect 15936 23248 15988 23254
rect 15936 23190 15988 23196
rect 16304 23248 16356 23254
rect 16304 23190 16356 23196
rect 15292 23180 15344 23186
rect 15292 23122 15344 23128
rect 14648 22568 14700 22574
rect 14648 22510 14700 22516
rect 14096 22500 14148 22506
rect 14096 22442 14148 22448
rect 13924 22222 14044 22250
rect 14660 22234 14688 22510
rect 15304 22234 15332 23122
rect 16408 22234 16436 23258
rect 16592 22794 16620 23462
rect 17236 23322 17264 24006
rect 17224 23316 17276 23322
rect 17224 23258 17276 23264
rect 17040 23112 17092 23118
rect 17040 23054 17092 23060
rect 16500 22766 16620 22794
rect 16500 22710 16528 22766
rect 16488 22704 16540 22710
rect 16488 22646 16540 22652
rect 17052 22642 17080 23054
rect 17236 22778 17264 23258
rect 17420 23118 17448 34886
rect 17880 34762 17908 35022
rect 17880 34746 18000 34762
rect 18064 34746 18092 36071
rect 18142 35456 18198 35465
rect 18142 35391 18198 35400
rect 18156 34921 18184 35391
rect 18340 35154 18368 39520
rect 18328 35148 18380 35154
rect 18328 35090 18380 35096
rect 18512 34944 18564 34950
rect 18142 34912 18198 34921
rect 18512 34886 18564 34892
rect 19154 34912 19210 34921
rect 18142 34847 18198 34856
rect 17868 34740 18000 34746
rect 17920 34734 18000 34740
rect 17868 34682 17920 34688
rect 17868 34604 17920 34610
rect 17868 34546 17920 34552
rect 17776 34128 17828 34134
rect 17776 34070 17828 34076
rect 17788 33318 17816 34070
rect 17776 33312 17828 33318
rect 17774 33280 17776 33289
rect 17828 33280 17830 33289
rect 17774 33215 17830 33224
rect 17776 32972 17828 32978
rect 17776 32914 17828 32920
rect 17500 32768 17552 32774
rect 17500 32710 17552 32716
rect 17512 32570 17540 32710
rect 17500 32564 17552 32570
rect 17500 32506 17552 32512
rect 17512 32026 17540 32506
rect 17788 32298 17816 32914
rect 17776 32292 17828 32298
rect 17776 32234 17828 32240
rect 17880 32026 17908 34546
rect 17972 34542 18000 34734
rect 18052 34740 18104 34746
rect 18052 34682 18104 34688
rect 18064 34649 18092 34682
rect 18050 34640 18106 34649
rect 18524 34610 18552 34886
rect 19154 34847 19210 34856
rect 18050 34575 18106 34584
rect 18512 34604 18564 34610
rect 18512 34546 18564 34552
rect 17960 34536 18012 34542
rect 17960 34478 18012 34484
rect 18052 34060 18104 34066
rect 18052 34002 18104 34008
rect 18064 33454 18092 34002
rect 18788 33856 18840 33862
rect 18788 33798 18840 33804
rect 18800 33454 18828 33798
rect 18052 33448 18104 33454
rect 18052 33390 18104 33396
rect 18788 33448 18840 33454
rect 18788 33390 18840 33396
rect 17960 33380 18012 33386
rect 17960 33322 18012 33328
rect 17972 33114 18000 33322
rect 17960 33108 18012 33114
rect 17960 33050 18012 33056
rect 17500 32020 17552 32026
rect 17500 31962 17552 31968
rect 17868 32020 17920 32026
rect 17868 31962 17920 31968
rect 17972 31754 18000 33050
rect 18064 32722 18092 33390
rect 18144 32768 18196 32774
rect 18064 32716 18144 32722
rect 18064 32710 18196 32716
rect 18064 32694 18184 32710
rect 18064 32570 18092 32694
rect 18052 32564 18104 32570
rect 18052 32506 18104 32512
rect 19064 32564 19116 32570
rect 19064 32506 19116 32512
rect 18604 32360 18656 32366
rect 18604 32302 18656 32308
rect 18616 32026 18644 32302
rect 19076 32026 19104 32506
rect 18604 32020 18656 32026
rect 18604 31962 18656 31968
rect 19064 32020 19116 32026
rect 19064 31962 19116 31968
rect 18052 31952 18104 31958
rect 18052 31894 18104 31900
rect 17684 31748 17736 31754
rect 17684 31690 17736 31696
rect 17960 31748 18012 31754
rect 17960 31690 18012 31696
rect 17696 31414 17724 31690
rect 17972 31482 18000 31690
rect 17960 31476 18012 31482
rect 17960 31418 18012 31424
rect 17684 31408 17736 31414
rect 17684 31350 17736 31356
rect 17592 31136 17644 31142
rect 17592 31078 17644 31084
rect 17604 30734 17632 31078
rect 17696 30938 17724 31350
rect 18064 31142 18092 31894
rect 18052 31136 18104 31142
rect 18052 31078 18104 31084
rect 17684 30932 17736 30938
rect 17684 30874 17736 30880
rect 18972 30932 19024 30938
rect 18972 30874 19024 30880
rect 17500 30728 17552 30734
rect 17500 30670 17552 30676
rect 17592 30728 17644 30734
rect 17592 30670 17644 30676
rect 17512 30394 17540 30670
rect 17500 30388 17552 30394
rect 17500 30330 17552 30336
rect 17512 30122 17540 30330
rect 17500 30116 17552 30122
rect 17500 30058 17552 30064
rect 17604 29782 17632 30670
rect 17776 30592 17828 30598
rect 17776 30534 17828 30540
rect 17592 29776 17644 29782
rect 17592 29718 17644 29724
rect 17788 29034 17816 30534
rect 18510 30424 18566 30433
rect 18510 30359 18566 30368
rect 18524 30258 18552 30359
rect 18512 30252 18564 30258
rect 18512 30194 18564 30200
rect 18696 30252 18748 30258
rect 18696 30194 18748 30200
rect 17960 30116 18012 30122
rect 17960 30058 18012 30064
rect 17776 29028 17828 29034
rect 17776 28970 17828 28976
rect 17972 27878 18000 30058
rect 18052 30048 18104 30054
rect 18052 29990 18104 29996
rect 18064 29073 18092 29990
rect 18708 29850 18736 30194
rect 18696 29844 18748 29850
rect 18696 29786 18748 29792
rect 18144 29640 18196 29646
rect 18144 29582 18196 29588
rect 18156 29209 18184 29582
rect 18236 29300 18288 29306
rect 18236 29242 18288 29248
rect 18142 29200 18198 29209
rect 18142 29135 18198 29144
rect 18050 29064 18106 29073
rect 18050 28999 18106 29008
rect 18248 28762 18276 29242
rect 18708 29238 18736 29786
rect 18880 29572 18932 29578
rect 18880 29514 18932 29520
rect 18892 29238 18920 29514
rect 18696 29232 18748 29238
rect 18696 29174 18748 29180
rect 18880 29232 18932 29238
rect 18880 29174 18932 29180
rect 18880 28960 18932 28966
rect 18880 28902 18932 28908
rect 18236 28756 18288 28762
rect 18236 28698 18288 28704
rect 18892 28014 18920 28902
rect 18984 28762 19012 30874
rect 19064 29504 19116 29510
rect 19064 29446 19116 29452
rect 18972 28756 19024 28762
rect 18972 28698 19024 28704
rect 18970 28520 19026 28529
rect 18970 28455 19026 28464
rect 18880 28008 18932 28014
rect 18880 27950 18932 27956
rect 17960 27872 18012 27878
rect 17960 27814 18012 27820
rect 18892 27402 18920 27950
rect 18984 27606 19012 28455
rect 19076 28014 19104 29446
rect 19064 28008 19116 28014
rect 19064 27950 19116 27956
rect 18972 27600 19024 27606
rect 18972 27542 19024 27548
rect 18880 27396 18932 27402
rect 18880 27338 18932 27344
rect 18694 27160 18750 27169
rect 18694 27095 18696 27104
rect 18748 27095 18750 27104
rect 18696 27066 18748 27072
rect 18708 26926 18736 27066
rect 18696 26920 18748 26926
rect 18696 26862 18748 26868
rect 17960 26784 18012 26790
rect 17960 26726 18012 26732
rect 17972 26330 18000 26726
rect 19168 26586 19196 34847
rect 19248 34604 19300 34610
rect 19248 34546 19300 34552
rect 19260 33640 19288 34546
rect 19340 33652 19392 33658
rect 19260 33612 19340 33640
rect 19260 32366 19288 33612
rect 19340 33594 19392 33600
rect 19338 33280 19394 33289
rect 19338 33215 19394 33224
rect 19352 33114 19380 33215
rect 19340 33108 19392 33114
rect 19340 33050 19392 33056
rect 19248 32360 19300 32366
rect 19248 32302 19300 32308
rect 19340 32224 19392 32230
rect 19340 32166 19392 32172
rect 19352 30274 19380 32166
rect 19260 30258 19380 30274
rect 19248 30252 19380 30258
rect 19300 30246 19380 30252
rect 19248 30194 19300 30200
rect 19248 29640 19300 29646
rect 19248 29582 19300 29588
rect 19260 29034 19288 29582
rect 19248 29028 19300 29034
rect 19248 28970 19300 28976
rect 19260 28762 19288 28970
rect 19248 28756 19300 28762
rect 19248 28698 19300 28704
rect 19340 28008 19392 28014
rect 19340 27950 19392 27956
rect 19352 27674 19380 27950
rect 19340 27668 19392 27674
rect 19340 27610 19392 27616
rect 19444 26874 19472 39520
rect 19580 37564 19876 37584
rect 19636 37562 19660 37564
rect 19716 37562 19740 37564
rect 19796 37562 19820 37564
rect 19658 37510 19660 37562
rect 19722 37510 19734 37562
rect 19796 37510 19798 37562
rect 19636 37508 19660 37510
rect 19716 37508 19740 37510
rect 19796 37508 19820 37510
rect 19580 37488 19876 37508
rect 19580 36476 19876 36496
rect 19636 36474 19660 36476
rect 19716 36474 19740 36476
rect 19796 36474 19820 36476
rect 19658 36422 19660 36474
rect 19722 36422 19734 36474
rect 19796 36422 19798 36474
rect 19636 36420 19660 36422
rect 19716 36420 19740 36422
rect 19796 36420 19820 36422
rect 19580 36400 19876 36420
rect 19580 35388 19876 35408
rect 19636 35386 19660 35388
rect 19716 35386 19740 35388
rect 19796 35386 19820 35388
rect 19658 35334 19660 35386
rect 19722 35334 19734 35386
rect 19796 35334 19798 35386
rect 19636 35332 19660 35334
rect 19716 35332 19740 35334
rect 19796 35332 19820 35334
rect 19580 35312 19876 35332
rect 20168 34400 20220 34406
rect 20168 34342 20220 34348
rect 19580 34300 19876 34320
rect 19636 34298 19660 34300
rect 19716 34298 19740 34300
rect 19796 34298 19820 34300
rect 19658 34246 19660 34298
rect 19722 34246 19734 34298
rect 19796 34246 19798 34298
rect 19636 34244 19660 34246
rect 19716 34244 19740 34246
rect 19796 34244 19820 34246
rect 19580 34224 19876 34244
rect 19580 33212 19876 33232
rect 19636 33210 19660 33212
rect 19716 33210 19740 33212
rect 19796 33210 19820 33212
rect 19658 33158 19660 33210
rect 19722 33158 19734 33210
rect 19796 33158 19798 33210
rect 19636 33156 19660 33158
rect 19716 33156 19740 33158
rect 19796 33156 19820 33158
rect 19580 33136 19876 33156
rect 20180 33017 20208 34342
rect 20166 33008 20222 33017
rect 20166 32943 20222 32952
rect 19580 32124 19876 32144
rect 19636 32122 19660 32124
rect 19716 32122 19740 32124
rect 19796 32122 19820 32124
rect 19658 32070 19660 32122
rect 19722 32070 19734 32122
rect 19796 32070 19798 32122
rect 19636 32068 19660 32070
rect 19716 32068 19740 32070
rect 19796 32068 19820 32070
rect 19580 32048 19876 32068
rect 19580 31036 19876 31056
rect 19636 31034 19660 31036
rect 19716 31034 19740 31036
rect 19796 31034 19820 31036
rect 19658 30982 19660 31034
rect 19722 30982 19734 31034
rect 19796 30982 19798 31034
rect 19636 30980 19660 30982
rect 19716 30980 19740 30982
rect 19796 30980 19820 30982
rect 19580 30960 19876 30980
rect 20168 30796 20220 30802
rect 20168 30738 20220 30744
rect 20180 30258 20208 30738
rect 20168 30252 20220 30258
rect 20168 30194 20220 30200
rect 19984 30048 20036 30054
rect 19984 29990 20036 29996
rect 19580 29948 19876 29968
rect 19636 29946 19660 29948
rect 19716 29946 19740 29948
rect 19796 29946 19820 29948
rect 19658 29894 19660 29946
rect 19722 29894 19734 29946
rect 19796 29894 19798 29946
rect 19636 29892 19660 29894
rect 19716 29892 19740 29894
rect 19796 29892 19820 29894
rect 19580 29872 19876 29892
rect 19524 29708 19576 29714
rect 19524 29650 19576 29656
rect 19536 29306 19564 29650
rect 19996 29646 20024 29990
rect 19984 29640 20036 29646
rect 19984 29582 20036 29588
rect 19892 29504 19944 29510
rect 19892 29446 19944 29452
rect 19524 29300 19576 29306
rect 19524 29242 19576 29248
rect 19904 29034 19932 29446
rect 19996 29306 20024 29582
rect 19984 29300 20036 29306
rect 19984 29242 20036 29248
rect 20180 29102 20208 30194
rect 20168 29096 20220 29102
rect 20168 29038 20220 29044
rect 19892 29028 19944 29034
rect 19892 28970 19944 28976
rect 19580 28860 19876 28880
rect 19636 28858 19660 28860
rect 19716 28858 19740 28860
rect 19796 28858 19820 28860
rect 19658 28806 19660 28858
rect 19722 28806 19734 28858
rect 19796 28806 19798 28858
rect 19636 28804 19660 28806
rect 19716 28804 19740 28806
rect 19796 28804 19820 28806
rect 19580 28784 19876 28804
rect 19708 28688 19760 28694
rect 19708 28630 19760 28636
rect 19720 28082 19748 28630
rect 19904 28558 19932 28970
rect 20180 28762 20208 29038
rect 20168 28756 20220 28762
rect 20168 28698 20220 28704
rect 19892 28552 19944 28558
rect 19890 28520 19892 28529
rect 19944 28520 19946 28529
rect 19890 28455 19946 28464
rect 19984 28484 20036 28490
rect 19984 28426 20036 28432
rect 19708 28076 19760 28082
rect 19708 28018 19760 28024
rect 19580 27772 19876 27792
rect 19636 27770 19660 27772
rect 19716 27770 19740 27772
rect 19796 27770 19820 27772
rect 19658 27718 19660 27770
rect 19722 27718 19734 27770
rect 19796 27718 19798 27770
rect 19636 27716 19660 27718
rect 19716 27716 19740 27718
rect 19796 27716 19820 27718
rect 19580 27696 19876 27716
rect 19996 27334 20024 28426
rect 20352 27396 20404 27402
rect 20352 27338 20404 27344
rect 19984 27328 20036 27334
rect 19984 27270 20036 27276
rect 19260 26846 19472 26874
rect 19156 26580 19208 26586
rect 19156 26522 19208 26528
rect 19260 26450 19288 26846
rect 19340 26784 19392 26790
rect 19340 26726 19392 26732
rect 19352 26586 19380 26726
rect 19580 26684 19876 26704
rect 19636 26682 19660 26684
rect 19716 26682 19740 26684
rect 19796 26682 19820 26684
rect 19658 26630 19660 26682
rect 19722 26630 19734 26682
rect 19796 26630 19798 26682
rect 19636 26628 19660 26630
rect 19716 26628 19740 26630
rect 19796 26628 19820 26630
rect 19580 26608 19876 26628
rect 19340 26580 19392 26586
rect 19340 26522 19392 26528
rect 18328 26444 18380 26450
rect 18328 26386 18380 26392
rect 19248 26444 19300 26450
rect 19248 26386 19300 26392
rect 17880 26302 18000 26330
rect 17880 26042 17908 26302
rect 17960 26240 18012 26246
rect 17960 26182 18012 26188
rect 17868 26036 17920 26042
rect 17868 25978 17920 25984
rect 17972 25294 18000 26182
rect 18340 26042 18368 26386
rect 19352 26330 19380 26522
rect 19432 26512 19484 26518
rect 19432 26454 19484 26460
rect 19168 26302 19380 26330
rect 19168 26042 19196 26302
rect 18328 26036 18380 26042
rect 18328 25978 18380 25984
rect 19156 26036 19208 26042
rect 19156 25978 19208 25984
rect 19444 25922 19472 26454
rect 19800 26240 19852 26246
rect 19800 26182 19852 26188
rect 19260 25906 19472 25922
rect 19812 25906 19840 26182
rect 19248 25900 19472 25906
rect 19300 25894 19472 25900
rect 19800 25900 19852 25906
rect 19248 25842 19300 25848
rect 19800 25842 19852 25848
rect 19812 25786 19840 25842
rect 19996 25838 20024 27270
rect 20168 26784 20220 26790
rect 20168 26726 20220 26732
rect 20180 26518 20208 26726
rect 20168 26512 20220 26518
rect 20168 26454 20220 26460
rect 20076 26444 20128 26450
rect 20076 26386 20128 26392
rect 19984 25832 20036 25838
rect 19340 25764 19392 25770
rect 19812 25758 19932 25786
rect 19984 25774 20036 25780
rect 19340 25706 19392 25712
rect 18418 25528 18474 25537
rect 19352 25498 19380 25706
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 18418 25463 18420 25472
rect 18472 25463 18474 25472
rect 19340 25492 19392 25498
rect 18420 25434 18472 25440
rect 19340 25434 19392 25440
rect 17960 25288 18012 25294
rect 17788 25236 17960 25242
rect 17788 25230 18012 25236
rect 17788 25214 18000 25230
rect 17788 24614 17816 25214
rect 17868 25152 17920 25158
rect 17868 25094 17920 25100
rect 17776 24608 17828 24614
rect 17776 24550 17828 24556
rect 17408 23112 17460 23118
rect 17408 23054 17460 23060
rect 17224 22772 17276 22778
rect 17224 22714 17276 22720
rect 17040 22636 17092 22642
rect 17040 22578 17092 22584
rect 17408 22636 17460 22642
rect 17408 22578 17460 22584
rect 17040 22500 17092 22506
rect 17040 22442 17092 22448
rect 16856 22432 16908 22438
rect 16856 22374 16908 22380
rect 16868 22273 16896 22374
rect 16854 22264 16910 22273
rect 13544 21966 13596 21972
rect 13634 21992 13690 22001
rect 13634 21927 13690 21936
rect 13728 21140 13780 21146
rect 13728 21082 13780 21088
rect 13266 20632 13322 20641
rect 12992 20596 13044 20602
rect 13266 20567 13322 20576
rect 12992 20538 13044 20544
rect 13740 20398 13768 21082
rect 13268 20392 13320 20398
rect 13268 20334 13320 20340
rect 13728 20392 13780 20398
rect 13728 20334 13780 20340
rect 12624 20256 12676 20262
rect 12624 20198 12676 20204
rect 2780 20052 2832 20058
rect 2780 19994 2832 20000
rect 12440 20052 12492 20058
rect 12440 19994 12492 20000
rect 12636 19922 12664 20198
rect 13280 20058 13308 20334
rect 14016 20330 14044 22222
rect 14096 22228 14148 22234
rect 14096 22170 14148 22176
rect 14648 22228 14700 22234
rect 14648 22170 14700 22176
rect 15292 22228 15344 22234
rect 15292 22170 15344 22176
rect 16396 22228 16448 22234
rect 17052 22234 17080 22442
rect 17420 22234 17448 22578
rect 16854 22199 16910 22208
rect 17040 22228 17092 22234
rect 16396 22170 16448 22176
rect 17040 22170 17092 22176
rect 17408 22228 17460 22234
rect 17408 22170 17460 22176
rect 14108 21350 14136 22170
rect 14648 22092 14700 22098
rect 14648 22034 14700 22040
rect 16856 22092 16908 22098
rect 16856 22034 16908 22040
rect 14660 21690 14688 22034
rect 15016 22024 15068 22030
rect 15752 22024 15804 22030
rect 15016 21966 15068 21972
rect 15750 21992 15752 22001
rect 16028 22024 16080 22030
rect 15804 21992 15806 22001
rect 14648 21684 14700 21690
rect 14648 21626 14700 21632
rect 14660 21418 14688 21626
rect 14648 21412 14700 21418
rect 14648 21354 14700 21360
rect 14096 21344 14148 21350
rect 14096 21286 14148 21292
rect 14108 21146 14136 21286
rect 14096 21140 14148 21146
rect 14096 21082 14148 21088
rect 15028 20466 15056 21966
rect 16028 21966 16080 21972
rect 15750 21927 15806 21936
rect 15844 21956 15896 21962
rect 15764 21690 15792 21927
rect 15844 21898 15896 21904
rect 15856 21690 15884 21898
rect 15752 21684 15804 21690
rect 15752 21626 15804 21632
rect 15844 21684 15896 21690
rect 15844 21626 15896 21632
rect 15292 21140 15344 21146
rect 15292 21082 15344 21088
rect 15304 21049 15332 21082
rect 15290 21040 15346 21049
rect 15290 20975 15346 20984
rect 16040 20942 16068 21966
rect 16868 21690 16896 22034
rect 16856 21684 16908 21690
rect 16856 21626 16908 21632
rect 17788 21554 17816 24550
rect 17880 24274 17908 25094
rect 18432 24954 18460 25434
rect 19904 25430 19932 25758
rect 20088 25498 20116 26386
rect 20364 26314 20392 27338
rect 20548 27169 20576 39520
rect 21456 36032 21508 36038
rect 21456 35974 21508 35980
rect 21468 35630 21496 35974
rect 20996 35624 21048 35630
rect 20996 35566 21048 35572
rect 21456 35624 21508 35630
rect 21456 35566 21508 35572
rect 20626 34776 20682 34785
rect 21008 34746 21036 35566
rect 21180 35488 21232 35494
rect 21180 35430 21232 35436
rect 21364 35488 21416 35494
rect 21364 35430 21416 35436
rect 21088 35216 21140 35222
rect 21088 35158 21140 35164
rect 20626 34711 20628 34720
rect 20680 34711 20682 34720
rect 20996 34740 21048 34746
rect 20628 34682 20680 34688
rect 20996 34682 21048 34688
rect 20640 34542 20668 34682
rect 21100 34542 21128 35158
rect 20628 34536 20680 34542
rect 20628 34478 20680 34484
rect 21088 34536 21140 34542
rect 21088 34478 21140 34484
rect 21100 34134 21128 34478
rect 21088 34128 21140 34134
rect 21088 34070 21140 34076
rect 21192 34066 21220 35430
rect 20720 34060 20772 34066
rect 20720 34002 20772 34008
rect 21180 34060 21232 34066
rect 21180 34002 21232 34008
rect 20732 33522 20760 34002
rect 21192 33640 21220 34002
rect 21376 33833 21404 35430
rect 21456 34944 21508 34950
rect 21456 34886 21508 34892
rect 21362 33824 21418 33833
rect 21362 33759 21418 33768
rect 21364 33652 21416 33658
rect 21192 33612 21364 33640
rect 20720 33516 20772 33522
rect 20720 33458 20772 33464
rect 20732 33114 20760 33458
rect 21192 33114 21220 33612
rect 21364 33594 21416 33600
rect 21468 33153 21496 34886
rect 21454 33144 21510 33153
rect 20720 33108 20772 33114
rect 20720 33050 20772 33056
rect 21180 33108 21232 33114
rect 21454 33079 21510 33088
rect 21180 33050 21232 33056
rect 20732 32570 20760 33050
rect 20720 32564 20772 32570
rect 20720 32506 20772 32512
rect 21548 31884 21600 31890
rect 21548 31826 21600 31832
rect 20996 31816 21048 31822
rect 20996 31758 21048 31764
rect 21008 31346 21036 31758
rect 20996 31340 21048 31346
rect 20996 31282 21048 31288
rect 21008 30802 21036 31282
rect 21560 31278 21588 31826
rect 21548 31272 21600 31278
rect 21548 31214 21600 31220
rect 21088 31204 21140 31210
rect 21088 31146 21140 31152
rect 21100 30870 21128 31146
rect 21560 30938 21588 31214
rect 21548 30932 21600 30938
rect 21548 30874 21600 30880
rect 21088 30864 21140 30870
rect 21088 30806 21140 30812
rect 20996 30796 21048 30802
rect 20996 30738 21048 30744
rect 21008 29782 21036 30738
rect 21100 30394 21128 30806
rect 21088 30388 21140 30394
rect 21088 30330 21140 30336
rect 21100 29850 21128 30330
rect 21088 29844 21140 29850
rect 21088 29786 21140 29792
rect 20996 29776 21048 29782
rect 20996 29718 21048 29724
rect 20720 28620 20772 28626
rect 20720 28562 20772 28568
rect 21180 28620 21232 28626
rect 21180 28562 21232 28568
rect 20628 27872 20680 27878
rect 20628 27814 20680 27820
rect 20640 27418 20668 27814
rect 20732 27606 20760 28562
rect 21192 28082 21220 28562
rect 21652 28370 21680 39520
rect 22468 36236 22520 36242
rect 22468 36178 22520 36184
rect 22480 35834 22508 36178
rect 22560 36032 22612 36038
rect 22560 35974 22612 35980
rect 22468 35828 22520 35834
rect 22468 35770 22520 35776
rect 22100 35692 22152 35698
rect 22100 35634 22152 35640
rect 21916 35148 21968 35154
rect 21916 35090 21968 35096
rect 21928 34950 21956 35090
rect 21916 34944 21968 34950
rect 21916 34886 21968 34892
rect 21928 34513 21956 34886
rect 21914 34504 21970 34513
rect 21914 34439 21970 34448
rect 22112 33998 22140 35634
rect 22468 35148 22520 35154
rect 22468 35090 22520 35096
rect 22480 34746 22508 35090
rect 22468 34740 22520 34746
rect 22468 34682 22520 34688
rect 22192 34468 22244 34474
rect 22192 34410 22244 34416
rect 22204 34202 22232 34410
rect 22192 34196 22244 34202
rect 22192 34138 22244 34144
rect 22100 33992 22152 33998
rect 22100 33934 22152 33940
rect 21916 33584 21968 33590
rect 21916 33526 21968 33532
rect 21732 33380 21784 33386
rect 21732 33322 21784 33328
rect 21744 33046 21772 33322
rect 21732 33040 21784 33046
rect 21732 32982 21784 32988
rect 21744 32570 21772 32982
rect 21824 32972 21876 32978
rect 21824 32914 21876 32920
rect 21732 32564 21784 32570
rect 21732 32506 21784 32512
rect 21836 32366 21864 32914
rect 21928 32910 21956 33526
rect 22112 33522 22140 33934
rect 22100 33516 22152 33522
rect 22100 33458 22152 33464
rect 22572 33046 22600 35974
rect 22756 34785 22784 39520
rect 23860 36242 23888 39520
rect 23848 36236 23900 36242
rect 23848 36178 23900 36184
rect 24964 35850 24992 39520
rect 26068 39494 26188 39520
rect 24780 35834 24992 35850
rect 24768 35828 24992 35834
rect 24820 35822 24992 35828
rect 24768 35770 24820 35776
rect 25688 35624 25740 35630
rect 25134 35592 25190 35601
rect 25688 35566 25740 35572
rect 25134 35527 25190 35536
rect 25596 35556 25648 35562
rect 22928 35216 22980 35222
rect 22928 35158 22980 35164
rect 22742 34776 22798 34785
rect 22742 34711 22798 34720
rect 22940 34610 22968 35158
rect 24032 34944 24084 34950
rect 24032 34886 24084 34892
rect 24216 34944 24268 34950
rect 24216 34886 24268 34892
rect 23388 34740 23440 34746
rect 23388 34682 23440 34688
rect 22928 34604 22980 34610
rect 22928 34546 22980 34552
rect 22940 34202 22968 34546
rect 23400 34218 23428 34682
rect 23662 34504 23718 34513
rect 23662 34439 23718 34448
rect 23400 34202 23520 34218
rect 22928 34196 22980 34202
rect 23400 34196 23532 34202
rect 23400 34190 23480 34196
rect 22928 34138 22980 34144
rect 23480 34138 23532 34144
rect 23112 34060 23164 34066
rect 23112 34002 23164 34008
rect 23124 33658 23152 34002
rect 23388 33856 23440 33862
rect 23388 33798 23440 33804
rect 23112 33652 23164 33658
rect 23112 33594 23164 33600
rect 23400 33454 23428 33798
rect 23492 33658 23520 34138
rect 23676 33658 23704 34439
rect 24044 34406 24072 34886
rect 24228 34610 24256 34886
rect 25042 34776 25098 34785
rect 25042 34711 25098 34720
rect 24216 34604 24268 34610
rect 24216 34546 24268 34552
rect 24032 34400 24084 34406
rect 24032 34342 24084 34348
rect 24044 34066 24072 34342
rect 24032 34060 24084 34066
rect 24032 34002 24084 34008
rect 24400 33856 24452 33862
rect 24122 33824 24178 33833
rect 24400 33798 24452 33804
rect 24122 33759 24178 33768
rect 23480 33652 23532 33658
rect 23480 33594 23532 33600
rect 23664 33652 23716 33658
rect 23664 33594 23716 33600
rect 24136 33522 24164 33759
rect 24412 33522 24440 33798
rect 24124 33516 24176 33522
rect 24124 33458 24176 33464
rect 24400 33516 24452 33522
rect 24400 33458 24452 33464
rect 23388 33448 23440 33454
rect 23388 33390 23440 33396
rect 24308 33448 24360 33454
rect 24308 33390 24360 33396
rect 23572 33380 23624 33386
rect 23572 33322 23624 33328
rect 23296 33108 23348 33114
rect 23296 33050 23348 33056
rect 22560 33040 22612 33046
rect 22560 32982 22612 32988
rect 21916 32904 21968 32910
rect 21916 32846 21968 32852
rect 21824 32360 21876 32366
rect 21824 32302 21876 32308
rect 21836 32026 21864 32302
rect 21824 32020 21876 32026
rect 21824 31962 21876 31968
rect 21928 31958 21956 32846
rect 23308 31958 23336 33050
rect 23584 33046 23612 33322
rect 23938 33144 23994 33153
rect 24320 33114 24348 33390
rect 24768 33380 24820 33386
rect 24768 33322 24820 33328
rect 23938 33079 23940 33088
rect 23992 33079 23994 33088
rect 24308 33108 24360 33114
rect 23940 33050 23992 33056
rect 24308 33050 24360 33056
rect 23572 33040 23624 33046
rect 23572 32982 23624 32988
rect 23388 32904 23440 32910
rect 23388 32846 23440 32852
rect 23400 32026 23428 32846
rect 23480 32768 23532 32774
rect 23480 32710 23532 32716
rect 23388 32020 23440 32026
rect 23388 31962 23440 31968
rect 21916 31952 21968 31958
rect 21916 31894 21968 31900
rect 22008 31952 22060 31958
rect 22008 31894 22060 31900
rect 23296 31952 23348 31958
rect 23296 31894 23348 31900
rect 21928 31414 21956 31894
rect 22020 31482 22048 31894
rect 23492 31890 23520 32710
rect 23952 32366 23980 33050
rect 24674 33008 24730 33017
rect 24674 32943 24676 32952
rect 24728 32943 24730 32952
rect 24676 32914 24728 32920
rect 24216 32564 24268 32570
rect 24216 32506 24268 32512
rect 24124 32428 24176 32434
rect 24124 32370 24176 32376
rect 23940 32360 23992 32366
rect 23940 32302 23992 32308
rect 23572 32292 23624 32298
rect 23572 32234 23624 32240
rect 23584 32026 23612 32234
rect 24136 32026 24164 32370
rect 23572 32020 23624 32026
rect 23572 31962 23624 31968
rect 24124 32020 24176 32026
rect 24124 31962 24176 31968
rect 24228 31958 24256 32506
rect 24688 32434 24716 32914
rect 24676 32428 24728 32434
rect 24676 32370 24728 32376
rect 24216 31952 24268 31958
rect 24216 31894 24268 31900
rect 23480 31884 23532 31890
rect 23480 31826 23532 31832
rect 23492 31482 23520 31826
rect 24124 31816 24176 31822
rect 24124 31758 24176 31764
rect 22008 31476 22060 31482
rect 22008 31418 22060 31424
rect 23480 31476 23532 31482
rect 23480 31418 23532 31424
rect 21916 31408 21968 31414
rect 21916 31350 21968 31356
rect 24032 31340 24084 31346
rect 24032 31282 24084 31288
rect 24044 30938 24072 31282
rect 24032 30932 24084 30938
rect 24032 30874 24084 30880
rect 23480 30796 23532 30802
rect 23480 30738 23532 30744
rect 23492 30394 23520 30738
rect 23756 30592 23808 30598
rect 23756 30534 23808 30540
rect 23768 30394 23796 30534
rect 23480 30388 23532 30394
rect 23480 30330 23532 30336
rect 23756 30388 23808 30394
rect 23756 30330 23808 30336
rect 24044 30190 24072 30874
rect 24032 30184 24084 30190
rect 24032 30126 24084 30132
rect 24136 29850 24164 31758
rect 24228 31482 24256 31894
rect 24780 31890 24808 33322
rect 24860 32768 24912 32774
rect 24860 32710 24912 32716
rect 24872 32026 24900 32710
rect 24860 32020 24912 32026
rect 24860 31962 24912 31968
rect 24768 31884 24820 31890
rect 24768 31826 24820 31832
rect 24676 31680 24728 31686
rect 24676 31622 24728 31628
rect 24216 31476 24268 31482
rect 24216 31418 24268 31424
rect 24228 30802 24256 31418
rect 24688 31113 24716 31622
rect 24674 31104 24730 31113
rect 24674 31039 24730 31048
rect 24676 30932 24728 30938
rect 24676 30874 24728 30880
rect 24216 30796 24268 30802
rect 24216 30738 24268 30744
rect 24584 30796 24636 30802
rect 24584 30738 24636 30744
rect 24124 29844 24176 29850
rect 24124 29786 24176 29792
rect 23570 29744 23626 29753
rect 23570 29679 23572 29688
rect 23624 29679 23626 29688
rect 23572 29650 23624 29656
rect 23584 29306 23612 29650
rect 24492 29504 24544 29510
rect 24492 29446 24544 29452
rect 23572 29300 23624 29306
rect 23572 29242 23624 29248
rect 24032 29096 24084 29102
rect 24032 29038 24084 29044
rect 24044 28762 24072 29038
rect 24124 28960 24176 28966
rect 24124 28902 24176 28908
rect 24032 28756 24084 28762
rect 24032 28698 24084 28704
rect 22282 28520 22338 28529
rect 22282 28455 22284 28464
rect 22336 28455 22338 28464
rect 22284 28426 22336 28432
rect 21560 28342 21680 28370
rect 21180 28076 21232 28082
rect 21180 28018 21232 28024
rect 20812 27872 20864 27878
rect 20812 27814 20864 27820
rect 21456 27872 21508 27878
rect 21456 27814 21508 27820
rect 20720 27600 20772 27606
rect 20720 27542 20772 27548
rect 20640 27390 20760 27418
rect 20534 27160 20590 27169
rect 20534 27095 20590 27104
rect 20352 26308 20404 26314
rect 20352 26250 20404 26256
rect 20536 26308 20588 26314
rect 20536 26250 20588 26256
rect 20548 25906 20576 26250
rect 20536 25900 20588 25906
rect 20536 25842 20588 25848
rect 20628 25832 20680 25838
rect 20628 25774 20680 25780
rect 20260 25696 20312 25702
rect 20260 25638 20312 25644
rect 20076 25492 20128 25498
rect 20076 25434 20128 25440
rect 19892 25424 19944 25430
rect 19892 25366 19944 25372
rect 18604 25356 18656 25362
rect 18604 25298 18656 25304
rect 18420 24948 18472 24954
rect 18420 24890 18472 24896
rect 18616 24614 18644 25298
rect 20272 24954 20300 25638
rect 20640 25378 20668 25774
rect 20732 25702 20760 27390
rect 20824 25786 20852 27814
rect 21468 27674 21496 27814
rect 21456 27668 21508 27674
rect 21456 27610 21508 27616
rect 20904 27600 20956 27606
rect 20904 27542 20956 27548
rect 20916 26382 20944 27542
rect 21272 26784 21324 26790
rect 21272 26726 21324 26732
rect 20904 26376 20956 26382
rect 20904 26318 20956 26324
rect 21284 25906 21312 26726
rect 20996 25900 21048 25906
rect 20996 25842 21048 25848
rect 21272 25900 21324 25906
rect 21272 25842 21324 25848
rect 20904 25832 20956 25838
rect 20824 25780 20904 25786
rect 21008 25809 21036 25842
rect 20824 25774 20956 25780
rect 20994 25800 21050 25809
rect 20824 25758 20944 25774
rect 20720 25696 20772 25702
rect 20720 25638 20772 25644
rect 20824 25498 20852 25758
rect 20994 25735 21050 25744
rect 20812 25492 20864 25498
rect 20812 25434 20864 25440
rect 20640 25350 20852 25378
rect 20720 25288 20772 25294
rect 20720 25230 20772 25236
rect 20260 24948 20312 24954
rect 20260 24890 20312 24896
rect 18972 24744 19024 24750
rect 18972 24686 19024 24692
rect 19892 24744 19944 24750
rect 19892 24686 19944 24692
rect 18604 24608 18656 24614
rect 18602 24576 18604 24585
rect 18656 24576 18658 24585
rect 18602 24511 18658 24520
rect 18984 24274 19012 24686
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 17868 24268 17920 24274
rect 17868 24210 17920 24216
rect 18512 24268 18564 24274
rect 18512 24210 18564 24216
rect 18972 24268 19024 24274
rect 18972 24210 19024 24216
rect 18236 24132 18288 24138
rect 18236 24074 18288 24080
rect 18248 23322 18276 24074
rect 18420 24064 18472 24070
rect 18420 24006 18472 24012
rect 18432 23662 18460 24006
rect 18420 23656 18472 23662
rect 18420 23598 18472 23604
rect 18236 23316 18288 23322
rect 18236 23258 18288 23264
rect 18144 23180 18196 23186
rect 18144 23122 18196 23128
rect 18156 22234 18184 23122
rect 18432 22710 18460 23598
rect 18524 23526 18552 24210
rect 18788 24200 18840 24206
rect 18788 24142 18840 24148
rect 18604 24064 18656 24070
rect 18604 24006 18656 24012
rect 18512 23520 18564 23526
rect 18512 23462 18564 23468
rect 18420 22704 18472 22710
rect 18420 22646 18472 22652
rect 18144 22228 18196 22234
rect 18144 22170 18196 22176
rect 18616 22098 18644 24006
rect 18696 23520 18748 23526
rect 18696 23462 18748 23468
rect 18708 23186 18736 23462
rect 18800 23322 18828 24142
rect 19340 24132 19392 24138
rect 19340 24074 19392 24080
rect 19062 23896 19118 23905
rect 19062 23831 19064 23840
rect 19116 23831 19118 23840
rect 19064 23802 19116 23808
rect 19064 23656 19116 23662
rect 19064 23598 19116 23604
rect 19154 23624 19210 23633
rect 18788 23316 18840 23322
rect 18788 23258 18840 23264
rect 18696 23180 18748 23186
rect 18696 23122 18748 23128
rect 18800 23050 18828 23258
rect 18788 23044 18840 23050
rect 18788 22986 18840 22992
rect 18800 22642 18828 22986
rect 19076 22778 19104 23598
rect 19154 23559 19210 23568
rect 19168 23526 19196 23559
rect 19352 23526 19380 24074
rect 19524 24064 19576 24070
rect 19524 24006 19576 24012
rect 19800 24064 19852 24070
rect 19800 24006 19852 24012
rect 19432 23724 19484 23730
rect 19432 23666 19484 23672
rect 19156 23520 19208 23526
rect 19340 23520 19392 23526
rect 19156 23462 19208 23468
rect 19260 23480 19340 23508
rect 19156 23180 19208 23186
rect 19156 23122 19208 23128
rect 19064 22772 19116 22778
rect 19064 22714 19116 22720
rect 18788 22636 18840 22642
rect 18788 22578 18840 22584
rect 19168 22574 19196 23122
rect 19156 22568 19208 22574
rect 19156 22510 19208 22516
rect 18604 22092 18656 22098
rect 18604 22034 18656 22040
rect 17132 21548 17184 21554
rect 17132 21490 17184 21496
rect 17776 21548 17828 21554
rect 17776 21490 17828 21496
rect 16764 21344 16816 21350
rect 16764 21286 16816 21292
rect 16856 21344 16908 21350
rect 16856 21286 16908 21292
rect 16776 21146 16804 21286
rect 16764 21140 16816 21146
rect 16764 21082 16816 21088
rect 16488 21004 16540 21010
rect 16488 20946 16540 20952
rect 15752 20936 15804 20942
rect 15752 20878 15804 20884
rect 16028 20936 16080 20942
rect 16028 20878 16080 20884
rect 15764 20602 15792 20878
rect 16500 20618 16528 20946
rect 16868 20874 16896 21286
rect 17144 21078 17172 21490
rect 17960 21344 18012 21350
rect 17960 21286 18012 21292
rect 17132 21072 17184 21078
rect 17132 21014 17184 21020
rect 17972 21010 18000 21286
rect 18616 21146 18644 22034
rect 19168 21894 19196 22510
rect 19260 21962 19288 23480
rect 19340 23462 19392 23468
rect 19444 23254 19472 23666
rect 19536 23662 19564 24006
rect 19812 23730 19840 24006
rect 19800 23724 19852 23730
rect 19800 23666 19852 23672
rect 19524 23656 19576 23662
rect 19524 23598 19576 23604
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 19580 23344 19876 23364
rect 19432 23248 19484 23254
rect 19432 23190 19484 23196
rect 19444 22778 19472 23190
rect 19904 23186 19932 24686
rect 20260 24676 20312 24682
rect 20260 24618 20312 24624
rect 20074 24304 20130 24313
rect 20074 24239 20130 24248
rect 19892 23180 19944 23186
rect 19892 23122 19944 23128
rect 19432 22772 19484 22778
rect 19432 22714 19484 22720
rect 19338 22264 19394 22273
rect 19338 22199 19394 22208
rect 19248 21956 19300 21962
rect 19248 21898 19300 21904
rect 19156 21888 19208 21894
rect 19156 21830 19208 21836
rect 19168 21486 19196 21830
rect 19156 21480 19208 21486
rect 19156 21422 19208 21428
rect 19248 21412 19300 21418
rect 19248 21354 19300 21360
rect 18604 21140 18656 21146
rect 18604 21082 18656 21088
rect 19154 21040 19210 21049
rect 17960 21004 18012 21010
rect 17960 20946 18012 20952
rect 18328 21004 18380 21010
rect 19154 20975 19156 20984
rect 18328 20946 18380 20952
rect 19208 20975 19210 20984
rect 19156 20946 19208 20952
rect 16856 20868 16908 20874
rect 16856 20810 16908 20816
rect 17868 20868 17920 20874
rect 17868 20810 17920 20816
rect 16672 20800 16724 20806
rect 16672 20742 16724 20748
rect 16500 20602 16620 20618
rect 15752 20596 15804 20602
rect 15752 20538 15804 20544
rect 16500 20596 16632 20602
rect 16500 20590 16580 20596
rect 15016 20460 15068 20466
rect 15016 20402 15068 20408
rect 16396 20460 16448 20466
rect 16396 20402 16448 20408
rect 14004 20324 14056 20330
rect 14004 20266 14056 20272
rect 13728 20256 13780 20262
rect 13728 20198 13780 20204
rect 13268 20052 13320 20058
rect 13268 19994 13320 20000
rect 13452 20052 13504 20058
rect 13452 19994 13504 20000
rect 1952 19916 2004 19922
rect 1952 19858 2004 19864
rect 12624 19916 12676 19922
rect 12624 19858 12676 19864
rect 1964 19514 1992 19858
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 1584 19508 1636 19514
rect 1584 19450 1636 19456
rect 1952 19508 2004 19514
rect 1952 19450 2004 19456
rect 13464 19378 13492 19994
rect 13544 19916 13596 19922
rect 13544 19858 13596 19864
rect 13452 19372 13504 19378
rect 13452 19314 13504 19320
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 13464 18222 13492 19314
rect 13556 18970 13584 19858
rect 13740 19310 13768 20198
rect 14016 20058 14044 20266
rect 15028 20058 15056 20402
rect 15752 20256 15804 20262
rect 15752 20198 15804 20204
rect 15764 20058 15792 20198
rect 14004 20052 14056 20058
rect 14004 19994 14056 20000
rect 15016 20052 15068 20058
rect 15016 19994 15068 20000
rect 15752 20052 15804 20058
rect 15752 19994 15804 20000
rect 15764 19514 15792 19994
rect 16212 19916 16264 19922
rect 16212 19858 16264 19864
rect 14832 19508 14884 19514
rect 14832 19450 14884 19456
rect 15752 19508 15804 19514
rect 15752 19450 15804 19456
rect 13728 19304 13780 19310
rect 13728 19246 13780 19252
rect 13544 18964 13596 18970
rect 13544 18906 13596 18912
rect 14004 18760 14056 18766
rect 14004 18702 14056 18708
rect 14016 18222 14044 18702
rect 14844 18222 14872 19450
rect 16224 19310 16252 19858
rect 16408 19378 16436 20402
rect 16396 19372 16448 19378
rect 16396 19314 16448 19320
rect 16212 19304 16264 19310
rect 16212 19246 16264 19252
rect 15844 19236 15896 19242
rect 15844 19178 15896 19184
rect 15856 18902 15884 19178
rect 16224 18970 16252 19246
rect 16500 19174 16528 20590
rect 16580 20538 16632 20544
rect 16684 19990 16712 20742
rect 17880 20482 17908 20810
rect 17972 20602 18000 20946
rect 18236 20936 18288 20942
rect 18236 20878 18288 20884
rect 17960 20596 18012 20602
rect 17960 20538 18012 20544
rect 17880 20454 18000 20482
rect 17972 20058 18000 20454
rect 18052 20392 18104 20398
rect 18052 20334 18104 20340
rect 17960 20052 18012 20058
rect 17960 19994 18012 20000
rect 16672 19984 16724 19990
rect 16672 19926 16724 19932
rect 17868 19848 17920 19854
rect 17868 19790 17920 19796
rect 17880 19514 17908 19790
rect 17960 19712 18012 19718
rect 17960 19654 18012 19660
rect 17868 19508 17920 19514
rect 17868 19450 17920 19456
rect 16488 19168 16540 19174
rect 16488 19110 16540 19116
rect 16212 18964 16264 18970
rect 16212 18906 16264 18912
rect 15844 18896 15896 18902
rect 15844 18838 15896 18844
rect 15856 18426 15884 18838
rect 16304 18624 16356 18630
rect 16304 18566 16356 18572
rect 15844 18420 15896 18426
rect 15844 18362 15896 18368
rect 13452 18216 13504 18222
rect 13452 18158 13504 18164
rect 14004 18216 14056 18222
rect 14004 18158 14056 18164
rect 14832 18216 14884 18222
rect 14832 18158 14884 18164
rect 14016 17882 14044 18158
rect 16316 18086 16344 18566
rect 17880 18426 17908 19450
rect 17972 19378 18000 19654
rect 17960 19372 18012 19378
rect 17960 19314 18012 19320
rect 18064 19310 18092 20334
rect 18248 19718 18276 20878
rect 18340 20330 18368 20946
rect 19260 20618 19288 21354
rect 19352 21146 19380 22199
rect 19444 22166 19472 22714
rect 19984 22568 20036 22574
rect 19984 22510 20036 22516
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 19432 22160 19484 22166
rect 19432 22102 19484 22108
rect 19996 21690 20024 22510
rect 19984 21684 20036 21690
rect 19984 21626 20036 21632
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 19340 21140 19392 21146
rect 19340 21082 19392 21088
rect 19524 21004 19576 21010
rect 19524 20946 19576 20952
rect 19260 20602 19380 20618
rect 19536 20602 19564 20946
rect 19260 20596 19392 20602
rect 19260 20590 19340 20596
rect 19340 20538 19392 20544
rect 19524 20596 19576 20602
rect 19524 20538 19576 20544
rect 18328 20324 18380 20330
rect 18328 20266 18380 20272
rect 18236 19712 18288 19718
rect 18236 19654 18288 19660
rect 18340 19514 18368 20266
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 19580 20080 19876 20100
rect 18788 19916 18840 19922
rect 18788 19858 18840 19864
rect 18328 19508 18380 19514
rect 18328 19450 18380 19456
rect 18052 19304 18104 19310
rect 18052 19246 18104 19252
rect 18064 18630 18092 19246
rect 18800 19242 18828 19858
rect 18144 19236 18196 19242
rect 18144 19178 18196 19184
rect 18788 19236 18840 19242
rect 18788 19178 18840 19184
rect 18156 18970 18184 19178
rect 19984 19168 20036 19174
rect 19984 19110 20036 19116
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 18144 18964 18196 18970
rect 18144 18906 18196 18912
rect 18420 18828 18472 18834
rect 18420 18770 18472 18776
rect 18052 18624 18104 18630
rect 18052 18566 18104 18572
rect 17868 18420 17920 18426
rect 17868 18362 17920 18368
rect 18064 18222 18092 18566
rect 18052 18216 18104 18222
rect 18052 18158 18104 18164
rect 16304 18080 16356 18086
rect 16304 18022 16356 18028
rect 16316 17882 16344 18022
rect 18064 17882 18092 18158
rect 14004 17876 14056 17882
rect 14004 17818 14056 17824
rect 16304 17876 16356 17882
rect 16304 17818 16356 17824
rect 18052 17876 18104 17882
rect 18052 17818 18104 17824
rect 18432 17542 18460 18770
rect 19996 18358 20024 19110
rect 20088 18766 20116 24239
rect 20272 24138 20300 24618
rect 20732 24342 20760 25230
rect 20824 24410 20852 25350
rect 20904 25288 20956 25294
rect 20904 25230 20956 25236
rect 20916 24750 20944 25230
rect 21284 24954 21312 25842
rect 21456 25424 21508 25430
rect 21456 25366 21508 25372
rect 21468 24954 21496 25366
rect 21272 24948 21324 24954
rect 21272 24890 21324 24896
rect 21456 24948 21508 24954
rect 21456 24890 21508 24896
rect 20904 24744 20956 24750
rect 20904 24686 20956 24692
rect 20812 24404 20864 24410
rect 20812 24346 20864 24352
rect 20720 24336 20772 24342
rect 20720 24278 20772 24284
rect 20260 24132 20312 24138
rect 20260 24074 20312 24080
rect 20272 23866 20300 24074
rect 20732 23866 20760 24278
rect 20916 24274 20944 24686
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 21088 24200 21140 24206
rect 21088 24142 21140 24148
rect 20260 23860 20312 23866
rect 20260 23802 20312 23808
rect 20720 23860 20772 23866
rect 20720 23802 20772 23808
rect 20272 23322 20300 23802
rect 21100 23633 21128 24142
rect 21560 23905 21588 28342
rect 21638 28248 21694 28257
rect 21638 28183 21640 28192
rect 21692 28183 21694 28192
rect 21640 28154 21692 28160
rect 22468 28076 22520 28082
rect 22468 28018 22520 28024
rect 21640 27872 21692 27878
rect 21640 27814 21692 27820
rect 21652 27130 21680 27814
rect 22480 27674 22508 28018
rect 24136 27713 24164 28902
rect 24504 27860 24532 29446
rect 24596 29102 24624 30738
rect 24688 30326 24716 30874
rect 24872 30818 24900 31962
rect 25056 30954 25084 34711
rect 24780 30802 24900 30818
rect 24768 30796 24900 30802
rect 24820 30790 24900 30796
rect 24964 30926 25084 30954
rect 24768 30738 24820 30744
rect 24768 30592 24820 30598
rect 24768 30534 24820 30540
rect 24676 30320 24728 30326
rect 24676 30262 24728 30268
rect 24780 29594 24808 30534
rect 24860 29640 24912 29646
rect 24780 29588 24860 29594
rect 24780 29582 24912 29588
rect 24780 29566 24900 29582
rect 24584 29096 24636 29102
rect 24584 29038 24636 29044
rect 24676 29028 24728 29034
rect 24676 28970 24728 28976
rect 24688 28694 24716 28970
rect 24780 28762 24808 29566
rect 24860 28960 24912 28966
rect 24860 28902 24912 28908
rect 24768 28756 24820 28762
rect 24768 28698 24820 28704
rect 24676 28688 24728 28694
rect 24676 28630 24728 28636
rect 24584 28552 24636 28558
rect 24584 28494 24636 28500
rect 24596 28218 24624 28494
rect 24584 28212 24636 28218
rect 24584 28154 24636 28160
rect 24872 28082 24900 28902
rect 24860 28076 24912 28082
rect 24860 28018 24912 28024
rect 24872 27962 24900 28018
rect 24780 27934 24900 27962
rect 24584 27872 24636 27878
rect 24504 27832 24584 27860
rect 24584 27814 24636 27820
rect 24122 27704 24178 27713
rect 22468 27668 22520 27674
rect 24122 27639 24178 27648
rect 22468 27610 22520 27616
rect 21732 27532 21784 27538
rect 21732 27474 21784 27480
rect 21640 27124 21692 27130
rect 21640 27066 21692 27072
rect 21744 26994 21772 27474
rect 24596 27334 24624 27814
rect 24780 27606 24808 27934
rect 24768 27600 24820 27606
rect 24768 27542 24820 27548
rect 24964 27402 24992 30926
rect 25044 30796 25096 30802
rect 25044 30738 25096 30744
rect 25056 30394 25084 30738
rect 25044 30388 25096 30394
rect 25044 30330 25096 30336
rect 25044 29708 25096 29714
rect 25044 29650 25096 29656
rect 25056 29238 25084 29650
rect 25044 29232 25096 29238
rect 25044 29174 25096 29180
rect 25044 29096 25096 29102
rect 25044 29038 25096 29044
rect 25056 28422 25084 29038
rect 25148 28762 25176 35527
rect 25596 35498 25648 35504
rect 25608 34746 25636 35498
rect 25700 34950 25728 35566
rect 25688 34944 25740 34950
rect 25688 34886 25740 34892
rect 25596 34740 25648 34746
rect 25596 34682 25648 34688
rect 25320 34060 25372 34066
rect 25320 34002 25372 34008
rect 25332 33318 25360 34002
rect 25504 33856 25556 33862
rect 25504 33798 25556 33804
rect 25320 33312 25372 33318
rect 25320 33254 25372 33260
rect 25516 33114 25544 33798
rect 25608 33658 25636 34682
rect 25964 34060 26016 34066
rect 25964 34002 26016 34008
rect 25780 33924 25832 33930
rect 25780 33866 25832 33872
rect 25596 33652 25648 33658
rect 25596 33594 25648 33600
rect 25504 33108 25556 33114
rect 25504 33050 25556 33056
rect 25228 33040 25280 33046
rect 25228 32982 25280 32988
rect 25240 32502 25268 32982
rect 25516 32570 25544 33050
rect 25792 33046 25820 33866
rect 25872 33448 25924 33454
rect 25872 33390 25924 33396
rect 25884 33114 25912 33390
rect 25872 33108 25924 33114
rect 25872 33050 25924 33056
rect 25780 33040 25832 33046
rect 25780 32982 25832 32988
rect 25976 32570 26004 34002
rect 26160 32994 26188 39494
rect 27264 35737 27292 39520
rect 27250 35728 27306 35737
rect 27250 35663 27306 35672
rect 26976 35488 27028 35494
rect 26976 35430 27028 35436
rect 26700 34944 26752 34950
rect 26700 34886 26752 34892
rect 26712 34610 26740 34886
rect 26700 34604 26752 34610
rect 26700 34546 26752 34552
rect 26988 34542 27016 35430
rect 29472 35193 29500 39520
rect 29458 35184 29514 35193
rect 28080 35148 28132 35154
rect 29458 35119 29514 35128
rect 28080 35090 28132 35096
rect 28092 34746 28120 35090
rect 30576 35057 30604 39520
rect 30562 35048 30618 35057
rect 30562 34983 30618 34992
rect 28356 34944 28408 34950
rect 28356 34886 28408 34892
rect 28816 34944 28868 34950
rect 28816 34886 28868 34892
rect 28080 34740 28132 34746
rect 28080 34682 28132 34688
rect 26976 34536 27028 34542
rect 26976 34478 27028 34484
rect 26608 34468 26660 34474
rect 26608 34410 26660 34416
rect 26424 33992 26476 33998
rect 26424 33934 26476 33940
rect 26240 33584 26292 33590
rect 26292 33544 26372 33572
rect 26240 33526 26292 33532
rect 26240 33312 26292 33318
rect 26240 33254 26292 33260
rect 26252 33114 26280 33254
rect 26240 33108 26292 33114
rect 26240 33050 26292 33056
rect 26344 33046 26372 33544
rect 26436 33522 26464 33934
rect 26424 33516 26476 33522
rect 26424 33458 26476 33464
rect 26620 33454 26648 34410
rect 28092 34202 28120 34682
rect 28368 34406 28396 34886
rect 28356 34400 28408 34406
rect 28356 34342 28408 34348
rect 28080 34196 28132 34202
rect 28080 34138 28132 34144
rect 27620 33516 27672 33522
rect 27620 33458 27672 33464
rect 26608 33448 26660 33454
rect 26608 33390 26660 33396
rect 26884 33312 26936 33318
rect 26884 33254 26936 33260
rect 26896 33114 26924 33254
rect 27632 33114 27660 33458
rect 28092 33454 28120 34138
rect 28368 34082 28396 34342
rect 28828 34134 28856 34886
rect 31680 34649 31708 39520
rect 31666 34640 31722 34649
rect 31666 34575 31722 34584
rect 30104 34400 30156 34406
rect 30104 34342 30156 34348
rect 28816 34128 28868 34134
rect 28368 34066 28488 34082
rect 28816 34070 28868 34076
rect 28368 34060 28500 34066
rect 28368 34054 28448 34060
rect 28080 33448 28132 33454
rect 28080 33390 28132 33396
rect 28368 33318 28396 34054
rect 28448 34002 28500 34008
rect 28828 33658 28856 34070
rect 29092 33856 29144 33862
rect 29092 33798 29144 33804
rect 28816 33652 28868 33658
rect 28816 33594 28868 33600
rect 28356 33312 28408 33318
rect 28356 33254 28408 33260
rect 26884 33108 26936 33114
rect 26884 33050 26936 33056
rect 27620 33108 27672 33114
rect 27620 33050 27672 33056
rect 28172 33108 28224 33114
rect 28172 33050 28224 33056
rect 26332 33040 26384 33046
rect 26160 32966 26280 32994
rect 26332 32982 26384 32988
rect 25504 32564 25556 32570
rect 25504 32506 25556 32512
rect 25964 32564 26016 32570
rect 25964 32506 26016 32512
rect 25228 32496 25280 32502
rect 25228 32438 25280 32444
rect 26148 32428 26200 32434
rect 26148 32370 26200 32376
rect 26160 32026 26188 32370
rect 26148 32020 26200 32026
rect 26148 31962 26200 31968
rect 26252 31890 26280 32966
rect 26608 32904 26660 32910
rect 26608 32846 26660 32852
rect 26332 32768 26384 32774
rect 26332 32710 26384 32716
rect 26344 32298 26372 32710
rect 26620 32434 26648 32846
rect 26608 32428 26660 32434
rect 26608 32370 26660 32376
rect 26332 32292 26384 32298
rect 26332 32234 26384 32240
rect 26620 31958 26648 32370
rect 26896 32366 26924 33050
rect 27068 33040 27120 33046
rect 27068 32982 27120 32988
rect 27080 32570 27108 32982
rect 27068 32564 27120 32570
rect 27068 32506 27120 32512
rect 28184 32434 28212 33050
rect 28368 32910 28396 33254
rect 28632 32972 28684 32978
rect 28632 32914 28684 32920
rect 28356 32904 28408 32910
rect 28356 32846 28408 32852
rect 28172 32428 28224 32434
rect 28172 32370 28224 32376
rect 26884 32360 26936 32366
rect 27712 32360 27764 32366
rect 26884 32302 26936 32308
rect 27540 32298 27660 32314
rect 27712 32302 27764 32308
rect 27528 32292 27660 32298
rect 27580 32286 27660 32292
rect 27528 32234 27580 32240
rect 27068 32020 27120 32026
rect 27068 31962 27120 31968
rect 26608 31952 26660 31958
rect 26608 31894 26660 31900
rect 26240 31884 26292 31890
rect 26240 31826 26292 31832
rect 26252 31482 26280 31826
rect 26884 31816 26936 31822
rect 26884 31758 26936 31764
rect 26240 31476 26292 31482
rect 26240 31418 26292 31424
rect 25320 31136 25372 31142
rect 25320 31078 25372 31084
rect 26514 31104 26570 31113
rect 25332 30734 25360 31078
rect 26514 31039 26570 31048
rect 26528 30802 26556 31039
rect 26516 30796 26568 30802
rect 26516 30738 26568 30744
rect 25320 30728 25372 30734
rect 25320 30670 25372 30676
rect 25332 30190 25360 30670
rect 26528 30394 26556 30738
rect 26516 30388 26568 30394
rect 26516 30330 26568 30336
rect 25320 30184 25372 30190
rect 25320 30126 25372 30132
rect 25332 29850 25360 30126
rect 25780 30048 25832 30054
rect 25780 29990 25832 29996
rect 25792 29850 25820 29990
rect 25320 29844 25372 29850
rect 25320 29786 25372 29792
rect 25780 29844 25832 29850
rect 25780 29786 25832 29792
rect 25792 29646 25820 29786
rect 26896 29753 26924 31758
rect 27080 31482 27108 31962
rect 27632 31482 27660 32286
rect 27724 31958 27752 32302
rect 27712 31952 27764 31958
rect 27712 31894 27764 31900
rect 27068 31476 27120 31482
rect 27068 31418 27120 31424
rect 27620 31476 27672 31482
rect 27620 31418 27672 31424
rect 27080 31278 27108 31418
rect 28184 31346 28212 32370
rect 28368 31686 28396 32846
rect 28644 32570 28672 32914
rect 29000 32768 29052 32774
rect 29000 32710 29052 32716
rect 28632 32564 28684 32570
rect 28632 32506 28684 32512
rect 28644 32366 28672 32506
rect 28632 32360 28684 32366
rect 28632 32302 28684 32308
rect 28724 31884 28776 31890
rect 28724 31826 28776 31832
rect 28356 31680 28408 31686
rect 28356 31622 28408 31628
rect 28172 31340 28224 31346
rect 28172 31282 28224 31288
rect 27068 31272 27120 31278
rect 27068 31214 27120 31220
rect 28080 31136 28132 31142
rect 28080 31078 28132 31084
rect 28092 30802 28120 31078
rect 28184 30938 28212 31282
rect 28736 31142 28764 31826
rect 28816 31680 28868 31686
rect 28816 31622 28868 31628
rect 28828 31142 28856 31622
rect 28724 31136 28776 31142
rect 28724 31078 28776 31084
rect 28816 31136 28868 31142
rect 28816 31078 28868 31084
rect 28736 30938 28764 31078
rect 28172 30932 28224 30938
rect 28172 30874 28224 30880
rect 28724 30932 28776 30938
rect 28724 30874 28776 30880
rect 28828 30818 28856 31078
rect 29012 30818 29040 32710
rect 29104 32502 29132 33798
rect 30116 32609 30144 34342
rect 32784 33969 32812 39520
rect 33888 35329 33916 39520
rect 34992 37754 35020 39520
rect 35622 39400 35678 39409
rect 35622 39335 35678 39344
rect 34808 37726 35020 37754
rect 33874 35320 33930 35329
rect 33874 35255 33930 35264
rect 34808 34921 34836 37726
rect 34940 37020 35236 37040
rect 34996 37018 35020 37020
rect 35076 37018 35100 37020
rect 35156 37018 35180 37020
rect 35018 36966 35020 37018
rect 35082 36966 35094 37018
rect 35156 36966 35158 37018
rect 34996 36964 35020 36966
rect 35076 36964 35100 36966
rect 35156 36964 35180 36966
rect 34940 36944 35236 36964
rect 34940 35932 35236 35952
rect 34996 35930 35020 35932
rect 35076 35930 35100 35932
rect 35156 35930 35180 35932
rect 35018 35878 35020 35930
rect 35082 35878 35094 35930
rect 35156 35878 35158 35930
rect 34996 35876 35020 35878
rect 35076 35876 35100 35878
rect 35156 35876 35180 35878
rect 34940 35856 35236 35876
rect 35636 35834 35664 39335
rect 35806 36952 35862 36961
rect 35806 36887 35862 36896
rect 35624 35828 35676 35834
rect 35624 35770 35676 35776
rect 35624 35624 35676 35630
rect 35624 35566 35676 35572
rect 35530 35320 35586 35329
rect 35530 35255 35532 35264
rect 35584 35255 35586 35264
rect 35532 35226 35584 35232
rect 35636 35170 35664 35566
rect 35714 35456 35770 35465
rect 35714 35391 35770 35400
rect 35348 35148 35400 35154
rect 35348 35090 35400 35096
rect 35544 35142 35664 35170
rect 34794 34912 34850 34921
rect 34794 34847 34850 34856
rect 34940 34844 35236 34864
rect 34996 34842 35020 34844
rect 35076 34842 35100 34844
rect 35156 34842 35180 34844
rect 35018 34790 35020 34842
rect 35082 34790 35094 34842
rect 35156 34790 35158 34842
rect 34996 34788 35020 34790
rect 35076 34788 35100 34790
rect 35156 34788 35180 34790
rect 34940 34768 35236 34788
rect 35256 34536 35308 34542
rect 35256 34478 35308 34484
rect 32770 33960 32826 33969
rect 32770 33895 32826 33904
rect 34940 33756 35236 33776
rect 34996 33754 35020 33756
rect 35076 33754 35100 33756
rect 35156 33754 35180 33756
rect 35018 33702 35020 33754
rect 35082 33702 35094 33754
rect 35156 33702 35158 33754
rect 34996 33700 35020 33702
rect 35076 33700 35100 33702
rect 35156 33700 35180 33702
rect 34940 33680 35236 33700
rect 34940 32668 35236 32688
rect 34996 32666 35020 32668
rect 35076 32666 35100 32668
rect 35156 32666 35180 32668
rect 35018 32614 35020 32666
rect 35082 32614 35094 32666
rect 35156 32614 35158 32666
rect 34996 32612 35020 32614
rect 35076 32612 35100 32614
rect 35156 32612 35180 32614
rect 30102 32600 30158 32609
rect 34940 32592 35236 32612
rect 30102 32535 30158 32544
rect 29092 32496 29144 32502
rect 29092 32438 29144 32444
rect 29276 32360 29328 32366
rect 29276 32302 29328 32308
rect 29288 31686 29316 32302
rect 29276 31680 29328 31686
rect 29276 31622 29328 31628
rect 28080 30796 28132 30802
rect 28080 30738 28132 30744
rect 28736 30790 28856 30818
rect 28920 30802 29040 30818
rect 28908 30796 29040 30802
rect 28092 30394 28120 30738
rect 28736 30598 28764 30790
rect 28960 30790 29040 30796
rect 28908 30738 28960 30744
rect 28724 30592 28776 30598
rect 28724 30534 28776 30540
rect 28080 30388 28132 30394
rect 28080 30330 28132 30336
rect 28736 30054 28764 30534
rect 28724 30048 28776 30054
rect 28724 29990 28776 29996
rect 26882 29744 26938 29753
rect 26882 29679 26938 29688
rect 27712 29708 27764 29714
rect 27712 29650 27764 29656
rect 25320 29640 25372 29646
rect 25320 29582 25372 29588
rect 25780 29640 25832 29646
rect 25780 29582 25832 29588
rect 26148 29640 26200 29646
rect 26148 29582 26200 29588
rect 25332 29034 25360 29582
rect 25320 29028 25372 29034
rect 25320 28970 25372 28976
rect 26160 28762 26188 29582
rect 26516 29504 26568 29510
rect 26516 29446 26568 29452
rect 26424 28960 26476 28966
rect 26424 28902 26476 28908
rect 25136 28756 25188 28762
rect 25136 28698 25188 28704
rect 25688 28756 25740 28762
rect 25688 28698 25740 28704
rect 26148 28756 26200 28762
rect 26148 28698 26200 28704
rect 25504 28552 25556 28558
rect 25504 28494 25556 28500
rect 25044 28416 25096 28422
rect 25044 28358 25096 28364
rect 25516 28082 25544 28494
rect 25700 28218 25728 28698
rect 26436 28694 26464 28902
rect 26424 28688 26476 28694
rect 26424 28630 26476 28636
rect 26148 28416 26200 28422
rect 26148 28358 26200 28364
rect 25688 28212 25740 28218
rect 25688 28154 25740 28160
rect 25504 28076 25556 28082
rect 25504 28018 25556 28024
rect 26160 28014 26188 28358
rect 26436 28218 26464 28630
rect 26528 28558 26556 29446
rect 27724 29306 27752 29650
rect 28736 29510 28764 29990
rect 28724 29504 28776 29510
rect 28724 29446 28776 29452
rect 27712 29300 27764 29306
rect 27712 29242 27764 29248
rect 26516 28552 26568 28558
rect 26516 28494 26568 28500
rect 26424 28212 26476 28218
rect 26424 28154 26476 28160
rect 26148 28008 26200 28014
rect 26148 27950 26200 27956
rect 26160 27674 26188 27950
rect 26332 27940 26384 27946
rect 26332 27882 26384 27888
rect 26344 27690 26372 27882
rect 27252 27872 27304 27878
rect 27252 27814 27304 27820
rect 26974 27704 27030 27713
rect 26148 27668 26200 27674
rect 26344 27662 26464 27690
rect 26148 27610 26200 27616
rect 25136 27532 25188 27538
rect 25136 27474 25188 27480
rect 25412 27532 25464 27538
rect 25412 27474 25464 27480
rect 26148 27532 26200 27538
rect 26200 27492 26372 27520
rect 26148 27474 26200 27480
rect 24952 27396 25004 27402
rect 24952 27338 25004 27344
rect 24584 27328 24636 27334
rect 24584 27270 24636 27276
rect 21732 26988 21784 26994
rect 21732 26930 21784 26936
rect 22284 26988 22336 26994
rect 22284 26930 22336 26936
rect 21916 26852 21968 26858
rect 21916 26794 21968 26800
rect 21928 26042 21956 26794
rect 22296 26790 22324 26930
rect 22284 26784 22336 26790
rect 22284 26726 22336 26732
rect 22296 26586 22324 26726
rect 22284 26580 22336 26586
rect 22284 26522 22336 26528
rect 22008 26444 22060 26450
rect 22008 26386 22060 26392
rect 22020 26330 22048 26386
rect 24596 26382 24624 27270
rect 25148 26994 25176 27474
rect 25228 27328 25280 27334
rect 25228 27270 25280 27276
rect 25136 26988 25188 26994
rect 25136 26930 25188 26936
rect 25240 26926 25268 27270
rect 25424 27130 25452 27474
rect 25504 27464 25556 27470
rect 25502 27432 25504 27441
rect 25556 27432 25558 27441
rect 25502 27367 25558 27376
rect 25412 27124 25464 27130
rect 25412 27066 25464 27072
rect 25228 26920 25280 26926
rect 25228 26862 25280 26868
rect 24952 26444 25004 26450
rect 24952 26386 25004 26392
rect 24124 26376 24176 26382
rect 22020 26302 22140 26330
rect 24124 26318 24176 26324
rect 24584 26376 24636 26382
rect 24584 26318 24636 26324
rect 21916 26036 21968 26042
rect 21916 25978 21968 25984
rect 22006 25800 22062 25809
rect 22006 25735 22062 25744
rect 21546 23896 21602 23905
rect 22020 23866 22048 25735
rect 22112 25498 22140 26302
rect 22928 26240 22980 26246
rect 22928 26182 22980 26188
rect 22940 26042 22968 26182
rect 22928 26036 22980 26042
rect 22928 25978 22980 25984
rect 23480 25832 23532 25838
rect 23478 25800 23480 25809
rect 23532 25800 23534 25809
rect 23478 25735 23534 25744
rect 24136 25498 24164 26318
rect 24584 26240 24636 26246
rect 24398 26208 24454 26217
rect 24584 26182 24636 26188
rect 24398 26143 24454 26152
rect 24308 25968 24360 25974
rect 24308 25910 24360 25916
rect 24320 25498 24348 25910
rect 24412 25838 24440 26143
rect 24596 25906 24624 26182
rect 24584 25900 24636 25906
rect 24584 25842 24636 25848
rect 24400 25832 24452 25838
rect 24400 25774 24452 25780
rect 24596 25498 24624 25842
rect 24964 25838 24992 26386
rect 25044 26240 25096 26246
rect 25044 26182 25096 26188
rect 24952 25832 25004 25838
rect 24952 25774 25004 25780
rect 22100 25492 22152 25498
rect 22100 25434 22152 25440
rect 24124 25492 24176 25498
rect 24124 25434 24176 25440
rect 24308 25492 24360 25498
rect 24308 25434 24360 25440
rect 24584 25492 24636 25498
rect 24584 25434 24636 25440
rect 24768 25356 24820 25362
rect 24768 25298 24820 25304
rect 24780 24818 24808 25298
rect 25056 25294 25084 26182
rect 25240 25498 25268 26862
rect 25516 26858 25544 27367
rect 25504 26852 25556 26858
rect 25504 26794 25556 26800
rect 25320 26784 25372 26790
rect 25320 26726 25372 26732
rect 25332 26518 25360 26726
rect 25516 26586 25544 26794
rect 25504 26580 25556 26586
rect 25504 26522 25556 26528
rect 25320 26512 25372 26518
rect 25320 26454 25372 26460
rect 25332 26382 25360 26454
rect 25320 26376 25372 26382
rect 25320 26318 25372 26324
rect 25228 25492 25280 25498
rect 25148 25452 25228 25480
rect 25044 25288 25096 25294
rect 25044 25230 25096 25236
rect 24860 25220 24912 25226
rect 24860 25162 24912 25168
rect 24768 24812 24820 24818
rect 24768 24754 24820 24760
rect 22376 24608 22428 24614
rect 22376 24550 22428 24556
rect 22388 24274 22416 24550
rect 24780 24410 24808 24754
rect 24872 24750 24900 25162
rect 25056 24886 25084 25230
rect 25044 24880 25096 24886
rect 25044 24822 25096 24828
rect 25148 24750 25176 25452
rect 25228 25434 25280 25440
rect 25332 24750 25360 26318
rect 26240 26308 26292 26314
rect 26240 26250 26292 26256
rect 26252 26217 26280 26250
rect 26238 26208 26294 26217
rect 26238 26143 26294 26152
rect 26344 26042 26372 27492
rect 26436 26450 26464 27662
rect 26974 27639 27030 27648
rect 26516 27464 26568 27470
rect 26516 27406 26568 27412
rect 26528 27062 26556 27406
rect 26516 27056 26568 27062
rect 26516 26998 26568 27004
rect 26424 26444 26476 26450
rect 26424 26386 26476 26392
rect 26332 26036 26384 26042
rect 26332 25978 26384 25984
rect 26436 25974 26464 26386
rect 26988 26382 27016 27639
rect 27264 27538 27292 27814
rect 27252 27532 27304 27538
rect 27252 27474 27304 27480
rect 27264 26790 27292 27474
rect 27252 26784 27304 26790
rect 27252 26726 27304 26732
rect 26700 26376 26752 26382
rect 26620 26324 26700 26330
rect 26620 26318 26752 26324
rect 26976 26376 27028 26382
rect 26976 26318 27028 26324
rect 26620 26302 26740 26318
rect 26424 25968 26476 25974
rect 26424 25910 26476 25916
rect 26620 25702 26648 26302
rect 26988 25820 27016 26318
rect 27264 25906 27292 26726
rect 27724 26024 27752 29242
rect 27896 28416 27948 28422
rect 30012 28416 30064 28422
rect 27896 28358 27948 28364
rect 30010 28384 30012 28393
rect 30064 28384 30066 28393
rect 27908 28014 27936 28358
rect 30010 28319 30066 28328
rect 30024 28082 30052 28319
rect 30012 28076 30064 28082
rect 30012 28018 30064 28024
rect 27896 28008 27948 28014
rect 27896 27950 27948 27956
rect 30024 27674 30052 28018
rect 29828 27668 29880 27674
rect 29828 27610 29880 27616
rect 30012 27668 30064 27674
rect 30012 27610 30064 27616
rect 29092 27532 29144 27538
rect 29092 27474 29144 27480
rect 27894 27432 27950 27441
rect 27894 27367 27896 27376
rect 27948 27367 27950 27376
rect 27896 27338 27948 27344
rect 29104 27130 29132 27474
rect 29552 27464 29604 27470
rect 29552 27406 29604 27412
rect 29092 27124 29144 27130
rect 29092 27066 29144 27072
rect 29564 27062 29592 27406
rect 29552 27056 29604 27062
rect 29552 26998 29604 27004
rect 29182 26616 29238 26625
rect 29564 26586 29592 26998
rect 29840 26994 29868 27610
rect 29828 26988 29880 26994
rect 29828 26930 29880 26936
rect 29736 26852 29788 26858
rect 29736 26794 29788 26800
rect 29182 26551 29238 26560
rect 29368 26580 29420 26586
rect 29196 26450 29224 26551
rect 29368 26522 29420 26528
rect 29552 26580 29604 26586
rect 29552 26522 29604 26528
rect 29380 26489 29408 26522
rect 29366 26480 29422 26489
rect 28908 26444 28960 26450
rect 28908 26386 28960 26392
rect 29184 26444 29236 26450
rect 29366 26415 29422 26424
rect 29184 26386 29236 26392
rect 28264 26308 28316 26314
rect 28264 26250 28316 26256
rect 27540 25996 27752 26024
rect 27252 25900 27304 25906
rect 27252 25842 27304 25848
rect 27068 25832 27120 25838
rect 26988 25792 27068 25820
rect 26608 25696 26660 25702
rect 26608 25638 26660 25644
rect 26620 25537 26648 25638
rect 26606 25528 26662 25537
rect 26988 25498 27016 25792
rect 27068 25774 27120 25780
rect 27540 25498 27568 25996
rect 27712 25900 27764 25906
rect 27712 25842 27764 25848
rect 27724 25498 27752 25842
rect 28276 25770 28304 26250
rect 28920 26042 28948 26386
rect 28908 26036 28960 26042
rect 28908 25978 28960 25984
rect 29184 25832 29236 25838
rect 29184 25774 29236 25780
rect 28264 25764 28316 25770
rect 28264 25706 28316 25712
rect 26606 25463 26662 25472
rect 26976 25492 27028 25498
rect 26976 25434 27028 25440
rect 27528 25492 27580 25498
rect 27528 25434 27580 25440
rect 27712 25492 27764 25498
rect 27712 25434 27764 25440
rect 26240 25356 26292 25362
rect 26240 25298 26292 25304
rect 27344 25356 27396 25362
rect 27344 25298 27396 25304
rect 26148 25288 26200 25294
rect 26148 25230 26200 25236
rect 24860 24744 24912 24750
rect 24860 24686 24912 24692
rect 25136 24744 25188 24750
rect 25136 24686 25188 24692
rect 25320 24744 25372 24750
rect 25320 24686 25372 24692
rect 25148 24410 25176 24686
rect 24768 24404 24820 24410
rect 24768 24346 24820 24352
rect 25136 24404 25188 24410
rect 25136 24346 25188 24352
rect 22376 24268 22428 24274
rect 22376 24210 22428 24216
rect 21546 23831 21602 23840
rect 22008 23860 22060 23866
rect 22008 23802 22060 23808
rect 21086 23624 21142 23633
rect 21086 23559 21142 23568
rect 21548 23588 21600 23594
rect 21100 23322 21128 23559
rect 21548 23530 21600 23536
rect 20260 23316 20312 23322
rect 20260 23258 20312 23264
rect 21088 23316 21140 23322
rect 21088 23258 21140 23264
rect 21560 22982 21588 23530
rect 25148 23322 25176 24346
rect 25332 24342 25360 24686
rect 26160 24614 26188 25230
rect 26148 24608 26200 24614
rect 26148 24550 26200 24556
rect 26252 24410 26280 25298
rect 27356 24954 27384 25298
rect 27344 24948 27396 24954
rect 27344 24890 27396 24896
rect 26424 24608 26476 24614
rect 26424 24550 26476 24556
rect 26240 24404 26292 24410
rect 26240 24346 26292 24352
rect 25320 24336 25372 24342
rect 25320 24278 25372 24284
rect 25136 23316 25188 23322
rect 25136 23258 25188 23264
rect 21548 22976 21600 22982
rect 21548 22918 21600 22924
rect 21560 22137 21588 22918
rect 25148 22642 25176 23258
rect 26148 22976 26200 22982
rect 26148 22918 26200 22924
rect 25136 22636 25188 22642
rect 25136 22578 25188 22584
rect 22376 22432 22428 22438
rect 22376 22374 22428 22380
rect 21546 22128 21602 22137
rect 21546 22063 21602 22072
rect 22284 22092 22336 22098
rect 22284 22034 22336 22040
rect 22296 21894 22324 22034
rect 22388 22030 22416 22374
rect 23112 22092 23164 22098
rect 23112 22034 23164 22040
rect 24032 22092 24084 22098
rect 24032 22034 24084 22040
rect 22376 22024 22428 22030
rect 22376 21966 22428 21972
rect 23020 22024 23072 22030
rect 23020 21966 23072 21972
rect 21088 21888 21140 21894
rect 21088 21830 21140 21836
rect 22284 21888 22336 21894
rect 22284 21830 22336 21836
rect 21100 21486 21128 21830
rect 22296 21690 22324 21830
rect 22284 21684 22336 21690
rect 22284 21626 22336 21632
rect 21088 21480 21140 21486
rect 21088 21422 21140 21428
rect 21100 21146 21128 21422
rect 21088 21140 21140 21146
rect 21088 21082 21140 21088
rect 21730 21040 21786 21049
rect 21730 20975 21732 20984
rect 21784 20975 21786 20984
rect 22008 21004 22060 21010
rect 21732 20946 21784 20952
rect 22008 20946 22060 20952
rect 20536 20800 20588 20806
rect 20536 20742 20588 20748
rect 20168 19236 20220 19242
rect 20168 19178 20220 19184
rect 20076 18760 20128 18766
rect 20076 18702 20128 18708
rect 19984 18352 20036 18358
rect 19984 18294 20036 18300
rect 20180 18086 20208 19178
rect 20548 18970 20576 20742
rect 21456 20256 21508 20262
rect 21456 20198 21508 20204
rect 21468 19922 21496 20198
rect 21744 20058 21772 20946
rect 22020 20618 22048 20946
rect 23032 20806 23060 21966
rect 23124 21350 23152 22034
rect 23480 21888 23532 21894
rect 23480 21830 23532 21836
rect 23664 21888 23716 21894
rect 23664 21830 23716 21836
rect 23112 21344 23164 21350
rect 23112 21286 23164 21292
rect 23124 21146 23152 21286
rect 23112 21140 23164 21146
rect 23112 21082 23164 21088
rect 23020 20800 23072 20806
rect 23020 20742 23072 20748
rect 23032 20641 23060 20742
rect 23018 20632 23074 20641
rect 22020 20590 22140 20618
rect 22112 20398 22140 20590
rect 23018 20567 23074 20576
rect 23032 20466 23060 20567
rect 23388 20528 23440 20534
rect 23388 20470 23440 20476
rect 23020 20460 23072 20466
rect 23020 20402 23072 20408
rect 22100 20392 22152 20398
rect 22100 20334 22152 20340
rect 22112 20262 22140 20334
rect 21916 20256 21968 20262
rect 21916 20198 21968 20204
rect 22100 20256 22152 20262
rect 22100 20198 22152 20204
rect 21732 20052 21784 20058
rect 21732 19994 21784 20000
rect 21456 19916 21508 19922
rect 21456 19858 21508 19864
rect 20628 19304 20680 19310
rect 20628 19246 20680 19252
rect 20536 18964 20588 18970
rect 20536 18906 20588 18912
rect 20260 18760 20312 18766
rect 20260 18702 20312 18708
rect 20168 18080 20220 18086
rect 20168 18022 20220 18028
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 20180 17882 20208 18022
rect 20168 17876 20220 17882
rect 20168 17818 20220 17824
rect 19616 17808 19668 17814
rect 19616 17750 19668 17756
rect 18970 17640 19026 17649
rect 18970 17575 19026 17584
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 16670 7576 16726 7585
rect 16670 7511 16726 7520
rect 570 6760 626 6769
rect 570 6695 626 6704
rect 584 5681 612 6695
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 570 5672 626 5681
rect 570 5607 626 5616
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 3330 3496 3386 3505
rect 3330 3431 3386 3440
rect 3344 480 3372 3431
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 9956 2304 10008 2310
rect 9956 2246 10008 2252
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 9968 480 9996 2246
rect 16684 480 16712 7511
rect 18432 5681 18460 17478
rect 18984 17338 19012 17575
rect 18972 17332 19024 17338
rect 18972 17274 19024 17280
rect 19628 17202 19656 17750
rect 20272 17377 20300 18702
rect 20548 18358 20576 18906
rect 20536 18352 20588 18358
rect 20536 18294 20588 18300
rect 20640 18306 20668 19246
rect 21468 19174 21496 19858
rect 21744 19310 21772 19994
rect 21928 19394 21956 20198
rect 22112 20058 22140 20198
rect 23400 20058 23428 20470
rect 23492 20466 23520 21830
rect 23676 21486 23704 21830
rect 23664 21480 23716 21486
rect 23664 21422 23716 21428
rect 23676 21049 23704 21422
rect 24044 21350 24072 22034
rect 25148 21894 25176 22578
rect 25320 22500 25372 22506
rect 25320 22442 25372 22448
rect 25332 21894 25360 22442
rect 25502 22128 25558 22137
rect 25502 22063 25558 22072
rect 25136 21888 25188 21894
rect 25136 21830 25188 21836
rect 25320 21888 25372 21894
rect 25320 21830 25372 21836
rect 25148 21418 25176 21830
rect 25136 21412 25188 21418
rect 25136 21354 25188 21360
rect 24032 21344 24084 21350
rect 24032 21286 24084 21292
rect 24952 21344 25004 21350
rect 24952 21286 25004 21292
rect 24044 21146 24072 21286
rect 24032 21140 24084 21146
rect 24032 21082 24084 21088
rect 23662 21040 23718 21049
rect 23662 20975 23718 20984
rect 24216 21004 24268 21010
rect 24216 20946 24268 20952
rect 23480 20460 23532 20466
rect 23480 20402 23532 20408
rect 23492 20058 23520 20402
rect 23664 20256 23716 20262
rect 23664 20198 23716 20204
rect 22100 20052 22152 20058
rect 22100 19994 22152 20000
rect 23388 20052 23440 20058
rect 23388 19994 23440 20000
rect 23480 20052 23532 20058
rect 23480 19994 23532 20000
rect 21928 19366 22140 19394
rect 21732 19304 21784 19310
rect 21732 19246 21784 19252
rect 21456 19168 21508 19174
rect 21456 19110 21508 19116
rect 21468 18970 21496 19110
rect 21456 18964 21508 18970
rect 21456 18906 21508 18912
rect 22112 18902 22140 19366
rect 22100 18896 22152 18902
rect 22100 18838 22152 18844
rect 23676 18834 23704 20198
rect 23848 19848 23900 19854
rect 23848 19790 23900 19796
rect 23860 19281 23888 19790
rect 24228 19718 24256 20946
rect 24492 20528 24544 20534
rect 24492 20470 24544 20476
rect 24216 19712 24268 19718
rect 24216 19654 24268 19660
rect 23846 19272 23902 19281
rect 23846 19207 23902 19216
rect 24124 19168 24176 19174
rect 24124 19110 24176 19116
rect 24136 18873 24164 19110
rect 24122 18864 24178 18873
rect 22928 18828 22980 18834
rect 22928 18770 22980 18776
rect 23664 18828 23716 18834
rect 24122 18799 24178 18808
rect 23664 18770 23716 18776
rect 22376 18760 22428 18766
rect 22376 18702 22428 18708
rect 22388 18426 22416 18702
rect 22940 18426 22968 18770
rect 23388 18624 23440 18630
rect 23388 18566 23440 18572
rect 22376 18420 22428 18426
rect 22376 18362 22428 18368
rect 22928 18420 22980 18426
rect 22928 18362 22980 18368
rect 20548 17814 20576 18294
rect 20640 18290 20852 18306
rect 20628 18284 20852 18290
rect 20680 18278 20852 18284
rect 20628 18226 20680 18232
rect 20720 18148 20772 18154
rect 20720 18090 20772 18096
rect 20536 17808 20588 17814
rect 20536 17750 20588 17756
rect 20732 17542 20760 18090
rect 20824 17882 20852 18278
rect 20812 17876 20864 17882
rect 20812 17818 20864 17824
rect 23400 17746 23428 18566
rect 23676 18426 23704 18770
rect 23664 18420 23716 18426
rect 23664 18362 23716 18368
rect 23848 18352 23900 18358
rect 23848 18294 23900 18300
rect 22192 17740 22244 17746
rect 22192 17682 22244 17688
rect 22468 17740 22520 17746
rect 22468 17682 22520 17688
rect 23388 17740 23440 17746
rect 23388 17682 23440 17688
rect 22204 17649 22232 17682
rect 22190 17640 22246 17649
rect 22190 17575 22246 17584
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 21824 17536 21876 17542
rect 21824 17478 21876 17484
rect 20258 17368 20314 17377
rect 20732 17338 20760 17478
rect 20258 17303 20314 17312
rect 20720 17332 20772 17338
rect 20720 17274 20772 17280
rect 21836 17241 21864 17478
rect 22204 17338 22232 17575
rect 22192 17332 22244 17338
rect 22192 17274 22244 17280
rect 21822 17232 21878 17241
rect 19616 17196 19668 17202
rect 19616 17138 19668 17144
rect 19892 17196 19944 17202
rect 21822 17167 21878 17176
rect 19892 17138 19944 17144
rect 19246 17096 19302 17105
rect 19064 17060 19116 17066
rect 19246 17031 19302 17040
rect 19064 17002 19116 17008
rect 19076 16794 19104 17002
rect 19260 16794 19288 17031
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 19064 16788 19116 16794
rect 19064 16730 19116 16736
rect 19248 16788 19300 16794
rect 19248 16730 19300 16736
rect 19616 16652 19668 16658
rect 19616 16594 19668 16600
rect 19628 15978 19656 16594
rect 19904 16590 19932 17138
rect 22480 17134 22508 17682
rect 23400 17338 23428 17682
rect 23860 17338 23888 18294
rect 23388 17332 23440 17338
rect 23388 17274 23440 17280
rect 23848 17332 23900 17338
rect 23848 17274 23900 17280
rect 23662 17232 23718 17241
rect 23662 17167 23718 17176
rect 23676 17134 23704 17167
rect 20628 17128 20680 17134
rect 22468 17128 22520 17134
rect 22466 17096 22468 17105
rect 23664 17128 23716 17134
rect 22520 17096 22522 17105
rect 20680 17076 20760 17082
rect 20628 17070 20760 17076
rect 20640 17054 20760 17070
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 20180 16726 20208 16934
rect 20168 16720 20220 16726
rect 20168 16662 20220 16668
rect 19708 16584 19760 16590
rect 19708 16526 19760 16532
rect 19892 16584 19944 16590
rect 19892 16526 19944 16532
rect 19720 16114 19748 16526
rect 19904 16250 19932 16526
rect 20180 16250 20208 16662
rect 20732 16658 20760 17054
rect 22284 17060 22336 17066
rect 23664 17070 23716 17076
rect 22466 17031 22522 17040
rect 22284 17002 22336 17008
rect 22296 16794 22324 17002
rect 23676 16794 23704 17070
rect 24124 17060 24176 17066
rect 24124 17002 24176 17008
rect 22284 16788 22336 16794
rect 22284 16730 22336 16736
rect 23664 16788 23716 16794
rect 23664 16730 23716 16736
rect 24136 16726 24164 17002
rect 22100 16720 22152 16726
rect 22100 16662 22152 16668
rect 24124 16720 24176 16726
rect 24124 16662 24176 16668
rect 20720 16652 20772 16658
rect 20720 16594 20772 16600
rect 19892 16244 19944 16250
rect 19892 16186 19944 16192
rect 20168 16244 20220 16250
rect 20168 16186 20220 16192
rect 19708 16108 19760 16114
rect 19708 16050 19760 16056
rect 20628 16108 20680 16114
rect 20628 16050 20680 16056
rect 19616 15972 19668 15978
rect 19616 15914 19668 15920
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19580 15728 19876 15748
rect 20640 15570 20668 16050
rect 20732 16046 20760 16594
rect 22112 16250 22140 16662
rect 24136 16250 24164 16662
rect 22100 16244 22152 16250
rect 22100 16186 22152 16192
rect 24124 16244 24176 16250
rect 24124 16186 24176 16192
rect 20720 16040 20772 16046
rect 20720 15982 20772 15988
rect 20628 15564 20680 15570
rect 20628 15506 20680 15512
rect 20640 15162 20668 15506
rect 20732 15502 20760 15982
rect 22284 15972 22336 15978
rect 22284 15914 22336 15920
rect 22296 15706 22324 15914
rect 22284 15700 22336 15706
rect 22284 15642 22336 15648
rect 22008 15564 22060 15570
rect 22008 15506 22060 15512
rect 20720 15496 20772 15502
rect 20720 15438 20772 15444
rect 20904 15496 20956 15502
rect 20904 15438 20956 15444
rect 22020 15450 22048 15506
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20916 14958 20944 15438
rect 22020 15422 22140 15450
rect 21362 15192 21418 15201
rect 22112 15162 22140 15422
rect 21362 15127 21418 15136
rect 22100 15156 22152 15162
rect 21376 14958 21404 15127
rect 22100 15098 22152 15104
rect 20904 14952 20956 14958
rect 20904 14894 20956 14900
rect 21364 14952 21416 14958
rect 21364 14894 21416 14900
rect 21180 14884 21232 14890
rect 21180 14826 21232 14832
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19580 14640 19876 14660
rect 21192 14278 21220 14826
rect 23848 14476 23900 14482
rect 23848 14418 23900 14424
rect 23112 14340 23164 14346
rect 23112 14282 23164 14288
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 21192 12782 21220 14214
rect 23124 14074 23152 14282
rect 23860 14074 23888 14418
rect 23940 14408 23992 14414
rect 23940 14350 23992 14356
rect 23112 14068 23164 14074
rect 23112 14010 23164 14016
rect 23848 14068 23900 14074
rect 23848 14010 23900 14016
rect 23020 13728 23072 13734
rect 23020 13670 23072 13676
rect 22836 13320 22888 13326
rect 22836 13262 22888 13268
rect 22376 13184 22428 13190
rect 22376 13126 22428 13132
rect 22388 12850 22416 13126
rect 22376 12844 22428 12850
rect 22376 12786 22428 12792
rect 21180 12776 21232 12782
rect 21180 12718 21232 12724
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19580 12464 19876 12484
rect 21192 12238 21220 12718
rect 22848 12714 22876 13262
rect 23032 12986 23060 13670
rect 23124 13326 23152 14010
rect 23664 13864 23716 13870
rect 23716 13812 23796 13818
rect 23664 13806 23796 13812
rect 23676 13790 23796 13806
rect 23768 13512 23796 13790
rect 23860 13530 23888 14010
rect 23952 13870 23980 14350
rect 24032 14272 24084 14278
rect 24032 14214 24084 14220
rect 23940 13864 23992 13870
rect 23940 13806 23992 13812
rect 23584 13484 23796 13512
rect 23112 13320 23164 13326
rect 23112 13262 23164 13268
rect 23020 12980 23072 12986
rect 23020 12922 23072 12928
rect 22376 12708 22428 12714
rect 22376 12650 22428 12656
rect 22836 12708 22888 12714
rect 22836 12650 22888 12656
rect 22388 12374 22416 12650
rect 22376 12368 22428 12374
rect 22376 12310 22428 12316
rect 21180 12232 21232 12238
rect 21180 12174 21232 12180
rect 22284 12232 22336 12238
rect 22284 12174 22336 12180
rect 22296 11830 22324 12174
rect 22284 11824 22336 11830
rect 22284 11766 22336 11772
rect 22388 11558 22416 12310
rect 23388 11824 23440 11830
rect 23584 11778 23612 13484
rect 23768 13394 23796 13484
rect 23848 13524 23900 13530
rect 23848 13466 23900 13472
rect 23664 13388 23716 13394
rect 23664 13330 23716 13336
rect 23756 13388 23808 13394
rect 23756 13330 23808 13336
rect 23676 12646 23704 13330
rect 24044 12782 24072 14214
rect 24124 12844 24176 12850
rect 24124 12786 24176 12792
rect 24032 12776 24084 12782
rect 24032 12718 24084 12724
rect 23664 12640 23716 12646
rect 23664 12582 23716 12588
rect 23676 12442 23704 12582
rect 24136 12442 24164 12786
rect 23664 12436 23716 12442
rect 23664 12378 23716 12384
rect 24124 12436 24176 12442
rect 24124 12378 24176 12384
rect 23440 11772 23612 11778
rect 23388 11766 23612 11772
rect 23400 11750 23612 11766
rect 23664 11756 23716 11762
rect 23664 11698 23716 11704
rect 22560 11688 22612 11694
rect 22560 11630 22612 11636
rect 22376 11552 22428 11558
rect 22376 11494 22428 11500
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 22388 11354 22416 11494
rect 22376 11348 22428 11354
rect 22376 11290 22428 11296
rect 22468 11212 22520 11218
rect 22468 11154 22520 11160
rect 22284 10600 22336 10606
rect 22284 10542 22336 10548
rect 22296 10470 22324 10542
rect 22284 10464 22336 10470
rect 22284 10406 22336 10412
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 22480 9926 22508 11154
rect 22572 11014 22600 11630
rect 23480 11620 23532 11626
rect 23480 11562 23532 11568
rect 22652 11212 22704 11218
rect 22652 11154 22704 11160
rect 22560 11008 22612 11014
rect 22560 10950 22612 10956
rect 22572 10674 22600 10950
rect 22560 10668 22612 10674
rect 22560 10610 22612 10616
rect 22664 10606 22692 11154
rect 22652 10600 22704 10606
rect 22652 10542 22704 10548
rect 23112 10600 23164 10606
rect 23112 10542 23164 10548
rect 23124 10470 23152 10542
rect 22928 10464 22980 10470
rect 23112 10464 23164 10470
rect 22980 10412 23060 10418
rect 22928 10406 23060 10412
rect 23112 10406 23164 10412
rect 22940 10390 23060 10406
rect 23032 10130 23060 10390
rect 23124 10266 23152 10406
rect 23112 10260 23164 10266
rect 23112 10202 23164 10208
rect 23020 10124 23072 10130
rect 23020 10066 23072 10072
rect 22468 9920 22520 9926
rect 22468 9862 22520 9868
rect 22480 9450 22508 9862
rect 23032 9722 23060 10066
rect 23020 9716 23072 9722
rect 23020 9658 23072 9664
rect 23492 9654 23520 11562
rect 23676 10690 23704 11698
rect 23756 11552 23808 11558
rect 23756 11494 23808 11500
rect 23768 10810 23796 11494
rect 23756 10804 23808 10810
rect 23756 10746 23808 10752
rect 23676 10662 23796 10690
rect 23480 9648 23532 9654
rect 23480 9590 23532 9596
rect 22468 9444 22520 9450
rect 22468 9386 22520 9392
rect 23480 9444 23532 9450
rect 23480 9386 23532 9392
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 23492 9042 23520 9386
rect 23768 9042 23796 10662
rect 23480 9036 23532 9042
rect 23480 8978 23532 8984
rect 23756 9036 23808 9042
rect 23756 8978 23808 8984
rect 23768 8634 23796 8978
rect 23756 8628 23808 8634
rect 23756 8570 23808 8576
rect 24124 8424 24176 8430
rect 24124 8366 24176 8372
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 24136 8090 24164 8366
rect 24124 8084 24176 8090
rect 24124 8026 24176 8032
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19580 7024 19876 7044
rect 19580 6012 19876 6032
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 18418 5672 18474 5681
rect 18418 5607 18474 5616
rect 19580 4924 19876 4944
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 24228 4049 24256 19654
rect 24308 19168 24360 19174
rect 24308 19110 24360 19116
rect 24320 17882 24348 19110
rect 24504 18766 24532 20470
rect 24964 20466 24992 21286
rect 25134 20632 25190 20641
rect 25134 20567 25190 20576
rect 25148 20466 25176 20567
rect 24952 20460 25004 20466
rect 24952 20402 25004 20408
rect 25136 20460 25188 20466
rect 25136 20402 25188 20408
rect 24964 20058 24992 20402
rect 25332 20398 25360 21830
rect 25516 21146 25544 22063
rect 26160 21690 26188 22918
rect 26148 21684 26200 21690
rect 26148 21626 26200 21632
rect 26160 21486 26188 21626
rect 26332 21616 26384 21622
rect 26332 21558 26384 21564
rect 26148 21480 26200 21486
rect 26148 21422 26200 21428
rect 26240 21344 26292 21350
rect 26240 21286 26292 21292
rect 25504 21140 25556 21146
rect 25556 21100 25636 21128
rect 25504 21082 25556 21088
rect 25320 20392 25372 20398
rect 25320 20334 25372 20340
rect 25410 20360 25466 20369
rect 25410 20295 25466 20304
rect 25424 20058 25452 20295
rect 24952 20052 25004 20058
rect 24952 19994 25004 20000
rect 25412 20052 25464 20058
rect 25412 19994 25464 20000
rect 25320 19916 25372 19922
rect 25320 19858 25372 19864
rect 24768 19780 24820 19786
rect 24768 19722 24820 19728
rect 24780 19310 24808 19722
rect 24860 19508 24912 19514
rect 24860 19450 24912 19456
rect 24768 19304 24820 19310
rect 24768 19246 24820 19252
rect 24584 19168 24636 19174
rect 24584 19110 24636 19116
rect 24676 19168 24728 19174
rect 24676 19110 24728 19116
rect 24596 18873 24624 19110
rect 24688 18970 24716 19110
rect 24872 18970 24900 19450
rect 24676 18964 24728 18970
rect 24676 18906 24728 18912
rect 24860 18964 24912 18970
rect 24860 18906 24912 18912
rect 25332 18873 25360 19858
rect 25424 19514 25452 19994
rect 25412 19508 25464 19514
rect 25412 19450 25464 19456
rect 25412 19372 25464 19378
rect 25412 19314 25464 19320
rect 24582 18864 24638 18873
rect 25318 18864 25374 18873
rect 24582 18799 24638 18808
rect 25228 18828 25280 18834
rect 25318 18799 25374 18808
rect 25228 18770 25280 18776
rect 24492 18760 24544 18766
rect 24398 18728 24454 18737
rect 24492 18702 24544 18708
rect 24398 18663 24454 18672
rect 24412 18426 24440 18663
rect 24400 18420 24452 18426
rect 24400 18362 24452 18368
rect 24504 18290 24532 18702
rect 25240 18358 25268 18770
rect 25424 18766 25452 19314
rect 25504 18964 25556 18970
rect 25504 18906 25556 18912
rect 25412 18760 25464 18766
rect 25412 18702 25464 18708
rect 25228 18352 25280 18358
rect 25228 18294 25280 18300
rect 24492 18284 24544 18290
rect 24492 18226 24544 18232
rect 24308 17876 24360 17882
rect 24308 17818 24360 17824
rect 24504 17746 24532 18226
rect 24860 18148 24912 18154
rect 24860 18090 24912 18096
rect 24768 18080 24820 18086
rect 24768 18022 24820 18028
rect 24780 17921 24808 18022
rect 24766 17912 24822 17921
rect 24872 17882 24900 18090
rect 25424 17882 25452 18702
rect 25516 18426 25544 18906
rect 25608 18902 25636 21100
rect 26146 20496 26202 20505
rect 26146 20431 26148 20440
rect 26200 20431 26202 20440
rect 26148 20402 26200 20408
rect 25872 20324 25924 20330
rect 25872 20266 25924 20272
rect 25884 19718 25912 20266
rect 26148 19848 26200 19854
rect 26252 19836 26280 21286
rect 26344 20330 26372 21558
rect 26332 20324 26384 20330
rect 26332 20266 26384 20272
rect 26200 19808 26280 19836
rect 26148 19790 26200 19796
rect 25780 19712 25832 19718
rect 25780 19654 25832 19660
rect 25872 19712 25924 19718
rect 25872 19654 25924 19660
rect 26056 19712 26108 19718
rect 26056 19654 26108 19660
rect 25596 18896 25648 18902
rect 25596 18838 25648 18844
rect 25792 18834 25820 19654
rect 25780 18828 25832 18834
rect 25780 18770 25832 18776
rect 25792 18426 25820 18770
rect 25504 18420 25556 18426
rect 25504 18362 25556 18368
rect 25780 18420 25832 18426
rect 25780 18362 25832 18368
rect 24766 17847 24822 17856
rect 24860 17876 24912 17882
rect 24780 17814 24808 17847
rect 24860 17818 24912 17824
rect 25412 17876 25464 17882
rect 25412 17818 25464 17824
rect 24768 17808 24820 17814
rect 24768 17750 24820 17756
rect 24492 17740 24544 17746
rect 24492 17682 24544 17688
rect 25228 17740 25280 17746
rect 25228 17682 25280 17688
rect 25136 17604 25188 17610
rect 25136 17546 25188 17552
rect 24952 17536 25004 17542
rect 24952 17478 25004 17484
rect 24964 17134 24992 17478
rect 24860 17128 24912 17134
rect 24860 17070 24912 17076
rect 24952 17128 25004 17134
rect 24952 17070 25004 17076
rect 24872 16726 24900 17070
rect 24860 16720 24912 16726
rect 24860 16662 24912 16668
rect 24872 16046 24900 16662
rect 25148 16182 25176 17546
rect 25240 16998 25268 17682
rect 25320 17672 25372 17678
rect 25320 17614 25372 17620
rect 25332 17066 25360 17614
rect 25884 17542 25912 19654
rect 26068 19514 26096 19654
rect 26056 19508 26108 19514
rect 26056 19450 26108 19456
rect 25964 18896 26016 18902
rect 25964 18838 26016 18844
rect 25976 18222 26004 18838
rect 25964 18216 26016 18222
rect 25964 18158 26016 18164
rect 25872 17536 25924 17542
rect 25872 17478 25924 17484
rect 26436 17218 26464 24550
rect 27160 23248 27212 23254
rect 27160 23190 27212 23196
rect 26792 23180 26844 23186
rect 26792 23122 26844 23128
rect 26804 22710 26832 23122
rect 27172 23089 27200 23190
rect 27158 23080 27214 23089
rect 27158 23015 27214 23024
rect 27172 22778 27200 23015
rect 27160 22772 27212 22778
rect 27160 22714 27212 22720
rect 26792 22704 26844 22710
rect 26792 22646 26844 22652
rect 26804 22166 26832 22646
rect 26792 22160 26844 22166
rect 26792 22102 26844 22108
rect 26516 22024 26568 22030
rect 26516 21966 26568 21972
rect 26528 21418 26556 21966
rect 26804 21690 26832 22102
rect 27894 21992 27950 22001
rect 27894 21927 27950 21936
rect 27160 21888 27212 21894
rect 27160 21830 27212 21836
rect 26792 21684 26844 21690
rect 26792 21626 26844 21632
rect 26516 21412 26568 21418
rect 26516 21354 26568 21360
rect 26608 21140 26660 21146
rect 26608 21082 26660 21088
rect 26516 20800 26568 20806
rect 26516 20742 26568 20748
rect 26528 19310 26556 20742
rect 26620 20602 26648 21082
rect 27172 20942 27200 21830
rect 27908 21690 27936 21927
rect 27896 21684 27948 21690
rect 27896 21626 27948 21632
rect 27908 21486 27936 21626
rect 27896 21480 27948 21486
rect 27896 21422 27948 21428
rect 27620 21412 27672 21418
rect 27620 21354 27672 21360
rect 26976 20936 27028 20942
rect 26976 20878 27028 20884
rect 27160 20936 27212 20942
rect 27160 20878 27212 20884
rect 26608 20596 26660 20602
rect 26608 20538 26660 20544
rect 26606 20088 26662 20097
rect 26988 20058 27016 20878
rect 27172 20330 27200 20878
rect 27632 20806 27660 21354
rect 28080 21004 28132 21010
rect 28080 20946 28132 20952
rect 27620 20800 27672 20806
rect 27620 20742 27672 20748
rect 27632 20330 27660 20742
rect 28092 20602 28120 20946
rect 28080 20596 28132 20602
rect 28080 20538 28132 20544
rect 28092 20369 28120 20538
rect 28078 20360 28134 20369
rect 27160 20324 27212 20330
rect 27160 20266 27212 20272
rect 27620 20324 27672 20330
rect 28078 20295 28134 20304
rect 27620 20266 27672 20272
rect 26606 20023 26662 20032
rect 26976 20052 27028 20058
rect 26620 19922 26648 20023
rect 27172 20040 27200 20266
rect 27252 20052 27304 20058
rect 27172 20012 27252 20040
rect 26976 19994 27028 20000
rect 27252 19994 27304 20000
rect 26608 19916 26660 19922
rect 26608 19858 26660 19864
rect 26620 19514 26648 19858
rect 26608 19508 26660 19514
rect 26608 19450 26660 19456
rect 26516 19304 26568 19310
rect 26516 19246 26568 19252
rect 26882 19272 26938 19281
rect 26882 19207 26884 19216
rect 26936 19207 26938 19216
rect 26884 19178 26936 19184
rect 26884 18828 26936 18834
rect 26884 18770 26936 18776
rect 26896 18737 26924 18770
rect 26882 18728 26938 18737
rect 26988 18698 27016 19994
rect 27632 19922 27660 20266
rect 28080 20256 28132 20262
rect 28080 20198 28132 20204
rect 28092 19990 28120 20198
rect 28080 19984 28132 19990
rect 28080 19926 28132 19932
rect 27620 19916 27672 19922
rect 27620 19858 27672 19864
rect 28092 19514 28120 19926
rect 28080 19508 28132 19514
rect 28080 19450 28132 19456
rect 27804 19304 27856 19310
rect 27804 19246 27856 19252
rect 27816 18970 27844 19246
rect 27804 18964 27856 18970
rect 27804 18906 27856 18912
rect 27802 18864 27858 18873
rect 27802 18799 27858 18808
rect 26882 18663 26938 18672
rect 26976 18692 27028 18698
rect 26976 18634 27028 18640
rect 27816 18222 27844 18799
rect 27804 18216 27856 18222
rect 27804 18158 27856 18164
rect 26514 17912 26570 17921
rect 27816 17882 27844 18158
rect 26514 17847 26516 17856
rect 26568 17847 26570 17856
rect 27804 17876 27856 17882
rect 26516 17818 26568 17824
rect 27804 17818 27856 17824
rect 26884 17740 26936 17746
rect 26884 17682 26936 17688
rect 26436 17190 26832 17218
rect 25320 17060 25372 17066
rect 25320 17002 25372 17008
rect 25228 16992 25280 16998
rect 25228 16934 25280 16940
rect 26240 16992 26292 16998
rect 26240 16934 26292 16940
rect 25240 16794 25268 16934
rect 25228 16788 25280 16794
rect 25228 16730 25280 16736
rect 25136 16176 25188 16182
rect 25136 16118 25188 16124
rect 24584 16040 24636 16046
rect 24584 15982 24636 15988
rect 24860 16040 24912 16046
rect 24860 15982 24912 15988
rect 24596 14618 24624 15982
rect 25780 15972 25832 15978
rect 25780 15914 25832 15920
rect 25792 15881 25820 15914
rect 25778 15872 25834 15881
rect 25778 15807 25834 15816
rect 26252 15201 26280 16934
rect 26516 16584 26568 16590
rect 26516 16526 26568 16532
rect 26528 16046 26556 16526
rect 26516 16040 26568 16046
rect 26516 15982 26568 15988
rect 26528 15366 26556 15982
rect 26516 15360 26568 15366
rect 26516 15302 26568 15308
rect 26238 15192 26294 15201
rect 26238 15127 26294 15136
rect 26516 14884 26568 14890
rect 26516 14826 26568 14832
rect 26528 14618 26556 14826
rect 26608 14816 26660 14822
rect 26608 14758 26660 14764
rect 24584 14612 24636 14618
rect 24584 14554 24636 14560
rect 26516 14612 26568 14618
rect 26516 14554 26568 14560
rect 24596 13394 24624 14554
rect 26148 14068 26200 14074
rect 26148 14010 26200 14016
rect 26160 13530 26188 14010
rect 25596 13524 25648 13530
rect 25596 13466 25648 13472
rect 26148 13524 26200 13530
rect 26148 13466 26200 13472
rect 24676 13456 24728 13462
rect 24676 13398 24728 13404
rect 24584 13388 24636 13394
rect 24584 13330 24636 13336
rect 24688 12986 24716 13398
rect 25608 12986 25636 13466
rect 26620 13394 26648 14758
rect 26700 13864 26752 13870
rect 26700 13806 26752 13812
rect 26608 13388 26660 13394
rect 26608 13330 26660 13336
rect 24676 12980 24728 12986
rect 24676 12922 24728 12928
rect 25596 12980 25648 12986
rect 25596 12922 25648 12928
rect 24860 12912 24912 12918
rect 24860 12854 24912 12860
rect 24584 12844 24636 12850
rect 24584 12786 24636 12792
rect 24596 12102 24624 12786
rect 24872 12306 24900 12854
rect 25688 12776 25740 12782
rect 25688 12718 25740 12724
rect 24860 12300 24912 12306
rect 24860 12242 24912 12248
rect 24584 12096 24636 12102
rect 24584 12038 24636 12044
rect 24308 11008 24360 11014
rect 24308 10950 24360 10956
rect 24320 10538 24348 10950
rect 24596 10674 24624 12038
rect 24872 11898 24900 12242
rect 25700 12102 25728 12718
rect 26620 12442 26648 13330
rect 26608 12436 26660 12442
rect 26608 12378 26660 12384
rect 26608 12232 26660 12238
rect 26608 12174 26660 12180
rect 25504 12096 25556 12102
rect 25504 12038 25556 12044
rect 25688 12096 25740 12102
rect 25688 12038 25740 12044
rect 25516 11898 25544 12038
rect 24860 11892 24912 11898
rect 24860 11834 24912 11840
rect 25504 11892 25556 11898
rect 25504 11834 25556 11840
rect 25320 11212 25372 11218
rect 25320 11154 25372 11160
rect 25332 10742 25360 11154
rect 25320 10736 25372 10742
rect 25320 10678 25372 10684
rect 24584 10668 24636 10674
rect 24584 10610 24636 10616
rect 24308 10532 24360 10538
rect 24308 10474 24360 10480
rect 25700 9518 25728 12038
rect 26620 11830 26648 12174
rect 26712 11898 26740 13806
rect 26700 11892 26752 11898
rect 26700 11834 26752 11840
rect 26608 11824 26660 11830
rect 26608 11766 26660 11772
rect 26240 11552 26292 11558
rect 26240 11494 26292 11500
rect 26252 9636 26280 11494
rect 26424 11212 26476 11218
rect 26424 11154 26476 11160
rect 26436 10470 26464 11154
rect 26424 10464 26476 10470
rect 26424 10406 26476 10412
rect 26608 10464 26660 10470
rect 26608 10406 26660 10412
rect 26436 10266 26464 10406
rect 26424 10260 26476 10266
rect 26424 10202 26476 10208
rect 26332 9920 26384 9926
rect 26332 9862 26384 9868
rect 26160 9608 26280 9636
rect 24860 9512 24912 9518
rect 24860 9454 24912 9460
rect 25688 9512 25740 9518
rect 25688 9454 25740 9460
rect 24492 9444 24544 9450
rect 24492 9386 24544 9392
rect 24504 8906 24532 9386
rect 24872 9178 24900 9454
rect 26056 9444 26108 9450
rect 26056 9386 26108 9392
rect 24860 9172 24912 9178
rect 24860 9114 24912 9120
rect 24492 8900 24544 8906
rect 24492 8842 24544 8848
rect 24504 8090 24532 8842
rect 26068 8634 26096 9386
rect 26160 9042 26188 9608
rect 26240 9512 26292 9518
rect 26344 9466 26372 9862
rect 26292 9460 26372 9466
rect 26240 9454 26372 9460
rect 26252 9438 26372 9454
rect 26148 9036 26200 9042
rect 26148 8978 26200 8984
rect 26056 8628 26108 8634
rect 26056 8570 26108 8576
rect 26160 8090 26188 8978
rect 26252 8974 26280 9438
rect 26436 9042 26464 10202
rect 26620 9926 26648 10406
rect 26608 9920 26660 9926
rect 26608 9862 26660 9868
rect 26424 9036 26476 9042
rect 26424 8978 26476 8984
rect 26240 8968 26292 8974
rect 26240 8910 26292 8916
rect 26436 8634 26464 8978
rect 26516 8968 26568 8974
rect 26516 8910 26568 8916
rect 26424 8628 26476 8634
rect 26424 8570 26476 8576
rect 24492 8084 24544 8090
rect 24492 8026 24544 8032
rect 26148 8084 26200 8090
rect 26148 8026 26200 8032
rect 26528 6798 26556 8910
rect 26620 8634 26648 9862
rect 26608 8628 26660 8634
rect 26608 8570 26660 8576
rect 26804 6866 26832 17190
rect 26896 16998 26924 17682
rect 26976 17672 27028 17678
rect 26976 17614 27028 17620
rect 26988 17134 27016 17614
rect 27896 17536 27948 17542
rect 27434 17504 27490 17513
rect 27434 17439 27490 17448
rect 27710 17504 27766 17513
rect 27896 17478 27948 17484
rect 27710 17439 27766 17448
rect 27448 17338 27476 17439
rect 27618 17368 27674 17377
rect 27436 17332 27488 17338
rect 27618 17303 27674 17312
rect 27436 17274 27488 17280
rect 27632 17134 27660 17303
rect 26976 17128 27028 17134
rect 26976 17070 27028 17076
rect 27620 17128 27672 17134
rect 27620 17070 27672 17076
rect 26884 16992 26936 16998
rect 26884 16934 26936 16940
rect 26988 16794 27016 17070
rect 26976 16788 27028 16794
rect 26976 16730 27028 16736
rect 27068 16652 27120 16658
rect 27068 16594 27120 16600
rect 27080 16250 27108 16594
rect 27068 16244 27120 16250
rect 27068 16186 27120 16192
rect 27160 15904 27212 15910
rect 27160 15846 27212 15852
rect 27172 15434 27200 15846
rect 27160 15428 27212 15434
rect 27160 15370 27212 15376
rect 27068 15360 27120 15366
rect 27068 15302 27120 15308
rect 27080 15094 27108 15302
rect 27068 15088 27120 15094
rect 27068 15030 27120 15036
rect 27172 15026 27200 15370
rect 27344 15360 27396 15366
rect 27344 15302 27396 15308
rect 27160 15020 27212 15026
rect 27160 14962 27212 14968
rect 27068 14544 27120 14550
rect 27068 14486 27120 14492
rect 26976 14408 27028 14414
rect 26976 14350 27028 14356
rect 26988 14074 27016 14350
rect 26976 14068 27028 14074
rect 26976 14010 27028 14016
rect 27080 13802 27108 14486
rect 27068 13796 27120 13802
rect 27068 13738 27120 13744
rect 27080 12986 27108 13738
rect 27068 12980 27120 12986
rect 27068 12922 27120 12928
rect 27172 11354 27200 14962
rect 27356 14958 27384 15302
rect 27344 14952 27396 14958
rect 27344 14894 27396 14900
rect 27344 14408 27396 14414
rect 27344 14350 27396 14356
rect 27356 13530 27384 14350
rect 27344 13524 27396 13530
rect 27344 13466 27396 13472
rect 27356 11778 27384 13466
rect 27620 13184 27672 13190
rect 27620 13126 27672 13132
rect 27436 12436 27488 12442
rect 27436 12378 27488 12384
rect 27448 12345 27476 12378
rect 27434 12336 27490 12345
rect 27632 12306 27660 13126
rect 27434 12271 27490 12280
rect 27620 12300 27672 12306
rect 27620 12242 27672 12248
rect 27356 11762 27476 11778
rect 27356 11756 27488 11762
rect 27356 11750 27436 11756
rect 27436 11698 27488 11704
rect 27344 11688 27396 11694
rect 27344 11630 27396 11636
rect 27160 11348 27212 11354
rect 27160 11290 27212 11296
rect 26976 11008 27028 11014
rect 26976 10950 27028 10956
rect 26988 10674 27016 10950
rect 27172 10674 27200 11290
rect 27356 10810 27384 11630
rect 27448 11150 27476 11698
rect 27528 11280 27580 11286
rect 27528 11222 27580 11228
rect 27436 11144 27488 11150
rect 27436 11086 27488 11092
rect 27344 10804 27396 10810
rect 27344 10746 27396 10752
rect 26976 10668 27028 10674
rect 26976 10610 27028 10616
rect 27160 10668 27212 10674
rect 27160 10610 27212 10616
rect 27448 10538 27476 11086
rect 27540 10962 27568 11222
rect 27540 10934 27660 10962
rect 27160 10532 27212 10538
rect 27160 10474 27212 10480
rect 27436 10532 27488 10538
rect 27436 10474 27488 10480
rect 27172 8498 27200 10474
rect 27632 10470 27660 10934
rect 27620 10464 27672 10470
rect 27620 10406 27672 10412
rect 27632 10130 27660 10406
rect 27620 10124 27672 10130
rect 27620 10066 27672 10072
rect 27632 9382 27660 10066
rect 27528 9376 27580 9382
rect 27528 9318 27580 9324
rect 27620 9376 27672 9382
rect 27620 9318 27672 9324
rect 27160 8492 27212 8498
rect 27160 8434 27212 8440
rect 26884 8424 26936 8430
rect 26884 8366 26936 8372
rect 26896 8090 26924 8366
rect 27172 8090 27200 8434
rect 27540 8430 27568 9318
rect 27724 9042 27752 17439
rect 27908 17338 27936 17478
rect 27896 17332 27948 17338
rect 27896 17274 27948 17280
rect 27988 15564 28040 15570
rect 27988 15506 28040 15512
rect 27804 15496 27856 15502
rect 27804 15438 27856 15444
rect 27896 15496 27948 15502
rect 27896 15438 27948 15444
rect 27816 15162 27844 15438
rect 27804 15156 27856 15162
rect 27804 15098 27856 15104
rect 27816 14074 27844 15098
rect 27908 14618 27936 15438
rect 28000 15162 28028 15506
rect 27988 15156 28040 15162
rect 27988 15098 28040 15104
rect 27896 14612 27948 14618
rect 27896 14554 27948 14560
rect 28000 14550 28028 15098
rect 28080 15088 28132 15094
rect 28080 15030 28132 15036
rect 27988 14544 28040 14550
rect 27988 14486 28040 14492
rect 28092 14414 28120 15030
rect 28080 14408 28132 14414
rect 28080 14350 28132 14356
rect 27804 14068 27856 14074
rect 27804 14010 27856 14016
rect 27816 13462 27844 14010
rect 28092 13870 28120 14350
rect 28080 13864 28132 13870
rect 28080 13806 28132 13812
rect 28092 13462 28120 13806
rect 27804 13456 27856 13462
rect 27804 13398 27856 13404
rect 28080 13456 28132 13462
rect 28080 13398 28132 13404
rect 27816 12986 27844 13398
rect 28092 12986 28120 13398
rect 27804 12980 27856 12986
rect 27804 12922 27856 12928
rect 28080 12980 28132 12986
rect 28080 12922 28132 12928
rect 27804 12300 27856 12306
rect 27804 12242 27856 12248
rect 27816 11898 27844 12242
rect 28080 12232 28132 12238
rect 28078 12200 28080 12209
rect 28132 12200 28134 12209
rect 28078 12135 28134 12144
rect 27804 11892 27856 11898
rect 27804 11834 27856 11840
rect 28092 11762 28120 12135
rect 28080 11756 28132 11762
rect 28080 11698 28132 11704
rect 27896 11552 27948 11558
rect 27896 11494 27948 11500
rect 27908 11082 27936 11494
rect 28092 11354 28120 11698
rect 28080 11348 28132 11354
rect 28080 11290 28132 11296
rect 27896 11076 27948 11082
rect 27896 11018 27948 11024
rect 28276 10810 28304 25706
rect 28908 25696 28960 25702
rect 28906 25664 28908 25673
rect 28960 25664 28962 25673
rect 28906 25599 28962 25608
rect 28920 25362 28948 25599
rect 28908 25356 28960 25362
rect 28908 25298 28960 25304
rect 29196 25158 29224 25774
rect 29366 25528 29422 25537
rect 29748 25498 29776 26794
rect 29840 25838 29868 26930
rect 29828 25832 29880 25838
rect 29828 25774 29880 25780
rect 29366 25463 29422 25472
rect 29736 25492 29788 25498
rect 29184 25152 29236 25158
rect 29184 25094 29236 25100
rect 29092 24268 29144 24274
rect 29092 24210 29144 24216
rect 29104 23866 29132 24210
rect 29092 23860 29144 23866
rect 29092 23802 29144 23808
rect 28724 23520 28776 23526
rect 28724 23462 28776 23468
rect 28736 22574 28764 23462
rect 28724 22568 28776 22574
rect 28724 22510 28776 22516
rect 29092 20868 29144 20874
rect 29092 20810 29144 20816
rect 29104 20602 29132 20810
rect 29092 20596 29144 20602
rect 29092 20538 29144 20544
rect 28724 19916 28776 19922
rect 28724 19858 28776 19864
rect 28736 19802 28764 19858
rect 29092 19848 29144 19854
rect 28736 19774 28856 19802
rect 29092 19790 29144 19796
rect 28356 19168 28408 19174
rect 28356 19110 28408 19116
rect 28632 19168 28684 19174
rect 28632 19110 28684 19116
rect 28368 18970 28396 19110
rect 28356 18964 28408 18970
rect 28356 18906 28408 18912
rect 28448 18760 28500 18766
rect 28448 18702 28500 18708
rect 28460 18465 28488 18702
rect 28446 18456 28502 18465
rect 28446 18391 28448 18400
rect 28500 18391 28502 18400
rect 28448 18362 28500 18368
rect 28644 18290 28672 19110
rect 28724 18964 28776 18970
rect 28724 18906 28776 18912
rect 28736 18426 28764 18906
rect 28828 18902 28856 19774
rect 29000 19712 29052 19718
rect 29000 19654 29052 19660
rect 28816 18896 28868 18902
rect 29012 18850 29040 19654
rect 29104 18970 29132 19790
rect 29092 18964 29144 18970
rect 29092 18906 29144 18912
rect 28816 18838 28868 18844
rect 28920 18822 29040 18850
rect 28920 18766 28948 18822
rect 28908 18760 28960 18766
rect 28908 18702 28960 18708
rect 29092 18760 29144 18766
rect 29092 18702 29144 18708
rect 28816 18624 28868 18630
rect 28816 18566 28868 18572
rect 28724 18420 28776 18426
rect 28724 18362 28776 18368
rect 28632 18284 28684 18290
rect 28632 18226 28684 18232
rect 28828 16810 28856 18566
rect 28920 17814 28948 18702
rect 28908 17808 28960 17814
rect 28908 17750 28960 17756
rect 29104 17542 29132 18702
rect 29092 17536 29144 17542
rect 29196 17513 29224 25094
rect 29380 19174 29408 25463
rect 29736 25434 29788 25440
rect 29840 25362 29868 25774
rect 30012 25764 30064 25770
rect 30012 25706 30064 25712
rect 30024 25362 30052 25706
rect 29828 25356 29880 25362
rect 29828 25298 29880 25304
rect 30012 25356 30064 25362
rect 30012 25298 30064 25304
rect 29736 24744 29788 24750
rect 29736 24686 29788 24692
rect 29748 24070 29776 24686
rect 29736 24064 29788 24070
rect 29736 24006 29788 24012
rect 29748 23662 29776 24006
rect 29736 23656 29788 23662
rect 29736 23598 29788 23604
rect 29748 23254 29776 23598
rect 29736 23248 29788 23254
rect 29736 23190 29788 23196
rect 29644 23180 29696 23186
rect 29644 23122 29696 23128
rect 29552 22500 29604 22506
rect 29552 22442 29604 22448
rect 29564 21690 29592 22442
rect 29656 22234 29684 23122
rect 29748 22574 29776 23190
rect 29736 22568 29788 22574
rect 29736 22510 29788 22516
rect 29644 22228 29696 22234
rect 29644 22170 29696 22176
rect 29748 21894 29776 22510
rect 29736 21888 29788 21894
rect 29736 21830 29788 21836
rect 29552 21684 29604 21690
rect 29552 21626 29604 21632
rect 29564 20874 29592 21626
rect 29828 21004 29880 21010
rect 29828 20946 29880 20952
rect 29552 20868 29604 20874
rect 29552 20810 29604 20816
rect 29460 20800 29512 20806
rect 29460 20742 29512 20748
rect 29472 20058 29500 20742
rect 29840 20602 29868 20946
rect 29828 20596 29880 20602
rect 29828 20538 29880 20544
rect 29460 20052 29512 20058
rect 29460 19994 29512 20000
rect 29472 19378 29500 19994
rect 29460 19372 29512 19378
rect 29460 19314 29512 19320
rect 29368 19168 29420 19174
rect 29368 19110 29420 19116
rect 30116 18136 30144 32535
rect 34940 31580 35236 31600
rect 34996 31578 35020 31580
rect 35076 31578 35100 31580
rect 35156 31578 35180 31580
rect 35018 31526 35020 31578
rect 35082 31526 35094 31578
rect 35156 31526 35158 31578
rect 34996 31524 35020 31526
rect 35076 31524 35100 31526
rect 35156 31524 35180 31526
rect 34940 31504 35236 31524
rect 34704 31136 34756 31142
rect 34704 31078 34756 31084
rect 34612 30320 34664 30326
rect 34612 30262 34664 30268
rect 32680 29776 32732 29782
rect 32680 29718 32732 29724
rect 31300 29640 31352 29646
rect 31300 29582 31352 29588
rect 31312 29170 31340 29582
rect 32692 29238 32720 29718
rect 34520 29708 34572 29714
rect 34520 29650 34572 29656
rect 33140 29504 33192 29510
rect 33060 29464 33140 29492
rect 32680 29232 32732 29238
rect 32680 29174 32732 29180
rect 31300 29164 31352 29170
rect 31300 29106 31352 29112
rect 31944 29096 31996 29102
rect 31944 29038 31996 29044
rect 31576 29028 31628 29034
rect 31576 28970 31628 28976
rect 30840 28960 30892 28966
rect 31588 28937 31616 28970
rect 30840 28902 30892 28908
rect 31574 28928 31630 28937
rect 30852 28490 30880 28902
rect 31574 28863 31630 28872
rect 31588 28762 31616 28863
rect 31576 28756 31628 28762
rect 31576 28698 31628 28704
rect 30932 28552 30984 28558
rect 30932 28494 30984 28500
rect 30840 28484 30892 28490
rect 30840 28426 30892 28432
rect 30472 28416 30524 28422
rect 30472 28358 30524 28364
rect 30484 27674 30512 28358
rect 30472 27668 30524 27674
rect 30472 27610 30524 27616
rect 30748 27532 30800 27538
rect 30748 27474 30800 27480
rect 30760 26790 30788 27474
rect 30748 26784 30800 26790
rect 30748 26726 30800 26732
rect 30760 26586 30788 26726
rect 30852 26586 30880 28426
rect 30944 28218 30972 28494
rect 31956 28422 31984 29038
rect 32220 28620 32272 28626
rect 32220 28562 32272 28568
rect 31944 28416 31996 28422
rect 31942 28384 31944 28393
rect 31996 28384 31998 28393
rect 31942 28319 31998 28328
rect 32232 28218 32260 28562
rect 30932 28212 30984 28218
rect 30932 28154 30984 28160
rect 32220 28212 32272 28218
rect 32220 28154 32272 28160
rect 30932 27940 30984 27946
rect 30932 27882 30984 27888
rect 30944 27334 30972 27882
rect 32588 27600 32640 27606
rect 32588 27542 32640 27548
rect 32496 27532 32548 27538
rect 32496 27474 32548 27480
rect 30932 27328 30984 27334
rect 30932 27270 30984 27276
rect 31576 27328 31628 27334
rect 31576 27270 31628 27276
rect 32128 27328 32180 27334
rect 32128 27270 32180 27276
rect 30748 26580 30800 26586
rect 30748 26522 30800 26528
rect 30840 26580 30892 26586
rect 30840 26522 30892 26528
rect 30852 26382 30880 26522
rect 30944 26450 30972 27270
rect 30932 26444 30984 26450
rect 30932 26386 30984 26392
rect 31484 26444 31536 26450
rect 31484 26386 31536 26392
rect 30840 26376 30892 26382
rect 30194 26344 30250 26353
rect 30840 26318 30892 26324
rect 30194 26279 30250 26288
rect 30208 25498 30236 26279
rect 30196 25492 30248 25498
rect 30196 25434 30248 25440
rect 30656 25356 30708 25362
rect 30656 25298 30708 25304
rect 30668 24954 30696 25298
rect 30852 25294 30880 26318
rect 31496 25906 31524 26386
rect 31588 26246 31616 27270
rect 31668 26784 31720 26790
rect 31720 26732 31800 26738
rect 31668 26726 31800 26732
rect 31680 26710 31800 26726
rect 31668 26376 31720 26382
rect 31668 26318 31720 26324
rect 31576 26240 31628 26246
rect 31576 26182 31628 26188
rect 31484 25900 31536 25906
rect 31484 25842 31536 25848
rect 31116 25696 31168 25702
rect 31116 25638 31168 25644
rect 31128 25430 31156 25638
rect 31588 25430 31616 26182
rect 31680 25498 31708 26318
rect 31772 26042 31800 26710
rect 32140 26625 32168 27270
rect 32508 27062 32536 27474
rect 32600 27130 32628 27542
rect 32588 27124 32640 27130
rect 32588 27066 32640 27072
rect 32496 27056 32548 27062
rect 32496 26998 32548 27004
rect 32692 26994 32720 29174
rect 32956 28076 33008 28082
rect 32956 28018 33008 28024
rect 32968 27878 32996 28018
rect 32956 27872 33008 27878
rect 32956 27814 33008 27820
rect 32968 26994 32996 27814
rect 32680 26988 32732 26994
rect 32680 26930 32732 26936
rect 32956 26988 33008 26994
rect 32956 26930 33008 26936
rect 32126 26616 32182 26625
rect 32968 26586 32996 26930
rect 33060 26858 33088 29464
rect 33140 29446 33192 29452
rect 34532 29034 34560 29650
rect 34520 29028 34572 29034
rect 34520 28970 34572 28976
rect 34336 28960 34388 28966
rect 33506 28928 33562 28937
rect 34336 28902 34388 28908
rect 33506 28863 33562 28872
rect 33520 28762 33548 28863
rect 33508 28756 33560 28762
rect 33508 28698 33560 28704
rect 34348 28422 34376 28902
rect 34336 28416 34388 28422
rect 34336 28358 34388 28364
rect 33968 28212 34020 28218
rect 33968 28154 34020 28160
rect 33324 27940 33376 27946
rect 33324 27882 33376 27888
rect 33336 27674 33364 27882
rect 33324 27668 33376 27674
rect 33324 27610 33376 27616
rect 33048 26852 33100 26858
rect 33048 26794 33100 26800
rect 32126 26551 32182 26560
rect 32680 26580 32732 26586
rect 32680 26522 32732 26528
rect 32956 26580 33008 26586
rect 32956 26522 33008 26528
rect 31944 26512 31996 26518
rect 31944 26454 31996 26460
rect 31956 26353 31984 26454
rect 31942 26344 31998 26353
rect 31942 26279 31998 26288
rect 32312 26308 32364 26314
rect 32312 26250 32364 26256
rect 31760 26036 31812 26042
rect 31760 25978 31812 25984
rect 31760 25832 31812 25838
rect 31760 25774 31812 25780
rect 31772 25498 31800 25774
rect 31942 25664 31998 25673
rect 31942 25599 31998 25608
rect 31668 25492 31720 25498
rect 31668 25434 31720 25440
rect 31760 25492 31812 25498
rect 31760 25434 31812 25440
rect 31116 25424 31168 25430
rect 31116 25366 31168 25372
rect 31576 25424 31628 25430
rect 31576 25366 31628 25372
rect 30840 25288 30892 25294
rect 30840 25230 30892 25236
rect 30656 24948 30708 24954
rect 30656 24890 30708 24896
rect 30852 24614 30880 25230
rect 31588 25226 31616 25366
rect 31956 25362 31984 25599
rect 31944 25356 31996 25362
rect 31996 25316 32076 25344
rect 31944 25298 31996 25304
rect 31576 25220 31628 25226
rect 31576 25162 31628 25168
rect 31944 24948 31996 24954
rect 31944 24890 31996 24896
rect 30932 24676 30984 24682
rect 30932 24618 30984 24624
rect 30840 24608 30892 24614
rect 30840 24550 30892 24556
rect 30944 24410 30972 24618
rect 31116 24608 31168 24614
rect 31116 24550 31168 24556
rect 30932 24404 30984 24410
rect 30932 24346 30984 24352
rect 31128 24274 31156 24550
rect 31956 24410 31984 24890
rect 31944 24404 31996 24410
rect 31944 24346 31996 24352
rect 32048 24342 32076 25316
rect 32128 25288 32180 25294
rect 32128 25230 32180 25236
rect 32140 24614 32168 25230
rect 32220 25152 32272 25158
rect 32220 25094 32272 25100
rect 32128 24608 32180 24614
rect 32128 24550 32180 24556
rect 32140 24410 32168 24550
rect 32128 24404 32180 24410
rect 32128 24346 32180 24352
rect 32036 24336 32088 24342
rect 32036 24278 32088 24284
rect 31116 24268 31168 24274
rect 31116 24210 31168 24216
rect 32128 24268 32180 24274
rect 32128 24210 32180 24216
rect 31128 23866 31156 24210
rect 32140 23866 32168 24210
rect 31116 23860 31168 23866
rect 31116 23802 31168 23808
rect 32128 23860 32180 23866
rect 32128 23802 32180 23808
rect 30932 23588 30984 23594
rect 30932 23530 30984 23536
rect 30944 23322 30972 23530
rect 31760 23520 31812 23526
rect 31760 23462 31812 23468
rect 30932 23316 30984 23322
rect 30932 23258 30984 23264
rect 31024 23180 31076 23186
rect 31024 23122 31076 23128
rect 31036 22778 31064 23122
rect 31772 22794 31800 23462
rect 32140 23322 32168 23802
rect 32128 23316 32180 23322
rect 32128 23258 32180 23264
rect 32232 23186 32260 25094
rect 32324 23662 32352 26250
rect 32496 25356 32548 25362
rect 32496 25298 32548 25304
rect 32508 24954 32536 25298
rect 32496 24948 32548 24954
rect 32496 24890 32548 24896
rect 32692 24818 32720 26522
rect 33048 26376 33100 26382
rect 33048 26318 33100 26324
rect 33060 25838 33088 26318
rect 33324 25968 33376 25974
rect 33324 25910 33376 25916
rect 33048 25832 33100 25838
rect 33048 25774 33100 25780
rect 32864 25696 32916 25702
rect 32864 25638 32916 25644
rect 32680 24812 32732 24818
rect 32680 24754 32732 24760
rect 32692 24206 32720 24754
rect 32588 24200 32640 24206
rect 32588 24142 32640 24148
rect 32680 24200 32732 24206
rect 32680 24142 32732 24148
rect 32312 23656 32364 23662
rect 32312 23598 32364 23604
rect 32600 23594 32628 24142
rect 32692 23798 32720 24142
rect 32680 23792 32732 23798
rect 32680 23734 32732 23740
rect 32588 23588 32640 23594
rect 32588 23530 32640 23536
rect 32876 23322 32904 25638
rect 33060 25106 33088 25774
rect 33140 25696 33192 25702
rect 33140 25638 33192 25644
rect 33152 25158 33180 25638
rect 32968 25078 33088 25106
rect 33140 25152 33192 25158
rect 33140 25094 33192 25100
rect 32864 23316 32916 23322
rect 32864 23258 32916 23264
rect 32220 23180 32272 23186
rect 32220 23122 32272 23128
rect 31680 22778 31800 22794
rect 32232 22778 32260 23122
rect 32968 22778 32996 25078
rect 33152 24970 33180 25094
rect 33060 24942 33180 24970
rect 33060 23866 33088 24942
rect 33336 24138 33364 25910
rect 33692 25900 33744 25906
rect 33692 25842 33744 25848
rect 33704 25226 33732 25842
rect 33876 25424 33928 25430
rect 33876 25366 33928 25372
rect 33692 25220 33744 25226
rect 33692 25162 33744 25168
rect 33784 24744 33836 24750
rect 33784 24686 33836 24692
rect 33796 24410 33824 24686
rect 33784 24404 33836 24410
rect 33784 24346 33836 24352
rect 33324 24132 33376 24138
rect 33324 24074 33376 24080
rect 33048 23860 33100 23866
rect 33048 23802 33100 23808
rect 33336 23186 33364 24074
rect 33324 23180 33376 23186
rect 33324 23122 33376 23128
rect 33336 22778 33364 23122
rect 31024 22772 31076 22778
rect 31024 22714 31076 22720
rect 31668 22772 31800 22778
rect 31720 22766 31800 22772
rect 32220 22772 32272 22778
rect 31668 22714 31720 22720
rect 32220 22714 32272 22720
rect 32956 22772 33008 22778
rect 32956 22714 33008 22720
rect 33324 22772 33376 22778
rect 33324 22714 33376 22720
rect 32968 22574 32996 22714
rect 33888 22574 33916 25366
rect 32956 22568 33008 22574
rect 32956 22510 33008 22516
rect 33876 22568 33928 22574
rect 33876 22510 33928 22516
rect 32128 22432 32180 22438
rect 32128 22374 32180 22380
rect 32140 22030 32168 22374
rect 33888 22234 33916 22510
rect 33876 22228 33928 22234
rect 33876 22170 33928 22176
rect 32128 22024 32180 22030
rect 32128 21966 32180 21972
rect 30564 21888 30616 21894
rect 30564 21830 30616 21836
rect 30576 21486 30604 21830
rect 30564 21480 30616 21486
rect 30564 21422 30616 21428
rect 30196 21412 30248 21418
rect 30196 21354 30248 21360
rect 30208 19990 30236 21354
rect 30576 21146 30604 21422
rect 32140 21146 32168 21966
rect 33324 21412 33376 21418
rect 33324 21354 33376 21360
rect 33336 21146 33364 21354
rect 30564 21140 30616 21146
rect 30564 21082 30616 21088
rect 32128 21140 32180 21146
rect 32128 21082 32180 21088
rect 33324 21140 33376 21146
rect 33324 21082 33376 21088
rect 30288 21004 30340 21010
rect 30340 20964 30420 20992
rect 30288 20946 30340 20952
rect 30392 20058 30420 20964
rect 30576 20466 30604 21082
rect 33336 20466 33364 21082
rect 33692 20936 33744 20942
rect 33692 20878 33744 20884
rect 30564 20460 30616 20466
rect 30564 20402 30616 20408
rect 33324 20460 33376 20466
rect 33324 20402 33376 20408
rect 30380 20052 30432 20058
rect 30380 19994 30432 20000
rect 30196 19984 30248 19990
rect 30196 19926 30248 19932
rect 30576 19378 30604 20402
rect 33416 20392 33468 20398
rect 33416 20334 33468 20340
rect 30932 20324 30984 20330
rect 30932 20266 30984 20272
rect 30748 19916 30800 19922
rect 30748 19858 30800 19864
rect 30196 19372 30248 19378
rect 30196 19314 30248 19320
rect 30564 19372 30616 19378
rect 30564 19314 30616 19320
rect 30208 18834 30236 19314
rect 30760 19310 30788 19858
rect 30944 19718 30972 20266
rect 31944 20256 31996 20262
rect 31944 20198 31996 20204
rect 31956 19854 31984 20198
rect 33428 20058 33456 20334
rect 33416 20052 33468 20058
rect 33416 19994 33468 20000
rect 31944 19848 31996 19854
rect 31944 19790 31996 19796
rect 30932 19712 30984 19718
rect 30932 19654 30984 19660
rect 32404 19712 32456 19718
rect 32404 19654 32456 19660
rect 30748 19304 30800 19310
rect 30748 19246 30800 19252
rect 30380 19168 30432 19174
rect 30380 19110 30432 19116
rect 30288 18896 30340 18902
rect 30392 18873 30420 19110
rect 30944 18970 30972 19654
rect 32416 19378 32444 19654
rect 32404 19372 32456 19378
rect 32404 19314 32456 19320
rect 33048 19304 33100 19310
rect 32310 19272 32366 19281
rect 32128 19236 32180 19242
rect 33048 19246 33100 19252
rect 32310 19207 32366 19216
rect 32128 19178 32180 19184
rect 31300 19168 31352 19174
rect 31300 19110 31352 19116
rect 30932 18964 30984 18970
rect 30932 18906 30984 18912
rect 30288 18838 30340 18844
rect 30378 18864 30434 18873
rect 30196 18828 30248 18834
rect 30196 18770 30248 18776
rect 30085 18108 30144 18136
rect 29552 18080 29604 18086
rect 30085 18068 30113 18108
rect 30085 18040 30144 18068
rect 29552 18022 29604 18028
rect 29460 17808 29512 17814
rect 29460 17750 29512 17756
rect 29092 17478 29144 17484
rect 29182 17504 29238 17513
rect 29104 17338 29132 17478
rect 29182 17439 29238 17448
rect 29472 17338 29500 17750
rect 29092 17332 29144 17338
rect 29092 17274 29144 17280
rect 29460 17332 29512 17338
rect 29460 17274 29512 17280
rect 28828 16782 29040 16810
rect 29012 16658 29040 16782
rect 29564 16726 29592 18022
rect 29920 16788 29972 16794
rect 29920 16730 29972 16736
rect 29552 16720 29604 16726
rect 29932 16697 29960 16730
rect 29552 16662 29604 16668
rect 29918 16688 29974 16697
rect 29000 16652 29052 16658
rect 29918 16623 29974 16632
rect 29000 16594 29052 16600
rect 29918 16280 29974 16289
rect 29918 16215 29920 16224
rect 29972 16215 29974 16224
rect 29920 16186 29972 16192
rect 28630 16144 28686 16153
rect 28630 16079 28632 16088
rect 28684 16079 28686 16088
rect 28632 16050 28684 16056
rect 29932 16046 29960 16186
rect 29920 16040 29972 16046
rect 29920 15982 29972 15988
rect 29460 15904 29512 15910
rect 29460 15846 29512 15852
rect 29472 15502 29500 15846
rect 29736 15564 29788 15570
rect 29736 15506 29788 15512
rect 29460 15496 29512 15502
rect 29460 15438 29512 15444
rect 29748 15162 29776 15506
rect 29736 15156 29788 15162
rect 29736 15098 29788 15104
rect 30012 14952 30064 14958
rect 30012 14894 30064 14900
rect 30024 14618 30052 14894
rect 30012 14612 30064 14618
rect 30012 14554 30064 14560
rect 28724 14544 28776 14550
rect 28724 14486 28776 14492
rect 28736 14074 28764 14486
rect 30024 14074 30052 14554
rect 28724 14068 28776 14074
rect 28724 14010 28776 14016
rect 29000 14068 29052 14074
rect 29000 14010 29052 14016
rect 30012 14068 30064 14074
rect 30012 14010 30064 14016
rect 29012 13530 29040 14010
rect 30024 13870 30052 14010
rect 30012 13864 30064 13870
rect 30012 13806 30064 13812
rect 29000 13524 29052 13530
rect 29000 13466 29052 13472
rect 30012 13184 30064 13190
rect 30012 13126 30064 13132
rect 30024 12782 30052 13126
rect 29644 12776 29696 12782
rect 29644 12718 29696 12724
rect 30012 12776 30064 12782
rect 30012 12718 30064 12724
rect 29656 12442 29684 12718
rect 30116 12628 30144 18040
rect 30300 17354 30328 18838
rect 30378 18799 30434 18808
rect 30392 18426 30420 18799
rect 30564 18692 30616 18698
rect 30564 18634 30616 18640
rect 30380 18420 30432 18426
rect 30380 18362 30432 18368
rect 30392 18154 30420 18362
rect 30576 18222 30604 18634
rect 31312 18465 31340 19110
rect 32140 18970 32168 19178
rect 32324 19174 32352 19207
rect 32312 19168 32364 19174
rect 32312 19110 32364 19116
rect 32772 19168 32824 19174
rect 32772 19110 32824 19116
rect 32128 18964 32180 18970
rect 32128 18906 32180 18912
rect 32128 18624 32180 18630
rect 32128 18566 32180 18572
rect 31298 18456 31354 18465
rect 31298 18391 31354 18400
rect 31312 18222 31340 18391
rect 30564 18216 30616 18222
rect 30564 18158 30616 18164
rect 31300 18216 31352 18222
rect 31300 18158 31352 18164
rect 31760 18216 31812 18222
rect 31760 18158 31812 18164
rect 30380 18148 30432 18154
rect 30380 18090 30432 18096
rect 31312 17882 31340 18158
rect 31772 17882 31800 18158
rect 31300 17876 31352 17882
rect 31300 17818 31352 17824
rect 31760 17876 31812 17882
rect 31760 17818 31812 17824
rect 32140 17610 32168 18566
rect 32324 18057 32352 19110
rect 32784 18630 32812 19110
rect 32772 18624 32824 18630
rect 32772 18566 32824 18572
rect 32588 18080 32640 18086
rect 32310 18048 32366 18057
rect 32588 18022 32640 18028
rect 32310 17983 32366 17992
rect 32600 17882 32628 18022
rect 32496 17876 32548 17882
rect 32496 17818 32548 17824
rect 32588 17876 32640 17882
rect 32588 17818 32640 17824
rect 32128 17604 32180 17610
rect 32128 17546 32180 17552
rect 30472 17536 30524 17542
rect 30472 17478 30524 17484
rect 30300 17338 30420 17354
rect 30300 17332 30432 17338
rect 30300 17326 30380 17332
rect 30380 17274 30432 17280
rect 30484 17134 30512 17478
rect 32508 17270 32536 17818
rect 32496 17264 32548 17270
rect 32496 17206 32548 17212
rect 32600 17202 32628 17818
rect 32772 17672 32824 17678
rect 32772 17614 32824 17620
rect 32784 17338 32812 17614
rect 32772 17332 32824 17338
rect 32772 17274 32824 17280
rect 32588 17196 32640 17202
rect 32588 17138 32640 17144
rect 30288 17128 30340 17134
rect 30472 17128 30524 17134
rect 30340 17076 30420 17082
rect 30288 17070 30420 17076
rect 30472 17070 30524 17076
rect 30300 17054 30420 17070
rect 30392 16794 30420 17054
rect 30380 16788 30432 16794
rect 30380 16730 30432 16736
rect 30196 16720 30248 16726
rect 30392 16674 30420 16730
rect 30196 16662 30248 16668
rect 30208 16250 30236 16662
rect 30300 16646 30420 16674
rect 30196 16244 30248 16250
rect 30196 16186 30248 16192
rect 30196 15360 30248 15366
rect 30196 15302 30248 15308
rect 30208 13410 30236 15302
rect 30300 14482 30328 16646
rect 30484 16590 30512 17070
rect 30380 16584 30432 16590
rect 30380 16526 30432 16532
rect 30472 16584 30524 16590
rect 30472 16526 30524 16532
rect 30392 15706 30420 16526
rect 30484 16250 30512 16526
rect 30472 16244 30524 16250
rect 30472 16186 30524 16192
rect 33060 16182 33088 19246
rect 33428 18154 33456 19994
rect 33704 18834 33732 20878
rect 33876 20528 33928 20534
rect 33876 20470 33928 20476
rect 33782 20360 33838 20369
rect 33782 20295 33838 20304
rect 33796 19854 33824 20295
rect 33784 19848 33836 19854
rect 33784 19790 33836 19796
rect 33796 19174 33824 19790
rect 33784 19168 33836 19174
rect 33784 19110 33836 19116
rect 33888 18873 33916 20470
rect 33980 19281 34008 28154
rect 34348 27878 34376 28358
rect 34532 28234 34560 28970
rect 34440 28206 34560 28234
rect 34624 28218 34652 30262
rect 34612 28212 34664 28218
rect 34336 27872 34388 27878
rect 34336 27814 34388 27820
rect 34152 27532 34204 27538
rect 34152 27474 34204 27480
rect 34164 27130 34192 27474
rect 34244 27328 34296 27334
rect 34244 27270 34296 27276
rect 34152 27124 34204 27130
rect 34152 27066 34204 27072
rect 34058 27024 34114 27033
rect 34058 26959 34114 26968
rect 34072 26450 34100 26959
rect 34256 26897 34284 27270
rect 34440 27010 34468 28206
rect 34612 28154 34664 28160
rect 34520 28144 34572 28150
rect 34520 28086 34572 28092
rect 34610 28112 34666 28121
rect 34532 27130 34560 28086
rect 34610 28047 34666 28056
rect 34624 27538 34652 28047
rect 34716 27554 34744 31078
rect 34940 30492 35236 30512
rect 34996 30490 35020 30492
rect 35076 30490 35100 30492
rect 35156 30490 35180 30492
rect 35018 30438 35020 30490
rect 35082 30438 35094 30490
rect 35156 30438 35158 30490
rect 34996 30436 35020 30438
rect 35076 30436 35100 30438
rect 35156 30436 35180 30438
rect 34940 30416 35236 30436
rect 34796 29504 34848 29510
rect 34796 29446 34848 29452
rect 34808 29034 34836 29446
rect 34940 29404 35236 29424
rect 34996 29402 35020 29404
rect 35076 29402 35100 29404
rect 35156 29402 35180 29404
rect 35018 29350 35020 29402
rect 35082 29350 35094 29402
rect 35156 29350 35158 29402
rect 34996 29348 35020 29350
rect 35076 29348 35100 29350
rect 35156 29348 35180 29350
rect 34940 29328 35236 29348
rect 34796 29028 34848 29034
rect 34796 28970 34848 28976
rect 34888 28960 34940 28966
rect 34888 28902 34940 28908
rect 34900 28694 34928 28902
rect 34888 28688 34940 28694
rect 34888 28630 34940 28636
rect 34900 28506 34928 28630
rect 34808 28478 34928 28506
rect 34808 28218 34836 28478
rect 34940 28316 35236 28336
rect 34996 28314 35020 28316
rect 35076 28314 35100 28316
rect 35156 28314 35180 28316
rect 35018 28262 35020 28314
rect 35082 28262 35094 28314
rect 35156 28262 35158 28314
rect 34996 28260 35020 28262
rect 35076 28260 35100 28262
rect 35156 28260 35180 28262
rect 34940 28240 35236 28260
rect 34796 28212 34848 28218
rect 34796 28154 34848 28160
rect 34980 28008 35032 28014
rect 34980 27950 35032 27956
rect 35072 28008 35124 28014
rect 35072 27950 35124 27956
rect 34992 27878 35020 27950
rect 34980 27872 35032 27878
rect 34980 27814 35032 27820
rect 34612 27532 34664 27538
rect 34716 27526 34836 27554
rect 34612 27474 34664 27480
rect 34704 27464 34756 27470
rect 34704 27406 34756 27412
rect 34520 27124 34572 27130
rect 34520 27066 34572 27072
rect 34440 26982 34652 27010
rect 34716 26994 34744 27406
rect 34242 26888 34298 26897
rect 34624 26874 34652 26982
rect 34704 26988 34756 26994
rect 34704 26930 34756 26936
rect 34624 26846 34744 26874
rect 34242 26823 34298 26832
rect 34256 26586 34284 26823
rect 34428 26784 34480 26790
rect 34428 26726 34480 26732
rect 34244 26580 34296 26586
rect 34244 26522 34296 26528
rect 34242 26480 34298 26489
rect 34060 26444 34112 26450
rect 34242 26415 34298 26424
rect 34060 26386 34112 26392
rect 34072 26042 34100 26386
rect 34060 26036 34112 26042
rect 34060 25978 34112 25984
rect 34256 25498 34284 26415
rect 34244 25492 34296 25498
rect 34244 25434 34296 25440
rect 34060 25356 34112 25362
rect 34060 25298 34112 25304
rect 34072 24954 34100 25298
rect 34256 24954 34284 25434
rect 34336 25288 34388 25294
rect 34336 25230 34388 25236
rect 34060 24948 34112 24954
rect 34060 24890 34112 24896
rect 34244 24948 34296 24954
rect 34244 24890 34296 24896
rect 34348 24410 34376 25230
rect 34440 24750 34468 26726
rect 34612 26444 34664 26450
rect 34612 26386 34664 26392
rect 34624 26042 34652 26386
rect 34612 26036 34664 26042
rect 34612 25978 34664 25984
rect 34624 25498 34652 25978
rect 34612 25492 34664 25498
rect 34612 25434 34664 25440
rect 34520 25220 34572 25226
rect 34520 25162 34572 25168
rect 34428 24744 34480 24750
rect 34428 24686 34480 24692
rect 34336 24404 34388 24410
rect 34336 24346 34388 24352
rect 34532 24290 34560 25162
rect 34624 24818 34652 25434
rect 34612 24812 34664 24818
rect 34612 24754 34664 24760
rect 34348 24262 34560 24290
rect 34612 24268 34664 24274
rect 34244 23860 34296 23866
rect 34244 23802 34296 23808
rect 34150 23624 34206 23633
rect 34150 23559 34206 23568
rect 34164 22001 34192 23559
rect 34256 23322 34284 23802
rect 34348 23798 34376 24262
rect 34612 24210 34664 24216
rect 34428 24200 34480 24206
rect 34428 24142 34480 24148
rect 34336 23792 34388 23798
rect 34336 23734 34388 23740
rect 34336 23588 34388 23594
rect 34336 23530 34388 23536
rect 34244 23316 34296 23322
rect 34244 23258 34296 23264
rect 34348 23254 34376 23530
rect 34440 23526 34468 24142
rect 34520 24064 34572 24070
rect 34520 24006 34572 24012
rect 34428 23520 34480 23526
rect 34428 23462 34480 23468
rect 34440 23322 34468 23462
rect 34532 23322 34560 24006
rect 34624 23866 34652 24210
rect 34612 23860 34664 23866
rect 34612 23802 34664 23808
rect 34716 23361 34744 26846
rect 34702 23352 34758 23361
rect 34428 23316 34480 23322
rect 34428 23258 34480 23264
rect 34520 23316 34572 23322
rect 34572 23276 34652 23304
rect 34702 23287 34758 23296
rect 34520 23258 34572 23264
rect 34336 23248 34388 23254
rect 34336 23190 34388 23196
rect 34520 22976 34572 22982
rect 34520 22918 34572 22924
rect 34532 22522 34560 22918
rect 34256 22494 34560 22522
rect 34150 21992 34206 22001
rect 34150 21927 34206 21936
rect 34152 20936 34204 20942
rect 34152 20878 34204 20884
rect 34164 20534 34192 20878
rect 34152 20528 34204 20534
rect 34152 20470 34204 20476
rect 34256 20398 34284 22494
rect 34428 22432 34480 22438
rect 34428 22374 34480 22380
rect 34518 22400 34574 22409
rect 34336 22160 34388 22166
rect 34336 22102 34388 22108
rect 34348 20602 34376 22102
rect 34440 20942 34468 22374
rect 34518 22335 34574 22344
rect 34428 20936 34480 20942
rect 34428 20878 34480 20884
rect 34440 20602 34468 20878
rect 34336 20596 34388 20602
rect 34336 20538 34388 20544
rect 34428 20596 34480 20602
rect 34428 20538 34480 20544
rect 34244 20392 34296 20398
rect 34244 20334 34296 20340
rect 34440 19990 34468 20538
rect 34060 19984 34112 19990
rect 34428 19984 34480 19990
rect 34060 19926 34112 19932
rect 34150 19952 34206 19961
rect 34072 19514 34100 19926
rect 34428 19926 34480 19932
rect 34150 19887 34206 19896
rect 34060 19508 34112 19514
rect 34060 19450 34112 19456
rect 33966 19272 34022 19281
rect 33966 19207 34022 19216
rect 33968 19168 34020 19174
rect 33968 19110 34020 19116
rect 33874 18864 33930 18873
rect 33692 18828 33744 18834
rect 33874 18799 33876 18808
rect 33692 18770 33744 18776
rect 33928 18799 33930 18808
rect 33876 18770 33928 18776
rect 33600 18216 33652 18222
rect 33600 18158 33652 18164
rect 33416 18148 33468 18154
rect 33416 18090 33468 18096
rect 33232 18080 33284 18086
rect 33232 18022 33284 18028
rect 33244 17338 33272 18022
rect 33428 17814 33456 18090
rect 33612 17882 33640 18158
rect 33600 17876 33652 17882
rect 33600 17818 33652 17824
rect 33416 17808 33468 17814
rect 33416 17750 33468 17756
rect 33232 17332 33284 17338
rect 33232 17274 33284 17280
rect 33704 17270 33732 18770
rect 33888 18358 33916 18770
rect 33876 18352 33928 18358
rect 33876 18294 33928 18300
rect 33692 17264 33744 17270
rect 33692 17206 33744 17212
rect 33048 16176 33100 16182
rect 33048 16118 33100 16124
rect 33048 15904 33100 15910
rect 31758 15872 31814 15881
rect 33048 15846 33100 15852
rect 31758 15807 31814 15816
rect 30380 15700 30432 15706
rect 30380 15642 30432 15648
rect 31772 15502 31800 15807
rect 33060 15570 33088 15846
rect 32220 15564 32272 15570
rect 32220 15506 32272 15512
rect 33048 15564 33100 15570
rect 33048 15506 33100 15512
rect 31760 15496 31812 15502
rect 31760 15438 31812 15444
rect 31772 15162 31800 15438
rect 32232 15162 32260 15506
rect 32956 15496 33008 15502
rect 32956 15438 33008 15444
rect 32404 15360 32456 15366
rect 32404 15302 32456 15308
rect 31760 15156 31812 15162
rect 31760 15098 31812 15104
rect 32220 15156 32272 15162
rect 32220 15098 32272 15104
rect 30562 15056 30618 15065
rect 30562 14991 30564 15000
rect 30616 14991 30618 15000
rect 30564 14962 30616 14968
rect 30748 14952 30800 14958
rect 30748 14894 30800 14900
rect 30288 14476 30340 14482
rect 30288 14418 30340 14424
rect 30300 13802 30328 14418
rect 30288 13796 30340 13802
rect 30288 13738 30340 13744
rect 30300 13530 30328 13738
rect 30760 13530 30788 14894
rect 32232 14618 32260 15098
rect 32312 14952 32364 14958
rect 32312 14894 32364 14900
rect 32220 14612 32272 14618
rect 32220 14554 32272 14560
rect 32324 14278 32352 14894
rect 32312 14272 32364 14278
rect 32312 14214 32364 14220
rect 32324 13870 32352 14214
rect 32312 13864 32364 13870
rect 32312 13806 32364 13812
rect 30932 13728 30984 13734
rect 30932 13670 30984 13676
rect 32128 13728 32180 13734
rect 32128 13670 32180 13676
rect 30288 13524 30340 13530
rect 30288 13466 30340 13472
rect 30472 13524 30524 13530
rect 30472 13466 30524 13472
rect 30748 13524 30800 13530
rect 30748 13466 30800 13472
rect 30208 13394 30420 13410
rect 30208 13388 30432 13394
rect 30208 13382 30380 13388
rect 30196 12980 30248 12986
rect 30196 12922 30248 12928
rect 29932 12600 30144 12628
rect 29644 12436 29696 12442
rect 29644 12378 29696 12384
rect 29932 12322 29960 12600
rect 30208 12374 30236 12922
rect 30300 12442 30328 13382
rect 30380 13330 30432 13336
rect 30484 12918 30512 13466
rect 30656 13456 30708 13462
rect 30656 13398 30708 13404
rect 30564 13320 30616 13326
rect 30564 13262 30616 13268
rect 30576 12986 30604 13262
rect 30564 12980 30616 12986
rect 30564 12922 30616 12928
rect 30380 12912 30432 12918
rect 30380 12854 30432 12860
rect 30472 12912 30524 12918
rect 30524 12860 30604 12866
rect 30472 12854 30604 12860
rect 30392 12442 30420 12854
rect 30484 12838 30604 12854
rect 30668 12850 30696 13398
rect 30288 12436 30340 12442
rect 30288 12378 30340 12384
rect 30380 12436 30432 12442
rect 30380 12378 30432 12384
rect 30196 12368 30248 12374
rect 29000 12300 29052 12306
rect 29932 12294 30052 12322
rect 30196 12310 30248 12316
rect 29000 12242 29052 12248
rect 29012 11898 29040 12242
rect 29184 12096 29236 12102
rect 29184 12038 29236 12044
rect 29196 11898 29224 12038
rect 29000 11892 29052 11898
rect 29000 11834 29052 11840
rect 29184 11892 29236 11898
rect 29184 11834 29236 11840
rect 28724 11620 28776 11626
rect 28724 11562 28776 11568
rect 28736 11354 28764 11562
rect 28724 11348 28776 11354
rect 28724 11290 28776 11296
rect 28540 11212 28592 11218
rect 28540 11154 28592 11160
rect 28264 10804 28316 10810
rect 28264 10746 28316 10752
rect 28552 10742 28580 11154
rect 29184 11076 29236 11082
rect 29184 11018 29236 11024
rect 28540 10736 28592 10742
rect 28540 10678 28592 10684
rect 28908 10600 28960 10606
rect 29196 10554 29224 11018
rect 28960 10548 29224 10554
rect 28908 10542 29224 10548
rect 28920 10526 29224 10542
rect 29092 10124 29144 10130
rect 29092 10066 29144 10072
rect 29104 9722 29132 10066
rect 29092 9716 29144 9722
rect 29092 9658 29144 9664
rect 28724 9648 28776 9654
rect 28724 9590 28776 9596
rect 27712 9036 27764 9042
rect 27712 8978 27764 8984
rect 27724 8634 27752 8978
rect 27896 8832 27948 8838
rect 27896 8774 27948 8780
rect 27712 8628 27764 8634
rect 27712 8570 27764 8576
rect 27908 8566 27936 8774
rect 27896 8560 27948 8566
rect 27896 8502 27948 8508
rect 27528 8424 27580 8430
rect 27528 8366 27580 8372
rect 28356 8288 28408 8294
rect 28356 8230 28408 8236
rect 26884 8084 26936 8090
rect 26884 8026 26936 8032
rect 27160 8084 27212 8090
rect 27160 8026 27212 8032
rect 28368 7886 28396 8230
rect 28736 8022 28764 9590
rect 28908 9376 28960 9382
rect 28960 9324 29040 9330
rect 28908 9318 29040 9324
rect 28920 9302 29040 9318
rect 29012 8090 29040 9302
rect 29000 8084 29052 8090
rect 29000 8026 29052 8032
rect 28724 8016 28776 8022
rect 28724 7958 28776 7964
rect 28356 7880 28408 7886
rect 28356 7822 28408 7828
rect 28368 7206 28396 7822
rect 28736 7546 28764 7958
rect 28724 7540 28776 7546
rect 28724 7482 28776 7488
rect 29104 7410 29132 9658
rect 29196 8838 29224 10526
rect 29920 10464 29972 10470
rect 29920 10406 29972 10412
rect 29932 10062 29960 10406
rect 29920 10056 29972 10062
rect 29920 9998 29972 10004
rect 29828 9988 29880 9994
rect 29828 9930 29880 9936
rect 29460 9920 29512 9926
rect 29460 9862 29512 9868
rect 29472 9586 29500 9862
rect 29840 9761 29868 9930
rect 29826 9752 29882 9761
rect 29826 9687 29882 9696
rect 29460 9580 29512 9586
rect 29460 9522 29512 9528
rect 29840 9518 29868 9687
rect 29828 9512 29880 9518
rect 29828 9454 29880 9460
rect 29644 9376 29696 9382
rect 29644 9318 29696 9324
rect 29368 8968 29420 8974
rect 29368 8910 29420 8916
rect 29184 8832 29236 8838
rect 29184 8774 29236 8780
rect 29380 8498 29408 8910
rect 29368 8492 29420 8498
rect 29368 8434 29420 8440
rect 29656 7585 29684 9318
rect 29826 9208 29882 9217
rect 29932 9178 29960 9998
rect 29826 9143 29882 9152
rect 29920 9172 29972 9178
rect 29840 9110 29868 9143
rect 29920 9114 29972 9120
rect 29828 9104 29880 9110
rect 29828 9046 29880 9052
rect 29736 8628 29788 8634
rect 29840 8616 29868 9046
rect 29788 8588 29868 8616
rect 29736 8570 29788 8576
rect 29642 7576 29698 7585
rect 29642 7511 29698 7520
rect 29092 7404 29144 7410
rect 29092 7346 29144 7352
rect 27620 7200 27672 7206
rect 27540 7148 27620 7154
rect 27540 7142 27672 7148
rect 28356 7200 28408 7206
rect 28356 7142 28408 7148
rect 27540 7126 27660 7142
rect 26792 6860 26844 6866
rect 26792 6802 26844 6808
rect 26516 6792 26568 6798
rect 26516 6734 26568 6740
rect 26528 6662 26556 6734
rect 26516 6656 26568 6662
rect 26516 6598 26568 6604
rect 26528 6118 26556 6598
rect 26804 6458 26832 6802
rect 27540 6662 27568 7126
rect 27528 6656 27580 6662
rect 27528 6598 27580 6604
rect 27896 6656 27948 6662
rect 27896 6598 27948 6604
rect 29828 6656 29880 6662
rect 29828 6598 29880 6604
rect 26792 6452 26844 6458
rect 26792 6394 26844 6400
rect 27908 6322 27936 6598
rect 29840 6322 29868 6598
rect 27896 6316 27948 6322
rect 27896 6258 27948 6264
rect 28724 6316 28776 6322
rect 28724 6258 28776 6264
rect 29828 6316 29880 6322
rect 29828 6258 29880 6264
rect 26516 6112 26568 6118
rect 26516 6054 26568 6060
rect 26700 6112 26752 6118
rect 26700 6054 26752 6060
rect 26712 5710 26740 6054
rect 27908 5846 27936 6258
rect 28736 6118 28764 6258
rect 27988 6112 28040 6118
rect 27988 6054 28040 6060
rect 28724 6112 28776 6118
rect 28724 6054 28776 6060
rect 29000 6112 29052 6118
rect 29000 6054 29052 6060
rect 28000 5914 28028 6054
rect 27988 5908 28040 5914
rect 27988 5850 28040 5856
rect 27436 5840 27488 5846
rect 27436 5782 27488 5788
rect 27896 5840 27948 5846
rect 27896 5782 27948 5788
rect 26700 5704 26752 5710
rect 26700 5646 26752 5652
rect 26712 5030 26740 5646
rect 27448 5370 27476 5782
rect 27436 5364 27488 5370
rect 27436 5306 27488 5312
rect 26700 5024 26752 5030
rect 27896 5024 27948 5030
rect 26700 4966 26752 4972
rect 27342 4992 27398 5001
rect 26712 4690 26740 4966
rect 27896 4966 27948 4972
rect 27342 4927 27398 4936
rect 26700 4684 26752 4690
rect 26700 4626 26752 4632
rect 23294 4040 23350 4049
rect 23294 3975 23350 3984
rect 24214 4040 24270 4049
rect 24214 3975 24270 3984
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19580 3760 19876 3780
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 23308 480 23336 3975
rect 26792 3936 26844 3942
rect 26792 3878 26844 3884
rect 26804 3670 26832 3878
rect 27356 3738 27384 4927
rect 27618 4856 27674 4865
rect 27618 4791 27674 4800
rect 27344 3732 27396 3738
rect 27344 3674 27396 3680
rect 26792 3664 26844 3670
rect 26792 3606 26844 3612
rect 27632 2854 27660 4791
rect 27908 4214 27936 4966
rect 28000 4758 28028 5850
rect 28736 5234 28764 6054
rect 29012 5574 29040 6054
rect 29840 5846 29868 6258
rect 29828 5840 29880 5846
rect 29828 5782 29880 5788
rect 29000 5568 29052 5574
rect 28920 5528 29000 5556
rect 28920 5370 28948 5528
rect 29000 5510 29052 5516
rect 29828 5568 29880 5574
rect 29828 5510 29880 5516
rect 28908 5364 28960 5370
rect 28908 5306 28960 5312
rect 28724 5228 28776 5234
rect 28724 5170 28776 5176
rect 28736 5030 28764 5170
rect 29276 5160 29328 5166
rect 29276 5102 29328 5108
rect 28080 5024 28132 5030
rect 28080 4966 28132 4972
rect 28724 5024 28776 5030
rect 28724 4966 28776 4972
rect 28092 4826 28120 4966
rect 28080 4820 28132 4826
rect 28080 4762 28132 4768
rect 27988 4752 28040 4758
rect 27988 4694 28040 4700
rect 28000 4282 28028 4694
rect 28448 4684 28500 4690
rect 28448 4626 28500 4632
rect 27988 4276 28040 4282
rect 27988 4218 28040 4224
rect 27896 4208 27948 4214
rect 27896 4150 27948 4156
rect 27988 4140 28040 4146
rect 27988 4082 28040 4088
rect 28172 4140 28224 4146
rect 28172 4082 28224 4088
rect 28000 3942 28028 4082
rect 27988 3936 28040 3942
rect 27988 3878 28040 3884
rect 27712 3596 27764 3602
rect 27712 3538 27764 3544
rect 27724 3126 27752 3538
rect 28184 3534 28212 4082
rect 28460 3738 28488 4626
rect 28736 4593 28764 4966
rect 28722 4584 28778 4593
rect 28722 4519 28778 4528
rect 28736 4146 28764 4519
rect 29000 4480 29052 4486
rect 28920 4428 29000 4434
rect 28920 4422 29052 4428
rect 28920 4406 29040 4422
rect 28724 4140 28776 4146
rect 28724 4082 28776 4088
rect 28920 4010 28948 4406
rect 29288 4078 29316 5102
rect 29840 4729 29868 5510
rect 29826 4720 29882 4729
rect 29826 4655 29882 4664
rect 30024 4570 30052 12294
rect 30104 12300 30156 12306
rect 30104 12242 30156 12248
rect 30116 11898 30144 12242
rect 30392 11898 30420 12378
rect 30576 12345 30604 12838
rect 30656 12844 30708 12850
rect 30656 12786 30708 12792
rect 30944 12782 30972 13670
rect 30932 12776 30984 12782
rect 30932 12718 30984 12724
rect 30562 12336 30618 12345
rect 30562 12271 30618 12280
rect 30944 12238 30972 12718
rect 32140 12646 32168 13670
rect 32324 13530 32352 13806
rect 32416 13530 32444 15302
rect 32968 15162 32996 15438
rect 32956 15156 33008 15162
rect 32956 15098 33008 15104
rect 32772 14884 32824 14890
rect 32772 14826 32824 14832
rect 32784 14278 32812 14826
rect 32772 14272 32824 14278
rect 32772 14214 32824 14220
rect 32680 14068 32732 14074
rect 32680 14010 32732 14016
rect 32312 13524 32364 13530
rect 32312 13466 32364 13472
rect 32404 13524 32456 13530
rect 32404 13466 32456 13472
rect 32692 13326 32720 14010
rect 32784 13841 32812 14214
rect 32770 13832 32826 13841
rect 32770 13767 32826 13776
rect 32772 13524 32824 13530
rect 32772 13466 32824 13472
rect 32680 13320 32732 13326
rect 32680 13262 32732 13268
rect 31760 12640 31812 12646
rect 31588 12588 31760 12594
rect 31588 12582 31812 12588
rect 32128 12640 32180 12646
rect 32128 12582 32180 12588
rect 31588 12566 31800 12582
rect 30656 12232 30708 12238
rect 30656 12174 30708 12180
rect 30932 12232 30984 12238
rect 30932 12174 30984 12180
rect 30104 11892 30156 11898
rect 30104 11834 30156 11840
rect 30380 11892 30432 11898
rect 30380 11834 30432 11840
rect 30668 11830 30696 12174
rect 31484 12164 31536 12170
rect 31484 12106 31536 12112
rect 30656 11824 30708 11830
rect 30656 11766 30708 11772
rect 31496 11762 31524 12106
rect 31484 11756 31536 11762
rect 31484 11698 31536 11704
rect 31588 11694 31616 12566
rect 32692 12170 32720 13262
rect 32784 12986 32812 13466
rect 33060 12986 33088 15506
rect 33704 14634 33732 17206
rect 33784 14816 33836 14822
rect 33784 14758 33836 14764
rect 33612 14606 33732 14634
rect 33612 14414 33640 14606
rect 33796 14414 33824 14758
rect 33888 14618 33916 18294
rect 33876 14612 33928 14618
rect 33876 14554 33928 14560
rect 33600 14408 33652 14414
rect 33600 14350 33652 14356
rect 33784 14408 33836 14414
rect 33784 14350 33836 14356
rect 33232 14272 33284 14278
rect 33232 14214 33284 14220
rect 32772 12980 32824 12986
rect 32772 12922 32824 12928
rect 33048 12980 33100 12986
rect 33048 12922 33100 12928
rect 32784 12866 32812 12922
rect 32784 12838 32996 12866
rect 32680 12164 32732 12170
rect 32680 12106 32732 12112
rect 31944 12096 31996 12102
rect 31944 12038 31996 12044
rect 32772 12096 32824 12102
rect 32772 12038 32824 12044
rect 31392 11688 31444 11694
rect 31392 11630 31444 11636
rect 31576 11688 31628 11694
rect 31576 11630 31628 11636
rect 31404 11354 31432 11630
rect 31392 11348 31444 11354
rect 31392 11290 31444 11296
rect 30288 11008 30340 11014
rect 30288 10950 30340 10956
rect 30104 10804 30156 10810
rect 30104 10746 30156 10752
rect 30116 10538 30144 10746
rect 30196 10668 30248 10674
rect 30196 10610 30248 10616
rect 30104 10532 30156 10538
rect 30104 10474 30156 10480
rect 30116 10266 30144 10474
rect 30104 10260 30156 10266
rect 30104 10202 30156 10208
rect 30104 10056 30156 10062
rect 30104 9998 30156 10004
rect 30116 9722 30144 9998
rect 30104 9716 30156 9722
rect 30104 9658 30156 9664
rect 30208 9178 30236 10610
rect 30300 10470 30328 10950
rect 30288 10464 30340 10470
rect 30288 10406 30340 10412
rect 30300 10305 30328 10406
rect 30286 10296 30342 10305
rect 30286 10231 30342 10240
rect 30564 10260 30616 10266
rect 30564 10202 30616 10208
rect 30288 9716 30340 9722
rect 30288 9658 30340 9664
rect 30196 9172 30248 9178
rect 30196 9114 30248 9120
rect 30208 8362 30236 9114
rect 30300 8616 30328 9658
rect 30576 9586 30604 10202
rect 31956 9761 31984 12038
rect 32784 11801 32812 12038
rect 32770 11792 32826 11801
rect 32770 11727 32826 11736
rect 32128 11620 32180 11626
rect 32128 11562 32180 11568
rect 32140 11354 32168 11562
rect 32128 11348 32180 11354
rect 32128 11290 32180 11296
rect 32494 10296 32550 10305
rect 32494 10231 32496 10240
rect 32548 10231 32550 10240
rect 32496 10202 32548 10208
rect 31942 9752 31998 9761
rect 31942 9687 31998 9696
rect 31852 9648 31904 9654
rect 31852 9590 31904 9596
rect 30564 9580 30616 9586
rect 30564 9522 30616 9528
rect 31864 8634 31892 9590
rect 31956 8974 31984 9687
rect 32508 9518 32536 10202
rect 32496 9512 32548 9518
rect 32416 9460 32496 9466
rect 32416 9454 32548 9460
rect 32416 9438 32536 9454
rect 31944 8968 31996 8974
rect 31944 8910 31996 8916
rect 30380 8628 30432 8634
rect 30300 8588 30380 8616
rect 30380 8570 30432 8576
rect 31852 8628 31904 8634
rect 31852 8570 31904 8576
rect 30196 8356 30248 8362
rect 30196 8298 30248 8304
rect 30380 8356 30432 8362
rect 30380 8298 30432 8304
rect 30392 8090 30420 8298
rect 31760 8288 31812 8294
rect 31760 8230 31812 8236
rect 31772 8090 31800 8230
rect 30380 8084 30432 8090
rect 30380 8026 30432 8032
rect 31760 8084 31812 8090
rect 31760 8026 31812 8032
rect 31208 7268 31260 7274
rect 31208 7210 31260 7216
rect 30288 6860 30340 6866
rect 30288 6802 30340 6808
rect 30300 6390 30328 6802
rect 31220 6746 31248 7210
rect 31300 7200 31352 7206
rect 31300 7142 31352 7148
rect 31312 6934 31340 7142
rect 31300 6928 31352 6934
rect 31300 6870 31352 6876
rect 31864 6866 31892 8570
rect 31956 8022 31984 8910
rect 32036 8832 32088 8838
rect 32036 8774 32088 8780
rect 32048 8430 32076 8774
rect 32036 8424 32088 8430
rect 32036 8366 32088 8372
rect 31944 8016 31996 8022
rect 31944 7958 31996 7964
rect 32128 7948 32180 7954
rect 32128 7890 32180 7896
rect 32036 7880 32088 7886
rect 32036 7822 32088 7828
rect 32048 7546 32076 7822
rect 32036 7540 32088 7546
rect 32036 7482 32088 7488
rect 32048 7342 32076 7482
rect 32036 7336 32088 7342
rect 32036 7278 32088 7284
rect 32140 7002 32168 7890
rect 32416 7546 32444 9438
rect 32496 9376 32548 9382
rect 32496 9318 32548 9324
rect 32508 8634 32536 9318
rect 32968 9178 32996 12838
rect 33140 12708 33192 12714
rect 33140 12650 33192 12656
rect 33152 12442 33180 12650
rect 33140 12436 33192 12442
rect 33140 12378 33192 12384
rect 33140 12300 33192 12306
rect 33140 12242 33192 12248
rect 33152 11762 33180 12242
rect 33244 12238 33272 14214
rect 33612 14074 33640 14350
rect 33600 14068 33652 14074
rect 33600 14010 33652 14016
rect 33796 13938 33824 14350
rect 33888 14074 33916 14554
rect 33876 14068 33928 14074
rect 33876 14010 33928 14016
rect 33784 13932 33836 13938
rect 33784 13874 33836 13880
rect 33782 13832 33838 13841
rect 33782 13767 33838 13776
rect 33692 13728 33744 13734
rect 33692 13670 33744 13676
rect 33416 13320 33468 13326
rect 33416 13262 33468 13268
rect 33428 12714 33456 13262
rect 33416 12708 33468 12714
rect 33416 12650 33468 12656
rect 33600 12640 33652 12646
rect 33600 12582 33652 12588
rect 33324 12436 33376 12442
rect 33324 12378 33376 12384
rect 33232 12232 33284 12238
rect 33232 12174 33284 12180
rect 33244 11898 33272 12174
rect 33232 11892 33284 11898
rect 33232 11834 33284 11840
rect 33140 11756 33192 11762
rect 33140 11698 33192 11704
rect 33140 10192 33192 10198
rect 33140 10134 33192 10140
rect 33048 10124 33100 10130
rect 33048 10066 33100 10072
rect 33060 9722 33088 10066
rect 33048 9716 33100 9722
rect 33048 9658 33100 9664
rect 33152 9450 33180 10134
rect 33336 9466 33364 12378
rect 33612 12306 33640 12582
rect 33600 12300 33652 12306
rect 33600 12242 33652 12248
rect 33704 12238 33732 13670
rect 33796 12850 33824 13767
rect 33888 13530 33916 14010
rect 33876 13524 33928 13530
rect 33876 13466 33928 13472
rect 33876 12912 33928 12918
rect 33876 12854 33928 12860
rect 33784 12844 33836 12850
rect 33784 12786 33836 12792
rect 33796 12646 33824 12786
rect 33784 12640 33836 12646
rect 33784 12582 33836 12588
rect 33888 12306 33916 12854
rect 33980 12617 34008 19110
rect 34060 18760 34112 18766
rect 34060 18702 34112 18708
rect 34072 17882 34100 18702
rect 34060 17876 34112 17882
rect 34060 17818 34112 17824
rect 34060 17672 34112 17678
rect 34060 17614 34112 17620
rect 34072 17338 34100 17614
rect 34060 17332 34112 17338
rect 34060 17274 34112 17280
rect 34164 15065 34192 19887
rect 34244 19848 34296 19854
rect 34244 19790 34296 19796
rect 34256 19242 34284 19790
rect 34244 19236 34296 19242
rect 34244 19178 34296 19184
rect 34256 18970 34284 19178
rect 34244 18964 34296 18970
rect 34244 18906 34296 18912
rect 34336 18760 34388 18766
rect 34336 18702 34388 18708
rect 34348 18222 34376 18702
rect 34336 18216 34388 18222
rect 34336 18158 34388 18164
rect 34426 18048 34482 18057
rect 34426 17983 34482 17992
rect 34244 17604 34296 17610
rect 34244 17546 34296 17552
rect 34150 15056 34206 15065
rect 34150 14991 34206 15000
rect 34256 13258 34284 17546
rect 34440 17490 34468 17983
rect 34532 17610 34560 22335
rect 34624 22234 34652 23276
rect 34704 23180 34756 23186
rect 34704 23122 34756 23128
rect 34716 22778 34744 23122
rect 34704 22772 34756 22778
rect 34704 22714 34756 22720
rect 34702 22264 34758 22273
rect 34612 22228 34664 22234
rect 34702 22199 34758 22208
rect 34612 22170 34664 22176
rect 34612 22024 34664 22030
rect 34612 21966 34664 21972
rect 34624 21486 34652 21966
rect 34612 21480 34664 21486
rect 34612 21422 34664 21428
rect 34612 20936 34664 20942
rect 34612 20878 34664 20884
rect 34624 20330 34652 20878
rect 34612 20324 34664 20330
rect 34612 20266 34664 20272
rect 34624 19786 34652 20266
rect 34612 19780 34664 19786
rect 34612 19722 34664 19728
rect 34610 18728 34666 18737
rect 34610 18663 34666 18672
rect 34520 17604 34572 17610
rect 34520 17546 34572 17552
rect 34440 17462 34560 17490
rect 34532 15450 34560 17462
rect 34624 16289 34652 18663
rect 34610 16280 34666 16289
rect 34610 16215 34666 16224
rect 34612 16176 34664 16182
rect 34612 16118 34664 16124
rect 34348 15422 34560 15450
rect 34244 13252 34296 13258
rect 34244 13194 34296 13200
rect 34348 12850 34376 15422
rect 34520 15360 34572 15366
rect 34520 15302 34572 15308
rect 34428 14476 34480 14482
rect 34428 14418 34480 14424
rect 34440 13530 34468 14418
rect 34428 13524 34480 13530
rect 34428 13466 34480 13472
rect 34336 12844 34388 12850
rect 34336 12786 34388 12792
rect 34532 12730 34560 15302
rect 34624 14618 34652 16118
rect 34612 14612 34664 14618
rect 34612 14554 34664 14560
rect 34072 12702 34560 12730
rect 33966 12608 34022 12617
rect 33966 12543 34022 12552
rect 33876 12300 33928 12306
rect 33876 12242 33928 12248
rect 33692 12232 33744 12238
rect 33692 12174 33744 12180
rect 33704 12102 33732 12174
rect 33692 12096 33744 12102
rect 33692 12038 33744 12044
rect 33704 11898 33732 12038
rect 33888 11898 33916 12242
rect 34072 12209 34100 12702
rect 34152 12640 34204 12646
rect 34428 12640 34480 12646
rect 34334 12608 34390 12617
rect 34204 12588 34284 12594
rect 34152 12582 34284 12588
rect 34164 12566 34284 12582
rect 34256 12442 34284 12566
rect 34428 12582 34480 12588
rect 34520 12640 34572 12646
rect 34520 12582 34572 12588
rect 34334 12543 34390 12552
rect 34348 12442 34376 12543
rect 34244 12436 34296 12442
rect 34244 12378 34296 12384
rect 34336 12436 34388 12442
rect 34336 12378 34388 12384
rect 34440 12322 34468 12582
rect 34256 12294 34468 12322
rect 34058 12200 34114 12209
rect 34058 12135 34114 12144
rect 33692 11892 33744 11898
rect 33692 11834 33744 11840
rect 33876 11892 33928 11898
rect 33876 11834 33928 11840
rect 33888 11218 33916 11834
rect 33876 11212 33928 11218
rect 33876 11154 33928 11160
rect 33888 10198 33916 11154
rect 33876 10192 33928 10198
rect 33876 10134 33928 10140
rect 33508 10124 33560 10130
rect 33508 10066 33560 10072
rect 33520 9586 33548 10066
rect 33508 9580 33560 9586
rect 33508 9522 33560 9528
rect 33140 9444 33192 9450
rect 33140 9386 33192 9392
rect 33244 9438 33364 9466
rect 32956 9172 33008 9178
rect 32956 9114 33008 9120
rect 32864 8832 32916 8838
rect 32864 8774 32916 8780
rect 32496 8628 32548 8634
rect 32496 8570 32548 8576
rect 32876 8362 32904 8774
rect 32864 8356 32916 8362
rect 32864 8298 32916 8304
rect 32404 7540 32456 7546
rect 32404 7482 32456 7488
rect 32876 7449 32904 8298
rect 32968 8022 32996 9114
rect 33048 8968 33100 8974
rect 33048 8910 33100 8916
rect 33060 8090 33088 8910
rect 33152 8430 33180 9386
rect 33140 8424 33192 8430
rect 33140 8366 33192 8372
rect 33048 8084 33100 8090
rect 33048 8026 33100 8032
rect 32956 8016 33008 8022
rect 32956 7958 33008 7964
rect 32968 7585 32996 7958
rect 33152 7954 33180 8366
rect 33140 7948 33192 7954
rect 33140 7890 33192 7896
rect 32954 7576 33010 7585
rect 33152 7546 33180 7890
rect 32954 7511 33010 7520
rect 33140 7540 33192 7546
rect 33140 7482 33192 7488
rect 32862 7440 32918 7449
rect 32862 7375 32864 7384
rect 32916 7375 32918 7384
rect 32864 7346 32916 7352
rect 32680 7268 32732 7274
rect 32680 7210 32732 7216
rect 32692 7002 32720 7210
rect 32128 6996 32180 7002
rect 32128 6938 32180 6944
rect 32680 6996 32732 7002
rect 32680 6938 32732 6944
rect 31852 6860 31904 6866
rect 31852 6802 31904 6808
rect 31944 6860 31996 6866
rect 31944 6802 31996 6808
rect 31220 6718 31340 6746
rect 30840 6656 30892 6662
rect 30840 6598 30892 6604
rect 30852 6458 30880 6598
rect 30840 6452 30892 6458
rect 30840 6394 30892 6400
rect 30288 6384 30340 6390
rect 30288 6326 30340 6332
rect 31312 6118 31340 6718
rect 31392 6656 31444 6662
rect 31392 6598 31444 6604
rect 31404 6322 31432 6598
rect 31392 6316 31444 6322
rect 31392 6258 31444 6264
rect 31864 6186 31892 6802
rect 31852 6180 31904 6186
rect 31852 6122 31904 6128
rect 31116 6112 31168 6118
rect 31116 6054 31168 6060
rect 31300 6112 31352 6118
rect 31300 6054 31352 6060
rect 31668 6112 31720 6118
rect 31668 6054 31720 6060
rect 30288 5840 30340 5846
rect 30288 5782 30340 5788
rect 30196 5772 30248 5778
rect 30196 5714 30248 5720
rect 30104 5704 30156 5710
rect 30104 5646 30156 5652
rect 29748 4542 30052 4570
rect 29000 4072 29052 4078
rect 29000 4014 29052 4020
rect 29276 4072 29328 4078
rect 29276 4014 29328 4020
rect 28908 4004 28960 4010
rect 28908 3946 28960 3952
rect 28448 3732 28500 3738
rect 28448 3674 28500 3680
rect 29012 3670 29040 4014
rect 29288 3738 29316 4014
rect 29368 3936 29420 3942
rect 29368 3878 29420 3884
rect 29380 3738 29408 3878
rect 29276 3732 29328 3738
rect 29276 3674 29328 3680
rect 29368 3732 29420 3738
rect 29368 3674 29420 3680
rect 29000 3664 29052 3670
rect 29000 3606 29052 3612
rect 27804 3528 27856 3534
rect 27804 3470 27856 3476
rect 28172 3528 28224 3534
rect 28172 3470 28224 3476
rect 27816 3233 27844 3470
rect 27802 3224 27858 3233
rect 27802 3159 27804 3168
rect 27856 3159 27858 3168
rect 27804 3130 27856 3136
rect 27712 3120 27764 3126
rect 27816 3099 27844 3130
rect 27712 3062 27764 3068
rect 28078 3088 28134 3097
rect 27724 2961 27752 3062
rect 28184 3058 28212 3470
rect 29012 3194 29040 3606
rect 29000 3188 29052 3194
rect 29000 3130 29052 3136
rect 28078 3023 28080 3032
rect 28132 3023 28134 3032
rect 28172 3052 28224 3058
rect 28080 2994 28132 3000
rect 28172 2994 28224 3000
rect 27710 2952 27766 2961
rect 27710 2887 27766 2896
rect 28000 2854 28028 2885
rect 27620 2848 27672 2854
rect 27988 2848 28040 2854
rect 27620 2790 27672 2796
rect 27986 2816 27988 2825
rect 28040 2816 28042 2825
rect 27986 2751 28042 2760
rect 28000 2650 28028 2751
rect 28184 2650 28212 2994
rect 29288 2990 29316 3674
rect 29276 2984 29328 2990
rect 29276 2926 29328 2932
rect 27988 2644 28040 2650
rect 27988 2586 28040 2592
rect 28172 2644 28224 2650
rect 28172 2586 28224 2592
rect 29288 2514 29316 2926
rect 29380 2922 29408 3674
rect 29368 2916 29420 2922
rect 29368 2858 29420 2864
rect 29380 2650 29408 2858
rect 29368 2644 29420 2650
rect 29368 2586 29420 2592
rect 29276 2508 29328 2514
rect 29276 2450 29328 2456
rect 29748 626 29776 4542
rect 30116 4486 30144 5646
rect 30208 4826 30236 5714
rect 30300 5386 30328 5782
rect 31128 5642 31156 6054
rect 31312 5846 31340 6054
rect 31680 5914 31708 6054
rect 31668 5908 31720 5914
rect 31668 5850 31720 5856
rect 31300 5840 31352 5846
rect 31300 5782 31352 5788
rect 31116 5636 31168 5642
rect 31116 5578 31168 5584
rect 30300 5370 30420 5386
rect 30300 5364 30432 5370
rect 30300 5358 30380 5364
rect 30380 5306 30432 5312
rect 30380 5024 30432 5030
rect 30300 4972 30380 4978
rect 30300 4966 30432 4972
rect 30300 4950 30420 4966
rect 30196 4820 30248 4826
rect 30196 4762 30248 4768
rect 30104 4480 30156 4486
rect 30104 4422 30156 4428
rect 30300 4078 30328 4950
rect 30748 4684 30800 4690
rect 30748 4626 30800 4632
rect 30760 4078 30788 4626
rect 31024 4616 31076 4622
rect 31022 4584 31024 4593
rect 31076 4584 31078 4593
rect 31022 4519 31078 4528
rect 30288 4072 30340 4078
rect 30288 4014 30340 4020
rect 30748 4072 30800 4078
rect 30748 4014 30800 4020
rect 30656 3936 30708 3942
rect 30656 3878 30708 3884
rect 30668 3670 30696 3878
rect 30656 3664 30708 3670
rect 30656 3606 30708 3612
rect 30760 3398 30788 4014
rect 31036 3738 31064 4519
rect 31128 4146 31156 5578
rect 31680 5556 31708 5850
rect 31956 5846 31984 6802
rect 32140 6254 32168 6938
rect 32772 6928 32824 6934
rect 32772 6870 32824 6876
rect 32404 6724 32456 6730
rect 32404 6666 32456 6672
rect 32416 6458 32444 6666
rect 32784 6458 32812 6870
rect 32404 6452 32456 6458
rect 32404 6394 32456 6400
rect 32772 6452 32824 6458
rect 32772 6394 32824 6400
rect 32128 6248 32180 6254
rect 32128 6190 32180 6196
rect 33140 6248 33192 6254
rect 33140 6190 33192 6196
rect 32956 6112 33008 6118
rect 32402 6080 32458 6089
rect 32956 6054 33008 6060
rect 32402 6015 32458 6024
rect 31944 5840 31996 5846
rect 31944 5782 31996 5788
rect 31680 5528 31800 5556
rect 31772 4826 31800 5528
rect 32416 5370 32444 6015
rect 32968 5846 32996 6054
rect 32956 5840 33008 5846
rect 32956 5782 33008 5788
rect 33152 5642 33180 6190
rect 33140 5636 33192 5642
rect 33140 5578 33192 5584
rect 32772 5568 32824 5574
rect 32772 5510 32824 5516
rect 32404 5364 32456 5370
rect 32404 5306 32456 5312
rect 32784 5030 32812 5510
rect 33048 5228 33100 5234
rect 33048 5170 33100 5176
rect 32220 5024 32272 5030
rect 32218 4992 32220 5001
rect 32772 5024 32824 5030
rect 32272 4992 32274 5001
rect 32772 4966 32824 4972
rect 32218 4927 32274 4936
rect 32784 4865 32812 4966
rect 32770 4856 32826 4865
rect 31760 4820 31812 4826
rect 32770 4791 32826 4800
rect 31760 4762 31812 4768
rect 32126 4720 32182 4729
rect 31208 4684 31260 4690
rect 32126 4655 32128 4664
rect 31208 4626 31260 4632
rect 32180 4655 32182 4664
rect 32128 4626 32180 4632
rect 31116 4140 31168 4146
rect 31116 4082 31168 4088
rect 31220 4010 31248 4626
rect 33060 4622 33088 5170
rect 33048 4616 33100 4622
rect 33048 4558 33100 4564
rect 31760 4072 31812 4078
rect 33244 4026 33272 9438
rect 33324 9376 33376 9382
rect 33324 9318 33376 9324
rect 33336 8974 33364 9318
rect 33324 8968 33376 8974
rect 33324 8910 33376 8916
rect 33336 8090 33364 8910
rect 33520 8566 33548 9522
rect 34256 9178 34284 12294
rect 34336 12096 34388 12102
rect 34336 12038 34388 12044
rect 34348 11898 34376 12038
rect 34336 11892 34388 11898
rect 34336 11834 34388 11840
rect 34532 10554 34560 12582
rect 34612 12300 34664 12306
rect 34612 12242 34664 12248
rect 34624 12102 34652 12242
rect 34612 12096 34664 12102
rect 34612 12038 34664 12044
rect 34612 11892 34664 11898
rect 34612 11834 34664 11840
rect 34440 10526 34560 10554
rect 34244 9172 34296 9178
rect 34244 9114 34296 9120
rect 33508 8560 33560 8566
rect 33508 8502 33560 8508
rect 34440 8514 34468 10526
rect 34520 10464 34572 10470
rect 34520 10406 34572 10412
rect 34532 8634 34560 10406
rect 34520 8628 34572 8634
rect 34520 8570 34572 8576
rect 34440 8486 34560 8514
rect 33324 8084 33376 8090
rect 33324 8026 33376 8032
rect 33324 7948 33376 7954
rect 33324 7890 33376 7896
rect 33336 7342 33364 7890
rect 33324 7336 33376 7342
rect 33324 7278 33376 7284
rect 33336 6934 33364 7278
rect 33324 6928 33376 6934
rect 33324 6870 33376 6876
rect 34244 6860 34296 6866
rect 34244 6802 34296 6808
rect 33784 6656 33836 6662
rect 33784 6598 33836 6604
rect 33796 6361 33824 6598
rect 34256 6390 34284 6802
rect 34532 6644 34560 8486
rect 34624 8378 34652 11834
rect 34716 8566 34744 22199
rect 34808 13734 34836 27526
rect 34992 27470 35020 27814
rect 35084 27674 35112 27950
rect 35072 27668 35124 27674
rect 35072 27610 35124 27616
rect 34980 27464 35032 27470
rect 34980 27406 35032 27412
rect 34940 27228 35236 27248
rect 34996 27226 35020 27228
rect 35076 27226 35100 27228
rect 35156 27226 35180 27228
rect 35018 27174 35020 27226
rect 35082 27174 35094 27226
rect 35156 27174 35158 27226
rect 34996 27172 35020 27174
rect 35076 27172 35100 27174
rect 35156 27172 35180 27174
rect 34940 27152 35236 27172
rect 34980 26852 35032 26858
rect 34980 26794 35032 26800
rect 34992 26586 35020 26794
rect 35268 26625 35296 34478
rect 35360 34406 35388 35090
rect 35348 34400 35400 34406
rect 35348 34342 35400 34348
rect 35348 33312 35400 33318
rect 35348 33254 35400 33260
rect 35360 30326 35388 33254
rect 35440 31884 35492 31890
rect 35440 31826 35492 31832
rect 35452 31142 35480 31826
rect 35440 31136 35492 31142
rect 35440 31078 35492 31084
rect 35544 30954 35572 35142
rect 35622 34640 35678 34649
rect 35622 34575 35678 34584
rect 35636 34202 35664 34575
rect 35624 34196 35676 34202
rect 35624 34138 35676 34144
rect 35728 33658 35756 35391
rect 35820 34746 35848 36887
rect 36096 35873 36124 39520
rect 36726 38176 36782 38185
rect 36726 38111 36782 38120
rect 36082 35864 36138 35873
rect 36082 35799 36138 35808
rect 36740 34746 36768 38111
rect 37200 35601 37228 39520
rect 37186 35592 37242 35601
rect 37186 35527 37242 35536
rect 38304 35329 38332 39520
rect 38290 35320 38346 35329
rect 38290 35255 38346 35264
rect 35808 34740 35860 34746
rect 35808 34682 35860 34688
rect 36728 34740 36780 34746
rect 36728 34682 36780 34688
rect 39408 34649 39436 39520
rect 39394 34640 39450 34649
rect 39394 34575 39450 34584
rect 37096 34536 37148 34542
rect 35806 34504 35862 34513
rect 37096 34478 37148 34484
rect 35806 34439 35862 34448
rect 35716 33652 35768 33658
rect 35716 33594 35768 33600
rect 35622 33280 35678 33289
rect 35622 33215 35678 33224
rect 35452 30926 35572 30954
rect 35636 30938 35664 33215
rect 35714 32056 35770 32065
rect 35820 32026 35848 34439
rect 35900 34060 35952 34066
rect 35900 34002 35952 34008
rect 35912 33318 35940 34002
rect 35900 33312 35952 33318
rect 35900 33254 35952 33260
rect 35714 31991 35770 32000
rect 35808 32020 35860 32026
rect 35624 30932 35676 30938
rect 35348 30320 35400 30326
rect 35348 30262 35400 30268
rect 35348 30184 35400 30190
rect 35348 30126 35400 30132
rect 35360 27441 35388 30126
rect 35346 27432 35402 27441
rect 35346 27367 35402 27376
rect 35254 26616 35310 26625
rect 34980 26580 35032 26586
rect 35254 26551 35310 26560
rect 34980 26522 35032 26528
rect 35256 26444 35308 26450
rect 35256 26386 35308 26392
rect 34940 26140 35236 26160
rect 34996 26138 35020 26140
rect 35076 26138 35100 26140
rect 35156 26138 35180 26140
rect 35018 26086 35020 26138
rect 35082 26086 35094 26138
rect 35156 26086 35158 26138
rect 34996 26084 35020 26086
rect 35076 26084 35100 26086
rect 35156 26084 35180 26086
rect 34940 26064 35236 26084
rect 35268 25498 35296 26386
rect 35256 25492 35308 25498
rect 35256 25434 35308 25440
rect 34940 25052 35236 25072
rect 34996 25050 35020 25052
rect 35076 25050 35100 25052
rect 35156 25050 35180 25052
rect 35018 24998 35020 25050
rect 35082 24998 35094 25050
rect 35156 24998 35158 25050
rect 34996 24996 35020 24998
rect 35076 24996 35100 24998
rect 35156 24996 35180 24998
rect 34940 24976 35236 24996
rect 35164 24608 35216 24614
rect 35164 24550 35216 24556
rect 35176 24206 35204 24550
rect 35164 24200 35216 24206
rect 35216 24148 35296 24154
rect 35164 24142 35296 24148
rect 35176 24126 35296 24142
rect 34940 23964 35236 23984
rect 34996 23962 35020 23964
rect 35076 23962 35100 23964
rect 35156 23962 35180 23964
rect 35018 23910 35020 23962
rect 35082 23910 35094 23962
rect 35156 23910 35158 23962
rect 34996 23908 35020 23910
rect 35076 23908 35100 23910
rect 35156 23908 35180 23910
rect 34940 23888 35236 23908
rect 35268 23594 35296 24126
rect 35256 23588 35308 23594
rect 35256 23530 35308 23536
rect 35256 23112 35308 23118
rect 35256 23054 35308 23060
rect 34940 22876 35236 22896
rect 34996 22874 35020 22876
rect 35076 22874 35100 22876
rect 35156 22874 35180 22876
rect 35018 22822 35020 22874
rect 35082 22822 35094 22874
rect 35156 22822 35158 22874
rect 34996 22820 35020 22822
rect 35076 22820 35100 22822
rect 35156 22820 35180 22822
rect 34940 22800 35236 22820
rect 35164 22432 35216 22438
rect 35164 22374 35216 22380
rect 35176 22234 35204 22374
rect 35164 22228 35216 22234
rect 35164 22170 35216 22176
rect 35268 22166 35296 23054
rect 35452 22778 35480 30926
rect 35624 30874 35676 30880
rect 35622 30832 35678 30841
rect 35532 30796 35584 30802
rect 35622 30767 35678 30776
rect 35532 30738 35584 30744
rect 35544 30054 35572 30738
rect 35532 30048 35584 30054
rect 35532 29990 35584 29996
rect 35544 29730 35572 29990
rect 35636 29850 35664 30767
rect 35728 30326 35756 31991
rect 35808 31962 35860 31968
rect 35912 31906 35940 33254
rect 35820 31878 35940 31906
rect 35716 30320 35768 30326
rect 35716 30262 35768 30268
rect 35624 29844 35676 29850
rect 35624 29786 35676 29792
rect 35544 29702 35664 29730
rect 35532 27328 35584 27334
rect 35532 27270 35584 27276
rect 35544 26625 35572 27270
rect 35530 26616 35586 26625
rect 35530 26551 35586 26560
rect 35544 26518 35572 26551
rect 35532 26512 35584 26518
rect 35532 26454 35584 26460
rect 35532 26240 35584 26246
rect 35532 26182 35584 26188
rect 35544 25838 35572 26182
rect 35532 25832 35584 25838
rect 35532 25774 35584 25780
rect 35544 24682 35572 25774
rect 35532 24676 35584 24682
rect 35532 24618 35584 24624
rect 35530 24576 35586 24585
rect 35530 24511 35586 24520
rect 35544 23497 35572 24511
rect 35530 23488 35586 23497
rect 35530 23423 35586 23432
rect 35532 22976 35584 22982
rect 35532 22918 35584 22924
rect 35440 22772 35492 22778
rect 35440 22714 35492 22720
rect 35256 22160 35308 22166
rect 35256 22102 35308 22108
rect 34940 21788 35236 21808
rect 34996 21786 35020 21788
rect 35076 21786 35100 21788
rect 35156 21786 35180 21788
rect 35018 21734 35020 21786
rect 35082 21734 35094 21786
rect 35156 21734 35158 21786
rect 34996 21732 35020 21734
rect 35076 21732 35100 21734
rect 35156 21732 35180 21734
rect 34940 21712 35236 21732
rect 35268 21690 35296 22102
rect 35348 21888 35400 21894
rect 35348 21830 35400 21836
rect 35256 21684 35308 21690
rect 35256 21626 35308 21632
rect 34888 21480 34940 21486
rect 34888 21422 34940 21428
rect 34900 20942 34928 21422
rect 34888 20936 34940 20942
rect 34888 20878 34940 20884
rect 35360 20806 35388 21830
rect 35348 20800 35400 20806
rect 35348 20742 35400 20748
rect 34940 20700 35236 20720
rect 34996 20698 35020 20700
rect 35076 20698 35100 20700
rect 35156 20698 35180 20700
rect 35018 20646 35020 20698
rect 35082 20646 35094 20698
rect 35156 20646 35158 20698
rect 34996 20644 35020 20646
rect 35076 20644 35100 20646
rect 35156 20644 35180 20646
rect 34940 20624 35236 20644
rect 35072 20392 35124 20398
rect 35360 20369 35388 20742
rect 35072 20334 35124 20340
rect 35346 20360 35402 20369
rect 35084 19990 35112 20334
rect 35346 20295 35402 20304
rect 35072 19984 35124 19990
rect 35072 19926 35124 19932
rect 35346 19816 35402 19825
rect 35256 19780 35308 19786
rect 35346 19751 35402 19760
rect 35256 19722 35308 19728
rect 34940 19612 35236 19632
rect 34996 19610 35020 19612
rect 35076 19610 35100 19612
rect 35156 19610 35180 19612
rect 35018 19558 35020 19610
rect 35082 19558 35094 19610
rect 35156 19558 35158 19610
rect 34996 19556 35020 19558
rect 35076 19556 35100 19558
rect 35156 19556 35180 19558
rect 34940 19536 35236 19556
rect 35268 18970 35296 19722
rect 35360 19718 35388 19751
rect 35348 19712 35400 19718
rect 35348 19654 35400 19660
rect 35256 18964 35308 18970
rect 35256 18906 35308 18912
rect 34940 18524 35236 18544
rect 34996 18522 35020 18524
rect 35076 18522 35100 18524
rect 35156 18522 35180 18524
rect 35018 18470 35020 18522
rect 35082 18470 35094 18522
rect 35156 18470 35158 18522
rect 34996 18468 35020 18470
rect 35076 18468 35100 18470
rect 35156 18468 35180 18470
rect 34940 18448 35236 18468
rect 35360 17814 35388 19654
rect 35348 17808 35400 17814
rect 35348 17750 35400 17756
rect 35256 17740 35308 17746
rect 35256 17682 35308 17688
rect 34940 17436 35236 17456
rect 34996 17434 35020 17436
rect 35076 17434 35100 17436
rect 35156 17434 35180 17436
rect 35018 17382 35020 17434
rect 35082 17382 35094 17434
rect 35156 17382 35158 17434
rect 34996 17380 35020 17382
rect 35076 17380 35100 17382
rect 35156 17380 35180 17382
rect 34940 17360 35236 17380
rect 35268 17338 35296 17682
rect 35348 17672 35400 17678
rect 35348 17614 35400 17620
rect 35256 17332 35308 17338
rect 35256 17274 35308 17280
rect 35360 16998 35388 17614
rect 35348 16992 35400 16998
rect 35348 16934 35400 16940
rect 35452 16590 35480 22714
rect 35544 22574 35572 22918
rect 35532 22568 35584 22574
rect 35532 22510 35584 22516
rect 35530 22400 35586 22409
rect 35530 22335 35586 22344
rect 35544 20505 35572 22335
rect 35636 22166 35664 29702
rect 35714 29608 35770 29617
rect 35714 29543 35770 29552
rect 35728 26042 35756 29543
rect 35716 26036 35768 26042
rect 35716 25978 35768 25984
rect 35728 25770 35756 25978
rect 35716 25764 35768 25770
rect 35716 25706 35768 25712
rect 35716 25220 35768 25226
rect 35716 25162 35768 25168
rect 35728 24138 35756 25162
rect 35716 24132 35768 24138
rect 35716 24074 35768 24080
rect 35820 22166 35848 31878
rect 35992 28416 36044 28422
rect 35992 28358 36044 28364
rect 36004 28014 36032 28358
rect 35992 28008 36044 28014
rect 35992 27950 36044 27956
rect 36360 27872 36412 27878
rect 36360 27814 36412 27820
rect 36372 27538 36400 27814
rect 36360 27532 36412 27538
rect 36360 27474 36412 27480
rect 36372 27130 36400 27474
rect 36820 27328 36872 27334
rect 36820 27270 36872 27276
rect 36360 27124 36412 27130
rect 36360 27066 36412 27072
rect 36372 26926 36400 27066
rect 36360 26920 36412 26926
rect 36360 26862 36412 26868
rect 36832 26790 36860 27270
rect 37004 26988 37056 26994
rect 37004 26930 37056 26936
rect 37016 26897 37044 26930
rect 37002 26888 37058 26897
rect 37002 26823 37058 26832
rect 36820 26784 36872 26790
rect 36820 26726 36872 26732
rect 36832 26450 36860 26726
rect 37016 26586 37044 26823
rect 37004 26580 37056 26586
rect 37004 26522 37056 26528
rect 36820 26444 36872 26450
rect 36820 26386 36872 26392
rect 36910 26072 36966 26081
rect 36910 26007 36966 26016
rect 36820 25696 36872 25702
rect 36820 25638 36872 25644
rect 35900 25356 35952 25362
rect 35900 25298 35952 25304
rect 35912 24342 35940 25298
rect 36832 25294 36860 25638
rect 36820 25288 36872 25294
rect 36820 25230 36872 25236
rect 36832 24954 36860 25230
rect 36820 24948 36872 24954
rect 36820 24890 36872 24896
rect 35900 24336 35952 24342
rect 35900 24278 35952 24284
rect 36924 24274 36952 26007
rect 36912 24268 36964 24274
rect 36912 24210 36964 24216
rect 36924 23866 36952 24210
rect 36912 23860 36964 23866
rect 36912 23802 36964 23808
rect 36544 23656 36596 23662
rect 36544 23598 36596 23604
rect 35900 23588 35952 23594
rect 35900 23530 35952 23536
rect 35912 23322 35940 23530
rect 36268 23520 36320 23526
rect 36268 23462 36320 23468
rect 35900 23316 35952 23322
rect 35900 23258 35952 23264
rect 36280 23118 36308 23462
rect 36268 23112 36320 23118
rect 36268 23054 36320 23060
rect 36280 22778 36308 23054
rect 36556 22982 36584 23598
rect 36544 22976 36596 22982
rect 36544 22918 36596 22924
rect 36268 22772 36320 22778
rect 36268 22714 36320 22720
rect 36084 22636 36136 22642
rect 36084 22578 36136 22584
rect 35900 22568 35952 22574
rect 35900 22510 35952 22516
rect 35624 22160 35676 22166
rect 35624 22102 35676 22108
rect 35808 22160 35860 22166
rect 35808 22102 35860 22108
rect 35716 22092 35768 22098
rect 35716 22034 35768 22040
rect 35622 21176 35678 21185
rect 35622 21111 35678 21120
rect 35530 20496 35586 20505
rect 35530 20431 35586 20440
rect 35636 20097 35664 21111
rect 35622 20088 35678 20097
rect 35622 20023 35678 20032
rect 35728 19972 35756 22034
rect 35808 21684 35860 21690
rect 35808 21626 35860 21632
rect 35820 20398 35848 21626
rect 35912 21146 35940 22510
rect 35992 21888 36044 21894
rect 35992 21830 36044 21836
rect 36004 21486 36032 21830
rect 36096 21690 36124 22578
rect 36176 22160 36228 22166
rect 36176 22102 36228 22108
rect 36188 21962 36216 22102
rect 36176 21956 36228 21962
rect 36176 21898 36228 21904
rect 36084 21684 36136 21690
rect 36084 21626 36136 21632
rect 35992 21480 36044 21486
rect 35992 21422 36044 21428
rect 35900 21140 35952 21146
rect 35900 21082 35952 21088
rect 36556 20806 36584 22918
rect 35900 20800 35952 20806
rect 35900 20742 35952 20748
rect 36544 20800 36596 20806
rect 36544 20742 36596 20748
rect 35808 20392 35860 20398
rect 35808 20334 35860 20340
rect 35808 20256 35860 20262
rect 35912 20244 35940 20742
rect 35860 20216 35940 20244
rect 36176 20256 36228 20262
rect 35808 20198 35860 20204
rect 36176 20198 36228 20204
rect 35636 19944 35756 19972
rect 35532 19916 35584 19922
rect 35532 19858 35584 19864
rect 35544 19174 35572 19858
rect 35532 19168 35584 19174
rect 35532 19110 35584 19116
rect 35544 18970 35572 19110
rect 35532 18964 35584 18970
rect 35532 18906 35584 18912
rect 35636 17610 35664 19944
rect 35716 19848 35768 19854
rect 35716 19790 35768 19796
rect 35728 19174 35756 19790
rect 35820 19514 35848 20198
rect 35808 19508 35860 19514
rect 35808 19450 35860 19456
rect 35820 19242 35848 19450
rect 36188 19310 36216 20198
rect 37108 19825 37136 34478
rect 37832 26784 37884 26790
rect 37832 26726 37884 26732
rect 37844 26625 37872 26726
rect 37830 26616 37886 26625
rect 37830 26551 37886 26560
rect 37094 19816 37150 19825
rect 37094 19751 37150 19760
rect 36176 19304 36228 19310
rect 36176 19246 36228 19252
rect 35808 19236 35860 19242
rect 35808 19178 35860 19184
rect 35716 19168 35768 19174
rect 35716 19110 35768 19116
rect 35728 18630 35756 19110
rect 35716 18624 35768 18630
rect 35716 18566 35768 18572
rect 35820 18578 35848 19178
rect 36188 18902 36216 19246
rect 36176 18896 36228 18902
rect 36176 18838 36228 18844
rect 35728 18154 35756 18566
rect 35820 18550 35940 18578
rect 35808 18420 35860 18426
rect 35808 18362 35860 18368
rect 35716 18148 35768 18154
rect 35716 18090 35768 18096
rect 35624 17604 35676 17610
rect 35624 17546 35676 17552
rect 35716 17536 35768 17542
rect 35622 17504 35678 17513
rect 35716 17478 35768 17484
rect 35622 17439 35678 17448
rect 35440 16584 35492 16590
rect 35440 16526 35492 16532
rect 34940 16348 35236 16368
rect 34996 16346 35020 16348
rect 35076 16346 35100 16348
rect 35156 16346 35180 16348
rect 35018 16294 35020 16346
rect 35082 16294 35094 16346
rect 35156 16294 35158 16346
rect 34996 16292 35020 16294
rect 35076 16292 35100 16294
rect 35156 16292 35180 16294
rect 34940 16272 35236 16292
rect 35438 16280 35494 16289
rect 35438 16215 35494 16224
rect 35452 15570 35480 16215
rect 35636 16153 35664 17439
rect 35728 17338 35756 17478
rect 35716 17332 35768 17338
rect 35716 17274 35768 17280
rect 35622 16144 35678 16153
rect 35622 16079 35678 16088
rect 35728 15706 35756 17274
rect 35820 17066 35848 18362
rect 35912 18222 35940 18550
rect 35900 18216 35952 18222
rect 35900 18158 35952 18164
rect 35912 17882 35940 18158
rect 35900 17876 35952 17882
rect 35900 17818 35952 17824
rect 36268 17808 36320 17814
rect 36268 17750 36320 17756
rect 35900 17604 35952 17610
rect 35900 17546 35952 17552
rect 35808 17060 35860 17066
rect 35808 17002 35860 17008
rect 35820 16794 35848 17002
rect 35808 16788 35860 16794
rect 35808 16730 35860 16736
rect 35808 15904 35860 15910
rect 35808 15846 35860 15852
rect 35716 15700 35768 15706
rect 35716 15642 35768 15648
rect 35440 15564 35492 15570
rect 35440 15506 35492 15512
rect 34940 15260 35236 15280
rect 34996 15258 35020 15260
rect 35076 15258 35100 15260
rect 35156 15258 35180 15260
rect 35018 15206 35020 15258
rect 35082 15206 35094 15258
rect 35156 15206 35158 15258
rect 34996 15204 35020 15206
rect 35076 15204 35100 15206
rect 35156 15204 35180 15206
rect 34940 15184 35236 15204
rect 35452 15162 35480 15506
rect 35440 15156 35492 15162
rect 35440 15098 35492 15104
rect 35622 15056 35678 15065
rect 35622 14991 35678 15000
rect 35256 14952 35308 14958
rect 35256 14894 35308 14900
rect 34940 14172 35236 14192
rect 34996 14170 35020 14172
rect 35076 14170 35100 14172
rect 35156 14170 35180 14172
rect 35018 14118 35020 14170
rect 35082 14118 35094 14170
rect 35156 14118 35158 14170
rect 34996 14116 35020 14118
rect 35076 14116 35100 14118
rect 35156 14116 35180 14118
rect 34940 14096 35236 14116
rect 35268 13870 35296 14894
rect 35532 14816 35584 14822
rect 35532 14758 35584 14764
rect 35544 14618 35572 14758
rect 35532 14612 35584 14618
rect 35532 14554 35584 14560
rect 35544 13870 35572 14554
rect 35256 13864 35308 13870
rect 35256 13806 35308 13812
rect 35532 13864 35584 13870
rect 35532 13806 35584 13812
rect 34796 13728 34848 13734
rect 34796 13670 34848 13676
rect 35268 13530 35296 13806
rect 35348 13728 35400 13734
rect 35348 13670 35400 13676
rect 34796 13524 34848 13530
rect 34796 13466 34848 13472
rect 35256 13524 35308 13530
rect 35256 13466 35308 13472
rect 34808 12850 34836 13466
rect 35256 13184 35308 13190
rect 35256 13126 35308 13132
rect 34940 13084 35236 13104
rect 34996 13082 35020 13084
rect 35076 13082 35100 13084
rect 35156 13082 35180 13084
rect 35018 13030 35020 13082
rect 35082 13030 35094 13082
rect 35156 13030 35158 13082
rect 34996 13028 35020 13030
rect 35076 13028 35100 13030
rect 35156 13028 35180 13030
rect 34940 13008 35236 13028
rect 34796 12844 34848 12850
rect 34796 12786 34848 12792
rect 35268 12782 35296 13126
rect 35256 12776 35308 12782
rect 35256 12718 35308 12724
rect 35360 12594 35388 13670
rect 35544 13394 35572 13806
rect 35532 13388 35584 13394
rect 35532 13330 35584 13336
rect 35532 13252 35584 13258
rect 35532 13194 35584 13200
rect 35268 12566 35388 12594
rect 34940 11996 35236 12016
rect 34996 11994 35020 11996
rect 35076 11994 35100 11996
rect 35156 11994 35180 11996
rect 35018 11942 35020 11994
rect 35082 11942 35094 11994
rect 35156 11942 35158 11994
rect 34996 11940 35020 11942
rect 35076 11940 35100 11942
rect 35156 11940 35180 11942
rect 34940 11920 35236 11940
rect 35268 11830 35296 12566
rect 35346 12472 35402 12481
rect 35346 12407 35402 12416
rect 35360 11898 35388 12407
rect 35440 12096 35492 12102
rect 35440 12038 35492 12044
rect 35348 11892 35400 11898
rect 35348 11834 35400 11840
rect 35256 11824 35308 11830
rect 35256 11766 35308 11772
rect 35346 11792 35402 11801
rect 35452 11762 35480 12038
rect 35346 11727 35402 11736
rect 35440 11756 35492 11762
rect 35360 11694 35388 11727
rect 35440 11698 35492 11704
rect 35348 11688 35400 11694
rect 35348 11630 35400 11636
rect 35072 11620 35124 11626
rect 35072 11562 35124 11568
rect 35084 11354 35112 11562
rect 35072 11348 35124 11354
rect 35072 11290 35124 11296
rect 35452 11286 35480 11698
rect 35440 11280 35492 11286
rect 35440 11222 35492 11228
rect 35440 11144 35492 11150
rect 35440 11086 35492 11092
rect 34940 10908 35236 10928
rect 34996 10906 35020 10908
rect 35076 10906 35100 10908
rect 35156 10906 35180 10908
rect 35018 10854 35020 10906
rect 35082 10854 35094 10906
rect 35156 10854 35158 10906
rect 34996 10852 35020 10854
rect 35076 10852 35100 10854
rect 35156 10852 35180 10854
rect 34940 10832 35236 10852
rect 35452 10674 35480 11086
rect 35440 10668 35492 10674
rect 35440 10610 35492 10616
rect 35452 10266 35480 10610
rect 35544 10266 35572 13194
rect 35440 10260 35492 10266
rect 35440 10202 35492 10208
rect 35532 10260 35584 10266
rect 35532 10202 35584 10208
rect 34796 9920 34848 9926
rect 34796 9862 34848 9868
rect 34808 9450 34836 9862
rect 34940 9820 35236 9840
rect 34996 9818 35020 9820
rect 35076 9818 35100 9820
rect 35156 9818 35180 9820
rect 35018 9766 35020 9818
rect 35082 9766 35094 9818
rect 35156 9766 35158 9818
rect 34996 9764 35020 9766
rect 35076 9764 35100 9766
rect 35156 9764 35180 9766
rect 34940 9744 35236 9764
rect 34796 9444 34848 9450
rect 34796 9386 34848 9392
rect 35440 9444 35492 9450
rect 35440 9386 35492 9392
rect 34888 9376 34940 9382
rect 34808 9324 34888 9330
rect 34808 9318 34940 9324
rect 34808 9302 34928 9318
rect 34704 8560 34756 8566
rect 34704 8502 34756 8508
rect 34624 8350 34744 8378
rect 34612 7744 34664 7750
rect 34612 7686 34664 7692
rect 34624 7449 34652 7686
rect 34610 7440 34666 7449
rect 34610 7375 34666 7384
rect 34716 6769 34744 8350
rect 34808 7750 34836 9302
rect 35348 9036 35400 9042
rect 35348 8978 35400 8984
rect 34940 8732 35236 8752
rect 34996 8730 35020 8732
rect 35076 8730 35100 8732
rect 35156 8730 35180 8732
rect 35018 8678 35020 8730
rect 35082 8678 35094 8730
rect 35156 8678 35158 8730
rect 34996 8676 35020 8678
rect 35076 8676 35100 8678
rect 35156 8676 35180 8678
rect 34940 8656 35236 8676
rect 35164 8560 35216 8566
rect 35216 8508 35296 8514
rect 35164 8502 35296 8508
rect 35176 8486 35296 8502
rect 34796 7744 34848 7750
rect 34796 7686 34848 7692
rect 34940 7644 35236 7664
rect 34996 7642 35020 7644
rect 35076 7642 35100 7644
rect 35156 7642 35180 7644
rect 35018 7590 35020 7642
rect 35082 7590 35094 7642
rect 35156 7590 35158 7642
rect 34996 7588 35020 7590
rect 35076 7588 35100 7590
rect 35156 7588 35180 7590
rect 34940 7568 35236 7588
rect 34796 6996 34848 7002
rect 34796 6938 34848 6944
rect 34702 6760 34758 6769
rect 34702 6695 34758 6704
rect 34532 6616 34744 6644
rect 34244 6384 34296 6390
rect 33782 6352 33838 6361
rect 33416 6316 33468 6322
rect 34244 6326 34296 6332
rect 33782 6287 33784 6296
rect 33416 6258 33468 6264
rect 33836 6287 33838 6296
rect 33784 6258 33836 6264
rect 33428 5710 33456 6258
rect 33796 6227 33824 6258
rect 34612 6112 34664 6118
rect 34612 6054 34664 6060
rect 33876 5908 33928 5914
rect 33876 5850 33928 5856
rect 33600 5840 33652 5846
rect 33600 5782 33652 5788
rect 33416 5704 33468 5710
rect 33416 5646 33468 5652
rect 33612 5370 33640 5782
rect 33888 5370 33916 5850
rect 34256 5710 34284 5741
rect 34244 5704 34296 5710
rect 34242 5672 34244 5681
rect 34428 5704 34480 5710
rect 34296 5672 34298 5681
rect 34428 5646 34480 5652
rect 34242 5607 34298 5616
rect 34256 5370 34284 5607
rect 33600 5364 33652 5370
rect 33600 5306 33652 5312
rect 33876 5364 33928 5370
rect 33876 5306 33928 5312
rect 34244 5364 34296 5370
rect 34244 5306 34296 5312
rect 34440 5234 34468 5646
rect 34520 5636 34572 5642
rect 34520 5578 34572 5584
rect 34428 5228 34480 5234
rect 34428 5170 34480 5176
rect 34532 4842 34560 5578
rect 34440 4826 34560 4842
rect 33784 4820 33836 4826
rect 33784 4762 33836 4768
rect 34428 4820 34560 4826
rect 34480 4814 34560 4820
rect 34428 4762 34480 4768
rect 33796 4282 33824 4762
rect 34624 4758 34652 6054
rect 34716 5273 34744 6616
rect 34808 5896 34836 6938
rect 34940 6556 35236 6576
rect 34996 6554 35020 6556
rect 35076 6554 35100 6556
rect 35156 6554 35180 6556
rect 35018 6502 35020 6554
rect 35082 6502 35094 6554
rect 35156 6502 35158 6554
rect 34996 6500 35020 6502
rect 35076 6500 35100 6502
rect 35156 6500 35180 6502
rect 34940 6480 35236 6500
rect 35072 6112 35124 6118
rect 35072 6054 35124 6060
rect 35084 5914 35112 6054
rect 35072 5908 35124 5914
rect 34808 5868 34928 5896
rect 34796 5772 34848 5778
rect 34796 5714 34848 5720
rect 34702 5264 34758 5273
rect 34702 5199 34758 5208
rect 34704 5160 34756 5166
rect 34704 5102 34756 5108
rect 34716 4826 34744 5102
rect 34808 5030 34836 5714
rect 34900 5710 34928 5868
rect 35072 5850 35124 5856
rect 35268 5794 35296 8486
rect 35360 8090 35388 8978
rect 35452 8906 35480 9386
rect 35440 8900 35492 8906
rect 35440 8842 35492 8848
rect 35452 8498 35480 8842
rect 35440 8492 35492 8498
rect 35440 8434 35492 8440
rect 35348 8084 35400 8090
rect 35348 8026 35400 8032
rect 35544 7818 35572 10202
rect 35636 8022 35664 14991
rect 35820 13530 35848 15846
rect 35912 14804 35940 17546
rect 35992 15700 36044 15706
rect 35992 15642 36044 15648
rect 36004 14958 36032 15642
rect 35992 14952 36044 14958
rect 35992 14894 36044 14900
rect 35912 14776 36032 14804
rect 35900 14272 35952 14278
rect 35900 14214 35952 14220
rect 35808 13524 35860 13530
rect 35808 13466 35860 13472
rect 35820 12986 35848 13466
rect 35912 13326 35940 14214
rect 35900 13320 35952 13326
rect 35900 13262 35952 13268
rect 35912 12986 35940 13262
rect 36004 13190 36032 14776
rect 36176 14612 36228 14618
rect 36176 14554 36228 14560
rect 36084 14544 36136 14550
rect 36084 14486 36136 14492
rect 36096 14074 36124 14486
rect 36188 14414 36216 14554
rect 36176 14408 36228 14414
rect 36176 14350 36228 14356
rect 36084 14068 36136 14074
rect 36084 14010 36136 14016
rect 36188 13530 36216 14350
rect 36176 13524 36228 13530
rect 36176 13466 36228 13472
rect 36084 13320 36136 13326
rect 36084 13262 36136 13268
rect 35992 13184 36044 13190
rect 35992 13126 36044 13132
rect 35808 12980 35860 12986
rect 35808 12922 35860 12928
rect 35900 12980 35952 12986
rect 35900 12922 35952 12928
rect 35716 12776 35768 12782
rect 35716 12718 35768 12724
rect 35728 12102 35756 12718
rect 35716 12096 35768 12102
rect 35716 12038 35768 12044
rect 35716 11892 35768 11898
rect 35716 11834 35768 11840
rect 35624 8016 35676 8022
rect 35624 7958 35676 7964
rect 35532 7812 35584 7818
rect 35532 7754 35584 7760
rect 35636 7546 35664 7958
rect 35728 7857 35756 11834
rect 35808 10532 35860 10538
rect 35808 10474 35860 10480
rect 35820 9722 35848 10474
rect 35808 9716 35860 9722
rect 35808 9658 35860 9664
rect 35820 8974 35848 9658
rect 36004 9382 36032 13126
rect 36096 12442 36124 13262
rect 36084 12436 36136 12442
rect 36084 12378 36136 12384
rect 36280 11898 36308 17750
rect 36912 16992 36964 16998
rect 36912 16934 36964 16940
rect 36636 16584 36688 16590
rect 36636 16526 36688 16532
rect 36452 14884 36504 14890
rect 36452 14826 36504 14832
rect 36464 14414 36492 14826
rect 36452 14408 36504 14414
rect 36452 14350 36504 14356
rect 36464 14074 36492 14350
rect 36452 14068 36504 14074
rect 36452 14010 36504 14016
rect 36464 12918 36492 14010
rect 36452 12912 36504 12918
rect 36452 12854 36504 12860
rect 36542 12744 36598 12753
rect 36542 12679 36598 12688
rect 36268 11892 36320 11898
rect 36268 11834 36320 11840
rect 36084 11824 36136 11830
rect 36084 11766 36136 11772
rect 35992 9376 36044 9382
rect 35992 9318 36044 9324
rect 35808 8968 35860 8974
rect 35808 8910 35860 8916
rect 35820 8634 35848 8910
rect 35900 8900 35952 8906
rect 35900 8842 35952 8848
rect 35808 8628 35860 8634
rect 35808 8570 35860 8576
rect 35912 8566 35940 8842
rect 35900 8560 35952 8566
rect 35900 8502 35952 8508
rect 36096 8362 36124 11766
rect 36268 10124 36320 10130
rect 36268 10066 36320 10072
rect 36280 9518 36308 10066
rect 36360 10056 36412 10062
rect 36360 9998 36412 10004
rect 36268 9512 36320 9518
rect 36268 9454 36320 9460
rect 36280 9178 36308 9454
rect 36372 9178 36400 9998
rect 36268 9172 36320 9178
rect 36268 9114 36320 9120
rect 36360 9172 36412 9178
rect 36360 9114 36412 9120
rect 35808 8356 35860 8362
rect 35808 8298 35860 8304
rect 36084 8356 36136 8362
rect 36084 8298 36136 8304
rect 35714 7848 35770 7857
rect 35714 7783 35770 7792
rect 35716 7744 35768 7750
rect 35716 7686 35768 7692
rect 35624 7540 35676 7546
rect 35624 7482 35676 7488
rect 35440 7336 35492 7342
rect 35440 7278 35492 7284
rect 35452 7002 35480 7278
rect 35440 6996 35492 7002
rect 35440 6938 35492 6944
rect 35440 6860 35492 6866
rect 35440 6802 35492 6808
rect 35452 6118 35480 6802
rect 35532 6656 35584 6662
rect 35532 6598 35584 6604
rect 35440 6112 35492 6118
rect 35438 6080 35440 6089
rect 35492 6080 35494 6089
rect 35438 6015 35494 6024
rect 35544 5846 35572 6598
rect 35532 5840 35584 5846
rect 35268 5766 35388 5794
rect 35532 5782 35584 5788
rect 34888 5704 34940 5710
rect 34888 5646 34940 5652
rect 35256 5704 35308 5710
rect 35256 5646 35308 5652
rect 34940 5468 35236 5488
rect 34996 5466 35020 5468
rect 35076 5466 35100 5468
rect 35156 5466 35180 5468
rect 35018 5414 35020 5466
rect 35082 5414 35094 5466
rect 35156 5414 35158 5466
rect 34996 5412 35020 5414
rect 35076 5412 35100 5414
rect 35156 5412 35180 5414
rect 34940 5392 35236 5412
rect 35164 5228 35216 5234
rect 35164 5170 35216 5176
rect 34796 5024 34848 5030
rect 34796 4966 34848 4972
rect 34704 4820 34756 4826
rect 34704 4762 34756 4768
rect 34612 4752 34664 4758
rect 34242 4720 34298 4729
rect 34060 4684 34112 4690
rect 34612 4694 34664 4700
rect 34242 4655 34298 4664
rect 34704 4684 34756 4690
rect 34060 4626 34112 4632
rect 34072 4570 34100 4626
rect 34256 4622 34284 4655
rect 34704 4626 34756 4632
rect 34244 4616 34296 4622
rect 34072 4542 34192 4570
rect 34244 4558 34296 4564
rect 33784 4276 33836 4282
rect 33784 4218 33836 4224
rect 31760 4014 31812 4020
rect 31208 4004 31260 4010
rect 31208 3946 31260 3952
rect 31024 3732 31076 3738
rect 31024 3674 31076 3680
rect 30748 3392 30800 3398
rect 30748 3334 30800 3340
rect 30288 2848 30340 2854
rect 30288 2790 30340 2796
rect 30300 2582 30328 2790
rect 30760 2650 30788 3334
rect 31220 2854 31248 3946
rect 31772 3534 31800 4014
rect 33060 3998 33272 4026
rect 33060 3602 33088 3998
rect 34164 3942 34192 4542
rect 34716 4282 34744 4626
rect 34704 4276 34756 4282
rect 34704 4218 34756 4224
rect 33140 3936 33192 3942
rect 34152 3936 34204 3942
rect 33140 3878 33192 3884
rect 34150 3904 34152 3913
rect 34204 3904 34206 3913
rect 32404 3596 32456 3602
rect 32404 3538 32456 3544
rect 33048 3596 33100 3602
rect 33048 3538 33100 3544
rect 31760 3528 31812 3534
rect 31760 3470 31812 3476
rect 31574 3224 31630 3233
rect 31574 3159 31576 3168
rect 31628 3159 31630 3168
rect 31576 3130 31628 3136
rect 31772 3058 31800 3470
rect 32036 3188 32088 3194
rect 32036 3130 32088 3136
rect 31300 3052 31352 3058
rect 31300 2994 31352 3000
rect 31760 3052 31812 3058
rect 31760 2994 31812 3000
rect 31208 2848 31260 2854
rect 31208 2790 31260 2796
rect 30748 2644 30800 2650
rect 30748 2586 30800 2592
rect 30288 2576 30340 2582
rect 30288 2518 30340 2524
rect 31312 2514 31340 2994
rect 32048 2990 32076 3130
rect 32036 2984 32088 2990
rect 31942 2952 31998 2961
rect 32036 2926 32088 2932
rect 31942 2887 31998 2896
rect 31956 2650 31984 2887
rect 32416 2650 32444 3538
rect 33060 3505 33088 3538
rect 32494 3496 32550 3505
rect 32494 3431 32496 3440
rect 32548 3431 32550 3440
rect 33046 3496 33102 3505
rect 33046 3431 33102 3440
rect 32496 3402 32548 3408
rect 33152 2990 33180 3878
rect 34150 3839 34206 3848
rect 34716 3670 34744 4218
rect 34808 4010 34836 4966
rect 35176 4622 35204 5170
rect 35268 5030 35296 5646
rect 35256 5024 35308 5030
rect 35256 4966 35308 4972
rect 34980 4616 35032 4622
rect 34978 4584 34980 4593
rect 35164 4616 35216 4622
rect 35032 4584 35034 4593
rect 35164 4558 35216 4564
rect 34978 4519 35034 4528
rect 34940 4380 35236 4400
rect 34996 4378 35020 4380
rect 35076 4378 35100 4380
rect 35156 4378 35180 4380
rect 35018 4326 35020 4378
rect 35082 4326 35094 4378
rect 35156 4326 35158 4378
rect 34996 4324 35020 4326
rect 35076 4324 35100 4326
rect 35156 4324 35180 4326
rect 34940 4304 35236 4324
rect 34796 4004 34848 4010
rect 34796 3946 34848 3952
rect 34704 3664 34756 3670
rect 34704 3606 34756 3612
rect 33692 3596 33744 3602
rect 33692 3538 33744 3544
rect 33416 3528 33468 3534
rect 33416 3470 33468 3476
rect 33428 2990 33456 3470
rect 33704 3097 33732 3538
rect 34612 3392 34664 3398
rect 34612 3334 34664 3340
rect 33690 3088 33746 3097
rect 33690 3023 33692 3032
rect 33744 3023 33746 3032
rect 33692 2994 33744 3000
rect 33140 2984 33192 2990
rect 33140 2926 33192 2932
rect 33416 2984 33468 2990
rect 33416 2926 33468 2932
rect 33048 2848 33100 2854
rect 33048 2790 33100 2796
rect 31944 2644 31996 2650
rect 31944 2586 31996 2592
rect 32404 2644 32456 2650
rect 32404 2586 32456 2592
rect 33060 2582 33088 2790
rect 33048 2576 33100 2582
rect 33048 2518 33100 2524
rect 33428 2514 33456 2926
rect 33704 2650 33732 2994
rect 34520 2984 34572 2990
rect 34520 2926 34572 2932
rect 34532 2650 34560 2926
rect 34624 2854 34652 3334
rect 34940 3292 35236 3312
rect 34996 3290 35020 3292
rect 35076 3290 35100 3292
rect 35156 3290 35180 3292
rect 35018 3238 35020 3290
rect 35082 3238 35094 3290
rect 35156 3238 35158 3290
rect 34996 3236 35020 3238
rect 35076 3236 35100 3238
rect 35156 3236 35180 3238
rect 34940 3216 35236 3236
rect 34612 2848 34664 2854
rect 34610 2816 34612 2825
rect 34664 2816 34666 2825
rect 34610 2751 34666 2760
rect 35268 2650 35296 4966
rect 33692 2644 33744 2650
rect 33692 2586 33744 2592
rect 34520 2644 34572 2650
rect 34520 2586 34572 2592
rect 35256 2644 35308 2650
rect 35256 2586 35308 2592
rect 31300 2508 31352 2514
rect 31300 2450 31352 2456
rect 33416 2508 33468 2514
rect 33416 2450 33468 2456
rect 34940 2204 35236 2224
rect 34996 2202 35020 2204
rect 35076 2202 35100 2204
rect 35156 2202 35180 2204
rect 35018 2150 35020 2202
rect 35082 2150 35094 2202
rect 35156 2150 35158 2202
rect 34996 2148 35020 2150
rect 35076 2148 35100 2150
rect 35156 2148 35180 2150
rect 34940 2128 35236 2148
rect 35360 1737 35388 5766
rect 35532 5704 35584 5710
rect 35532 5646 35584 5652
rect 35544 4593 35572 5646
rect 35530 4584 35586 4593
rect 35530 4519 35586 4528
rect 35532 4480 35584 4486
rect 35532 4422 35584 4428
rect 35544 4078 35572 4422
rect 35532 4072 35584 4078
rect 35532 4014 35584 4020
rect 35544 3738 35572 4014
rect 35532 3732 35584 3738
rect 35532 3674 35584 3680
rect 35544 2990 35572 3674
rect 35532 2984 35584 2990
rect 35728 2961 35756 7686
rect 35820 4185 35848 8298
rect 36176 7948 36228 7954
rect 36176 7890 36228 7896
rect 36084 7744 36136 7750
rect 36084 7686 36136 7692
rect 36096 6254 36124 7686
rect 36188 7274 36216 7890
rect 36360 7812 36412 7818
rect 36360 7754 36412 7760
rect 36176 7268 36228 7274
rect 36176 7210 36228 7216
rect 36188 6662 36216 7210
rect 36176 6656 36228 6662
rect 36176 6598 36228 6604
rect 36084 6248 36136 6254
rect 36084 6190 36136 6196
rect 35900 6112 35952 6118
rect 35900 6054 35952 6060
rect 35912 4729 35940 6054
rect 36188 5370 36216 6598
rect 36268 5568 36320 5574
rect 36268 5510 36320 5516
rect 36176 5364 36228 5370
rect 36176 5306 36228 5312
rect 36280 5098 36308 5510
rect 36268 5092 36320 5098
rect 36268 5034 36320 5040
rect 35898 4720 35954 4729
rect 35898 4655 35954 4664
rect 36280 4486 36308 5034
rect 36268 4480 36320 4486
rect 36268 4422 36320 4428
rect 35806 4176 35862 4185
rect 35806 4111 35862 4120
rect 35808 4004 35860 4010
rect 35808 3946 35860 3952
rect 35820 3618 35848 3946
rect 35898 3904 35954 3913
rect 35898 3839 35954 3848
rect 35912 3738 35940 3839
rect 35900 3732 35952 3738
rect 35900 3674 35952 3680
rect 35820 3590 36032 3618
rect 36280 3602 36308 4422
rect 35532 2926 35584 2932
rect 35714 2952 35770 2961
rect 35544 2514 35572 2926
rect 35714 2887 35770 2896
rect 35808 2848 35860 2854
rect 35808 2790 35860 2796
rect 35820 2582 35848 2790
rect 36004 2650 36032 3590
rect 36268 3596 36320 3602
rect 36268 3538 36320 3544
rect 36280 3194 36308 3538
rect 36268 3188 36320 3194
rect 36268 3130 36320 3136
rect 35992 2644 36044 2650
rect 35992 2586 36044 2592
rect 35808 2576 35860 2582
rect 35808 2518 35860 2524
rect 35532 2508 35584 2514
rect 35532 2450 35584 2456
rect 35346 1728 35402 1737
rect 35346 1663 35402 1672
rect 36372 649 36400 7754
rect 36452 6656 36504 6662
rect 36452 6598 36504 6604
rect 36464 4593 36492 6598
rect 36556 6458 36584 12679
rect 36648 9081 36676 16526
rect 36820 14000 36872 14006
rect 36820 13942 36872 13948
rect 36832 13841 36860 13942
rect 36818 13832 36874 13841
rect 36818 13767 36874 13776
rect 36820 10464 36872 10470
rect 36820 10406 36872 10412
rect 36832 10062 36860 10406
rect 36924 10305 36952 16934
rect 37002 13968 37058 13977
rect 37002 13903 37058 13912
rect 36910 10296 36966 10305
rect 36910 10231 36966 10240
rect 36820 10056 36872 10062
rect 36820 9998 36872 10004
rect 36832 9382 36860 9998
rect 36820 9376 36872 9382
rect 36820 9318 36872 9324
rect 36832 9217 36860 9318
rect 36818 9208 36874 9217
rect 36818 9143 36874 9152
rect 36634 9072 36690 9081
rect 36634 9007 36690 9016
rect 36636 8288 36688 8294
rect 36636 8230 36688 8236
rect 36544 6452 36596 6458
rect 36544 6394 36596 6400
rect 36648 5681 36676 8230
rect 37016 6866 37044 13903
rect 37094 11520 37150 11529
rect 37094 11455 37150 11464
rect 37108 8634 37136 11455
rect 37096 8628 37148 8634
rect 37096 8570 37148 8576
rect 37108 8430 37136 8570
rect 37096 8424 37148 8430
rect 37096 8366 37148 8372
rect 37004 6860 37056 6866
rect 37004 6802 37056 6808
rect 37016 6458 37044 6802
rect 37004 6452 37056 6458
rect 37004 6394 37056 6400
rect 37280 6384 37332 6390
rect 37278 6352 37280 6361
rect 37332 6352 37334 6361
rect 37278 6287 37334 6296
rect 36634 5672 36690 5681
rect 36634 5607 36690 5616
rect 36450 4584 36506 4593
rect 36450 4519 36506 4528
rect 36464 3534 36492 4519
rect 36820 3936 36872 3942
rect 36820 3878 36872 3884
rect 36832 3670 36860 3878
rect 36820 3664 36872 3670
rect 36820 3606 36872 3612
rect 36452 3528 36504 3534
rect 36452 3470 36504 3476
rect 36634 3496 36690 3505
rect 36464 3058 36492 3470
rect 36634 3431 36690 3440
rect 36452 3052 36504 3058
rect 36452 2994 36504 3000
rect 36358 640 36414 649
rect 29748 598 30052 626
rect 30024 480 30052 598
rect 36358 575 36414 584
rect 36648 480 36676 3431
rect 36832 3126 36860 3606
rect 36820 3120 36872 3126
rect 36820 3062 36872 3068
rect 3330 0 3386 480
rect 9954 0 10010 480
rect 16670 0 16726 480
rect 23294 0 23350 480
rect 30010 0 30066 480
rect 36634 0 36690 480
<< via2 >>
rect 1398 35264 1454 35320
rect 2042 34992 2098 35048
rect 3146 36080 3202 36136
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 4986 35436 4988 35456
rect 4988 35436 5040 35456
rect 5040 35436 5042 35456
rect 4986 35400 5042 35436
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 4066 33904 4122 33960
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 7470 35828 7526 35864
rect 7470 35808 7472 35828
rect 7472 35808 7524 35828
rect 7524 35808 7526 35828
rect 6642 35708 6644 35728
rect 6644 35708 6696 35728
rect 6696 35708 6698 35728
rect 6642 35672 6698 35708
rect 6826 35672 6882 35728
rect 8574 35556 8630 35592
rect 8574 35536 8576 35556
rect 8576 35536 8628 35556
rect 8628 35536 8630 35556
rect 5538 35436 5540 35456
rect 5540 35436 5592 35456
rect 5592 35436 5594 35456
rect 5538 35400 5594 35436
rect 6826 35148 6882 35184
rect 6826 35128 6828 35148
rect 6828 35128 6880 35148
rect 6880 35128 6882 35148
rect 5078 34604 5134 34640
rect 5078 34584 5080 34604
rect 5080 34584 5132 34604
rect 5132 34584 5134 34604
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 2870 32020 2926 32056
rect 2870 32000 2872 32020
rect 2872 32000 2924 32020
rect 2924 32000 2926 32020
rect 4986 32020 5042 32056
rect 4986 32000 4988 32020
rect 4988 32000 5040 32020
rect 5040 32000 5042 32020
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 3330 31048 3386 31104
rect 1674 29708 1730 29744
rect 1674 29688 1676 29708
rect 1676 29688 1728 29708
rect 1728 29688 1730 29708
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 5814 31084 5816 31104
rect 5816 31084 5868 31104
rect 5868 31084 5870 31104
rect 5814 31048 5870 31084
rect 11610 35808 11666 35864
rect 11886 35828 11942 35864
rect 11886 35808 11888 35828
rect 11888 35808 11940 35828
rect 11940 35808 11942 35828
rect 10506 35672 10562 35728
rect 10874 35284 10930 35320
rect 10874 35264 10876 35284
rect 10876 35264 10928 35284
rect 10928 35264 10930 35284
rect 7470 34584 7526 34640
rect 8022 33088 8078 33144
rect 9402 35128 9458 35184
rect 8850 34740 8906 34776
rect 8850 34720 8852 34740
rect 8852 34720 8904 34740
rect 8904 34720 8906 34740
rect 4158 29688 4214 29744
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 7930 29144 7986 29200
rect 3974 27396 4030 27432
rect 3974 27376 3976 27396
rect 3976 27376 4028 27396
rect 4028 27376 4030 27396
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 8022 28600 8078 28656
rect 10874 34992 10930 35048
rect 10138 33108 10194 33144
rect 10138 33088 10140 33108
rect 10140 33088 10192 33108
rect 10192 33088 10194 33108
rect 9494 32444 9496 32464
rect 9496 32444 9548 32464
rect 9548 32444 9550 32464
rect 9494 32408 9550 32444
rect 10874 32680 10930 32736
rect 10414 31084 10416 31104
rect 10416 31084 10468 31104
rect 10468 31084 10470 31104
rect 10414 31048 10470 31084
rect 5722 27376 5778 27432
rect 6458 26696 6514 26752
rect 10414 29960 10470 30016
rect 9678 29144 9734 29200
rect 13910 35808 13966 35864
rect 14462 35672 14518 35728
rect 13634 35128 13690 35184
rect 12714 34720 12770 34776
rect 13634 34856 13690 34912
rect 11610 33108 11666 33144
rect 11610 33088 11612 33108
rect 11612 33088 11664 33108
rect 11664 33088 11666 33108
rect 12990 33224 13046 33280
rect 13358 33224 13414 33280
rect 12806 32716 12808 32736
rect 12808 32716 12860 32736
rect 12860 32716 12862 32736
rect 12806 32680 12862 32716
rect 11334 32308 11336 32328
rect 11336 32308 11388 32328
rect 11388 32308 11390 32328
rect 11334 32272 11390 32308
rect 13818 32444 13820 32464
rect 13820 32444 13872 32464
rect 13872 32444 13874 32464
rect 13818 32408 13874 32444
rect 13174 31592 13230 31648
rect 11886 30252 11942 30288
rect 11886 30232 11888 30252
rect 11888 30232 11940 30252
rect 11940 30232 11942 30252
rect 9678 28620 9734 28656
rect 9678 28600 9680 28620
rect 9680 28600 9732 28620
rect 9732 28600 9734 28620
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 1582 20032 1638 20088
rect 8850 26732 8852 26752
rect 8852 26732 8904 26752
rect 8904 26732 8906 26752
rect 8850 26696 8906 26732
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 12622 29996 12624 30016
rect 12624 29996 12676 30016
rect 12676 29996 12678 30016
rect 12622 29960 12678 29996
rect 12990 29280 13046 29336
rect 11886 25472 11942 25528
rect 14554 33088 14610 33144
rect 14462 32680 14518 32736
rect 14278 31476 14334 31512
rect 14278 31456 14280 31476
rect 14280 31456 14332 31476
rect 14332 31456 14334 31476
rect 13818 31084 13820 31104
rect 13820 31084 13872 31104
rect 13872 31084 13874 31104
rect 13818 31048 13874 31084
rect 15290 33224 15346 33280
rect 15106 32408 15162 32464
rect 15842 33924 15898 33960
rect 15842 33904 15844 33924
rect 15844 33904 15896 33924
rect 15896 33904 15898 33924
rect 16026 32544 16082 32600
rect 15014 30232 15070 30288
rect 15290 30232 15346 30288
rect 17130 32408 17186 32464
rect 16118 31456 16174 31512
rect 15934 30368 15990 30424
rect 18050 36080 18106 36136
rect 17038 31592 17094 31648
rect 16946 30232 17002 30288
rect 15750 29144 15806 29200
rect 16394 29280 16450 29336
rect 15842 29008 15898 29064
rect 13726 26968 13782 27024
rect 15382 26968 15438 27024
rect 13266 25608 13322 25664
rect 13174 25472 13230 25528
rect 7194 23704 7250 23760
rect 10138 24692 10140 24712
rect 10140 24692 10192 24712
rect 10192 24692 10194 24712
rect 10138 24656 10194 24692
rect 10506 23704 10562 23760
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 10046 20596 10102 20632
rect 10046 20576 10048 20596
rect 10048 20576 10100 20596
rect 10100 20576 10102 20596
rect 14554 25608 14610 25664
rect 13818 25472 13874 25528
rect 13818 24656 13874 24712
rect 15658 25472 15714 25528
rect 15474 24520 15530 24576
rect 14462 24248 14518 24304
rect 18142 35400 18198 35456
rect 18142 34856 18198 34912
rect 17774 33260 17776 33280
rect 17776 33260 17828 33280
rect 17828 33260 17830 33280
rect 17774 33224 17830 33260
rect 18050 34584 18106 34640
rect 19154 34856 19210 34912
rect 18510 30368 18566 30424
rect 18142 29144 18198 29200
rect 18050 29008 18106 29064
rect 18970 28464 19026 28520
rect 18694 27124 18750 27160
rect 18694 27104 18696 27124
rect 18696 27104 18748 27124
rect 18748 27104 18750 27124
rect 19338 33224 19394 33280
rect 19580 37562 19636 37564
rect 19660 37562 19716 37564
rect 19740 37562 19796 37564
rect 19820 37562 19876 37564
rect 19580 37510 19606 37562
rect 19606 37510 19636 37562
rect 19660 37510 19670 37562
rect 19670 37510 19716 37562
rect 19740 37510 19786 37562
rect 19786 37510 19796 37562
rect 19820 37510 19850 37562
rect 19850 37510 19876 37562
rect 19580 37508 19636 37510
rect 19660 37508 19716 37510
rect 19740 37508 19796 37510
rect 19820 37508 19876 37510
rect 19580 36474 19636 36476
rect 19660 36474 19716 36476
rect 19740 36474 19796 36476
rect 19820 36474 19876 36476
rect 19580 36422 19606 36474
rect 19606 36422 19636 36474
rect 19660 36422 19670 36474
rect 19670 36422 19716 36474
rect 19740 36422 19786 36474
rect 19786 36422 19796 36474
rect 19820 36422 19850 36474
rect 19850 36422 19876 36474
rect 19580 36420 19636 36422
rect 19660 36420 19716 36422
rect 19740 36420 19796 36422
rect 19820 36420 19876 36422
rect 19580 35386 19636 35388
rect 19660 35386 19716 35388
rect 19740 35386 19796 35388
rect 19820 35386 19876 35388
rect 19580 35334 19606 35386
rect 19606 35334 19636 35386
rect 19660 35334 19670 35386
rect 19670 35334 19716 35386
rect 19740 35334 19786 35386
rect 19786 35334 19796 35386
rect 19820 35334 19850 35386
rect 19850 35334 19876 35386
rect 19580 35332 19636 35334
rect 19660 35332 19716 35334
rect 19740 35332 19796 35334
rect 19820 35332 19876 35334
rect 19580 34298 19636 34300
rect 19660 34298 19716 34300
rect 19740 34298 19796 34300
rect 19820 34298 19876 34300
rect 19580 34246 19606 34298
rect 19606 34246 19636 34298
rect 19660 34246 19670 34298
rect 19670 34246 19716 34298
rect 19740 34246 19786 34298
rect 19786 34246 19796 34298
rect 19820 34246 19850 34298
rect 19850 34246 19876 34298
rect 19580 34244 19636 34246
rect 19660 34244 19716 34246
rect 19740 34244 19796 34246
rect 19820 34244 19876 34246
rect 19580 33210 19636 33212
rect 19660 33210 19716 33212
rect 19740 33210 19796 33212
rect 19820 33210 19876 33212
rect 19580 33158 19606 33210
rect 19606 33158 19636 33210
rect 19660 33158 19670 33210
rect 19670 33158 19716 33210
rect 19740 33158 19786 33210
rect 19786 33158 19796 33210
rect 19820 33158 19850 33210
rect 19850 33158 19876 33210
rect 19580 33156 19636 33158
rect 19660 33156 19716 33158
rect 19740 33156 19796 33158
rect 19820 33156 19876 33158
rect 20166 32952 20222 33008
rect 19580 32122 19636 32124
rect 19660 32122 19716 32124
rect 19740 32122 19796 32124
rect 19820 32122 19876 32124
rect 19580 32070 19606 32122
rect 19606 32070 19636 32122
rect 19660 32070 19670 32122
rect 19670 32070 19716 32122
rect 19740 32070 19786 32122
rect 19786 32070 19796 32122
rect 19820 32070 19850 32122
rect 19850 32070 19876 32122
rect 19580 32068 19636 32070
rect 19660 32068 19716 32070
rect 19740 32068 19796 32070
rect 19820 32068 19876 32070
rect 19580 31034 19636 31036
rect 19660 31034 19716 31036
rect 19740 31034 19796 31036
rect 19820 31034 19876 31036
rect 19580 30982 19606 31034
rect 19606 30982 19636 31034
rect 19660 30982 19670 31034
rect 19670 30982 19716 31034
rect 19740 30982 19786 31034
rect 19786 30982 19796 31034
rect 19820 30982 19850 31034
rect 19850 30982 19876 31034
rect 19580 30980 19636 30982
rect 19660 30980 19716 30982
rect 19740 30980 19796 30982
rect 19820 30980 19876 30982
rect 19580 29946 19636 29948
rect 19660 29946 19716 29948
rect 19740 29946 19796 29948
rect 19820 29946 19876 29948
rect 19580 29894 19606 29946
rect 19606 29894 19636 29946
rect 19660 29894 19670 29946
rect 19670 29894 19716 29946
rect 19740 29894 19786 29946
rect 19786 29894 19796 29946
rect 19820 29894 19850 29946
rect 19850 29894 19876 29946
rect 19580 29892 19636 29894
rect 19660 29892 19716 29894
rect 19740 29892 19796 29894
rect 19820 29892 19876 29894
rect 19580 28858 19636 28860
rect 19660 28858 19716 28860
rect 19740 28858 19796 28860
rect 19820 28858 19876 28860
rect 19580 28806 19606 28858
rect 19606 28806 19636 28858
rect 19660 28806 19670 28858
rect 19670 28806 19716 28858
rect 19740 28806 19786 28858
rect 19786 28806 19796 28858
rect 19820 28806 19850 28858
rect 19850 28806 19876 28858
rect 19580 28804 19636 28806
rect 19660 28804 19716 28806
rect 19740 28804 19796 28806
rect 19820 28804 19876 28806
rect 19890 28500 19892 28520
rect 19892 28500 19944 28520
rect 19944 28500 19946 28520
rect 19890 28464 19946 28500
rect 19580 27770 19636 27772
rect 19660 27770 19716 27772
rect 19740 27770 19796 27772
rect 19820 27770 19876 27772
rect 19580 27718 19606 27770
rect 19606 27718 19636 27770
rect 19660 27718 19670 27770
rect 19670 27718 19716 27770
rect 19740 27718 19786 27770
rect 19786 27718 19796 27770
rect 19820 27718 19850 27770
rect 19850 27718 19876 27770
rect 19580 27716 19636 27718
rect 19660 27716 19716 27718
rect 19740 27716 19796 27718
rect 19820 27716 19876 27718
rect 19580 26682 19636 26684
rect 19660 26682 19716 26684
rect 19740 26682 19796 26684
rect 19820 26682 19876 26684
rect 19580 26630 19606 26682
rect 19606 26630 19636 26682
rect 19660 26630 19670 26682
rect 19670 26630 19716 26682
rect 19740 26630 19786 26682
rect 19786 26630 19796 26682
rect 19820 26630 19850 26682
rect 19850 26630 19876 26682
rect 19580 26628 19636 26630
rect 19660 26628 19716 26630
rect 19740 26628 19796 26630
rect 19820 26628 19876 26630
rect 18418 25492 18474 25528
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 18418 25472 18420 25492
rect 18420 25472 18472 25492
rect 18472 25472 18474 25492
rect 13634 21936 13690 21992
rect 13266 20576 13322 20632
rect 16854 22208 16910 22264
rect 15750 21972 15752 21992
rect 15752 21972 15804 21992
rect 15804 21972 15806 21992
rect 15750 21936 15806 21972
rect 15290 20984 15346 21040
rect 20626 34740 20682 34776
rect 20626 34720 20628 34740
rect 20628 34720 20680 34740
rect 20680 34720 20682 34740
rect 21362 33768 21418 33824
rect 21454 33088 21510 33144
rect 21914 34448 21970 34504
rect 25134 35536 25190 35592
rect 22742 34720 22798 34776
rect 23662 34448 23718 34504
rect 25042 34720 25098 34776
rect 24122 33768 24178 33824
rect 23938 33108 23994 33144
rect 23938 33088 23940 33108
rect 23940 33088 23992 33108
rect 23992 33088 23994 33108
rect 24674 32972 24730 33008
rect 24674 32952 24676 32972
rect 24676 32952 24728 32972
rect 24728 32952 24730 32972
rect 24674 31048 24730 31104
rect 23570 29708 23626 29744
rect 23570 29688 23572 29708
rect 23572 29688 23624 29708
rect 23624 29688 23626 29708
rect 22282 28484 22338 28520
rect 22282 28464 22284 28484
rect 22284 28464 22336 28484
rect 22336 28464 22338 28484
rect 20534 27104 20590 27160
rect 20994 25744 21050 25800
rect 18602 24556 18604 24576
rect 18604 24556 18656 24576
rect 18656 24556 18658 24576
rect 18602 24520 18658 24556
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 19062 23860 19118 23896
rect 19062 23840 19064 23860
rect 19064 23840 19116 23860
rect 19116 23840 19118 23860
rect 19154 23568 19210 23624
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 20074 24248 20130 24304
rect 19338 22208 19394 22264
rect 19154 21004 19210 21040
rect 19154 20984 19156 21004
rect 19156 20984 19208 21004
rect 19208 20984 19210 21004
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 21638 28212 21694 28248
rect 21638 28192 21640 28212
rect 21640 28192 21692 28212
rect 21692 28192 21694 28212
rect 24122 27648 24178 27704
rect 27250 35672 27306 35728
rect 29458 35128 29514 35184
rect 30562 34992 30618 35048
rect 31666 34584 31722 34640
rect 26514 31048 26570 31104
rect 35622 39344 35678 39400
rect 33874 35264 33930 35320
rect 34940 37018 34996 37020
rect 35020 37018 35076 37020
rect 35100 37018 35156 37020
rect 35180 37018 35236 37020
rect 34940 36966 34966 37018
rect 34966 36966 34996 37018
rect 35020 36966 35030 37018
rect 35030 36966 35076 37018
rect 35100 36966 35146 37018
rect 35146 36966 35156 37018
rect 35180 36966 35210 37018
rect 35210 36966 35236 37018
rect 34940 36964 34996 36966
rect 35020 36964 35076 36966
rect 35100 36964 35156 36966
rect 35180 36964 35236 36966
rect 34940 35930 34996 35932
rect 35020 35930 35076 35932
rect 35100 35930 35156 35932
rect 35180 35930 35236 35932
rect 34940 35878 34966 35930
rect 34966 35878 34996 35930
rect 35020 35878 35030 35930
rect 35030 35878 35076 35930
rect 35100 35878 35146 35930
rect 35146 35878 35156 35930
rect 35180 35878 35210 35930
rect 35210 35878 35236 35930
rect 34940 35876 34996 35878
rect 35020 35876 35076 35878
rect 35100 35876 35156 35878
rect 35180 35876 35236 35878
rect 35806 36896 35862 36952
rect 35530 35284 35586 35320
rect 35530 35264 35532 35284
rect 35532 35264 35584 35284
rect 35584 35264 35586 35284
rect 35714 35400 35770 35456
rect 34794 34856 34850 34912
rect 34940 34842 34996 34844
rect 35020 34842 35076 34844
rect 35100 34842 35156 34844
rect 35180 34842 35236 34844
rect 34940 34790 34966 34842
rect 34966 34790 34996 34842
rect 35020 34790 35030 34842
rect 35030 34790 35076 34842
rect 35100 34790 35146 34842
rect 35146 34790 35156 34842
rect 35180 34790 35210 34842
rect 35210 34790 35236 34842
rect 34940 34788 34996 34790
rect 35020 34788 35076 34790
rect 35100 34788 35156 34790
rect 35180 34788 35236 34790
rect 32770 33904 32826 33960
rect 34940 33754 34996 33756
rect 35020 33754 35076 33756
rect 35100 33754 35156 33756
rect 35180 33754 35236 33756
rect 34940 33702 34966 33754
rect 34966 33702 34996 33754
rect 35020 33702 35030 33754
rect 35030 33702 35076 33754
rect 35100 33702 35146 33754
rect 35146 33702 35156 33754
rect 35180 33702 35210 33754
rect 35210 33702 35236 33754
rect 34940 33700 34996 33702
rect 35020 33700 35076 33702
rect 35100 33700 35156 33702
rect 35180 33700 35236 33702
rect 34940 32666 34996 32668
rect 35020 32666 35076 32668
rect 35100 32666 35156 32668
rect 35180 32666 35236 32668
rect 34940 32614 34966 32666
rect 34966 32614 34996 32666
rect 35020 32614 35030 32666
rect 35030 32614 35076 32666
rect 35100 32614 35146 32666
rect 35146 32614 35156 32666
rect 35180 32614 35210 32666
rect 35210 32614 35236 32666
rect 34940 32612 34996 32614
rect 35020 32612 35076 32614
rect 35100 32612 35156 32614
rect 35180 32612 35236 32614
rect 30102 32544 30158 32600
rect 26882 29688 26938 29744
rect 25502 27412 25504 27432
rect 25504 27412 25556 27432
rect 25556 27412 25558 27432
rect 25502 27376 25558 27412
rect 22006 25744 22062 25800
rect 21546 23840 21602 23896
rect 23478 25780 23480 25800
rect 23480 25780 23532 25800
rect 23532 25780 23534 25800
rect 23478 25744 23534 25780
rect 24398 26152 24454 26208
rect 26238 26152 26294 26208
rect 26974 27648 27030 27704
rect 30010 28364 30012 28384
rect 30012 28364 30064 28384
rect 30064 28364 30066 28384
rect 30010 28328 30066 28364
rect 27894 27396 27950 27432
rect 27894 27376 27896 27396
rect 27896 27376 27948 27396
rect 27948 27376 27950 27396
rect 29182 26560 29238 26616
rect 29366 26424 29422 26480
rect 26606 25472 26662 25528
rect 21086 23568 21142 23624
rect 21546 22072 21602 22128
rect 21730 21004 21786 21040
rect 21730 20984 21732 21004
rect 21732 20984 21784 21004
rect 21784 20984 21786 21004
rect 23018 20576 23074 20632
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 18970 17584 19026 17640
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 16670 7520 16726 7576
rect 570 6704 626 6760
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 570 5616 626 5672
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 3330 3440 3386 3496
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 25502 22072 25558 22128
rect 23662 20984 23718 21040
rect 23846 19216 23902 19272
rect 24122 18808 24178 18864
rect 22190 17584 22246 17640
rect 20258 17312 20314 17368
rect 21822 17176 21878 17232
rect 19246 17040 19302 17096
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 23662 17176 23718 17232
rect 22466 17076 22468 17096
rect 22468 17076 22520 17096
rect 22520 17076 22522 17096
rect 22466 17040 22522 17076
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 21362 15136 21418 15192
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 18418 5616 18474 5672
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 25134 20576 25190 20632
rect 25410 20304 25466 20360
rect 24582 18808 24638 18864
rect 25318 18808 25374 18864
rect 24398 18672 24454 18728
rect 24766 17856 24822 17912
rect 26146 20460 26202 20496
rect 26146 20440 26148 20460
rect 26148 20440 26200 20460
rect 26200 20440 26202 20460
rect 27158 23024 27214 23080
rect 27894 21936 27950 21992
rect 26606 20032 26662 20088
rect 28078 20304 28134 20360
rect 26882 19236 26938 19272
rect 26882 19216 26884 19236
rect 26884 19216 26936 19236
rect 26936 19216 26938 19236
rect 26882 18672 26938 18728
rect 27802 18808 27858 18864
rect 26514 17876 26570 17912
rect 26514 17856 26516 17876
rect 26516 17856 26568 17876
rect 26568 17856 26570 17876
rect 25778 15816 25834 15872
rect 26238 15136 26294 15192
rect 27434 17448 27490 17504
rect 27710 17448 27766 17504
rect 27618 17312 27674 17368
rect 27434 12280 27490 12336
rect 28078 12180 28080 12200
rect 28080 12180 28132 12200
rect 28132 12180 28134 12200
rect 28078 12144 28134 12180
rect 28906 25644 28908 25664
rect 28908 25644 28960 25664
rect 28960 25644 28962 25664
rect 28906 25608 28962 25644
rect 29366 25472 29422 25528
rect 28446 18420 28502 18456
rect 28446 18400 28448 18420
rect 28448 18400 28500 18420
rect 28500 18400 28502 18420
rect 34940 31578 34996 31580
rect 35020 31578 35076 31580
rect 35100 31578 35156 31580
rect 35180 31578 35236 31580
rect 34940 31526 34966 31578
rect 34966 31526 34996 31578
rect 35020 31526 35030 31578
rect 35030 31526 35076 31578
rect 35100 31526 35146 31578
rect 35146 31526 35156 31578
rect 35180 31526 35210 31578
rect 35210 31526 35236 31578
rect 34940 31524 34996 31526
rect 35020 31524 35076 31526
rect 35100 31524 35156 31526
rect 35180 31524 35236 31526
rect 31574 28872 31630 28928
rect 31942 28364 31944 28384
rect 31944 28364 31996 28384
rect 31996 28364 31998 28384
rect 31942 28328 31998 28364
rect 30194 26288 30250 26344
rect 32126 26560 32182 26616
rect 33506 28872 33562 28928
rect 31942 26288 31998 26344
rect 31942 25608 31998 25664
rect 32310 19216 32366 19272
rect 29182 17448 29238 17504
rect 29918 16632 29974 16688
rect 29918 16244 29974 16280
rect 29918 16224 29920 16244
rect 29920 16224 29972 16244
rect 29972 16224 29974 16244
rect 28630 16108 28686 16144
rect 28630 16088 28632 16108
rect 28632 16088 28684 16108
rect 28684 16088 28686 16108
rect 30378 18808 30434 18864
rect 31298 18400 31354 18456
rect 32310 17992 32366 18048
rect 33782 20304 33838 20360
rect 34058 26968 34114 27024
rect 34610 28056 34666 28112
rect 34940 30490 34996 30492
rect 35020 30490 35076 30492
rect 35100 30490 35156 30492
rect 35180 30490 35236 30492
rect 34940 30438 34966 30490
rect 34966 30438 34996 30490
rect 35020 30438 35030 30490
rect 35030 30438 35076 30490
rect 35100 30438 35146 30490
rect 35146 30438 35156 30490
rect 35180 30438 35210 30490
rect 35210 30438 35236 30490
rect 34940 30436 34996 30438
rect 35020 30436 35076 30438
rect 35100 30436 35156 30438
rect 35180 30436 35236 30438
rect 34940 29402 34996 29404
rect 35020 29402 35076 29404
rect 35100 29402 35156 29404
rect 35180 29402 35236 29404
rect 34940 29350 34966 29402
rect 34966 29350 34996 29402
rect 35020 29350 35030 29402
rect 35030 29350 35076 29402
rect 35100 29350 35146 29402
rect 35146 29350 35156 29402
rect 35180 29350 35210 29402
rect 35210 29350 35236 29402
rect 34940 29348 34996 29350
rect 35020 29348 35076 29350
rect 35100 29348 35156 29350
rect 35180 29348 35236 29350
rect 34940 28314 34996 28316
rect 35020 28314 35076 28316
rect 35100 28314 35156 28316
rect 35180 28314 35236 28316
rect 34940 28262 34966 28314
rect 34966 28262 34996 28314
rect 35020 28262 35030 28314
rect 35030 28262 35076 28314
rect 35100 28262 35146 28314
rect 35146 28262 35156 28314
rect 35180 28262 35210 28314
rect 35210 28262 35236 28314
rect 34940 28260 34996 28262
rect 35020 28260 35076 28262
rect 35100 28260 35156 28262
rect 35180 28260 35236 28262
rect 34242 26832 34298 26888
rect 34242 26424 34298 26480
rect 34150 23568 34206 23624
rect 34702 23296 34758 23352
rect 34150 21936 34206 21992
rect 34518 22344 34574 22400
rect 34150 19896 34206 19952
rect 33966 19216 34022 19272
rect 33874 18828 33930 18864
rect 33874 18808 33876 18828
rect 33876 18808 33928 18828
rect 33928 18808 33930 18828
rect 31758 15816 31814 15872
rect 30562 15020 30618 15056
rect 30562 15000 30564 15020
rect 30564 15000 30616 15020
rect 30616 15000 30618 15020
rect 29826 9696 29882 9752
rect 29826 9152 29882 9208
rect 29642 7520 29698 7576
rect 27342 4936 27398 4992
rect 23294 3984 23350 4040
rect 24214 3984 24270 4040
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 27618 4800 27674 4856
rect 28722 4528 28778 4584
rect 29826 4664 29882 4720
rect 30562 12280 30618 12336
rect 32770 13776 32826 13832
rect 30286 10240 30342 10296
rect 32770 11736 32826 11792
rect 32494 10260 32550 10296
rect 32494 10240 32496 10260
rect 32496 10240 32548 10260
rect 32548 10240 32550 10260
rect 31942 9696 31998 9752
rect 33782 13776 33838 13832
rect 34426 17992 34482 18048
rect 34150 15000 34206 15056
rect 34702 22208 34758 22264
rect 34610 18672 34666 18728
rect 34610 16224 34666 16280
rect 33966 12552 34022 12608
rect 34334 12552 34390 12608
rect 34058 12144 34114 12200
rect 32954 7520 33010 7576
rect 32862 7404 32918 7440
rect 32862 7384 32864 7404
rect 32864 7384 32916 7404
rect 32916 7384 32918 7404
rect 27802 3188 27858 3224
rect 27802 3168 27804 3188
rect 27804 3168 27856 3188
rect 27856 3168 27858 3188
rect 28078 3052 28134 3088
rect 28078 3032 28080 3052
rect 28080 3032 28132 3052
rect 28132 3032 28134 3052
rect 27710 2896 27766 2952
rect 27986 2796 27988 2816
rect 27988 2796 28040 2816
rect 28040 2796 28042 2816
rect 27986 2760 28042 2796
rect 31022 4564 31024 4584
rect 31024 4564 31076 4584
rect 31076 4564 31078 4584
rect 31022 4528 31078 4564
rect 32402 6024 32458 6080
rect 32218 4972 32220 4992
rect 32220 4972 32272 4992
rect 32272 4972 32274 4992
rect 32218 4936 32274 4972
rect 32770 4800 32826 4856
rect 32126 4684 32182 4720
rect 32126 4664 32128 4684
rect 32128 4664 32180 4684
rect 32180 4664 32182 4684
rect 34940 27226 34996 27228
rect 35020 27226 35076 27228
rect 35100 27226 35156 27228
rect 35180 27226 35236 27228
rect 34940 27174 34966 27226
rect 34966 27174 34996 27226
rect 35020 27174 35030 27226
rect 35030 27174 35076 27226
rect 35100 27174 35146 27226
rect 35146 27174 35156 27226
rect 35180 27174 35210 27226
rect 35210 27174 35236 27226
rect 34940 27172 34996 27174
rect 35020 27172 35076 27174
rect 35100 27172 35156 27174
rect 35180 27172 35236 27174
rect 35622 34584 35678 34640
rect 36726 38120 36782 38176
rect 36082 35808 36138 35864
rect 37186 35536 37242 35592
rect 38290 35264 38346 35320
rect 39394 34584 39450 34640
rect 35806 34448 35862 34504
rect 35622 33224 35678 33280
rect 35714 32000 35770 32056
rect 35346 27376 35402 27432
rect 35254 26560 35310 26616
rect 34940 26138 34996 26140
rect 35020 26138 35076 26140
rect 35100 26138 35156 26140
rect 35180 26138 35236 26140
rect 34940 26086 34966 26138
rect 34966 26086 34996 26138
rect 35020 26086 35030 26138
rect 35030 26086 35076 26138
rect 35100 26086 35146 26138
rect 35146 26086 35156 26138
rect 35180 26086 35210 26138
rect 35210 26086 35236 26138
rect 34940 26084 34996 26086
rect 35020 26084 35076 26086
rect 35100 26084 35156 26086
rect 35180 26084 35236 26086
rect 34940 25050 34996 25052
rect 35020 25050 35076 25052
rect 35100 25050 35156 25052
rect 35180 25050 35236 25052
rect 34940 24998 34966 25050
rect 34966 24998 34996 25050
rect 35020 24998 35030 25050
rect 35030 24998 35076 25050
rect 35100 24998 35146 25050
rect 35146 24998 35156 25050
rect 35180 24998 35210 25050
rect 35210 24998 35236 25050
rect 34940 24996 34996 24998
rect 35020 24996 35076 24998
rect 35100 24996 35156 24998
rect 35180 24996 35236 24998
rect 34940 23962 34996 23964
rect 35020 23962 35076 23964
rect 35100 23962 35156 23964
rect 35180 23962 35236 23964
rect 34940 23910 34966 23962
rect 34966 23910 34996 23962
rect 35020 23910 35030 23962
rect 35030 23910 35076 23962
rect 35100 23910 35146 23962
rect 35146 23910 35156 23962
rect 35180 23910 35210 23962
rect 35210 23910 35236 23962
rect 34940 23908 34996 23910
rect 35020 23908 35076 23910
rect 35100 23908 35156 23910
rect 35180 23908 35236 23910
rect 34940 22874 34996 22876
rect 35020 22874 35076 22876
rect 35100 22874 35156 22876
rect 35180 22874 35236 22876
rect 34940 22822 34966 22874
rect 34966 22822 34996 22874
rect 35020 22822 35030 22874
rect 35030 22822 35076 22874
rect 35100 22822 35146 22874
rect 35146 22822 35156 22874
rect 35180 22822 35210 22874
rect 35210 22822 35236 22874
rect 34940 22820 34996 22822
rect 35020 22820 35076 22822
rect 35100 22820 35156 22822
rect 35180 22820 35236 22822
rect 35622 30776 35678 30832
rect 35530 26560 35586 26616
rect 35530 24520 35586 24576
rect 35530 23432 35586 23488
rect 34940 21786 34996 21788
rect 35020 21786 35076 21788
rect 35100 21786 35156 21788
rect 35180 21786 35236 21788
rect 34940 21734 34966 21786
rect 34966 21734 34996 21786
rect 35020 21734 35030 21786
rect 35030 21734 35076 21786
rect 35100 21734 35146 21786
rect 35146 21734 35156 21786
rect 35180 21734 35210 21786
rect 35210 21734 35236 21786
rect 34940 21732 34996 21734
rect 35020 21732 35076 21734
rect 35100 21732 35156 21734
rect 35180 21732 35236 21734
rect 34940 20698 34996 20700
rect 35020 20698 35076 20700
rect 35100 20698 35156 20700
rect 35180 20698 35236 20700
rect 34940 20646 34966 20698
rect 34966 20646 34996 20698
rect 35020 20646 35030 20698
rect 35030 20646 35076 20698
rect 35100 20646 35146 20698
rect 35146 20646 35156 20698
rect 35180 20646 35210 20698
rect 35210 20646 35236 20698
rect 34940 20644 34996 20646
rect 35020 20644 35076 20646
rect 35100 20644 35156 20646
rect 35180 20644 35236 20646
rect 35346 20304 35402 20360
rect 35346 19760 35402 19816
rect 34940 19610 34996 19612
rect 35020 19610 35076 19612
rect 35100 19610 35156 19612
rect 35180 19610 35236 19612
rect 34940 19558 34966 19610
rect 34966 19558 34996 19610
rect 35020 19558 35030 19610
rect 35030 19558 35076 19610
rect 35100 19558 35146 19610
rect 35146 19558 35156 19610
rect 35180 19558 35210 19610
rect 35210 19558 35236 19610
rect 34940 19556 34996 19558
rect 35020 19556 35076 19558
rect 35100 19556 35156 19558
rect 35180 19556 35236 19558
rect 34940 18522 34996 18524
rect 35020 18522 35076 18524
rect 35100 18522 35156 18524
rect 35180 18522 35236 18524
rect 34940 18470 34966 18522
rect 34966 18470 34996 18522
rect 35020 18470 35030 18522
rect 35030 18470 35076 18522
rect 35100 18470 35146 18522
rect 35146 18470 35156 18522
rect 35180 18470 35210 18522
rect 35210 18470 35236 18522
rect 34940 18468 34996 18470
rect 35020 18468 35076 18470
rect 35100 18468 35156 18470
rect 35180 18468 35236 18470
rect 34940 17434 34996 17436
rect 35020 17434 35076 17436
rect 35100 17434 35156 17436
rect 35180 17434 35236 17436
rect 34940 17382 34966 17434
rect 34966 17382 34996 17434
rect 35020 17382 35030 17434
rect 35030 17382 35076 17434
rect 35100 17382 35146 17434
rect 35146 17382 35156 17434
rect 35180 17382 35210 17434
rect 35210 17382 35236 17434
rect 34940 17380 34996 17382
rect 35020 17380 35076 17382
rect 35100 17380 35156 17382
rect 35180 17380 35236 17382
rect 35530 22344 35586 22400
rect 35714 29552 35770 29608
rect 37002 26832 37058 26888
rect 36910 26016 36966 26072
rect 35622 21120 35678 21176
rect 35530 20440 35586 20496
rect 35622 20032 35678 20088
rect 37830 26560 37886 26616
rect 37094 19760 37150 19816
rect 35622 17448 35678 17504
rect 34940 16346 34996 16348
rect 35020 16346 35076 16348
rect 35100 16346 35156 16348
rect 35180 16346 35236 16348
rect 34940 16294 34966 16346
rect 34966 16294 34996 16346
rect 35020 16294 35030 16346
rect 35030 16294 35076 16346
rect 35100 16294 35146 16346
rect 35146 16294 35156 16346
rect 35180 16294 35210 16346
rect 35210 16294 35236 16346
rect 34940 16292 34996 16294
rect 35020 16292 35076 16294
rect 35100 16292 35156 16294
rect 35180 16292 35236 16294
rect 35438 16224 35494 16280
rect 35622 16088 35678 16144
rect 34940 15258 34996 15260
rect 35020 15258 35076 15260
rect 35100 15258 35156 15260
rect 35180 15258 35236 15260
rect 34940 15206 34966 15258
rect 34966 15206 34996 15258
rect 35020 15206 35030 15258
rect 35030 15206 35076 15258
rect 35100 15206 35146 15258
rect 35146 15206 35156 15258
rect 35180 15206 35210 15258
rect 35210 15206 35236 15258
rect 34940 15204 34996 15206
rect 35020 15204 35076 15206
rect 35100 15204 35156 15206
rect 35180 15204 35236 15206
rect 35622 15000 35678 15056
rect 34940 14170 34996 14172
rect 35020 14170 35076 14172
rect 35100 14170 35156 14172
rect 35180 14170 35236 14172
rect 34940 14118 34966 14170
rect 34966 14118 34996 14170
rect 35020 14118 35030 14170
rect 35030 14118 35076 14170
rect 35100 14118 35146 14170
rect 35146 14118 35156 14170
rect 35180 14118 35210 14170
rect 35210 14118 35236 14170
rect 34940 14116 34996 14118
rect 35020 14116 35076 14118
rect 35100 14116 35156 14118
rect 35180 14116 35236 14118
rect 34940 13082 34996 13084
rect 35020 13082 35076 13084
rect 35100 13082 35156 13084
rect 35180 13082 35236 13084
rect 34940 13030 34966 13082
rect 34966 13030 34996 13082
rect 35020 13030 35030 13082
rect 35030 13030 35076 13082
rect 35100 13030 35146 13082
rect 35146 13030 35156 13082
rect 35180 13030 35210 13082
rect 35210 13030 35236 13082
rect 34940 13028 34996 13030
rect 35020 13028 35076 13030
rect 35100 13028 35156 13030
rect 35180 13028 35236 13030
rect 34940 11994 34996 11996
rect 35020 11994 35076 11996
rect 35100 11994 35156 11996
rect 35180 11994 35236 11996
rect 34940 11942 34966 11994
rect 34966 11942 34996 11994
rect 35020 11942 35030 11994
rect 35030 11942 35076 11994
rect 35100 11942 35146 11994
rect 35146 11942 35156 11994
rect 35180 11942 35210 11994
rect 35210 11942 35236 11994
rect 34940 11940 34996 11942
rect 35020 11940 35076 11942
rect 35100 11940 35156 11942
rect 35180 11940 35236 11942
rect 35346 12416 35402 12472
rect 35346 11736 35402 11792
rect 34940 10906 34996 10908
rect 35020 10906 35076 10908
rect 35100 10906 35156 10908
rect 35180 10906 35236 10908
rect 34940 10854 34966 10906
rect 34966 10854 34996 10906
rect 35020 10854 35030 10906
rect 35030 10854 35076 10906
rect 35100 10854 35146 10906
rect 35146 10854 35156 10906
rect 35180 10854 35210 10906
rect 35210 10854 35236 10906
rect 34940 10852 34996 10854
rect 35020 10852 35076 10854
rect 35100 10852 35156 10854
rect 35180 10852 35236 10854
rect 34940 9818 34996 9820
rect 35020 9818 35076 9820
rect 35100 9818 35156 9820
rect 35180 9818 35236 9820
rect 34940 9766 34966 9818
rect 34966 9766 34996 9818
rect 35020 9766 35030 9818
rect 35030 9766 35076 9818
rect 35100 9766 35146 9818
rect 35146 9766 35156 9818
rect 35180 9766 35210 9818
rect 35210 9766 35236 9818
rect 34940 9764 34996 9766
rect 35020 9764 35076 9766
rect 35100 9764 35156 9766
rect 35180 9764 35236 9766
rect 34610 7384 34666 7440
rect 34940 8730 34996 8732
rect 35020 8730 35076 8732
rect 35100 8730 35156 8732
rect 35180 8730 35236 8732
rect 34940 8678 34966 8730
rect 34966 8678 34996 8730
rect 35020 8678 35030 8730
rect 35030 8678 35076 8730
rect 35100 8678 35146 8730
rect 35146 8678 35156 8730
rect 35180 8678 35210 8730
rect 35210 8678 35236 8730
rect 34940 8676 34996 8678
rect 35020 8676 35076 8678
rect 35100 8676 35156 8678
rect 35180 8676 35236 8678
rect 34940 7642 34996 7644
rect 35020 7642 35076 7644
rect 35100 7642 35156 7644
rect 35180 7642 35236 7644
rect 34940 7590 34966 7642
rect 34966 7590 34996 7642
rect 35020 7590 35030 7642
rect 35030 7590 35076 7642
rect 35100 7590 35146 7642
rect 35146 7590 35156 7642
rect 35180 7590 35210 7642
rect 35210 7590 35236 7642
rect 34940 7588 34996 7590
rect 35020 7588 35076 7590
rect 35100 7588 35156 7590
rect 35180 7588 35236 7590
rect 34702 6704 34758 6760
rect 33782 6316 33838 6352
rect 33782 6296 33784 6316
rect 33784 6296 33836 6316
rect 33836 6296 33838 6316
rect 34242 5652 34244 5672
rect 34244 5652 34296 5672
rect 34296 5652 34298 5672
rect 34242 5616 34298 5652
rect 34940 6554 34996 6556
rect 35020 6554 35076 6556
rect 35100 6554 35156 6556
rect 35180 6554 35236 6556
rect 34940 6502 34966 6554
rect 34966 6502 34996 6554
rect 35020 6502 35030 6554
rect 35030 6502 35076 6554
rect 35100 6502 35146 6554
rect 35146 6502 35156 6554
rect 35180 6502 35210 6554
rect 35210 6502 35236 6554
rect 34940 6500 34996 6502
rect 35020 6500 35076 6502
rect 35100 6500 35156 6502
rect 35180 6500 35236 6502
rect 34702 5208 34758 5264
rect 36542 12688 36598 12744
rect 35714 7792 35770 7848
rect 35438 6060 35440 6080
rect 35440 6060 35492 6080
rect 35492 6060 35494 6080
rect 35438 6024 35494 6060
rect 34940 5466 34996 5468
rect 35020 5466 35076 5468
rect 35100 5466 35156 5468
rect 35180 5466 35236 5468
rect 34940 5414 34966 5466
rect 34966 5414 34996 5466
rect 35020 5414 35030 5466
rect 35030 5414 35076 5466
rect 35100 5414 35146 5466
rect 35146 5414 35156 5466
rect 35180 5414 35210 5466
rect 35210 5414 35236 5466
rect 34940 5412 34996 5414
rect 35020 5412 35076 5414
rect 35100 5412 35156 5414
rect 35180 5412 35236 5414
rect 34242 4664 34298 4720
rect 34150 3884 34152 3904
rect 34152 3884 34204 3904
rect 34204 3884 34206 3904
rect 31574 3188 31630 3224
rect 31574 3168 31576 3188
rect 31576 3168 31628 3188
rect 31628 3168 31630 3188
rect 31942 2896 31998 2952
rect 32494 3460 32550 3496
rect 32494 3440 32496 3460
rect 32496 3440 32548 3460
rect 32548 3440 32550 3460
rect 33046 3440 33102 3496
rect 34150 3848 34206 3884
rect 34978 4564 34980 4584
rect 34980 4564 35032 4584
rect 35032 4564 35034 4584
rect 34978 4528 35034 4564
rect 34940 4378 34996 4380
rect 35020 4378 35076 4380
rect 35100 4378 35156 4380
rect 35180 4378 35236 4380
rect 34940 4326 34966 4378
rect 34966 4326 34996 4378
rect 35020 4326 35030 4378
rect 35030 4326 35076 4378
rect 35100 4326 35146 4378
rect 35146 4326 35156 4378
rect 35180 4326 35210 4378
rect 35210 4326 35236 4378
rect 34940 4324 34996 4326
rect 35020 4324 35076 4326
rect 35100 4324 35156 4326
rect 35180 4324 35236 4326
rect 33690 3052 33746 3088
rect 33690 3032 33692 3052
rect 33692 3032 33744 3052
rect 33744 3032 33746 3052
rect 34940 3290 34996 3292
rect 35020 3290 35076 3292
rect 35100 3290 35156 3292
rect 35180 3290 35236 3292
rect 34940 3238 34966 3290
rect 34966 3238 34996 3290
rect 35020 3238 35030 3290
rect 35030 3238 35076 3290
rect 35100 3238 35146 3290
rect 35146 3238 35156 3290
rect 35180 3238 35210 3290
rect 35210 3238 35236 3290
rect 34940 3236 34996 3238
rect 35020 3236 35076 3238
rect 35100 3236 35156 3238
rect 35180 3236 35236 3238
rect 34610 2796 34612 2816
rect 34612 2796 34664 2816
rect 34664 2796 34666 2816
rect 34610 2760 34666 2796
rect 34940 2202 34996 2204
rect 35020 2202 35076 2204
rect 35100 2202 35156 2204
rect 35180 2202 35236 2204
rect 34940 2150 34966 2202
rect 34966 2150 34996 2202
rect 35020 2150 35030 2202
rect 35030 2150 35076 2202
rect 35100 2150 35146 2202
rect 35146 2150 35156 2202
rect 35180 2150 35210 2202
rect 35210 2150 35236 2202
rect 34940 2148 34996 2150
rect 35020 2148 35076 2150
rect 35100 2148 35156 2150
rect 35180 2148 35236 2150
rect 35530 4528 35586 4584
rect 35898 4664 35954 4720
rect 35806 4120 35862 4176
rect 35898 3848 35954 3904
rect 35714 2896 35770 2952
rect 35346 1672 35402 1728
rect 36818 13776 36874 13832
rect 37002 13912 37058 13968
rect 36910 10240 36966 10296
rect 36818 9152 36874 9208
rect 36634 9016 36690 9072
rect 37094 11464 37150 11520
rect 37278 6332 37280 6352
rect 37280 6332 37332 6352
rect 37332 6332 37334 6352
rect 37278 6296 37334 6332
rect 36634 5616 36690 5672
rect 36450 4528 36506 4584
rect 36634 3440 36690 3496
rect 36358 584 36414 640
<< metal3 >>
rect 35617 39402 35683 39405
rect 39520 39402 40000 39432
rect 35617 39400 40000 39402
rect 35617 39344 35622 39400
rect 35678 39344 40000 39400
rect 35617 39342 40000 39344
rect 35617 39339 35683 39342
rect 39520 39312 40000 39342
rect 36721 38178 36787 38181
rect 39520 38178 40000 38208
rect 36721 38176 40000 38178
rect 36721 38120 36726 38176
rect 36782 38120 40000 38176
rect 36721 38118 40000 38120
rect 36721 38115 36787 38118
rect 39520 38088 40000 38118
rect 19568 37568 19888 37569
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 37503 19888 37504
rect 4208 37024 4528 37025
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 34928 37024 35248 37025
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36959 35248 36960
rect 35801 36954 35867 36957
rect 39520 36954 40000 36984
rect 35801 36952 40000 36954
rect 35801 36896 35806 36952
rect 35862 36896 40000 36952
rect 35801 36894 40000 36896
rect 35801 36891 35867 36894
rect 39520 36864 40000 36894
rect 19568 36480 19888 36481
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 36415 19888 36416
rect 3141 36138 3207 36141
rect 18045 36138 18111 36141
rect 3141 36136 18111 36138
rect 3141 36080 3146 36136
rect 3202 36080 18050 36136
rect 18106 36080 18111 36136
rect 3141 36078 18111 36080
rect 3141 36075 3207 36078
rect 18045 36075 18111 36078
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 34928 35936 35248 35937
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 35871 35248 35872
rect 7465 35866 7531 35869
rect 11605 35866 11671 35869
rect 7465 35864 11671 35866
rect 7465 35808 7470 35864
rect 7526 35808 11610 35864
rect 11666 35808 11671 35864
rect 7465 35806 11671 35808
rect 7465 35803 7531 35806
rect 11605 35803 11671 35806
rect 11881 35866 11947 35869
rect 13905 35866 13971 35869
rect 11881 35864 13971 35866
rect 11881 35808 11886 35864
rect 11942 35808 13910 35864
rect 13966 35808 13971 35864
rect 11881 35806 13971 35808
rect 11881 35803 11947 35806
rect 13905 35803 13971 35806
rect 24894 35804 24900 35868
rect 24964 35866 24970 35868
rect 36077 35866 36143 35869
rect 24964 35806 27538 35866
rect 24964 35804 24970 35806
rect 6637 35732 6703 35733
rect 6637 35730 6684 35732
rect 6592 35728 6684 35730
rect 6592 35672 6642 35728
rect 6592 35670 6684 35672
rect 6637 35668 6684 35670
rect 6748 35668 6754 35732
rect 6821 35730 6887 35733
rect 10501 35730 10567 35733
rect 6821 35728 10567 35730
rect 6821 35672 6826 35728
rect 6882 35672 10506 35728
rect 10562 35672 10567 35728
rect 6821 35670 10567 35672
rect 6637 35667 6703 35668
rect 6821 35667 6887 35670
rect 10501 35667 10567 35670
rect 14457 35730 14523 35733
rect 27245 35730 27311 35733
rect 14457 35728 27311 35730
rect 14457 35672 14462 35728
rect 14518 35672 27250 35728
rect 27306 35672 27311 35728
rect 14457 35670 27311 35672
rect 27478 35730 27538 35806
rect 35390 35864 36143 35866
rect 35390 35808 36082 35864
rect 36138 35808 36143 35864
rect 35390 35806 36143 35808
rect 35390 35730 35450 35806
rect 36077 35803 36143 35806
rect 39520 35730 40000 35760
rect 27478 35670 35450 35730
rect 37782 35670 40000 35730
rect 14457 35667 14523 35670
rect 27245 35667 27311 35670
rect 8569 35594 8635 35597
rect 25129 35594 25195 35597
rect 37181 35594 37247 35597
rect 8569 35592 37247 35594
rect 8569 35536 8574 35592
rect 8630 35536 25134 35592
rect 25190 35536 37186 35592
rect 37242 35536 37247 35592
rect 8569 35534 37247 35536
rect 8569 35531 8635 35534
rect 25129 35531 25195 35534
rect 37181 35531 37247 35534
rect 4981 35460 5047 35461
rect 4981 35458 5028 35460
rect 4936 35456 5028 35458
rect 4936 35400 4986 35456
rect 4936 35398 5028 35400
rect 4981 35396 5028 35398
rect 5092 35396 5098 35460
rect 5533 35458 5599 35461
rect 18137 35458 18203 35461
rect 5533 35456 18203 35458
rect 5533 35400 5538 35456
rect 5594 35400 18142 35456
rect 18198 35400 18203 35456
rect 5533 35398 18203 35400
rect 4981 35395 5047 35396
rect 5533 35395 5599 35398
rect 18137 35395 18203 35398
rect 35709 35458 35775 35461
rect 37782 35458 37842 35670
rect 39520 35640 40000 35670
rect 35709 35456 37842 35458
rect 35709 35400 35714 35456
rect 35770 35400 37842 35456
rect 35709 35398 37842 35400
rect 35709 35395 35775 35398
rect 19568 35392 19888 35393
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 35327 19888 35328
rect 1393 35322 1459 35325
rect 10869 35322 10935 35325
rect 1393 35320 10935 35322
rect 1393 35264 1398 35320
rect 1454 35264 10874 35320
rect 10930 35264 10935 35320
rect 1393 35262 10935 35264
rect 1393 35259 1459 35262
rect 10869 35259 10935 35262
rect 20662 35260 20668 35324
rect 20732 35322 20738 35324
rect 21398 35322 21404 35324
rect 20732 35262 21404 35322
rect 20732 35260 20738 35262
rect 21398 35260 21404 35262
rect 21468 35322 21474 35324
rect 33869 35322 33935 35325
rect 21468 35320 33935 35322
rect 21468 35264 33874 35320
rect 33930 35264 33935 35320
rect 21468 35262 33935 35264
rect 21468 35260 21474 35262
rect 33869 35259 33935 35262
rect 35525 35322 35591 35325
rect 38285 35322 38351 35325
rect 35525 35320 38351 35322
rect 35525 35264 35530 35320
rect 35586 35264 38290 35320
rect 38346 35264 38351 35320
rect 35525 35262 38351 35264
rect 35525 35259 35591 35262
rect 38285 35259 38351 35262
rect 6821 35186 6887 35189
rect 9397 35186 9463 35189
rect 6821 35184 9463 35186
rect 6821 35128 6826 35184
rect 6882 35128 9402 35184
rect 9458 35128 9463 35184
rect 6821 35126 9463 35128
rect 6821 35123 6887 35126
rect 9397 35123 9463 35126
rect 13629 35186 13695 35189
rect 29453 35186 29519 35189
rect 13629 35184 29519 35186
rect 13629 35128 13634 35184
rect 13690 35128 29458 35184
rect 29514 35128 29519 35184
rect 13629 35126 29519 35128
rect 13629 35123 13695 35126
rect 29453 35123 29519 35126
rect 2037 35050 2103 35053
rect 10869 35050 10935 35053
rect 30557 35050 30623 35053
rect 2037 35048 7666 35050
rect 2037 34992 2042 35048
rect 2098 34992 7666 35048
rect 2037 34990 7666 34992
rect 2037 34987 2103 34990
rect 7606 34914 7666 34990
rect 10869 35048 30623 35050
rect 10869 34992 10874 35048
rect 10930 34992 30562 35048
rect 30618 34992 30623 35048
rect 10869 34990 30623 34992
rect 10869 34987 10935 34990
rect 30557 34987 30623 34990
rect 13629 34914 13695 34917
rect 7606 34912 13695 34914
rect 7606 34856 13634 34912
rect 13690 34856 13695 34912
rect 7606 34854 13695 34856
rect 13629 34851 13695 34854
rect 18137 34914 18203 34917
rect 19149 34914 19215 34917
rect 34789 34914 34855 34917
rect 18137 34912 34855 34914
rect 18137 34856 18142 34912
rect 18198 34856 19154 34912
rect 19210 34856 34794 34912
rect 34850 34856 34855 34912
rect 18137 34854 34855 34856
rect 18137 34851 18203 34854
rect 19149 34851 19215 34854
rect 34789 34851 34855 34854
rect 4208 34848 4528 34849
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 34928 34848 35248 34849
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 34783 35248 34784
rect 8845 34778 8911 34781
rect 12709 34778 12775 34781
rect 8845 34776 12775 34778
rect 8845 34720 8850 34776
rect 8906 34720 12714 34776
rect 12770 34720 12775 34776
rect 8845 34718 12775 34720
rect 8845 34715 8911 34718
rect 12709 34715 12775 34718
rect 20621 34778 20687 34781
rect 22737 34778 22803 34781
rect 20621 34776 22803 34778
rect 20621 34720 20626 34776
rect 20682 34720 22742 34776
rect 22798 34720 22803 34776
rect 20621 34718 22803 34720
rect 20621 34715 20687 34718
rect 22737 34715 22803 34718
rect 24894 34716 24900 34780
rect 24964 34778 24970 34780
rect 25037 34778 25103 34781
rect 24964 34776 25103 34778
rect 24964 34720 25042 34776
rect 25098 34720 25103 34776
rect 24964 34718 25103 34720
rect 24964 34716 24970 34718
rect 25037 34715 25103 34718
rect 5073 34642 5139 34645
rect 7465 34642 7531 34645
rect 5073 34640 7531 34642
rect 5073 34584 5078 34640
rect 5134 34584 7470 34640
rect 7526 34584 7531 34640
rect 5073 34582 7531 34584
rect 5073 34579 5139 34582
rect 7465 34579 7531 34582
rect 18045 34642 18111 34645
rect 31661 34642 31727 34645
rect 18045 34640 31727 34642
rect 18045 34584 18050 34640
rect 18106 34584 31666 34640
rect 31722 34584 31727 34640
rect 18045 34582 31727 34584
rect 18045 34579 18111 34582
rect 31661 34579 31727 34582
rect 35617 34642 35683 34645
rect 39389 34642 39455 34645
rect 35617 34640 39455 34642
rect 35617 34584 35622 34640
rect 35678 34584 39394 34640
rect 39450 34584 39455 34640
rect 35617 34582 39455 34584
rect 35617 34579 35683 34582
rect 39389 34579 39455 34582
rect 21909 34506 21975 34509
rect 23657 34506 23723 34509
rect 21909 34504 23723 34506
rect 21909 34448 21914 34504
rect 21970 34448 23662 34504
rect 23718 34448 23723 34504
rect 21909 34446 23723 34448
rect 21909 34443 21975 34446
rect 23657 34443 23723 34446
rect 35801 34506 35867 34509
rect 39520 34506 40000 34536
rect 35801 34504 40000 34506
rect 35801 34448 35806 34504
rect 35862 34448 40000 34504
rect 35801 34446 40000 34448
rect 35801 34443 35867 34446
rect 39520 34416 40000 34446
rect 19568 34304 19888 34305
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 34239 19888 34240
rect 4061 33962 4127 33965
rect 15837 33962 15903 33965
rect 32765 33962 32831 33965
rect 4061 33960 32831 33962
rect 4061 33904 4066 33960
rect 4122 33904 15842 33960
rect 15898 33904 32770 33960
rect 32826 33904 32831 33960
rect 4061 33902 32831 33904
rect 4061 33899 4127 33902
rect 15837 33899 15903 33902
rect 32765 33899 32831 33902
rect 21357 33826 21423 33829
rect 24117 33826 24183 33829
rect 21357 33824 24183 33826
rect 21357 33768 21362 33824
rect 21418 33768 24122 33824
rect 24178 33768 24183 33824
rect 21357 33766 24183 33768
rect 21357 33763 21423 33766
rect 24117 33763 24183 33766
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 34928 33760 35248 33761
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 33695 35248 33696
rect 0 33328 480 33448
rect 12985 33282 13051 33285
rect 13353 33282 13419 33285
rect 15285 33282 15351 33285
rect 12985 33280 15351 33282
rect 12985 33224 12990 33280
rect 13046 33224 13358 33280
rect 13414 33224 15290 33280
rect 15346 33224 15351 33280
rect 12985 33222 15351 33224
rect 12985 33219 13051 33222
rect 13353 33219 13419 33222
rect 15285 33219 15351 33222
rect 17769 33282 17835 33285
rect 19333 33282 19399 33285
rect 17769 33280 19399 33282
rect 17769 33224 17774 33280
rect 17830 33224 19338 33280
rect 19394 33224 19399 33280
rect 17769 33222 19399 33224
rect 17769 33219 17835 33222
rect 19333 33219 19399 33222
rect 35617 33282 35683 33285
rect 39520 33282 40000 33312
rect 35617 33280 40000 33282
rect 35617 33224 35622 33280
rect 35678 33224 40000 33280
rect 35617 33222 40000 33224
rect 35617 33219 35683 33222
rect 19568 33216 19888 33217
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 39520 33192 40000 33222
rect 19568 33151 19888 33152
rect 8017 33146 8083 33149
rect 10133 33146 10199 33149
rect 8017 33144 10199 33146
rect 8017 33088 8022 33144
rect 8078 33088 10138 33144
rect 10194 33088 10199 33144
rect 8017 33086 10199 33088
rect 8017 33083 8083 33086
rect 10133 33083 10199 33086
rect 11605 33146 11671 33149
rect 14549 33146 14615 33149
rect 11605 33144 14615 33146
rect 11605 33088 11610 33144
rect 11666 33088 14554 33144
rect 14610 33088 14615 33144
rect 11605 33086 14615 33088
rect 11605 33083 11671 33086
rect 14549 33083 14615 33086
rect 21449 33146 21515 33149
rect 23933 33146 23999 33149
rect 21449 33144 23999 33146
rect 21449 33088 21454 33144
rect 21510 33088 23938 33144
rect 23994 33088 23999 33144
rect 21449 33086 23999 33088
rect 21449 33083 21515 33086
rect 23933 33083 23999 33086
rect 20161 33010 20227 33013
rect 24669 33010 24735 33013
rect 20161 33008 24735 33010
rect 20161 32952 20166 33008
rect 20222 32952 24674 33008
rect 24730 32952 24735 33008
rect 20161 32950 24735 32952
rect 20161 32947 20227 32950
rect 24669 32947 24735 32950
rect 10869 32738 10935 32741
rect 12801 32738 12867 32741
rect 14457 32738 14523 32741
rect 10869 32736 14523 32738
rect 10869 32680 10874 32736
rect 10930 32680 12806 32736
rect 12862 32680 14462 32736
rect 14518 32680 14523 32736
rect 10869 32678 14523 32680
rect 10869 32675 10935 32678
rect 12801 32675 12867 32678
rect 14457 32675 14523 32678
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 34928 32672 35248 32673
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 32607 35248 32608
rect 16021 32602 16087 32605
rect 30097 32602 30163 32605
rect 16021 32600 30163 32602
rect 16021 32544 16026 32600
rect 16082 32544 30102 32600
rect 30158 32544 30163 32600
rect 16021 32542 30163 32544
rect 16021 32539 16087 32542
rect 30097 32539 30163 32542
rect 9489 32466 9555 32469
rect 13813 32466 13879 32469
rect 15101 32466 15167 32469
rect 17125 32466 17191 32469
rect 9489 32464 13879 32466
rect 9489 32408 9494 32464
rect 9550 32408 13818 32464
rect 13874 32408 13879 32464
rect 9489 32406 13879 32408
rect 9489 32403 9555 32406
rect 13813 32403 13879 32406
rect 14782 32464 17191 32466
rect 14782 32408 15106 32464
rect 15162 32408 17130 32464
rect 17186 32408 17191 32464
rect 14782 32406 17191 32408
rect 11329 32330 11395 32333
rect 14782 32330 14842 32406
rect 15101 32403 15167 32406
rect 17125 32403 17191 32406
rect 11329 32328 14842 32330
rect 11329 32272 11334 32328
rect 11390 32272 14842 32328
rect 11329 32270 14842 32272
rect 11329 32267 11395 32270
rect 19568 32128 19888 32129
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 32063 19888 32064
rect 2865 32058 2931 32061
rect 4981 32058 5047 32061
rect 2865 32056 5047 32058
rect 2865 32000 2870 32056
rect 2926 32000 4986 32056
rect 5042 32000 5047 32056
rect 2865 31998 5047 32000
rect 2865 31995 2931 31998
rect 4981 31995 5047 31998
rect 35709 32058 35775 32061
rect 39520 32058 40000 32088
rect 35709 32056 40000 32058
rect 35709 32000 35714 32056
rect 35770 32000 40000 32056
rect 35709 31998 40000 32000
rect 35709 31995 35775 31998
rect 39520 31968 40000 31998
rect 13169 31650 13235 31653
rect 17033 31650 17099 31653
rect 13169 31648 17099 31650
rect 13169 31592 13174 31648
rect 13230 31592 17038 31648
rect 17094 31592 17099 31648
rect 13169 31590 17099 31592
rect 13169 31587 13235 31590
rect 17033 31587 17099 31590
rect 4208 31584 4528 31585
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 34928 31584 35248 31585
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 31519 35248 31520
rect 14273 31514 14339 31517
rect 16113 31514 16179 31517
rect 14273 31512 16179 31514
rect 14273 31456 14278 31512
rect 14334 31456 16118 31512
rect 16174 31456 16179 31512
rect 14273 31454 16179 31456
rect 14273 31451 14339 31454
rect 16113 31451 16179 31454
rect 3325 31106 3391 31109
rect 5809 31106 5875 31109
rect 3325 31104 5875 31106
rect 3325 31048 3330 31104
rect 3386 31048 5814 31104
rect 5870 31048 5875 31104
rect 3325 31046 5875 31048
rect 3325 31043 3391 31046
rect 5809 31043 5875 31046
rect 10409 31106 10475 31109
rect 13813 31106 13879 31109
rect 10409 31104 13879 31106
rect 10409 31048 10414 31104
rect 10470 31048 13818 31104
rect 13874 31048 13879 31104
rect 10409 31046 13879 31048
rect 10409 31043 10475 31046
rect 13813 31043 13879 31046
rect 24669 31106 24735 31109
rect 26509 31106 26575 31109
rect 24669 31104 26575 31106
rect 24669 31048 24674 31104
rect 24730 31048 26514 31104
rect 26570 31048 26575 31104
rect 24669 31046 26575 31048
rect 24669 31043 24735 31046
rect 26509 31043 26575 31046
rect 19568 31040 19888 31041
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 30975 19888 30976
rect 35617 30834 35683 30837
rect 39520 30834 40000 30864
rect 35617 30832 40000 30834
rect 35617 30776 35622 30832
rect 35678 30776 40000 30832
rect 35617 30774 40000 30776
rect 35617 30771 35683 30774
rect 39520 30744 40000 30774
rect 4208 30496 4528 30497
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 34928 30496 35248 30497
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 30431 35248 30432
rect 15929 30426 15995 30429
rect 18505 30426 18571 30429
rect 15929 30424 18571 30426
rect 15929 30368 15934 30424
rect 15990 30368 18510 30424
rect 18566 30368 18571 30424
rect 15929 30366 18571 30368
rect 15929 30363 15995 30366
rect 18505 30363 18571 30366
rect 11881 30290 11947 30293
rect 15009 30290 15075 30293
rect 11881 30288 15075 30290
rect 11881 30232 11886 30288
rect 11942 30232 15014 30288
rect 15070 30232 15075 30288
rect 11881 30230 15075 30232
rect 11881 30227 11947 30230
rect 15009 30227 15075 30230
rect 15285 30290 15351 30293
rect 16941 30290 17007 30293
rect 15285 30288 17007 30290
rect 15285 30232 15290 30288
rect 15346 30232 16946 30288
rect 17002 30232 17007 30288
rect 15285 30230 17007 30232
rect 15285 30227 15351 30230
rect 16941 30227 17007 30230
rect 10409 30018 10475 30021
rect 12617 30018 12683 30021
rect 10409 30016 12683 30018
rect 10409 29960 10414 30016
rect 10470 29960 12622 30016
rect 12678 29960 12683 30016
rect 10409 29958 12683 29960
rect 10409 29955 10475 29958
rect 12617 29955 12683 29958
rect 19568 29952 19888 29953
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 29887 19888 29888
rect 1669 29746 1735 29749
rect 4153 29746 4219 29749
rect 1669 29744 4219 29746
rect 1669 29688 1674 29744
rect 1730 29688 4158 29744
rect 4214 29688 4219 29744
rect 1669 29686 4219 29688
rect 1669 29683 1735 29686
rect 4153 29683 4219 29686
rect 23565 29746 23631 29749
rect 26877 29746 26943 29749
rect 23565 29744 26943 29746
rect 23565 29688 23570 29744
rect 23626 29688 26882 29744
rect 26938 29688 26943 29744
rect 23565 29686 26943 29688
rect 23565 29683 23631 29686
rect 26877 29683 26943 29686
rect 35709 29610 35775 29613
rect 39520 29610 40000 29640
rect 35709 29608 40000 29610
rect 35709 29552 35714 29608
rect 35770 29552 40000 29608
rect 35709 29550 40000 29552
rect 35709 29547 35775 29550
rect 39520 29520 40000 29550
rect 4208 29408 4528 29409
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 34928 29408 35248 29409
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 29343 35248 29344
rect 12985 29338 13051 29341
rect 16389 29338 16455 29341
rect 12985 29336 16455 29338
rect 12985 29280 12990 29336
rect 13046 29280 16394 29336
rect 16450 29280 16455 29336
rect 12985 29278 16455 29280
rect 12985 29275 13051 29278
rect 16389 29275 16455 29278
rect 7925 29202 7991 29205
rect 9673 29202 9739 29205
rect 7925 29200 9739 29202
rect 7925 29144 7930 29200
rect 7986 29144 9678 29200
rect 9734 29144 9739 29200
rect 7925 29142 9739 29144
rect 7925 29139 7991 29142
rect 9673 29139 9739 29142
rect 15745 29202 15811 29205
rect 18137 29202 18203 29205
rect 15745 29200 18203 29202
rect 15745 29144 15750 29200
rect 15806 29144 18142 29200
rect 18198 29144 18203 29200
rect 15745 29142 18203 29144
rect 15745 29139 15811 29142
rect 18137 29139 18203 29142
rect 15837 29066 15903 29069
rect 18045 29066 18111 29069
rect 15837 29064 18111 29066
rect 15837 29008 15842 29064
rect 15898 29008 18050 29064
rect 18106 29008 18111 29064
rect 15837 29006 18111 29008
rect 15837 29003 15903 29006
rect 18045 29003 18111 29006
rect 31569 28930 31635 28933
rect 33501 28930 33567 28933
rect 31569 28928 33567 28930
rect 31569 28872 31574 28928
rect 31630 28872 33506 28928
rect 33562 28872 33567 28928
rect 31569 28870 33567 28872
rect 31569 28867 31635 28870
rect 33501 28867 33567 28870
rect 19568 28864 19888 28865
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 28799 19888 28800
rect 8017 28658 8083 28661
rect 9673 28658 9739 28661
rect 8017 28656 9739 28658
rect 8017 28600 8022 28656
rect 8078 28600 9678 28656
rect 9734 28600 9739 28656
rect 8017 28598 9739 28600
rect 8017 28595 8083 28598
rect 9673 28595 9739 28598
rect 18965 28522 19031 28525
rect 19885 28522 19951 28525
rect 22277 28522 22343 28525
rect 18965 28520 22343 28522
rect 18965 28464 18970 28520
rect 19026 28464 19890 28520
rect 19946 28464 22282 28520
rect 22338 28464 22343 28520
rect 18965 28462 22343 28464
rect 18965 28459 19031 28462
rect 19885 28459 19951 28462
rect 22277 28459 22343 28462
rect 30005 28386 30071 28389
rect 31937 28386 32003 28389
rect 39520 28386 40000 28416
rect 30005 28384 32003 28386
rect 30005 28328 30010 28384
rect 30066 28328 31942 28384
rect 31998 28328 32003 28384
rect 30005 28326 32003 28328
rect 30005 28323 30071 28326
rect 31937 28323 32003 28326
rect 35574 28326 40000 28386
rect 4208 28320 4528 28321
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 34928 28320 35248 28321
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 28255 35248 28256
rect 21398 28188 21404 28252
rect 21468 28250 21474 28252
rect 21633 28250 21699 28253
rect 21468 28248 21699 28250
rect 21468 28192 21638 28248
rect 21694 28192 21699 28248
rect 21468 28190 21699 28192
rect 21468 28188 21474 28190
rect 21633 28187 21699 28190
rect 34605 28114 34671 28117
rect 35574 28114 35634 28326
rect 39520 28296 40000 28326
rect 34605 28112 35634 28114
rect 34605 28056 34610 28112
rect 34666 28056 35634 28112
rect 34605 28054 35634 28056
rect 34605 28051 34671 28054
rect 19568 27776 19888 27777
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 27711 19888 27712
rect 24117 27706 24183 27709
rect 26969 27706 27035 27709
rect 24117 27704 27035 27706
rect 24117 27648 24122 27704
rect 24178 27648 26974 27704
rect 27030 27648 27035 27704
rect 24117 27646 27035 27648
rect 24117 27643 24183 27646
rect 26969 27643 27035 27646
rect 3969 27434 4035 27437
rect 5717 27434 5783 27437
rect 3969 27432 5783 27434
rect 3969 27376 3974 27432
rect 4030 27376 5722 27432
rect 5778 27376 5783 27432
rect 3969 27374 5783 27376
rect 3969 27371 4035 27374
rect 5717 27371 5783 27374
rect 25497 27434 25563 27437
rect 27889 27434 27955 27437
rect 25497 27432 27955 27434
rect 25497 27376 25502 27432
rect 25558 27376 27894 27432
rect 27950 27376 27955 27432
rect 25497 27374 27955 27376
rect 25497 27371 25563 27374
rect 27889 27371 27955 27374
rect 34646 27372 34652 27436
rect 34716 27434 34722 27436
rect 35341 27434 35407 27437
rect 34716 27432 35407 27434
rect 34716 27376 35346 27432
rect 35402 27376 35407 27432
rect 34716 27374 35407 27376
rect 34716 27372 34722 27374
rect 35341 27371 35407 27374
rect 39520 27298 40000 27328
rect 35390 27238 40000 27298
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 34928 27232 35248 27233
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 27167 35248 27168
rect 18689 27162 18755 27165
rect 20529 27162 20595 27165
rect 18689 27160 20595 27162
rect 18689 27104 18694 27160
rect 18750 27104 20534 27160
rect 20590 27104 20595 27160
rect 18689 27102 20595 27104
rect 18689 27099 18755 27102
rect 20529 27099 20595 27102
rect 13721 27026 13787 27029
rect 15377 27026 15443 27029
rect 13721 27024 15443 27026
rect 13721 26968 13726 27024
rect 13782 26968 15382 27024
rect 15438 26968 15443 27024
rect 13721 26966 15443 26968
rect 13721 26963 13787 26966
rect 15377 26963 15443 26966
rect 34053 27026 34119 27029
rect 35390 27026 35450 27238
rect 39520 27208 40000 27238
rect 34053 27024 35450 27026
rect 34053 26968 34058 27024
rect 34114 26968 35450 27024
rect 34053 26966 35450 26968
rect 34053 26963 34119 26966
rect 34237 26890 34303 26893
rect 36997 26890 37063 26893
rect 34237 26888 37063 26890
rect 34237 26832 34242 26888
rect 34298 26832 37002 26888
rect 37058 26832 37063 26888
rect 34237 26830 37063 26832
rect 34237 26827 34303 26830
rect 36997 26827 37063 26830
rect 6453 26754 6519 26757
rect 8845 26754 8911 26757
rect 6453 26752 8911 26754
rect 6453 26696 6458 26752
rect 6514 26696 8850 26752
rect 8906 26696 8911 26752
rect 6453 26694 8911 26696
rect 6453 26691 6519 26694
rect 8845 26691 8911 26694
rect 19568 26688 19888 26689
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 26623 19888 26624
rect 29177 26618 29243 26621
rect 32121 26618 32187 26621
rect 29177 26616 32187 26618
rect 29177 26560 29182 26616
rect 29238 26560 32126 26616
rect 32182 26560 32187 26616
rect 29177 26558 32187 26560
rect 29177 26555 29243 26558
rect 32121 26555 32187 26558
rect 35249 26618 35315 26621
rect 35382 26618 35388 26620
rect 35249 26616 35388 26618
rect 35249 26560 35254 26616
rect 35310 26560 35388 26616
rect 35249 26558 35388 26560
rect 35249 26555 35315 26558
rect 35382 26556 35388 26558
rect 35452 26556 35458 26620
rect 35525 26618 35591 26621
rect 37825 26618 37891 26621
rect 35525 26616 37891 26618
rect 35525 26560 35530 26616
rect 35586 26560 37830 26616
rect 37886 26560 37891 26616
rect 35525 26558 37891 26560
rect 35525 26555 35591 26558
rect 37825 26555 37891 26558
rect 29361 26482 29427 26485
rect 34237 26482 34303 26485
rect 29361 26480 34303 26482
rect 29361 26424 29366 26480
rect 29422 26424 34242 26480
rect 34298 26424 34303 26480
rect 29361 26422 34303 26424
rect 29361 26419 29427 26422
rect 34237 26419 34303 26422
rect 30189 26346 30255 26349
rect 31937 26346 32003 26349
rect 30189 26344 32003 26346
rect 30189 26288 30194 26344
rect 30250 26288 31942 26344
rect 31998 26288 32003 26344
rect 30189 26286 32003 26288
rect 30189 26283 30255 26286
rect 31937 26283 32003 26286
rect 24393 26210 24459 26213
rect 26233 26210 26299 26213
rect 24393 26208 26299 26210
rect 24393 26152 24398 26208
rect 24454 26152 26238 26208
rect 26294 26152 26299 26208
rect 24393 26150 26299 26152
rect 24393 26147 24459 26150
rect 26233 26147 26299 26150
rect 4208 26144 4528 26145
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 34928 26144 35248 26145
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 26079 35248 26080
rect 36905 26074 36971 26077
rect 39520 26074 40000 26104
rect 36905 26072 40000 26074
rect 36905 26016 36910 26072
rect 36966 26016 40000 26072
rect 36905 26014 40000 26016
rect 36905 26011 36971 26014
rect 39520 25984 40000 26014
rect 20989 25802 21055 25805
rect 22001 25802 22067 25805
rect 23473 25802 23539 25805
rect 20989 25800 23539 25802
rect 20989 25744 20994 25800
rect 21050 25744 22006 25800
rect 22062 25744 23478 25800
rect 23534 25744 23539 25800
rect 20989 25742 23539 25744
rect 20989 25739 21055 25742
rect 22001 25739 22067 25742
rect 23473 25739 23539 25742
rect 13261 25666 13327 25669
rect 14549 25666 14615 25669
rect 13261 25664 14615 25666
rect 13261 25608 13266 25664
rect 13322 25608 14554 25664
rect 14610 25608 14615 25664
rect 13261 25606 14615 25608
rect 13261 25603 13327 25606
rect 14549 25603 14615 25606
rect 28901 25666 28967 25669
rect 31937 25666 32003 25669
rect 28901 25664 32003 25666
rect 28901 25608 28906 25664
rect 28962 25608 31942 25664
rect 31998 25608 32003 25664
rect 28901 25606 32003 25608
rect 28901 25603 28967 25606
rect 31937 25603 32003 25606
rect 19568 25600 19888 25601
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25535 19888 25536
rect 11881 25530 11947 25533
rect 13169 25530 13235 25533
rect 13813 25530 13879 25533
rect 11881 25528 13879 25530
rect 11881 25472 11886 25528
rect 11942 25472 13174 25528
rect 13230 25472 13818 25528
rect 13874 25472 13879 25528
rect 11881 25470 13879 25472
rect 11881 25467 11947 25470
rect 13169 25467 13235 25470
rect 13813 25467 13879 25470
rect 15653 25530 15719 25533
rect 18413 25530 18479 25533
rect 15653 25528 18479 25530
rect 15653 25472 15658 25528
rect 15714 25472 18418 25528
rect 18474 25472 18479 25528
rect 15653 25470 18479 25472
rect 15653 25467 15719 25470
rect 18413 25467 18479 25470
rect 26601 25530 26667 25533
rect 29361 25530 29427 25533
rect 26601 25528 29427 25530
rect 26601 25472 26606 25528
rect 26662 25472 29366 25528
rect 29422 25472 29427 25528
rect 26601 25470 29427 25472
rect 26601 25467 26667 25470
rect 29361 25467 29427 25470
rect 4208 25056 4528 25057
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 34928 25056 35248 25057
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 24991 35248 24992
rect 39520 24850 40000 24880
rect 35574 24790 40000 24850
rect 10133 24714 10199 24717
rect 13813 24714 13879 24717
rect 10133 24712 13879 24714
rect 10133 24656 10138 24712
rect 10194 24656 13818 24712
rect 13874 24656 13879 24712
rect 10133 24654 13879 24656
rect 10133 24651 10199 24654
rect 13813 24651 13879 24654
rect 35574 24581 35634 24790
rect 39520 24760 40000 24790
rect 15469 24578 15535 24581
rect 18597 24578 18663 24581
rect 15469 24576 18663 24578
rect 15469 24520 15474 24576
rect 15530 24520 18602 24576
rect 18658 24520 18663 24576
rect 15469 24518 18663 24520
rect 15469 24515 15535 24518
rect 18597 24515 18663 24518
rect 35525 24576 35634 24581
rect 35525 24520 35530 24576
rect 35586 24520 35634 24576
rect 35525 24518 35634 24520
rect 35525 24515 35591 24518
rect 19568 24512 19888 24513
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 24447 19888 24448
rect 14457 24306 14523 24309
rect 20069 24306 20135 24309
rect 14457 24304 20135 24306
rect 14457 24248 14462 24304
rect 14518 24248 20074 24304
rect 20130 24248 20135 24304
rect 14457 24246 20135 24248
rect 14457 24243 14523 24246
rect 20069 24243 20135 24246
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 34928 23968 35248 23969
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 23903 35248 23904
rect 19057 23898 19123 23901
rect 21541 23898 21607 23901
rect 19057 23896 21607 23898
rect 19057 23840 19062 23896
rect 19118 23840 21546 23896
rect 21602 23840 21607 23896
rect 19057 23838 21607 23840
rect 19057 23835 19123 23838
rect 21541 23835 21607 23838
rect 7189 23762 7255 23765
rect 10501 23762 10567 23765
rect 7189 23760 10567 23762
rect 7189 23704 7194 23760
rect 7250 23704 10506 23760
rect 10562 23704 10567 23760
rect 7189 23702 10567 23704
rect 7189 23699 7255 23702
rect 10501 23699 10567 23702
rect 19149 23626 19215 23629
rect 21081 23626 21147 23629
rect 19149 23624 21147 23626
rect 19149 23568 19154 23624
rect 19210 23568 21086 23624
rect 21142 23568 21147 23624
rect 19149 23566 21147 23568
rect 19149 23563 19215 23566
rect 21081 23563 21147 23566
rect 34145 23626 34211 23629
rect 39520 23626 40000 23656
rect 34145 23624 40000 23626
rect 34145 23568 34150 23624
rect 34206 23568 40000 23624
rect 34145 23566 40000 23568
rect 34145 23563 34211 23566
rect 39520 23536 40000 23566
rect 35525 23490 35591 23493
rect 34470 23488 35591 23490
rect 34470 23432 35530 23488
rect 35586 23432 35591 23488
rect 34470 23430 35591 23432
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 23359 19888 23360
rect 27153 23082 27219 23085
rect 34470 23082 34530 23430
rect 35525 23427 35591 23430
rect 34697 23354 34763 23357
rect 27153 23080 34530 23082
rect 27153 23024 27158 23080
rect 27214 23024 34530 23080
rect 27153 23022 34530 23024
rect 34654 23352 34763 23354
rect 34654 23296 34702 23352
rect 34758 23296 34763 23352
rect 34654 23291 34763 23296
rect 27153 23019 27219 23022
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 34513 22402 34579 22405
rect 34654 22402 34714 23291
rect 34928 22880 35248 22881
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 22815 35248 22816
rect 34513 22400 34714 22402
rect 34513 22344 34518 22400
rect 34574 22344 34714 22400
rect 34513 22342 34714 22344
rect 35525 22402 35591 22405
rect 39520 22402 40000 22432
rect 35525 22400 40000 22402
rect 35525 22344 35530 22400
rect 35586 22344 40000 22400
rect 35525 22342 40000 22344
rect 34513 22339 34579 22342
rect 35525 22339 35591 22342
rect 19568 22336 19888 22337
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 39520 22312 40000 22342
rect 19568 22271 19888 22272
rect 16849 22266 16915 22269
rect 19333 22266 19399 22269
rect 34697 22268 34763 22269
rect 16849 22264 19399 22266
rect 16849 22208 16854 22264
rect 16910 22208 19338 22264
rect 19394 22208 19399 22264
rect 16849 22206 19399 22208
rect 16849 22203 16915 22206
rect 19333 22203 19399 22206
rect 34646 22204 34652 22268
rect 34716 22266 34763 22268
rect 34716 22264 34808 22266
rect 34758 22208 34808 22264
rect 34716 22206 34808 22208
rect 34716 22204 34763 22206
rect 34697 22203 34763 22204
rect 21541 22130 21607 22133
rect 25497 22130 25563 22133
rect 21541 22128 25563 22130
rect 21541 22072 21546 22128
rect 21602 22072 25502 22128
rect 25558 22072 25563 22128
rect 21541 22070 25563 22072
rect 21541 22067 21607 22070
rect 25497 22067 25563 22070
rect 13629 21994 13695 21997
rect 15745 21994 15811 21997
rect 13629 21992 15811 21994
rect 13629 21936 13634 21992
rect 13690 21936 15750 21992
rect 15806 21936 15811 21992
rect 13629 21934 15811 21936
rect 13629 21931 13695 21934
rect 15745 21931 15811 21934
rect 27889 21994 27955 21997
rect 34145 21994 34211 21997
rect 27889 21992 34211 21994
rect 27889 21936 27894 21992
rect 27950 21936 34150 21992
rect 34206 21936 34211 21992
rect 27889 21934 34211 21936
rect 27889 21931 27955 21934
rect 34145 21931 34211 21934
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 34928 21792 35248 21793
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 21727 35248 21728
rect 19568 21248 19888 21249
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 21183 19888 21184
rect 35617 21178 35683 21181
rect 39520 21178 40000 21208
rect 35617 21176 40000 21178
rect 35617 21120 35622 21176
rect 35678 21120 40000 21176
rect 35617 21118 40000 21120
rect 35617 21115 35683 21118
rect 39520 21088 40000 21118
rect 15285 21042 15351 21045
rect 19149 21042 19215 21045
rect 15285 21040 19215 21042
rect 15285 20984 15290 21040
rect 15346 20984 19154 21040
rect 19210 20984 19215 21040
rect 15285 20982 19215 20984
rect 15285 20979 15351 20982
rect 19149 20979 19215 20982
rect 21725 21042 21791 21045
rect 23657 21042 23723 21045
rect 21725 21040 23723 21042
rect 21725 20984 21730 21040
rect 21786 20984 23662 21040
rect 23718 20984 23723 21040
rect 21725 20982 23723 20984
rect 21725 20979 21791 20982
rect 23657 20979 23723 20982
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 34928 20704 35248 20705
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 20639 35248 20640
rect 10041 20634 10107 20637
rect 13261 20634 13327 20637
rect 10041 20632 13327 20634
rect 10041 20576 10046 20632
rect 10102 20576 13266 20632
rect 13322 20576 13327 20632
rect 10041 20574 13327 20576
rect 10041 20571 10107 20574
rect 13261 20571 13327 20574
rect 23013 20634 23079 20637
rect 25129 20634 25195 20637
rect 23013 20632 25195 20634
rect 23013 20576 23018 20632
rect 23074 20576 25134 20632
rect 25190 20576 25195 20632
rect 23013 20574 25195 20576
rect 23013 20571 23079 20574
rect 25129 20571 25195 20574
rect 26141 20498 26207 20501
rect 35525 20498 35591 20501
rect 26141 20496 35591 20498
rect 26141 20440 26146 20496
rect 26202 20440 35530 20496
rect 35586 20440 35591 20496
rect 26141 20438 35591 20440
rect 26141 20435 26207 20438
rect 35525 20435 35591 20438
rect 25405 20362 25471 20365
rect 28073 20362 28139 20365
rect 25405 20360 28139 20362
rect 25405 20304 25410 20360
rect 25466 20304 28078 20360
rect 28134 20304 28139 20360
rect 25405 20302 28139 20304
rect 25405 20299 25471 20302
rect 28073 20299 28139 20302
rect 33777 20362 33843 20365
rect 35341 20362 35407 20365
rect 33777 20360 35407 20362
rect 33777 20304 33782 20360
rect 33838 20304 35346 20360
rect 35402 20304 35407 20360
rect 33777 20302 35407 20304
rect 33777 20299 33843 20302
rect 35341 20299 35407 20302
rect 19568 20160 19888 20161
rect 0 20090 480 20120
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 20095 19888 20096
rect 1577 20090 1643 20093
rect 0 20088 1643 20090
rect 0 20032 1582 20088
rect 1638 20032 1643 20088
rect 0 20030 1643 20032
rect 0 20000 480 20030
rect 1577 20027 1643 20030
rect 26601 20090 26667 20093
rect 35617 20090 35683 20093
rect 26601 20088 35683 20090
rect 26601 20032 26606 20088
rect 26662 20032 35622 20088
rect 35678 20032 35683 20088
rect 26601 20030 35683 20032
rect 26601 20027 26667 20030
rect 35617 20027 35683 20030
rect 34145 19954 34211 19957
rect 39520 19954 40000 19984
rect 34145 19952 40000 19954
rect 34145 19896 34150 19952
rect 34206 19896 40000 19952
rect 34145 19894 40000 19896
rect 34145 19891 34211 19894
rect 39520 19864 40000 19894
rect 35341 19818 35407 19821
rect 37089 19818 37155 19821
rect 35341 19816 37155 19818
rect 35341 19760 35346 19816
rect 35402 19760 37094 19816
rect 37150 19760 37155 19816
rect 35341 19758 37155 19760
rect 35341 19755 35407 19758
rect 37089 19755 37155 19758
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 34928 19616 35248 19617
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 19551 35248 19552
rect 23841 19274 23907 19277
rect 26877 19274 26943 19277
rect 23841 19272 26943 19274
rect 23841 19216 23846 19272
rect 23902 19216 26882 19272
rect 26938 19216 26943 19272
rect 23841 19214 26943 19216
rect 23841 19211 23907 19214
rect 26877 19211 26943 19214
rect 32305 19274 32371 19277
rect 33961 19274 34027 19277
rect 32305 19272 34027 19274
rect 32305 19216 32310 19272
rect 32366 19216 33966 19272
rect 34022 19216 34027 19272
rect 32305 19214 34027 19216
rect 32305 19211 32371 19214
rect 33961 19211 34027 19214
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 19007 19888 19008
rect 24117 18866 24183 18869
rect 24577 18866 24643 18869
rect 25313 18866 25379 18869
rect 27797 18866 27863 18869
rect 24117 18864 27863 18866
rect 24117 18808 24122 18864
rect 24178 18808 24582 18864
rect 24638 18808 25318 18864
rect 25374 18808 27802 18864
rect 27858 18808 27863 18864
rect 24117 18806 27863 18808
rect 24117 18803 24183 18806
rect 24577 18803 24643 18806
rect 25313 18803 25379 18806
rect 27797 18803 27863 18806
rect 30373 18866 30439 18869
rect 33869 18866 33935 18869
rect 30373 18864 33935 18866
rect 30373 18808 30378 18864
rect 30434 18808 33874 18864
rect 33930 18808 33935 18864
rect 30373 18806 33935 18808
rect 30373 18803 30439 18806
rect 33869 18803 33935 18806
rect 24393 18730 24459 18733
rect 26877 18730 26943 18733
rect 24393 18728 26943 18730
rect 24393 18672 24398 18728
rect 24454 18672 26882 18728
rect 26938 18672 26943 18728
rect 24393 18670 26943 18672
rect 24393 18667 24459 18670
rect 26877 18667 26943 18670
rect 34605 18730 34671 18733
rect 39520 18730 40000 18760
rect 34605 18728 40000 18730
rect 34605 18672 34610 18728
rect 34666 18672 40000 18728
rect 34605 18670 40000 18672
rect 34605 18667 34671 18670
rect 39520 18640 40000 18670
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 34928 18528 35248 18529
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 18463 35248 18464
rect 28441 18458 28507 18461
rect 31293 18458 31359 18461
rect 28441 18456 31359 18458
rect 28441 18400 28446 18456
rect 28502 18400 31298 18456
rect 31354 18400 31359 18456
rect 28441 18398 31359 18400
rect 28441 18395 28507 18398
rect 31293 18395 31359 18398
rect 32305 18050 32371 18053
rect 34421 18050 34487 18053
rect 32305 18048 34487 18050
rect 32305 17992 32310 18048
rect 32366 17992 34426 18048
rect 34482 17992 34487 18048
rect 32305 17990 34487 17992
rect 32305 17987 32371 17990
rect 34421 17987 34487 17990
rect 19568 17984 19888 17985
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 24761 17914 24827 17917
rect 26509 17914 26575 17917
rect 24761 17912 26575 17914
rect 24761 17856 24766 17912
rect 24822 17856 26514 17912
rect 26570 17856 26575 17912
rect 24761 17854 26575 17856
rect 24761 17851 24827 17854
rect 26509 17851 26575 17854
rect 18965 17642 19031 17645
rect 22185 17642 22251 17645
rect 18965 17640 22251 17642
rect 18965 17584 18970 17640
rect 19026 17584 22190 17640
rect 22246 17584 22251 17640
rect 18965 17582 22251 17584
rect 18965 17579 19031 17582
rect 22185 17579 22251 17582
rect 27429 17506 27495 17509
rect 27705 17506 27771 17509
rect 29177 17506 29243 17509
rect 27429 17504 29243 17506
rect 27429 17448 27434 17504
rect 27490 17448 27710 17504
rect 27766 17448 29182 17504
rect 29238 17448 29243 17504
rect 27429 17446 29243 17448
rect 27429 17443 27495 17446
rect 27705 17443 27771 17446
rect 29177 17443 29243 17446
rect 35617 17506 35683 17509
rect 39520 17506 40000 17536
rect 35617 17504 40000 17506
rect 35617 17448 35622 17504
rect 35678 17448 40000 17504
rect 35617 17446 40000 17448
rect 35617 17443 35683 17446
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 34928 17440 35248 17441
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 39520 17416 40000 17446
rect 34928 17375 35248 17376
rect 20253 17370 20319 17373
rect 27613 17370 27679 17373
rect 20253 17368 27679 17370
rect 20253 17312 20258 17368
rect 20314 17312 27618 17368
rect 27674 17312 27679 17368
rect 20253 17310 27679 17312
rect 20253 17307 20319 17310
rect 27613 17307 27679 17310
rect 21817 17234 21883 17237
rect 23657 17234 23723 17237
rect 21817 17232 23723 17234
rect 21817 17176 21822 17232
rect 21878 17176 23662 17232
rect 23718 17176 23723 17232
rect 21817 17174 23723 17176
rect 21817 17171 21883 17174
rect 23657 17171 23723 17174
rect 19241 17098 19307 17101
rect 22461 17098 22527 17101
rect 19241 17096 22527 17098
rect 19241 17040 19246 17096
rect 19302 17040 22466 17096
rect 22522 17040 22527 17096
rect 19241 17038 22527 17040
rect 19241 17035 19307 17038
rect 22461 17035 22527 17038
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 16831 19888 16832
rect 29913 16690 29979 16693
rect 35382 16690 35388 16692
rect 29913 16688 35388 16690
rect 29913 16632 29918 16688
rect 29974 16632 35388 16688
rect 29913 16630 35388 16632
rect 29913 16627 29979 16630
rect 35382 16628 35388 16630
rect 35452 16628 35458 16692
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 34928 16352 35248 16353
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 16287 35248 16288
rect 29913 16282 29979 16285
rect 34605 16282 34671 16285
rect 29913 16280 34671 16282
rect 29913 16224 29918 16280
rect 29974 16224 34610 16280
rect 34666 16224 34671 16280
rect 29913 16222 34671 16224
rect 29913 16219 29979 16222
rect 34605 16219 34671 16222
rect 35433 16282 35499 16285
rect 39520 16282 40000 16312
rect 35433 16280 40000 16282
rect 35433 16224 35438 16280
rect 35494 16224 40000 16280
rect 35433 16222 40000 16224
rect 35433 16219 35499 16222
rect 39520 16192 40000 16222
rect 28625 16146 28691 16149
rect 35617 16146 35683 16149
rect 28625 16144 35683 16146
rect 28625 16088 28630 16144
rect 28686 16088 35622 16144
rect 35678 16088 35683 16144
rect 28625 16086 35683 16088
rect 28625 16083 28691 16086
rect 35617 16083 35683 16086
rect 25773 15874 25839 15877
rect 31753 15874 31819 15877
rect 25773 15872 31819 15874
rect 25773 15816 25778 15872
rect 25834 15816 31758 15872
rect 31814 15816 31819 15872
rect 25773 15814 31819 15816
rect 25773 15811 25839 15814
rect 31753 15811 31819 15814
rect 19568 15808 19888 15809
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 15743 19888 15744
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 34928 15264 35248 15265
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 15199 35248 15200
rect 21357 15194 21423 15197
rect 26233 15194 26299 15197
rect 21357 15192 26299 15194
rect 21357 15136 21362 15192
rect 21418 15136 26238 15192
rect 26294 15136 26299 15192
rect 21357 15134 26299 15136
rect 21357 15131 21423 15134
rect 26233 15131 26299 15134
rect 30557 15058 30623 15061
rect 34145 15058 34211 15061
rect 30557 15056 34211 15058
rect 30557 15000 30562 15056
rect 30618 15000 34150 15056
rect 34206 15000 34211 15056
rect 30557 14998 34211 15000
rect 30557 14995 30623 14998
rect 34145 14995 34211 14998
rect 35617 15058 35683 15061
rect 39520 15058 40000 15088
rect 35617 15056 40000 15058
rect 35617 15000 35622 15056
rect 35678 15000 40000 15056
rect 35617 14998 40000 15000
rect 35617 14995 35683 14998
rect 39520 14968 40000 14998
rect 19568 14720 19888 14721
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 14655 19888 14656
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 34928 14176 35248 14177
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 14111 35248 14112
rect 36997 13970 37063 13973
rect 39520 13970 40000 14000
rect 36997 13968 40000 13970
rect 36997 13912 37002 13968
rect 37058 13912 40000 13968
rect 36997 13910 40000 13912
rect 36997 13907 37063 13910
rect 39520 13880 40000 13910
rect 32765 13834 32831 13837
rect 33777 13834 33843 13837
rect 36813 13834 36879 13837
rect 32765 13832 36879 13834
rect 32765 13776 32770 13832
rect 32826 13776 33782 13832
rect 33838 13776 36818 13832
rect 36874 13776 36879 13832
rect 32765 13774 36879 13776
rect 32765 13771 32831 13774
rect 33777 13771 33843 13774
rect 36813 13771 36879 13774
rect 19568 13632 19888 13633
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 13567 19888 13568
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 34928 13088 35248 13089
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 13023 35248 13024
rect 36537 12746 36603 12749
rect 39520 12746 40000 12776
rect 36537 12744 40000 12746
rect 36537 12688 36542 12744
rect 36598 12688 40000 12744
rect 36537 12686 40000 12688
rect 36537 12683 36603 12686
rect 39520 12656 40000 12686
rect 33961 12610 34027 12613
rect 34329 12610 34395 12613
rect 33961 12608 34395 12610
rect 33961 12552 33966 12608
rect 34022 12552 34334 12608
rect 34390 12552 34395 12608
rect 33961 12550 34395 12552
rect 33961 12547 34027 12550
rect 34329 12547 34395 12550
rect 19568 12544 19888 12545
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect 35341 12476 35407 12477
rect 35341 12474 35388 12476
rect 35296 12472 35388 12474
rect 35296 12416 35346 12472
rect 35296 12414 35388 12416
rect 35341 12412 35388 12414
rect 35452 12412 35458 12476
rect 35341 12411 35407 12412
rect 27429 12338 27495 12341
rect 30557 12338 30623 12341
rect 27429 12336 30623 12338
rect 27429 12280 27434 12336
rect 27490 12280 30562 12336
rect 30618 12280 30623 12336
rect 27429 12278 30623 12280
rect 27429 12275 27495 12278
rect 30557 12275 30623 12278
rect 28073 12202 28139 12205
rect 34053 12202 34119 12205
rect 28073 12200 34119 12202
rect 28073 12144 28078 12200
rect 28134 12144 34058 12200
rect 34114 12144 34119 12200
rect 28073 12142 34119 12144
rect 28073 12139 28139 12142
rect 34053 12139 34119 12142
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 34928 12000 35248 12001
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 11935 35248 11936
rect 32765 11794 32831 11797
rect 35341 11794 35407 11797
rect 32765 11792 35407 11794
rect 32765 11736 32770 11792
rect 32826 11736 35346 11792
rect 35402 11736 35407 11792
rect 32765 11734 35407 11736
rect 32765 11731 32831 11734
rect 35341 11731 35407 11734
rect 37089 11522 37155 11525
rect 39520 11522 40000 11552
rect 37089 11520 40000 11522
rect 37089 11464 37094 11520
rect 37150 11464 40000 11520
rect 37089 11462 40000 11464
rect 37089 11459 37155 11462
rect 19568 11456 19888 11457
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 39520 11432 40000 11462
rect 19568 11391 19888 11392
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 34928 10912 35248 10913
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 10847 35248 10848
rect 19568 10368 19888 10369
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 10303 19888 10304
rect 30281 10298 30347 10301
rect 32489 10298 32555 10301
rect 30281 10296 32555 10298
rect 30281 10240 30286 10296
rect 30342 10240 32494 10296
rect 32550 10240 32555 10296
rect 30281 10238 32555 10240
rect 30281 10235 30347 10238
rect 32489 10235 32555 10238
rect 36905 10298 36971 10301
rect 39520 10298 40000 10328
rect 36905 10296 40000 10298
rect 36905 10240 36910 10296
rect 36966 10240 40000 10296
rect 36905 10238 40000 10240
rect 36905 10235 36971 10238
rect 39520 10208 40000 10238
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 34928 9824 35248 9825
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 9759 35248 9760
rect 29821 9754 29887 9757
rect 31937 9754 32003 9757
rect 29821 9752 32003 9754
rect 29821 9696 29826 9752
rect 29882 9696 31942 9752
rect 31998 9696 32003 9752
rect 29821 9694 32003 9696
rect 29821 9691 29887 9694
rect 31937 9691 32003 9694
rect 19568 9280 19888 9281
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect 29821 9210 29887 9213
rect 36813 9210 36879 9213
rect 29821 9208 36879 9210
rect 29821 9152 29826 9208
rect 29882 9152 36818 9208
rect 36874 9152 36879 9208
rect 29821 9150 36879 9152
rect 29821 9147 29887 9150
rect 36813 9147 36879 9150
rect 36629 9074 36695 9077
rect 39520 9074 40000 9104
rect 36629 9072 40000 9074
rect 36629 9016 36634 9072
rect 36690 9016 40000 9072
rect 36629 9014 40000 9016
rect 36629 9011 36695 9014
rect 39520 8984 40000 9014
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 34928 8736 35248 8737
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 8671 35248 8672
rect 19568 8192 19888 8193
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 8127 19888 8128
rect 35709 7850 35775 7853
rect 39520 7850 40000 7880
rect 35709 7848 40000 7850
rect 35709 7792 35714 7848
rect 35770 7792 40000 7848
rect 35709 7790 40000 7792
rect 35709 7787 35775 7790
rect 39520 7760 40000 7790
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 34928 7648 35248 7649
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 7583 35248 7584
rect 16665 7578 16731 7581
rect 29637 7578 29703 7581
rect 32949 7578 33015 7581
rect 16665 7576 33015 7578
rect 16665 7520 16670 7576
rect 16726 7520 29642 7576
rect 29698 7520 32954 7576
rect 33010 7520 33015 7576
rect 16665 7518 33015 7520
rect 16665 7515 16731 7518
rect 29637 7515 29703 7518
rect 32949 7515 33015 7518
rect 32857 7442 32923 7445
rect 34605 7442 34671 7445
rect 32857 7440 34671 7442
rect 32857 7384 32862 7440
rect 32918 7384 34610 7440
rect 34666 7384 34671 7440
rect 32857 7382 34671 7384
rect 32857 7379 32923 7382
rect 34605 7379 34671 7382
rect 19568 7104 19888 7105
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 7039 19888 7040
rect 0 6762 480 6792
rect 565 6762 631 6765
rect 0 6760 631 6762
rect 0 6704 570 6760
rect 626 6704 631 6760
rect 0 6702 631 6704
rect 0 6672 480 6702
rect 565 6699 631 6702
rect 34697 6762 34763 6765
rect 34697 6760 35404 6762
rect 34697 6704 34702 6760
rect 34758 6704 35404 6760
rect 34697 6702 35404 6704
rect 34697 6699 34763 6702
rect 35344 6626 35404 6702
rect 39520 6626 40000 6656
rect 35344 6566 40000 6626
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 34928 6560 35248 6561
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 39520 6536 40000 6566
rect 34928 6495 35248 6496
rect 33777 6354 33843 6357
rect 37273 6354 37339 6357
rect 33777 6352 37339 6354
rect 33777 6296 33782 6352
rect 33838 6296 37278 6352
rect 37334 6296 37339 6352
rect 33777 6294 37339 6296
rect 33777 6291 33843 6294
rect 37273 6291 37339 6294
rect 32397 6082 32463 6085
rect 35433 6082 35499 6085
rect 32397 6080 35499 6082
rect 32397 6024 32402 6080
rect 32458 6024 35438 6080
rect 35494 6024 35499 6080
rect 32397 6022 35499 6024
rect 32397 6019 32463 6022
rect 35433 6019 35499 6022
rect 19568 6016 19888 6017
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 5951 19888 5952
rect 565 5674 631 5677
rect 18413 5674 18479 5677
rect 565 5672 18479 5674
rect 565 5616 570 5672
rect 626 5616 18418 5672
rect 18474 5616 18479 5672
rect 565 5614 18479 5616
rect 565 5611 631 5614
rect 18413 5611 18479 5614
rect 34237 5674 34303 5677
rect 36629 5674 36695 5677
rect 34237 5672 36695 5674
rect 34237 5616 34242 5672
rect 34298 5616 36634 5672
rect 36690 5616 36695 5672
rect 34237 5614 36695 5616
rect 34237 5611 34303 5614
rect 36629 5611 36695 5614
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 34928 5472 35248 5473
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 5407 35248 5408
rect 39520 5402 40000 5432
rect 35344 5342 40000 5402
rect 34697 5266 34763 5269
rect 35344 5266 35404 5342
rect 39520 5312 40000 5342
rect 34697 5264 35404 5266
rect 34697 5208 34702 5264
rect 34758 5208 35404 5264
rect 34697 5206 35404 5208
rect 34697 5203 34763 5206
rect 27337 4994 27403 4997
rect 32213 4994 32279 4997
rect 27337 4992 32279 4994
rect 27337 4936 27342 4992
rect 27398 4936 32218 4992
rect 32274 4936 32279 4992
rect 27337 4934 32279 4936
rect 27337 4931 27403 4934
rect 32213 4931 32279 4934
rect 19568 4928 19888 4929
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 4863 19888 4864
rect 27613 4858 27679 4861
rect 32765 4858 32831 4861
rect 27613 4856 32831 4858
rect 27613 4800 27618 4856
rect 27674 4800 32770 4856
rect 32826 4800 32831 4856
rect 27613 4798 32831 4800
rect 27613 4795 27679 4798
rect 32765 4795 32831 4798
rect 29821 4722 29887 4725
rect 32121 4722 32187 4725
rect 29821 4720 32187 4722
rect 29821 4664 29826 4720
rect 29882 4664 32126 4720
rect 32182 4664 32187 4720
rect 29821 4662 32187 4664
rect 29821 4659 29887 4662
rect 32121 4659 32187 4662
rect 34237 4722 34303 4725
rect 35893 4722 35959 4725
rect 34237 4720 35959 4722
rect 34237 4664 34242 4720
rect 34298 4664 35898 4720
rect 35954 4664 35959 4720
rect 34237 4662 35959 4664
rect 34237 4659 34303 4662
rect 35893 4659 35959 4662
rect 28717 4586 28783 4589
rect 31017 4586 31083 4589
rect 34973 4586 35039 4589
rect 35525 4586 35591 4589
rect 36445 4586 36511 4589
rect 28717 4584 36511 4586
rect 28717 4528 28722 4584
rect 28778 4528 31022 4584
rect 31078 4528 34978 4584
rect 35034 4528 35530 4584
rect 35586 4528 36450 4584
rect 36506 4528 36511 4584
rect 28717 4526 36511 4528
rect 28717 4523 28783 4526
rect 31017 4523 31083 4526
rect 34973 4523 35039 4526
rect 35525 4523 35591 4526
rect 36445 4523 36511 4526
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 34928 4384 35248 4385
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 4319 35248 4320
rect 35801 4178 35867 4181
rect 39520 4178 40000 4208
rect 35801 4176 40000 4178
rect 35801 4120 35806 4176
rect 35862 4120 40000 4176
rect 35801 4118 40000 4120
rect 35801 4115 35867 4118
rect 39520 4088 40000 4118
rect 23289 4042 23355 4045
rect 24209 4042 24275 4045
rect 23289 4040 24275 4042
rect 23289 3984 23294 4040
rect 23350 3984 24214 4040
rect 24270 3984 24275 4040
rect 23289 3982 24275 3984
rect 23289 3979 23355 3982
rect 24209 3979 24275 3982
rect 34145 3906 34211 3909
rect 35893 3906 35959 3909
rect 34145 3904 35959 3906
rect 34145 3848 34150 3904
rect 34206 3848 35898 3904
rect 35954 3848 35959 3904
rect 34145 3846 35959 3848
rect 34145 3843 34211 3846
rect 35893 3843 35959 3846
rect 19568 3840 19888 3841
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 3325 3498 3391 3501
rect 32489 3498 32555 3501
rect 3325 3496 32555 3498
rect 3325 3440 3330 3496
rect 3386 3440 32494 3496
rect 32550 3440 32555 3496
rect 3325 3438 32555 3440
rect 3325 3435 3391 3438
rect 32489 3435 32555 3438
rect 33041 3498 33107 3501
rect 36629 3498 36695 3501
rect 33041 3496 36695 3498
rect 33041 3440 33046 3496
rect 33102 3440 36634 3496
rect 36690 3440 36695 3496
rect 33041 3438 36695 3440
rect 33041 3435 33107 3438
rect 36629 3435 36695 3438
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 34928 3296 35248 3297
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 3231 35248 3232
rect 27797 3226 27863 3229
rect 31569 3226 31635 3229
rect 27797 3224 31635 3226
rect 27797 3168 27802 3224
rect 27858 3168 31574 3224
rect 31630 3168 31635 3224
rect 27797 3166 31635 3168
rect 27797 3163 27863 3166
rect 31569 3163 31635 3166
rect 28073 3090 28139 3093
rect 33685 3090 33751 3093
rect 28073 3088 33751 3090
rect 28073 3032 28078 3088
rect 28134 3032 33690 3088
rect 33746 3032 33751 3088
rect 28073 3030 33751 3032
rect 28073 3027 28139 3030
rect 33685 3027 33751 3030
rect 27705 2954 27771 2957
rect 31937 2954 32003 2957
rect 27705 2952 32003 2954
rect 27705 2896 27710 2952
rect 27766 2896 31942 2952
rect 31998 2896 32003 2952
rect 27705 2894 32003 2896
rect 27705 2891 27771 2894
rect 31937 2891 32003 2894
rect 35709 2954 35775 2957
rect 39520 2954 40000 2984
rect 35709 2952 40000 2954
rect 35709 2896 35714 2952
rect 35770 2896 40000 2952
rect 35709 2894 40000 2896
rect 35709 2891 35775 2894
rect 39520 2864 40000 2894
rect 27981 2818 28047 2821
rect 34605 2818 34671 2821
rect 27981 2816 34671 2818
rect 27981 2760 27986 2816
rect 28042 2760 34610 2816
rect 34666 2760 34671 2816
rect 27981 2758 34671 2760
rect 27981 2755 28047 2758
rect 34605 2755 34671 2758
rect 19568 2752 19888 2753
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2687 19888 2688
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 34928 2208 35248 2209
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2143 35248 2144
rect 35341 1730 35407 1733
rect 39520 1730 40000 1760
rect 35341 1728 40000 1730
rect 35341 1672 35346 1728
rect 35402 1672 40000 1728
rect 35341 1670 40000 1672
rect 35341 1667 35407 1670
rect 39520 1640 40000 1670
rect 36353 642 36419 645
rect 39520 642 40000 672
rect 36353 640 40000 642
rect 36353 584 36358 640
rect 36414 584 40000 640
rect 36353 582 40000 584
rect 36353 579 36419 582
rect 39520 552 40000 582
<< via3 >>
rect 19576 37564 19640 37568
rect 19576 37508 19580 37564
rect 19580 37508 19636 37564
rect 19636 37508 19640 37564
rect 19576 37504 19640 37508
rect 19656 37564 19720 37568
rect 19656 37508 19660 37564
rect 19660 37508 19716 37564
rect 19716 37508 19720 37564
rect 19656 37504 19720 37508
rect 19736 37564 19800 37568
rect 19736 37508 19740 37564
rect 19740 37508 19796 37564
rect 19796 37508 19800 37564
rect 19736 37504 19800 37508
rect 19816 37564 19880 37568
rect 19816 37508 19820 37564
rect 19820 37508 19876 37564
rect 19876 37508 19880 37564
rect 19816 37504 19880 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 34936 37020 35000 37024
rect 34936 36964 34940 37020
rect 34940 36964 34996 37020
rect 34996 36964 35000 37020
rect 34936 36960 35000 36964
rect 35016 37020 35080 37024
rect 35016 36964 35020 37020
rect 35020 36964 35076 37020
rect 35076 36964 35080 37020
rect 35016 36960 35080 36964
rect 35096 37020 35160 37024
rect 35096 36964 35100 37020
rect 35100 36964 35156 37020
rect 35156 36964 35160 37020
rect 35096 36960 35160 36964
rect 35176 37020 35240 37024
rect 35176 36964 35180 37020
rect 35180 36964 35236 37020
rect 35236 36964 35240 37020
rect 35176 36960 35240 36964
rect 19576 36476 19640 36480
rect 19576 36420 19580 36476
rect 19580 36420 19636 36476
rect 19636 36420 19640 36476
rect 19576 36416 19640 36420
rect 19656 36476 19720 36480
rect 19656 36420 19660 36476
rect 19660 36420 19716 36476
rect 19716 36420 19720 36476
rect 19656 36416 19720 36420
rect 19736 36476 19800 36480
rect 19736 36420 19740 36476
rect 19740 36420 19796 36476
rect 19796 36420 19800 36476
rect 19736 36416 19800 36420
rect 19816 36476 19880 36480
rect 19816 36420 19820 36476
rect 19820 36420 19876 36476
rect 19876 36420 19880 36476
rect 19816 36416 19880 36420
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 34936 35932 35000 35936
rect 34936 35876 34940 35932
rect 34940 35876 34996 35932
rect 34996 35876 35000 35932
rect 34936 35872 35000 35876
rect 35016 35932 35080 35936
rect 35016 35876 35020 35932
rect 35020 35876 35076 35932
rect 35076 35876 35080 35932
rect 35016 35872 35080 35876
rect 35096 35932 35160 35936
rect 35096 35876 35100 35932
rect 35100 35876 35156 35932
rect 35156 35876 35160 35932
rect 35096 35872 35160 35876
rect 35176 35932 35240 35936
rect 35176 35876 35180 35932
rect 35180 35876 35236 35932
rect 35236 35876 35240 35932
rect 35176 35872 35240 35876
rect 24900 35804 24964 35868
rect 6684 35728 6748 35732
rect 6684 35672 6698 35728
rect 6698 35672 6748 35728
rect 6684 35668 6748 35672
rect 5028 35456 5092 35460
rect 5028 35400 5042 35456
rect 5042 35400 5092 35456
rect 5028 35396 5092 35400
rect 19576 35388 19640 35392
rect 19576 35332 19580 35388
rect 19580 35332 19636 35388
rect 19636 35332 19640 35388
rect 19576 35328 19640 35332
rect 19656 35388 19720 35392
rect 19656 35332 19660 35388
rect 19660 35332 19716 35388
rect 19716 35332 19720 35388
rect 19656 35328 19720 35332
rect 19736 35388 19800 35392
rect 19736 35332 19740 35388
rect 19740 35332 19796 35388
rect 19796 35332 19800 35388
rect 19736 35328 19800 35332
rect 19816 35388 19880 35392
rect 19816 35332 19820 35388
rect 19820 35332 19876 35388
rect 19876 35332 19880 35388
rect 19816 35328 19880 35332
rect 20668 35260 20732 35324
rect 21404 35260 21468 35324
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 34936 34844 35000 34848
rect 34936 34788 34940 34844
rect 34940 34788 34996 34844
rect 34996 34788 35000 34844
rect 34936 34784 35000 34788
rect 35016 34844 35080 34848
rect 35016 34788 35020 34844
rect 35020 34788 35076 34844
rect 35076 34788 35080 34844
rect 35016 34784 35080 34788
rect 35096 34844 35160 34848
rect 35096 34788 35100 34844
rect 35100 34788 35156 34844
rect 35156 34788 35160 34844
rect 35096 34784 35160 34788
rect 35176 34844 35240 34848
rect 35176 34788 35180 34844
rect 35180 34788 35236 34844
rect 35236 34788 35240 34844
rect 35176 34784 35240 34788
rect 24900 34716 24964 34780
rect 19576 34300 19640 34304
rect 19576 34244 19580 34300
rect 19580 34244 19636 34300
rect 19636 34244 19640 34300
rect 19576 34240 19640 34244
rect 19656 34300 19720 34304
rect 19656 34244 19660 34300
rect 19660 34244 19716 34300
rect 19716 34244 19720 34300
rect 19656 34240 19720 34244
rect 19736 34300 19800 34304
rect 19736 34244 19740 34300
rect 19740 34244 19796 34300
rect 19796 34244 19800 34300
rect 19736 34240 19800 34244
rect 19816 34300 19880 34304
rect 19816 34244 19820 34300
rect 19820 34244 19876 34300
rect 19876 34244 19880 34300
rect 19816 34240 19880 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 34936 33756 35000 33760
rect 34936 33700 34940 33756
rect 34940 33700 34996 33756
rect 34996 33700 35000 33756
rect 34936 33696 35000 33700
rect 35016 33756 35080 33760
rect 35016 33700 35020 33756
rect 35020 33700 35076 33756
rect 35076 33700 35080 33756
rect 35016 33696 35080 33700
rect 35096 33756 35160 33760
rect 35096 33700 35100 33756
rect 35100 33700 35156 33756
rect 35156 33700 35160 33756
rect 35096 33696 35160 33700
rect 35176 33756 35240 33760
rect 35176 33700 35180 33756
rect 35180 33700 35236 33756
rect 35236 33700 35240 33756
rect 35176 33696 35240 33700
rect 19576 33212 19640 33216
rect 19576 33156 19580 33212
rect 19580 33156 19636 33212
rect 19636 33156 19640 33212
rect 19576 33152 19640 33156
rect 19656 33212 19720 33216
rect 19656 33156 19660 33212
rect 19660 33156 19716 33212
rect 19716 33156 19720 33212
rect 19656 33152 19720 33156
rect 19736 33212 19800 33216
rect 19736 33156 19740 33212
rect 19740 33156 19796 33212
rect 19796 33156 19800 33212
rect 19736 33152 19800 33156
rect 19816 33212 19880 33216
rect 19816 33156 19820 33212
rect 19820 33156 19876 33212
rect 19876 33156 19880 33212
rect 19816 33152 19880 33156
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 34936 32668 35000 32672
rect 34936 32612 34940 32668
rect 34940 32612 34996 32668
rect 34996 32612 35000 32668
rect 34936 32608 35000 32612
rect 35016 32668 35080 32672
rect 35016 32612 35020 32668
rect 35020 32612 35076 32668
rect 35076 32612 35080 32668
rect 35016 32608 35080 32612
rect 35096 32668 35160 32672
rect 35096 32612 35100 32668
rect 35100 32612 35156 32668
rect 35156 32612 35160 32668
rect 35096 32608 35160 32612
rect 35176 32668 35240 32672
rect 35176 32612 35180 32668
rect 35180 32612 35236 32668
rect 35236 32612 35240 32668
rect 35176 32608 35240 32612
rect 19576 32124 19640 32128
rect 19576 32068 19580 32124
rect 19580 32068 19636 32124
rect 19636 32068 19640 32124
rect 19576 32064 19640 32068
rect 19656 32124 19720 32128
rect 19656 32068 19660 32124
rect 19660 32068 19716 32124
rect 19716 32068 19720 32124
rect 19656 32064 19720 32068
rect 19736 32124 19800 32128
rect 19736 32068 19740 32124
rect 19740 32068 19796 32124
rect 19796 32068 19800 32124
rect 19736 32064 19800 32068
rect 19816 32124 19880 32128
rect 19816 32068 19820 32124
rect 19820 32068 19876 32124
rect 19876 32068 19880 32124
rect 19816 32064 19880 32068
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 34936 31580 35000 31584
rect 34936 31524 34940 31580
rect 34940 31524 34996 31580
rect 34996 31524 35000 31580
rect 34936 31520 35000 31524
rect 35016 31580 35080 31584
rect 35016 31524 35020 31580
rect 35020 31524 35076 31580
rect 35076 31524 35080 31580
rect 35016 31520 35080 31524
rect 35096 31580 35160 31584
rect 35096 31524 35100 31580
rect 35100 31524 35156 31580
rect 35156 31524 35160 31580
rect 35096 31520 35160 31524
rect 35176 31580 35240 31584
rect 35176 31524 35180 31580
rect 35180 31524 35236 31580
rect 35236 31524 35240 31580
rect 35176 31520 35240 31524
rect 19576 31036 19640 31040
rect 19576 30980 19580 31036
rect 19580 30980 19636 31036
rect 19636 30980 19640 31036
rect 19576 30976 19640 30980
rect 19656 31036 19720 31040
rect 19656 30980 19660 31036
rect 19660 30980 19716 31036
rect 19716 30980 19720 31036
rect 19656 30976 19720 30980
rect 19736 31036 19800 31040
rect 19736 30980 19740 31036
rect 19740 30980 19796 31036
rect 19796 30980 19800 31036
rect 19736 30976 19800 30980
rect 19816 31036 19880 31040
rect 19816 30980 19820 31036
rect 19820 30980 19876 31036
rect 19876 30980 19880 31036
rect 19816 30976 19880 30980
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 34936 30492 35000 30496
rect 34936 30436 34940 30492
rect 34940 30436 34996 30492
rect 34996 30436 35000 30492
rect 34936 30432 35000 30436
rect 35016 30492 35080 30496
rect 35016 30436 35020 30492
rect 35020 30436 35076 30492
rect 35076 30436 35080 30492
rect 35016 30432 35080 30436
rect 35096 30492 35160 30496
rect 35096 30436 35100 30492
rect 35100 30436 35156 30492
rect 35156 30436 35160 30492
rect 35096 30432 35160 30436
rect 35176 30492 35240 30496
rect 35176 30436 35180 30492
rect 35180 30436 35236 30492
rect 35236 30436 35240 30492
rect 35176 30432 35240 30436
rect 19576 29948 19640 29952
rect 19576 29892 19580 29948
rect 19580 29892 19636 29948
rect 19636 29892 19640 29948
rect 19576 29888 19640 29892
rect 19656 29948 19720 29952
rect 19656 29892 19660 29948
rect 19660 29892 19716 29948
rect 19716 29892 19720 29948
rect 19656 29888 19720 29892
rect 19736 29948 19800 29952
rect 19736 29892 19740 29948
rect 19740 29892 19796 29948
rect 19796 29892 19800 29948
rect 19736 29888 19800 29892
rect 19816 29948 19880 29952
rect 19816 29892 19820 29948
rect 19820 29892 19876 29948
rect 19876 29892 19880 29948
rect 19816 29888 19880 29892
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 34936 29404 35000 29408
rect 34936 29348 34940 29404
rect 34940 29348 34996 29404
rect 34996 29348 35000 29404
rect 34936 29344 35000 29348
rect 35016 29404 35080 29408
rect 35016 29348 35020 29404
rect 35020 29348 35076 29404
rect 35076 29348 35080 29404
rect 35016 29344 35080 29348
rect 35096 29404 35160 29408
rect 35096 29348 35100 29404
rect 35100 29348 35156 29404
rect 35156 29348 35160 29404
rect 35096 29344 35160 29348
rect 35176 29404 35240 29408
rect 35176 29348 35180 29404
rect 35180 29348 35236 29404
rect 35236 29348 35240 29404
rect 35176 29344 35240 29348
rect 19576 28860 19640 28864
rect 19576 28804 19580 28860
rect 19580 28804 19636 28860
rect 19636 28804 19640 28860
rect 19576 28800 19640 28804
rect 19656 28860 19720 28864
rect 19656 28804 19660 28860
rect 19660 28804 19716 28860
rect 19716 28804 19720 28860
rect 19656 28800 19720 28804
rect 19736 28860 19800 28864
rect 19736 28804 19740 28860
rect 19740 28804 19796 28860
rect 19796 28804 19800 28860
rect 19736 28800 19800 28804
rect 19816 28860 19880 28864
rect 19816 28804 19820 28860
rect 19820 28804 19876 28860
rect 19876 28804 19880 28860
rect 19816 28800 19880 28804
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 34936 28316 35000 28320
rect 34936 28260 34940 28316
rect 34940 28260 34996 28316
rect 34996 28260 35000 28316
rect 34936 28256 35000 28260
rect 35016 28316 35080 28320
rect 35016 28260 35020 28316
rect 35020 28260 35076 28316
rect 35076 28260 35080 28316
rect 35016 28256 35080 28260
rect 35096 28316 35160 28320
rect 35096 28260 35100 28316
rect 35100 28260 35156 28316
rect 35156 28260 35160 28316
rect 35096 28256 35160 28260
rect 35176 28316 35240 28320
rect 35176 28260 35180 28316
rect 35180 28260 35236 28316
rect 35236 28260 35240 28316
rect 35176 28256 35240 28260
rect 21404 28188 21468 28252
rect 19576 27772 19640 27776
rect 19576 27716 19580 27772
rect 19580 27716 19636 27772
rect 19636 27716 19640 27772
rect 19576 27712 19640 27716
rect 19656 27772 19720 27776
rect 19656 27716 19660 27772
rect 19660 27716 19716 27772
rect 19716 27716 19720 27772
rect 19656 27712 19720 27716
rect 19736 27772 19800 27776
rect 19736 27716 19740 27772
rect 19740 27716 19796 27772
rect 19796 27716 19800 27772
rect 19736 27712 19800 27716
rect 19816 27772 19880 27776
rect 19816 27716 19820 27772
rect 19820 27716 19876 27772
rect 19876 27716 19880 27772
rect 19816 27712 19880 27716
rect 34652 27372 34716 27436
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 34936 27228 35000 27232
rect 34936 27172 34940 27228
rect 34940 27172 34996 27228
rect 34996 27172 35000 27228
rect 34936 27168 35000 27172
rect 35016 27228 35080 27232
rect 35016 27172 35020 27228
rect 35020 27172 35076 27228
rect 35076 27172 35080 27228
rect 35016 27168 35080 27172
rect 35096 27228 35160 27232
rect 35096 27172 35100 27228
rect 35100 27172 35156 27228
rect 35156 27172 35160 27228
rect 35096 27168 35160 27172
rect 35176 27228 35240 27232
rect 35176 27172 35180 27228
rect 35180 27172 35236 27228
rect 35236 27172 35240 27228
rect 35176 27168 35240 27172
rect 19576 26684 19640 26688
rect 19576 26628 19580 26684
rect 19580 26628 19636 26684
rect 19636 26628 19640 26684
rect 19576 26624 19640 26628
rect 19656 26684 19720 26688
rect 19656 26628 19660 26684
rect 19660 26628 19716 26684
rect 19716 26628 19720 26684
rect 19656 26624 19720 26628
rect 19736 26684 19800 26688
rect 19736 26628 19740 26684
rect 19740 26628 19796 26684
rect 19796 26628 19800 26684
rect 19736 26624 19800 26628
rect 19816 26684 19880 26688
rect 19816 26628 19820 26684
rect 19820 26628 19876 26684
rect 19876 26628 19880 26684
rect 19816 26624 19880 26628
rect 35388 26556 35452 26620
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 34936 26140 35000 26144
rect 34936 26084 34940 26140
rect 34940 26084 34996 26140
rect 34996 26084 35000 26140
rect 34936 26080 35000 26084
rect 35016 26140 35080 26144
rect 35016 26084 35020 26140
rect 35020 26084 35076 26140
rect 35076 26084 35080 26140
rect 35016 26080 35080 26084
rect 35096 26140 35160 26144
rect 35096 26084 35100 26140
rect 35100 26084 35156 26140
rect 35156 26084 35160 26140
rect 35096 26080 35160 26084
rect 35176 26140 35240 26144
rect 35176 26084 35180 26140
rect 35180 26084 35236 26140
rect 35236 26084 35240 26140
rect 35176 26080 35240 26084
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 34936 25052 35000 25056
rect 34936 24996 34940 25052
rect 34940 24996 34996 25052
rect 34996 24996 35000 25052
rect 34936 24992 35000 24996
rect 35016 25052 35080 25056
rect 35016 24996 35020 25052
rect 35020 24996 35076 25052
rect 35076 24996 35080 25052
rect 35016 24992 35080 24996
rect 35096 25052 35160 25056
rect 35096 24996 35100 25052
rect 35100 24996 35156 25052
rect 35156 24996 35160 25052
rect 35096 24992 35160 24996
rect 35176 25052 35240 25056
rect 35176 24996 35180 25052
rect 35180 24996 35236 25052
rect 35236 24996 35240 25052
rect 35176 24992 35240 24996
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 34936 23964 35000 23968
rect 34936 23908 34940 23964
rect 34940 23908 34996 23964
rect 34996 23908 35000 23964
rect 34936 23904 35000 23908
rect 35016 23964 35080 23968
rect 35016 23908 35020 23964
rect 35020 23908 35076 23964
rect 35076 23908 35080 23964
rect 35016 23904 35080 23908
rect 35096 23964 35160 23968
rect 35096 23908 35100 23964
rect 35100 23908 35156 23964
rect 35156 23908 35160 23964
rect 35096 23904 35160 23908
rect 35176 23964 35240 23968
rect 35176 23908 35180 23964
rect 35180 23908 35236 23964
rect 35236 23908 35240 23964
rect 35176 23904 35240 23908
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 34936 22876 35000 22880
rect 34936 22820 34940 22876
rect 34940 22820 34996 22876
rect 34996 22820 35000 22876
rect 34936 22816 35000 22820
rect 35016 22876 35080 22880
rect 35016 22820 35020 22876
rect 35020 22820 35076 22876
rect 35076 22820 35080 22876
rect 35016 22816 35080 22820
rect 35096 22876 35160 22880
rect 35096 22820 35100 22876
rect 35100 22820 35156 22876
rect 35156 22820 35160 22876
rect 35096 22816 35160 22820
rect 35176 22876 35240 22880
rect 35176 22820 35180 22876
rect 35180 22820 35236 22876
rect 35236 22820 35240 22876
rect 35176 22816 35240 22820
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 34652 22264 34716 22268
rect 34652 22208 34702 22264
rect 34702 22208 34716 22264
rect 34652 22204 34716 22208
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 34936 21788 35000 21792
rect 34936 21732 34940 21788
rect 34940 21732 34996 21788
rect 34996 21732 35000 21788
rect 34936 21728 35000 21732
rect 35016 21788 35080 21792
rect 35016 21732 35020 21788
rect 35020 21732 35076 21788
rect 35076 21732 35080 21788
rect 35016 21728 35080 21732
rect 35096 21788 35160 21792
rect 35096 21732 35100 21788
rect 35100 21732 35156 21788
rect 35156 21732 35160 21788
rect 35096 21728 35160 21732
rect 35176 21788 35240 21792
rect 35176 21732 35180 21788
rect 35180 21732 35236 21788
rect 35236 21732 35240 21788
rect 35176 21728 35240 21732
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 34936 20700 35000 20704
rect 34936 20644 34940 20700
rect 34940 20644 34996 20700
rect 34996 20644 35000 20700
rect 34936 20640 35000 20644
rect 35016 20700 35080 20704
rect 35016 20644 35020 20700
rect 35020 20644 35076 20700
rect 35076 20644 35080 20700
rect 35016 20640 35080 20644
rect 35096 20700 35160 20704
rect 35096 20644 35100 20700
rect 35100 20644 35156 20700
rect 35156 20644 35160 20700
rect 35096 20640 35160 20644
rect 35176 20700 35240 20704
rect 35176 20644 35180 20700
rect 35180 20644 35236 20700
rect 35236 20644 35240 20700
rect 35176 20640 35240 20644
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 34936 19612 35000 19616
rect 34936 19556 34940 19612
rect 34940 19556 34996 19612
rect 34996 19556 35000 19612
rect 34936 19552 35000 19556
rect 35016 19612 35080 19616
rect 35016 19556 35020 19612
rect 35020 19556 35076 19612
rect 35076 19556 35080 19612
rect 35016 19552 35080 19556
rect 35096 19612 35160 19616
rect 35096 19556 35100 19612
rect 35100 19556 35156 19612
rect 35156 19556 35160 19612
rect 35096 19552 35160 19556
rect 35176 19612 35240 19616
rect 35176 19556 35180 19612
rect 35180 19556 35236 19612
rect 35236 19556 35240 19612
rect 35176 19552 35240 19556
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 34936 18524 35000 18528
rect 34936 18468 34940 18524
rect 34940 18468 34996 18524
rect 34996 18468 35000 18524
rect 34936 18464 35000 18468
rect 35016 18524 35080 18528
rect 35016 18468 35020 18524
rect 35020 18468 35076 18524
rect 35076 18468 35080 18524
rect 35016 18464 35080 18468
rect 35096 18524 35160 18528
rect 35096 18468 35100 18524
rect 35100 18468 35156 18524
rect 35156 18468 35160 18524
rect 35096 18464 35160 18468
rect 35176 18524 35240 18528
rect 35176 18468 35180 18524
rect 35180 18468 35236 18524
rect 35236 18468 35240 18524
rect 35176 18464 35240 18468
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 34936 17436 35000 17440
rect 34936 17380 34940 17436
rect 34940 17380 34996 17436
rect 34996 17380 35000 17436
rect 34936 17376 35000 17380
rect 35016 17436 35080 17440
rect 35016 17380 35020 17436
rect 35020 17380 35076 17436
rect 35076 17380 35080 17436
rect 35016 17376 35080 17380
rect 35096 17436 35160 17440
rect 35096 17380 35100 17436
rect 35100 17380 35156 17436
rect 35156 17380 35160 17436
rect 35096 17376 35160 17380
rect 35176 17436 35240 17440
rect 35176 17380 35180 17436
rect 35180 17380 35236 17436
rect 35236 17380 35240 17436
rect 35176 17376 35240 17380
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 35388 16628 35452 16692
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 34936 16348 35000 16352
rect 34936 16292 34940 16348
rect 34940 16292 34996 16348
rect 34996 16292 35000 16348
rect 34936 16288 35000 16292
rect 35016 16348 35080 16352
rect 35016 16292 35020 16348
rect 35020 16292 35076 16348
rect 35076 16292 35080 16348
rect 35016 16288 35080 16292
rect 35096 16348 35160 16352
rect 35096 16292 35100 16348
rect 35100 16292 35156 16348
rect 35156 16292 35160 16348
rect 35096 16288 35160 16292
rect 35176 16348 35240 16352
rect 35176 16292 35180 16348
rect 35180 16292 35236 16348
rect 35236 16292 35240 16348
rect 35176 16288 35240 16292
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 34936 15260 35000 15264
rect 34936 15204 34940 15260
rect 34940 15204 34996 15260
rect 34996 15204 35000 15260
rect 34936 15200 35000 15204
rect 35016 15260 35080 15264
rect 35016 15204 35020 15260
rect 35020 15204 35076 15260
rect 35076 15204 35080 15260
rect 35016 15200 35080 15204
rect 35096 15260 35160 15264
rect 35096 15204 35100 15260
rect 35100 15204 35156 15260
rect 35156 15204 35160 15260
rect 35096 15200 35160 15204
rect 35176 15260 35240 15264
rect 35176 15204 35180 15260
rect 35180 15204 35236 15260
rect 35236 15204 35240 15260
rect 35176 15200 35240 15204
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 34936 14172 35000 14176
rect 34936 14116 34940 14172
rect 34940 14116 34996 14172
rect 34996 14116 35000 14172
rect 34936 14112 35000 14116
rect 35016 14172 35080 14176
rect 35016 14116 35020 14172
rect 35020 14116 35076 14172
rect 35076 14116 35080 14172
rect 35016 14112 35080 14116
rect 35096 14172 35160 14176
rect 35096 14116 35100 14172
rect 35100 14116 35156 14172
rect 35156 14116 35160 14172
rect 35096 14112 35160 14116
rect 35176 14172 35240 14176
rect 35176 14116 35180 14172
rect 35180 14116 35236 14172
rect 35236 14116 35240 14172
rect 35176 14112 35240 14116
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 34936 13084 35000 13088
rect 34936 13028 34940 13084
rect 34940 13028 34996 13084
rect 34996 13028 35000 13084
rect 34936 13024 35000 13028
rect 35016 13084 35080 13088
rect 35016 13028 35020 13084
rect 35020 13028 35076 13084
rect 35076 13028 35080 13084
rect 35016 13024 35080 13028
rect 35096 13084 35160 13088
rect 35096 13028 35100 13084
rect 35100 13028 35156 13084
rect 35156 13028 35160 13084
rect 35096 13024 35160 13028
rect 35176 13084 35240 13088
rect 35176 13028 35180 13084
rect 35180 13028 35236 13084
rect 35236 13028 35240 13084
rect 35176 13024 35240 13028
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 35388 12472 35452 12476
rect 35388 12416 35402 12472
rect 35402 12416 35452 12472
rect 35388 12412 35452 12416
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 34936 11996 35000 12000
rect 34936 11940 34940 11996
rect 34940 11940 34996 11996
rect 34996 11940 35000 11996
rect 34936 11936 35000 11940
rect 35016 11996 35080 12000
rect 35016 11940 35020 11996
rect 35020 11940 35076 11996
rect 35076 11940 35080 11996
rect 35016 11936 35080 11940
rect 35096 11996 35160 12000
rect 35096 11940 35100 11996
rect 35100 11940 35156 11996
rect 35156 11940 35160 11996
rect 35096 11936 35160 11940
rect 35176 11996 35240 12000
rect 35176 11940 35180 11996
rect 35180 11940 35236 11996
rect 35236 11940 35240 11996
rect 35176 11936 35240 11940
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 34936 10908 35000 10912
rect 34936 10852 34940 10908
rect 34940 10852 34996 10908
rect 34996 10852 35000 10908
rect 34936 10848 35000 10852
rect 35016 10908 35080 10912
rect 35016 10852 35020 10908
rect 35020 10852 35076 10908
rect 35076 10852 35080 10908
rect 35016 10848 35080 10852
rect 35096 10908 35160 10912
rect 35096 10852 35100 10908
rect 35100 10852 35156 10908
rect 35156 10852 35160 10908
rect 35096 10848 35160 10852
rect 35176 10908 35240 10912
rect 35176 10852 35180 10908
rect 35180 10852 35236 10908
rect 35236 10852 35240 10908
rect 35176 10848 35240 10852
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 34936 9820 35000 9824
rect 34936 9764 34940 9820
rect 34940 9764 34996 9820
rect 34996 9764 35000 9820
rect 34936 9760 35000 9764
rect 35016 9820 35080 9824
rect 35016 9764 35020 9820
rect 35020 9764 35076 9820
rect 35076 9764 35080 9820
rect 35016 9760 35080 9764
rect 35096 9820 35160 9824
rect 35096 9764 35100 9820
rect 35100 9764 35156 9820
rect 35156 9764 35160 9820
rect 35096 9760 35160 9764
rect 35176 9820 35240 9824
rect 35176 9764 35180 9820
rect 35180 9764 35236 9820
rect 35236 9764 35240 9820
rect 35176 9760 35240 9764
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 34936 8732 35000 8736
rect 34936 8676 34940 8732
rect 34940 8676 34996 8732
rect 34996 8676 35000 8732
rect 34936 8672 35000 8676
rect 35016 8732 35080 8736
rect 35016 8676 35020 8732
rect 35020 8676 35076 8732
rect 35076 8676 35080 8732
rect 35016 8672 35080 8676
rect 35096 8732 35160 8736
rect 35096 8676 35100 8732
rect 35100 8676 35156 8732
rect 35156 8676 35160 8732
rect 35096 8672 35160 8676
rect 35176 8732 35240 8736
rect 35176 8676 35180 8732
rect 35180 8676 35236 8732
rect 35236 8676 35240 8732
rect 35176 8672 35240 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 34936 7644 35000 7648
rect 34936 7588 34940 7644
rect 34940 7588 34996 7644
rect 34996 7588 35000 7644
rect 34936 7584 35000 7588
rect 35016 7644 35080 7648
rect 35016 7588 35020 7644
rect 35020 7588 35076 7644
rect 35076 7588 35080 7644
rect 35016 7584 35080 7588
rect 35096 7644 35160 7648
rect 35096 7588 35100 7644
rect 35100 7588 35156 7644
rect 35156 7588 35160 7644
rect 35096 7584 35160 7588
rect 35176 7644 35240 7648
rect 35176 7588 35180 7644
rect 35180 7588 35236 7644
rect 35236 7588 35240 7644
rect 35176 7584 35240 7588
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 34936 6556 35000 6560
rect 34936 6500 34940 6556
rect 34940 6500 34996 6556
rect 34996 6500 35000 6556
rect 34936 6496 35000 6500
rect 35016 6556 35080 6560
rect 35016 6500 35020 6556
rect 35020 6500 35076 6556
rect 35076 6500 35080 6556
rect 35016 6496 35080 6500
rect 35096 6556 35160 6560
rect 35096 6500 35100 6556
rect 35100 6500 35156 6556
rect 35156 6500 35160 6556
rect 35096 6496 35160 6500
rect 35176 6556 35240 6560
rect 35176 6500 35180 6556
rect 35180 6500 35236 6556
rect 35236 6500 35240 6556
rect 35176 6496 35240 6500
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 34936 5468 35000 5472
rect 34936 5412 34940 5468
rect 34940 5412 34996 5468
rect 34996 5412 35000 5468
rect 34936 5408 35000 5412
rect 35016 5468 35080 5472
rect 35016 5412 35020 5468
rect 35020 5412 35076 5468
rect 35076 5412 35080 5468
rect 35016 5408 35080 5412
rect 35096 5468 35160 5472
rect 35096 5412 35100 5468
rect 35100 5412 35156 5468
rect 35156 5412 35160 5468
rect 35096 5408 35160 5412
rect 35176 5468 35240 5472
rect 35176 5412 35180 5468
rect 35180 5412 35236 5468
rect 35236 5412 35240 5468
rect 35176 5408 35240 5412
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 34936 4380 35000 4384
rect 34936 4324 34940 4380
rect 34940 4324 34996 4380
rect 34996 4324 35000 4380
rect 34936 4320 35000 4324
rect 35016 4380 35080 4384
rect 35016 4324 35020 4380
rect 35020 4324 35076 4380
rect 35076 4324 35080 4380
rect 35016 4320 35080 4324
rect 35096 4380 35160 4384
rect 35096 4324 35100 4380
rect 35100 4324 35156 4380
rect 35156 4324 35160 4380
rect 35096 4320 35160 4324
rect 35176 4380 35240 4384
rect 35176 4324 35180 4380
rect 35180 4324 35236 4380
rect 35236 4324 35240 4380
rect 35176 4320 35240 4324
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 34936 3292 35000 3296
rect 34936 3236 34940 3292
rect 34940 3236 34996 3292
rect 34996 3236 35000 3292
rect 34936 3232 35000 3236
rect 35016 3292 35080 3296
rect 35016 3236 35020 3292
rect 35020 3236 35076 3292
rect 35076 3236 35080 3292
rect 35016 3232 35080 3236
rect 35096 3292 35160 3296
rect 35096 3236 35100 3292
rect 35100 3236 35156 3292
rect 35156 3236 35160 3292
rect 35096 3232 35160 3236
rect 35176 3292 35240 3296
rect 35176 3236 35180 3292
rect 35180 3236 35236 3292
rect 35236 3236 35240 3292
rect 35176 3232 35240 3236
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 34936 2204 35000 2208
rect 34936 2148 34940 2204
rect 34940 2148 34996 2204
rect 34996 2148 35000 2204
rect 34936 2144 35000 2148
rect 35016 2204 35080 2208
rect 35016 2148 35020 2204
rect 35020 2148 35076 2204
rect 35076 2148 35080 2204
rect 35016 2144 35080 2148
rect 35096 2204 35160 2208
rect 35096 2148 35100 2204
rect 35100 2148 35156 2204
rect 35156 2148 35160 2204
rect 35096 2144 35160 2148
rect 35176 2204 35240 2208
rect 35176 2148 35180 2204
rect 35180 2148 35236 2204
rect 35236 2148 35240 2204
rect 35176 2144 35240 2148
<< metal4 >>
rect 4208 37024 4528 37584
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 35936 4528 36960
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 19568 37568 19888 37584
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 36480 19888 37504
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 5027 35460 5093 35461
rect 5027 35396 5028 35460
rect 5092 35396 5093 35460
rect 5027 35395 5093 35396
rect 5030 35138 5090 35395
rect 19568 35392 19888 36416
rect 34928 37024 35248 37584
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 35936 35248 36960
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 24899 35868 24965 35869
rect 24899 35818 24900 35868
rect 24964 35818 24965 35868
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5472 4528 6496
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2128 4528 2144
rect 19568 34304 19888 35328
rect 20667 35324 20733 35325
rect 20667 35260 20668 35324
rect 20732 35260 20733 35324
rect 20667 35259 20733 35260
rect 21403 35324 21469 35325
rect 21403 35260 21404 35324
rect 21468 35260 21469 35324
rect 21403 35259 21469 35260
rect 20670 35138 20730 35259
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 33216 19888 34240
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 32128 19888 33152
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 31040 19888 32064
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 29952 19888 30976
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 28864 19888 29888
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 27776 19888 28800
rect 21406 28253 21466 35259
rect 24902 34781 24962 35582
rect 34928 34848 35248 35872
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 24899 34780 24965 34781
rect 24899 34716 24900 34780
rect 24964 34716 24965 34780
rect 24899 34715 24965 34716
rect 34928 33760 35248 34784
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 32672 35248 33696
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 31584 35248 32608
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 30496 35248 31520
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 29408 35248 30432
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 28320 35248 29344
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 21403 28252 21469 28253
rect 21403 28188 21404 28252
rect 21468 28188 21469 28252
rect 21403 28187 21469 28188
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 26688 19888 27712
rect 34651 27436 34717 27437
rect 34651 27372 34652 27436
rect 34716 27372 34717 27436
rect 34651 27371 34717 27372
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 25600 19888 26624
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 24512 19888 25536
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 23424 19888 24448
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 22336 19888 23360
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 21248 19888 22272
rect 34654 22269 34714 27371
rect 34928 27232 35248 28256
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 26144 35248 27168
rect 35387 26620 35453 26621
rect 35387 26556 35388 26620
rect 35452 26556 35453 26620
rect 35387 26555 35453 26556
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 25056 35248 26080
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 23968 35248 24992
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 22880 35248 23904
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34651 22268 34717 22269
rect 34651 22204 34652 22268
rect 34716 22204 34717 22268
rect 34651 22203 34717 22204
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20160 19888 21184
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 19072 19888 20096
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 17984 19888 19008
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 16896 19888 17920
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 15808 19888 16832
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 13632 19888 14656
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 10368 19888 11392
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 9280 19888 10304
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 6016 19888 7040
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 4928 19888 5952
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 3840 19888 4864
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 2752 19888 3776
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2128 19888 2688
rect 34928 21792 35248 22816
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 20704 35248 21728
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 19616 35248 20640
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 18528 35248 19552
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 17440 35248 18464
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 16352 35248 17376
rect 35390 16693 35450 26555
rect 35387 16692 35453 16693
rect 35387 16628 35388 16692
rect 35452 16628 35453 16692
rect 35387 16627 35453 16628
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 15264 35248 16288
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 14176 35248 15200
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 13088 35248 14112
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 12000 35248 13024
rect 35390 12477 35450 16627
rect 35387 12476 35453 12477
rect 35387 12412 35388 12476
rect 35452 12412 35453 12476
rect 35387 12411 35453 12412
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 10912 35248 11936
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 9824 35248 10848
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 8736 35248 9760
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 7648 35248 8672
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 6560 35248 7584
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 5472 35248 6496
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 4384 35248 5408
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 3296 35248 4320
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 2208 35248 3232
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2128 35248 2144
<< via4 >>
rect 6598 35732 6834 35818
rect 6598 35668 6684 35732
rect 6684 35668 6748 35732
rect 6748 35668 6834 35732
rect 6598 35582 6834 35668
rect 24814 35804 24900 35818
rect 24900 35804 24964 35818
rect 24964 35804 25050 35818
rect 24814 35582 25050 35804
rect 4942 34902 5178 35138
rect 20582 34902 20818 35138
<< metal5 >>
rect 6556 35818 25092 35860
rect 6556 35582 6598 35818
rect 6834 35582 24814 35818
rect 25050 35582 25092 35818
rect 6556 35540 25092 35582
rect 4900 35138 20860 35180
rect 4900 34902 4942 35138
rect 5178 34902 20582 35138
rect 20818 34902 20860 35138
rect 4900 34860 20860 34902
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1604681595
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1604681595
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1604681595
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1604681595
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1604681595
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _67_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8188 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75
timestamp 1604681595
transform 1 0 8004 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_81
timestamp 1604681595
transform 1 0 8556 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1604681595
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1604681595
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1604681595
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1604681595
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1604681595
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1604681595
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1604681595
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1604681595
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1604681595
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1604681595
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1604681595
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1604681595
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1604681595
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1604681595
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1604681595
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1604681595
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1604681595
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_230
timestamp 1604681595
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_220
timestamp 1604681595
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_232
timestamp 1604681595
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_242
timestamp 1604681595
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_249
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_261
timestamp 1604681595
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_245
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_257
timestamp 1604681595
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 27048 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 26680 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__CLK
timestamp 1604681595
transform 1 0 26588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_273
timestamp 1604681595
transform 1 0 26220 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_280
timestamp 1604681595
transform 1 0 26864 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_269
timestamp 1604681595
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_277 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 26588 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_280
timestamp 1604681595
transform 1 0 26864 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_284
timestamp 1604681595
transform 1 0 27232 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_290
timestamp 1604681595
transform 1 0 27784 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_286
timestamp 1604681595
transform 1 0 27416 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 27232 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1604681595
transform 1 0 27968 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1604681595
transform 1 0 27600 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1604681595
transform 1 0 27416 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 27600 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_301
timestamp 1604681595
transform 1 0 28796 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_297
timestamp 1604681595
transform 1 0 28428 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_300
timestamp 1604681595
transform 1 0 28704 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_294
timestamp 1604681595
transform 1 0 28152 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__CLK
timestamp 1604681595
transform 1 0 28520 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__D
timestamp 1604681595
transform 1 0 28888 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__D
timestamp 1604681595
transform 1 0 28888 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_304
timestamp 1604681595
transform 1 0 29072 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_304
timestamp 1604681595
transform 1 0 29072 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 29256 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_
timestamp 1604681595
transform 1 0 29716 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__D
timestamp 1604681595
transform 1 0 29256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__CLK
timestamp 1604681595
transform 1 0 31188 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_308
timestamp 1604681595
transform 1 0 29440 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_325
timestamp 1604681595
transform 1 0 31004 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_329
timestamp 1604681595
transform 1 0 31372 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1604681595
transform 1 0 32108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_334
timestamp 1604681595
transform 1 0 31832 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_330
timestamp 1604681595
transform 1 0 31464 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__D
timestamp 1604681595
transform 1 0 31924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__D
timestamp 1604681595
transform 1 0 31556 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1604681595
transform 1 0 32292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_
timestamp 1604681595
transform 1 0 31740 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_
timestamp 1604681595
transform 1 0 32568 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_1_360
timestamp 1604681595
transform 1 0 34224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_356
timestamp 1604681595
transform 1 0 33856 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_352
timestamp 1604681595
transform 1 0 33488 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__CLK
timestamp 1604681595
transform 1 0 34040 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__D
timestamp 1604681595
transform 1 0 33672 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_369
timestamp 1604681595
transform 1 0 35052 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_365
timestamp 1604681595
transform 1 0 34684 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_361
timestamp 1604681595
transform 1 0 34316 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__CLK
timestamp 1604681595
transform 1 0 34500 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__D
timestamp 1604681595
transform 1 0 35144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__D
timestamp 1604681595
transform 1 0 34592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_
timestamp 1604681595
transform 1 0 34868 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_
timestamp 1604681595
transform 1 0 35420 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1604681595
transform 1 0 36800 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1604681595
transform 1 0 37168 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_392
timestamp 1604681595
transform 1 0 37168 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_386
timestamp 1604681595
transform 1 0 36616 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1604681595
transform 1 0 36984 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_398
timestamp 1604681595
transform 1 0 37720 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_394
timestamp 1604681595
transform 1 0 37352 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_396
timestamp 1604681595
transform 1 0 37536 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__CLK
timestamp 1604681595
transform 1 0 37352 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1604681595
transform 1 0 37536 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_406
timestamp 1604681595
transform 1 0 38456 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_404
timestamp 1604681595
transform 1 0 38272 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_402
timestamp 1604681595
transform 1 0 38088 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 38824 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 38824 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604681595
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1604681595
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1604681595
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1604681595
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1604681595
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1604681595
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1604681595
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1604681595
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1604681595
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1604681595
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1604681595
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1604681595
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1604681595
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1604681595
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1604681595
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_251
timestamp 1604681595
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_263
timestamp 1604681595
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_276
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604681595
transform 1 0 27324 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_
timestamp 1604681595
transform 1 0 28888 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 28336 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__CLK
timestamp 1604681595
transform 1 0 28704 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_284
timestamp 1604681595
transform 1 0 27232 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_294
timestamp 1604681595
transform 1 0 28152 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_298
timestamp 1604681595
transform 1 0 28520 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 30820 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 31188 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_321
timestamp 1604681595
transform 1 0 30636 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_325
timestamp 1604681595
transform 1 0 31004 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604681595
transform 1 0 32292 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__CLK
timestamp 1604681595
transform 1 0 31740 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__CLK
timestamp 1604681595
transform 1 0 32844 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_329
timestamp 1604681595
transform 1 0 31372 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_335
timestamp 1604681595
transform 1 0 31924 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_337
timestamp 1604681595
transform 1 0 32108 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_343
timestamp 1604681595
transform 1 0 32660 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_347
timestamp 1604681595
transform 1 0 33028 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_
timestamp 1604681595
transform 1 0 33396 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_2_370
timestamp 1604681595
transform 1 0 35144 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604681595
transform 1 0 35880 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__CLK
timestamp 1604681595
transform 1 0 35328 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__CLK
timestamp 1604681595
transform 1 0 35696 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_374
timestamp 1604681595
transform 1 0 35512 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_387
timestamp 1604681595
transform 1 0 36708 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 38824 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_395
timestamp 1604681595
transform 1 0 37444 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_398
timestamp 1604681595
transform 1 0 37720 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_406
timestamp 1604681595
transform 1 0 38456 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1604681595
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1604681595
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1604681595
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1604681595
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1604681595
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1604681595
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1604681595
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1604681595
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1604681595
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1604681595
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1604681595
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1604681595
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1604681595
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_220
timestamp 1604681595
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_232
timestamp 1604681595
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_245
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_257
timestamp 1604681595
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 27048 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 26680 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_269
timestamp 1604681595
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_277
timestamp 1604681595
transform 1 0 26588 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_280
timestamp 1604681595
transform 1 0 26864 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604681595
transform 1 0 27600 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 28612 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__D
timestamp 1604681595
transform 1 0 28980 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 27416 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_284
timestamp 1604681595
transform 1 0 27232 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_297
timestamp 1604681595
transform 1 0 28428 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_301
timestamp 1604681595
transform 1 0 28796 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_
timestamp 1604681595
transform 1 0 29256 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 31188 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_325
timestamp 1604681595
transform 1 0 31004 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_
timestamp 1604681595
transform 1 0 31740 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__D
timestamp 1604681595
transform 1 0 31556 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_329
timestamp 1604681595
transform 1 0 31372 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__D
timestamp 1604681595
transform 1 0 35236 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__D
timestamp 1604681595
transform 1 0 34592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 33672 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 34040 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_352
timestamp 1604681595
transform 1 0 33488 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_356
timestamp 1604681595
transform 1 0 33856 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_360
timestamp 1604681595
transform 1 0 34224 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_367
timestamp 1604681595
transform 1 0 34868 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_
timestamp 1604681595
transform 1 0 35420 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_3_392
timestamp 1604681595
transform 1 0 37168 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 38824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_404
timestamp 1604681595
transform 1 0 38272 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604681595
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1604681595
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1604681595
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1604681595
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1604681595
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1604681595
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1604681595
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1604681595
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1604681595
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1604681595
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1604681595
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1604681595
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1604681595
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1604681595
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_239
timestamp 1604681595
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_251
timestamp 1604681595
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_263
timestamp 1604681595
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_276
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 27876 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 27600 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_290
timestamp 1604681595
transform 1 0 27784 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604681595
transform 1 0 30360 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 29808 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 30176 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_310
timestamp 1604681595
transform 1 0 29624 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_314
timestamp 1604681595
transform 1 0 29992 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_327
timestamp 1604681595
transform 1 0 31188 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604681595
transform 1 0 32108 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
timestamp 1604681595
transform 1 0 32660 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_335
timestamp 1604681595
transform 1 0 31924 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_341
timestamp 1604681595
transform 1 0 32476 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_345
timestamp 1604681595
transform 1 0 32844 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604681595
transform 1 0 33580 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_
timestamp 1604681595
transform 1 0 35144 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1604681595
transform 1 0 34960 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 33396 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__CLK
timestamp 1604681595
transform 1 0 34592 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_362
timestamp 1604681595
transform 1 0 34408 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_366
timestamp 1604681595
transform 1 0 34776 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_389
timestamp 1604681595
transform 1 0 36892 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 38824 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_398
timestamp 1604681595
transform 1 0 37720 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_406
timestamp 1604681595
transform 1 0 38456 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1604681595
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1604681595
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1604681595
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1604681595
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1604681595
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1604681595
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1604681595
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1604681595
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1604681595
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1604681595
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1604681595
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1604681595
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1604681595
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1604681595
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_220
timestamp 1604681595
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_232
timestamp 1604681595
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_245
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_257
timestamp 1604681595
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 26956 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 26588 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_269
timestamp 1604681595
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_279
timestamp 1604681595
transform 1 0 26772 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_283
timestamp 1604681595
transform 1 0 27140 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604681595
transform 1 0 27600 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 27324 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 28980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 28612 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_287
timestamp 1604681595
transform 1 0 27508 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_297
timestamp 1604681595
transform 1 0 28428 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_301
timestamp 1604681595
transform 1 0 28796 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 29256 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 31188 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_325
timestamp 1604681595
transform 1 0 31004 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604681595
transform 1 0 32384 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 32200 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 31832 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_329
timestamp 1604681595
transform 1 0 31372 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_333
timestamp 1604681595
transform 1 0 31740 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_336
timestamp 1604681595
transform 1 0 32016 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_349
timestamp 1604681595
transform 1 0 33212 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_353
timestamp 1604681595
transform 1 0 33580 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 33396 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_357
timestamp 1604681595
transform 1 0 33948 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 33764 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 34132 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_361
timestamp 1604681595
transform 1 0 34316 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1604681595
transform 1 0 34592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_367
timestamp 1604681595
transform 1 0 34868 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_371
timestamp 1604681595
transform 1 0 35236 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1604681595
transform 1 0 35052 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_
timestamp 1604681595
transform 1 0 35420 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_5_392
timestamp 1604681595
transform 1 0 37168 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 38824 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_404
timestamp 1604681595
transform 1 0 38272 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1604681595
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604681595
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1604681595
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1604681595
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1604681595
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1604681595
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1604681595
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1604681595
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1604681595
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1604681595
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1604681595
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1604681595
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1604681595
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1604681595
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1604681595
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1604681595
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1604681595
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1604681595
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1604681595
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1604681595
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1604681595
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1604681595
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1604681595
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1604681595
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1604681595
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1604681595
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_202
timestamp 1604681595
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1604681595
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_227
timestamp 1604681595
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_239
timestamp 1604681595
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_220
timestamp 1604681595
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_232
timestamp 1604681595
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_251
timestamp 1604681595
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_257
timestamp 1604681595
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 26496 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 27048 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 26128 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_263
timestamp 1604681595
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_276
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_269
timestamp 1604681595
transform 1 0 25852 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_274
timestamp 1604681595
transform 1 0 26312 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_278
timestamp 1604681595
transform 1 0 26680 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_284
timestamp 1604681595
transform 1 0 27232 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_284
timestamp 1604681595
transform 1 0 27232 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 27416 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604681595
transform 1 0 27600 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_301
timestamp 1604681595
transform 1 0 28796 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_297
timestamp 1604681595
transform 1 0 28428 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_304
timestamp 1604681595
transform 1 0 29072 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 28612 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 28980 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 27324 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_315
timestamp 1604681595
transform 1 0 30084 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_308
timestamp 1604681595
transform 1 0 29440 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 29624 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 29256 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604681595
transform 1 0 29808 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604681595
transform 1 0 29256 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_7_319
timestamp 1604681595
transform 1 0 30452 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_321
timestamp 1604681595
transform 1 0 30636 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 30268 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 30820 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 31004 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_327
timestamp 1604681595
transform 1 0 31188 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_337
timestamp 1604681595
transform 1 0 32108 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_337
timestamp 1604681595
transform 1 0 32108 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_330
timestamp 1604681595
transform 1 0 31464 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 31832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 31280 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604681595
transform 1 0 31280 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_341
timestamp 1604681595
transform 1 0 32476 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_347
timestamp 1604681595
transform 1 0 33028 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_342
timestamp 1604681595
transform 1 0 32568 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 32384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 32844 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 32292 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 32660 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604681595
transform 1 0 32844 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604681595
transform 1 0 33120 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_358
timestamp 1604681595
transform 1 0 34040 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_354
timestamp 1604681595
transform 1 0 33672 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_357
timestamp 1604681595
transform 1 0 33948 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 33856 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_362
timestamp 1604681595
transform 1 0 34408 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_365
timestamp 1604681595
transform 1 0 34684 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__CLK
timestamp 1604681595
transform 1 0 34776 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 34224 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
timestamp 1604681595
transform 1 0 34592 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604681595
transform 1 0 34868 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604681595
transform 1 0 34960 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_371
timestamp 1604681595
transform 1 0 35236 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_375
timestamp 1604681595
transform 1 0 35604 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_377
timestamp 1604681595
transform 1 0 35788 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
timestamp 1604681595
transform 1 0 35420 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__D
timestamp 1604681595
transform 1 0 35972 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 35972 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_387
timestamp 1604681595
transform 1 0 36708 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_383
timestamp 1604681595
transform 1 0 36340 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_393
timestamp 1604681595
transform 1 0 37260 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 36892 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 36524 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 37076 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_381
timestamp 1604681595
transform 1 0 36156 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 38824 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 38824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 37628 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_398
timestamp 1604681595
transform 1 0 37720 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_406
timestamp 1604681595
transform 1 0 38456 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_395
timestamp 1604681595
transform 1 0 37444 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_399
timestamp 1604681595
transform 1 0 37812 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604681595
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1604681595
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1604681595
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1604681595
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1604681595
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1604681595
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1604681595
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1604681595
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1604681595
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1604681595
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1604681595
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1604681595
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_190
timestamp 1604681595
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_202
timestamp 1604681595
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_227
timestamp 1604681595
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_239
timestamp 1604681595
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_251
timestamp 1604681595
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_263
timestamp 1604681595
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_295
timestamp 1604681595
transform 1 0 28244 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_303
timestamp 1604681595
transform 1 0 28980 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 30268 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 29256 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_308
timestamp 1604681595
transform 1 0 29440 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_316
timestamp 1604681595
transform 1 0 30176 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_321
timestamp 1604681595
transform 1 0 30636 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_327
timestamp 1604681595
transform 1 0 31188 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 32660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 32292 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 31280 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_prog_clk_A
timestamp 1604681595
transform 1 0 31648 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_330
timestamp 1604681595
transform 1 0 31464 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_334
timestamp 1604681595
transform 1 0 31832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_337
timestamp 1604681595
transform 1 0 32108 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_341
timestamp 1604681595
transform 1 0 32476 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 34224 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 33672 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_352
timestamp 1604681595
transform 1 0 33488 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_356
timestamp 1604681595
transform 1 0 33856 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_364
timestamp 1604681595
transform 1 0 34592 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604681595
transform 1 0 35328 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 36432 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
timestamp 1604681595
transform 1 0 35880 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 36248 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_376
timestamp 1604681595
transform 1 0 35696 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_380
timestamp 1604681595
transform 1 0 36064 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_388
timestamp 1604681595
transform 1 0 36800 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 38824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_396
timestamp 1604681595
transform 1 0 37536 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_398
timestamp 1604681595
transform 1 0 37720 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_406
timestamp 1604681595
transform 1 0 38456 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1604681595
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1604681595
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1604681595
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1604681595
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1604681595
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_86
timestamp 1604681595
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_98
timestamp 1604681595
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_110
timestamp 1604681595
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1604681595
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_147
timestamp 1604681595
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_159
timestamp 1604681595
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_171
timestamp 1604681595
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1604681595
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1604681595
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_220
timestamp 1604681595
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_232
timestamp 1604681595
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1604681595
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_269
timestamp 1604681595
transform 1 0 25852 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1604681595
transform 1 0 26956 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 28336 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 28704 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_293
timestamp 1604681595
transform 1 0 28060 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_298
timestamp 1604681595
transform 1 0 28520 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_302
timestamp 1604681595
transform 1 0 28888 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _38_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 29440 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 31096 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 30912 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_306
timestamp 1604681595
transform 1 0 29256 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_311
timestamp 1604681595
transform 1 0 29716 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_323
timestamp 1604681595
transform 1 0 30820 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 32200 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 32016 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 31648 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 33212 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_330
timestamp 1604681595
transform 1 0 31464 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_334
timestamp 1604681595
transform 1 0 31832 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_347
timestamp 1604681595
transform 1 0 33028 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_351
timestamp 1604681595
transform 1 0 33396 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 33580 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_359
timestamp 1604681595
transform 1 0 34132 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_355
timestamp 1604681595
transform 1 0 33764 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 33948 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_363
timestamp 1604681595
transform 1 0 34500 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_367
timestamp 1604681595
transform 1 0 34868 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 34592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1604681595
transform 1 0 35236 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 35420 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_9_392
timestamp 1604681595
transform 1 0 37168 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 38824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_404
timestamp 1604681595
transform 1 0 38272 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1604681595
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1604681595
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1604681595
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1604681595
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1604681595
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_80
timestamp 1604681595
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1604681595
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1604681595
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1604681595
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1604681595
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_166
timestamp 1604681595
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_178
timestamp 1604681595
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_190
timestamp 1604681595
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_202
timestamp 1604681595
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1604681595
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_239
timestamp 1604681595
transform 1 0 23092 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__CLK
timestamp 1604681595
transform 1 0 24104 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_247
timestamp 1604681595
transform 1 0 23828 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_252
timestamp 1604681595
transform 1 0 24288 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 26680 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 27048 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_prog_clk_A
timestamp 1604681595
transform 1 0 25944 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_264
timestamp 1604681595
transform 1 0 25392 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_10_272
timestamp 1604681595
transform 1 0 26128 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_276
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_280
timestamp 1604681595
transform 1 0 26864 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 28336 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_10_284
timestamp 1604681595
transform 1 0 27232 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1604681595
transform 1 0 31004 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 30268 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_315
timestamp 1604681595
transform 1 0 30084 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_319
timestamp 1604681595
transform 1 0 30452 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 32108 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 33212 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 32660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 33028 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 31832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_328
timestamp 1604681595
transform 1 0 31280 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_341
timestamp 1604681595
transform 1 0 32476 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_345
timestamp 1604681595
transform 1 0 32844 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 35236 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_368
timestamp 1604681595
transform 1 0 34960 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 35696 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_10_373
timestamp 1604681595
transform 1 0 35420 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_381
timestamp 1604681595
transform 1 0 36156 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_393
timestamp 1604681595
transform 1 0 37260 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 38824 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_398
timestamp 1604681595
transform 1 0 37720 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_406
timestamp 1604681595
transform 1 0 38456 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1604681595
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1604681595
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1604681595
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1604681595
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_74
timestamp 1604681595
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_86
timestamp 1604681595
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_98
timestamp 1604681595
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_110
timestamp 1604681595
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1604681595
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_147
timestamp 1604681595
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_159
timestamp 1604681595
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_171
timestamp 1604681595
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1604681595
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1604681595
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__CLK
timestamp 1604681595
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_220
timestamp 1604681595
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_232
timestamp 1604681595
transform 1 0 22448 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_240
timestamp 1604681595
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_
timestamp 1604681595
transform 1 0 24104 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__D
timestamp 1604681595
transform 1 0 23920 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__D
timestamp 1604681595
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_245
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604681595
transform 1 0 26588 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 26404 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 26036 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_269
timestamp 1604681595
transform 1 0 25852 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_273
timestamp 1604681595
transform 1 0 26220 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_286
timestamp 1604681595
transform 1 0 27416 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 27600 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_290
timestamp 1604681595
transform 1 0 27784 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_297
timestamp 1604681595
transform 1 0 28428 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_294
timestamp 1604681595
transform 1 0 28152 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 28244 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_301
timestamp 1604681595
transform 1 0 28796 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 28612 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 28980 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 29348 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_11_306
timestamp 1604681595
transform 1 0 29256 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_326
timestamp 1604681595
transform 1 0 31096 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 32292 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 31832 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 31648 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 31280 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_330
timestamp 1604681595
transform 1 0 31464 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp 1604681595
transform 1 0 32108 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 34868 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 34592 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 34224 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_358
timestamp 1604681595
transform 1 0 34040 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_362
timestamp 1604681595
transform 1 0 34408 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 36432 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 36984 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 35880 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 36248 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_376
timestamp 1604681595
transform 1 0 35696 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_380
timestamp 1604681595
transform 1 0 36064 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_388
timestamp 1604681595
transform 1 0 36800 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_392
timestamp 1604681595
transform 1 0 37168 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 38824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_404
timestamp 1604681595
transform 1 0 38272 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1604681595
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1604681595
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1604681595
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1604681595
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1604681595
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_105
timestamp 1604681595
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_117
timestamp 1604681595
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_129
timestamp 1604681595
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1604681595
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1604681595
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1604681595
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1604681595
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1604681595
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1604681595
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_239
timestamp 1604681595
transform 1 0 23092 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_
timestamp 1604681595
transform 1 0 23460 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__CLK
timestamp 1604681595
transform 1 0 23276 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_262
timestamp 1604681595
transform 1 0 25208 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_prog_clk
timestamp 1604681595
transform 1 0 25944 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_273
timestamp 1604681595
transform 1 0 26220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 29072 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 28888 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 28520 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_295
timestamp 1604681595
transform 1 0 28244 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_300
timestamp 1604681595
transform 1 0 28704 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 29532 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_12_307
timestamp 1604681595
transform 1 0 29348 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 32568 0 -1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 32292 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 31832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_328
timestamp 1604681595
transform 1 0 31280 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_337
timestamp 1604681595
transform 1 0 32108 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_341
timestamp 1604681595
transform 1 0 32476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 35236 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 34868 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_363
timestamp 1604681595
transform 1 0 34500 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_369
timestamp 1604681595
transform 1 0 35052 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 36248 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 36616 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_380
timestamp 1604681595
transform 1 0 36064 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_384
timestamp 1604681595
transform 1 0 36432 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_388
timestamp 1604681595
transform 1 0 36800 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 38824 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_396
timestamp 1604681595
transform 1 0 37536 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_398
timestamp 1604681595
transform 1 0 37720 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_406
timestamp 1604681595
transform 1 0 38456 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1604681595
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1604681595
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1604681595
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1604681595
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1604681595
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1604681595
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1604681595
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_74
timestamp 1604681595
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_86
timestamp 1604681595
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1604681595
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1604681595
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_98
timestamp 1604681595
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_105
timestamp 1604681595
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_110
timestamp 1604681595
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_117
timestamp 1604681595
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_129
timestamp 1604681595
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_135
timestamp 1604681595
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_147
timestamp 1604681595
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1604681595
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_159
timestamp 1604681595
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_171
timestamp 1604681595
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_154
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_166
timestamp 1604681595
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1604681595
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_178
timestamp 1604681595
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_190
timestamp 1604681595
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1604681595
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_202
timestamp 1604681595
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_229
timestamp 1604681595
transform 1 0 22172 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_228
timestamp 1604681595
transform 1 0 22080 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_220
timestamp 1604681595
transform 1 0 21344 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 21988 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_233
timestamp 1604681595
transform 1 0 22540 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_237
timestamp 1604681595
transform 1 0 22908 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_233
timestamp 1604681595
transform 1 0 22540 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__CLK
timestamp 1604681595
transform 1 0 22356 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__CLK
timestamp 1604681595
transform 1 0 22356 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__D
timestamp 1604681595
transform 1 0 22724 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_
timestamp 1604681595
transform 1 0 22724 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__D
timestamp 1604681595
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_241
timestamp 1604681595
transform 1 0 23276 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_254
timestamp 1604681595
transform 1 0 24472 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_272
timestamp 1604681595
transform 1 0 26128 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_266
timestamp 1604681595
transform 1 0 25576 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_268
timestamp 1604681595
transform 1 0 25760 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_264
timestamp 1604681595
transform 1 0 25392 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 25576 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 25944 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_280
timestamp 1604681595
transform 1 0 26864 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_276
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 26220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 26680 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 26128 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 26956 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_13_291
timestamp 1604681595
transform 1 0 27876 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 28060 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_295
timestamp 1604681595
transform 1 0 28244 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_300
timestamp 1604681595
transform 1 0 28704 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_301
timestamp 1604681595
transform 1 0 28796 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 28888 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 28612 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 28980 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_304
timestamp 1604681595
transform 1 0 29072 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 29808 0 1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 29440 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 29624 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 30452 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 29256 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_306
timestamp 1604681595
transform 1 0 29256 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_317
timestamp 1604681595
transform 1 0 30268 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1604681595
transform 1 0 30636 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_337
timestamp 1604681595
transform 1 0 32108 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_333
timestamp 1604681595
transform 1 0 31740 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_337
timestamp 1604681595
transform 1 0 32108 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_333
timestamp 1604681595
transform 1 0 31740 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 31924 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_343
timestamp 1604681595
transform 1 0 32660 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 32476 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 32292 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_prog_clk
timestamp 1604681595
transform 1 0 32844 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 32476 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_14_348
timestamp 1604681595
transform 1 0 33120 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_358
timestamp 1604681595
transform 1 0 34040 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_354
timestamp 1604681595
transform 1 0 33672 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_350
timestamp 1604681595
transform 1 0 33304 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 34224 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_prog_clk_A
timestamp 1604681595
transform 1 0 33856 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 33488 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_370
timestamp 1604681595
transform 1 0 35144 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_362
timestamp 1604681595
transform 1 0 34408 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 34592 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 34868 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 33396 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 35880 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 36800 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 35328 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_386
timestamp 1604681595
transform 1 0 36616 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_390
timestamp 1604681595
transform 1 0 36984 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_374
timestamp 1604681595
transform 1 0 35512 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_387
timestamp 1604681595
transform 1 0 36708 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1604681595
transform 1 0 37352 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 38824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 38824 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_397
timestamp 1604681595
transform 1 0 37628 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1604681595
transform 1 0 38364 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_395
timestamp 1604681595
transform 1 0 37444 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_398
timestamp 1604681595
transform 1 0 37720 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_406
timestamp 1604681595
transform 1 0 38456 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1604681595
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1604681595
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1604681595
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1604681595
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1604681595
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_74
timestamp 1604681595
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_86
timestamp 1604681595
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_98
timestamp 1604681595
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_110
timestamp 1604681595
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_135
timestamp 1604681595
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_147
timestamp 1604681595
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_159
timestamp 1604681595
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_171
timestamp 1604681595
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1604681595
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1604681595
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604681595
transform 1 0 21988 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 21804 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__D
timestamp 1604681595
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_220
timestamp 1604681595
transform 1 0 21344 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_224
timestamp 1604681595
transform 1 0 21712 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_236
timestamp 1604681595
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_240
timestamp 1604681595
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604681595
transform 1 0 23920 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 24932 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_245
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_257
timestamp 1604681595
transform 1 0 24748 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_261
timestamp 1604681595
transform 1 0 25116 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604681595
transform 1 0 26496 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 26312 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 25944 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
timestamp 1604681595
transform 1 0 25300 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_265
timestamp 1604681595
transform 1 0 25484 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_269
timestamp 1604681595
transform 1 0 25852 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_272
timestamp 1604681595
transform 1 0 26128 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_285
timestamp 1604681595
transform 1 0 27324 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 27508 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_289
timestamp 1604681595
transform 1 0 27692 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 27876 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 28060 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_296
timestamp 1604681595
transform 1 0 28336 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 28520 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_300
timestamp 1604681595
transform 1 0 28704 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 28980 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 29808 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 29624 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_306
timestamp 1604681595
transform 1 0 29256 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_321
timestamp 1604681595
transform 1 0 30636 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_333
timestamp 1604681595
transform 1 0 31740 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_345
timestamp 1604681595
transform 1 0 32844 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1604681595
transform 1 0 33764 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 35236 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_353
timestamp 1604681595
transform 1 0 33580 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_358
timestamp 1604681595
transform 1 0 34040 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_367
timestamp 1604681595
transform 1 0 34868 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 35420 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_15_392
timestamp 1604681595
transform 1 0 37168 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 38824 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_404
timestamp 1604681595
transform 1 0 38272 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1604681595
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1604681595
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1604681595
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1604681595
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1604681595
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_80
timestamp 1604681595
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_105
timestamp 1604681595
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_117
timestamp 1604681595
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_129
timestamp 1604681595
transform 1 0 12972 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1604681595
transform 1 0 14076 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_154
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_166
timestamp 1604681595
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_178
timestamp 1604681595
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_190
timestamp 1604681595
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_202
timestamp 1604681595
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_
timestamp 1604681595
transform 1 0 22356 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 21988 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_229
timestamp 1604681595
transform 1 0 22172 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 24288 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1604681595
transform 1 0 24104 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_254
timestamp 1604681595
transform 1 0 24472 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_262
timestamp 1604681595
transform 1 0 25208 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604681595
transform 1 0 26956 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604681595
transform 1 0 25300 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 26680 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_267
timestamp 1604681595
transform 1 0 25668 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_276
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_280
timestamp 1604681595
transform 1 0 26864 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 28520 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 27968 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 28336 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 29072 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_290
timestamp 1604681595
transform 1 0 27784 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_294
timestamp 1604681595
transform 1 0 28152 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_302
timestamp 1604681595
transform 1 0 28888 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 29808 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_306
timestamp 1604681595
transform 1 0 29256 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_314
timestamp 1604681595
transform 1 0 29992 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_326
timestamp 1604681595
transform 1 0 31096 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1604681595
transform 1 0 32108 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 31280 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_330
timestamp 1604681595
transform 1 0 31464 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_340
timestamp 1604681595
transform 1 0 32384 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _40_
timestamp 1604681595
transform 1 0 35052 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 34868 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_352
timestamp 1604681595
transform 1 0 33488 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_364
timestamp 1604681595
transform 1 0 34592 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_4.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 35512 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_372
timestamp 1604681595
transform 1 0 35328 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_376
timestamp 1604681595
transform 1 0 35696 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_388
timestamp 1604681595
transform 1 0 36800 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 38824 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_396
timestamp 1604681595
transform 1 0 37536 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_398
timestamp 1604681595
transform 1 0 37720 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_406
timestamp 1604681595
transform 1 0 38456 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1604681595
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1604681595
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1604681595
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1604681595
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_74
timestamp 1604681595
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_86
timestamp 1604681595
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_98
timestamp 1604681595
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_110
timestamp 1604681595
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_135
timestamp 1604681595
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_147
timestamp 1604681595
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_159
timestamp 1604681595
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_171
timestamp 1604681595
transform 1 0 16836 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1604681595
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1604681595
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__D
timestamp 1604681595
transform 1 0 22264 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__CLK
timestamp 1604681595
transform 1 0 22632 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_220
timestamp 1604681595
transform 1 0 21344 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_228
timestamp 1604681595
transform 1 0 22080 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_232
timestamp 1604681595
transform 1 0 22448 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_236
timestamp 1604681595
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_240
timestamp 1604681595
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604681595
transform 1 0 23736 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
timestamp 1604681595
transform 1 0 25116 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 24748 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_245
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_255
timestamp 1604681595
transform 1 0 24564 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_259
timestamp 1604681595
transform 1 0 24932 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_prog_clk
timestamp 1604681595
transform 1 0 26680 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 26496 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_prog_clk_A
timestamp 1604681595
transform 1 0 26128 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_263
timestamp 1604681595
transform 1 0 25300 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_271
timestamp 1604681595
transform 1 0 26036 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_274
timestamp 1604681595
transform 1 0 26312 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_281
timestamp 1604681595
transform 1 0 26956 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604681595
transform 1 0 27508 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 27324 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 28520 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 28980 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_296
timestamp 1604681595
transform 1 0 28336 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_300
timestamp 1604681595
transform 1 0 28704 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_310
timestamp 1604681595
transform 1 0 29624 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_306
timestamp 1604681595
transform 1 0 29256 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_313
timestamp 1604681595
transform 1 0 29900 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 29716 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 30084 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_317
timestamp 1604681595
transform 1 0 30268 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 30452 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_325
timestamp 1604681595
transform 1 0 31004 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_321
timestamp 1604681595
transform 1 0 30636 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 31096 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 31280 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 32752 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 33120 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_337
timestamp 1604681595
transform 1 0 32108 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_343
timestamp 1604681595
transform 1 0 32660 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_346
timestamp 1604681595
transform 1 0 32936 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_358
timestamp 1604681595
transform 1 0 34040 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_354
timestamp 1604681595
transform 1 0 33672 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_350
timestamp 1604681595
transform 1 0 33304 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 33856 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 33488 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_362
timestamp 1604681595
transform 1 0 34408 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 34224 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 34592 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 34868 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 35880 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_376
timestamp 1604681595
transform 1 0 35696 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_380
timestamp 1604681595
transform 1 0 36064 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_392
timestamp 1604681595
transform 1 0 37168 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 38824 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_404
timestamp 1604681595
transform 1 0 38272 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1604681595
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1604681595
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1604681595
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1604681595
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_80
timestamp 1604681595
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1604681595
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_117
timestamp 1604681595
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_129
timestamp 1604681595
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1604681595
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_166
timestamp 1604681595
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_178
timestamp 1604681595
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_190
timestamp 1604681595
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__CLK
timestamp 1604681595
transform 1 0 21068 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_202
timestamp 1604681595
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_215
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_
timestamp 1604681595
transform 1 0 22264 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_18_219
timestamp 1604681595
transform 1 0 21252 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_227
timestamp 1604681595
transform 1 0 21988 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604681595
transform 1 0 25116 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 24196 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 24564 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__CLK
timestamp 1604681595
transform 1 0 24932 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_249
timestamp 1604681595
transform 1 0 24012 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1604681595
transform 1 0 24380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_257
timestamp 1604681595
transform 1 0 24748 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
timestamp 1604681595
transform 1 0 26680 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__CLK
timestamp 1604681595
transform 1 0 25668 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_265
timestamp 1604681595
transform 1 0 25484 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_269
timestamp 1604681595
transform 1 0 25852 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_276
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_280
timestamp 1604681595
transform 1 0 26864 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604681595
transform 1 0 27416 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 28980 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 27232 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_295
timestamp 1604681595
transform 1 0 28244 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 30084 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 29532 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 29900 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 31096 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_307
timestamp 1604681595
transform 1 0 29348 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_311
timestamp 1604681595
transform 1 0 29716 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_324
timestamp 1604681595
transform 1 0 30912 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 32752 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 32568 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 31464 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 31832 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_328
timestamp 1604681595
transform 1 0 31280 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_332
timestamp 1604681595
transform 1 0 31648 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_337
timestamp 1604681595
transform 1 0 32108 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_341
timestamp 1604681595
transform 1 0 32476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 34316 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 33764 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 34132 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_353
timestamp 1604681595
transform 1 0 33580 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_357
timestamp 1604681595
transform 1 0 33948 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 36248 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_380
timestamp 1604681595
transform 1 0 36064 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_384
timestamp 1604681595
transform 1 0 36432 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 38824 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_396
timestamp 1604681595
transform 1 0 37536 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_398
timestamp 1604681595
transform 1 0 37720 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_406
timestamp 1604681595
transform 1 0 38456 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1604681595
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1604681595
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1604681595
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1604681595
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1604681595
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1604681595
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1604681595
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1604681595
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_86
timestamp 1604681595
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1604681595
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1604681595
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_98
timestamp 1604681595
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1604681595
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_110
timestamp 1604681595
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1604681595
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1604681595
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1604681595
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_147
timestamp 1604681595
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1604681595
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_159
timestamp 1604681595
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_171
timestamp 1604681595
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1604681595
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1604681595
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1604681595
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_190
timestamp 1604681595
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_
timestamp 1604681595
transform 1 0 21068 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__D
timestamp 1604681595
transform 1 0 20884 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_208
timestamp 1604681595
transform 1 0 20240 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_214
timestamp 1604681595
transform 1 0 20792 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_202
timestamp 1604681595
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604681595
transform 1 0 22356 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 22172 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_236
timestamp 1604681595
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_240
timestamp 1604681595
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_227
timestamp 1604681595
transform 1 0 21988 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_240
timestamp 1604681595
transform 1 0 23184 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_245
timestamp 1604681595
transform 1 0 23644 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1604681595
transform 1 0 23460 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_19_262
timestamp 1604681595
transform 1 0 25208 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_258
timestamp 1604681595
transform 1 0 24840 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_254
timestamp 1604681595
transform 1 0 24472 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 25024 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__D
timestamp 1604681595
transform 1 0 24656 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_
timestamp 1604681595
transform 1 0 23920 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_
timestamp 1604681595
transform 1 0 25668 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__D
timestamp 1604681595
transform 1 0 25484 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1604681595
transform 1 0 27048 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_267
timestamp 1604681595
transform 1 0 25668 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_280
timestamp 1604681595
transform 1 0 26864 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_284
timestamp 1604681595
transform 1 0 27232 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_294
timestamp 1604681595
transform 1 0 28152 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_290
timestamp 1604681595
transform 1 0 27784 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_286
timestamp 1604681595
transform 1 0 27416 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__CLK
timestamp 1604681595
transform 1 0 27968 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__CLK
timestamp 1604681595
transform 1 0 27416 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__D
timestamp 1604681595
transform 1 0 27600 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_302
timestamp 1604681595
transform 1 0 28888 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604681595
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_
timestamp 1604681595
transform 1 0 27600 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_20_311
timestamp 1604681595
transform 1 0 29716 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_307
timestamp 1604681595
transform 1 0 29348 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_313
timestamp 1604681595
transform 1 0 29900 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_306
timestamp 1604681595
transform 1 0 29256 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 29900 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__CLK
timestamp 1604681595
transform 1 0 29532 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 30084 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 29532 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604681595
transform 1 0 30084 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_324
timestamp 1604681595
transform 1 0 30912 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_317
timestamp 1604681595
transform 1 0 30268 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 31096 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 30452 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 30636 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_20_337
timestamp 1604681595
transform 1 0 32108 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_328
timestamp 1604681595
transform 1 0 31280 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 31832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604681595
transform 1 0 32016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_345
timestamp 1604681595
transform 1 0 32844 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_340
timestamp 1604681595
transform 1 0 32384 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 32476 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 32660 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 33120 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 32660 0 -1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_19_357
timestamp 1604681595
transform 1 0 33948 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 34132 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_368
timestamp 1604681595
transform 1 0 34960 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_364
timestamp 1604681595
transform 1 0 34592 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_367
timestamp 1604681595
transform 1 0 34868 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_361
timestamp 1604681595
transform 1 0 34316 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 34776 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 35144 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 34592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604681595
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 35144 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_20_382
timestamp 1604681595
transform 1 0 36248 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_372
timestamp 1604681595
transform 1 0 35328 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 35420 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_20_390
timestamp 1604681595
transform 1 0 36984 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_386
timestamp 1604681595
transform 1 0 36616 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_389
timestamp 1604681595
transform 1 0 36892 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 36800 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 37076 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 36432 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1604681595
transform 1 0 37260 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 38824 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 38824 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604681595
transform 1 0 37628 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1604681595
transform 1 0 38364 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_396
timestamp 1604681595
transform 1 0 37536 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_398
timestamp 1604681595
transform 1 0 37720 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_406
timestamp 1604681595
transform 1 0 38456 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1604681595
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1604681595
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1604681595
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1604681595
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1604681595
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1604681595
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_98
timestamp 1604681595
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_110
timestamp 1604681595
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1604681595
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_147
timestamp 1604681595
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_159
timestamp 1604681595
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_171
timestamp 1604681595
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1604681595
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1604681595
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1604681595
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1604681595
transform 1 0 22632 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_220
timestamp 1604681595
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_232
timestamp 1604681595
transform 1 0 22448 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_236
timestamp 1604681595
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_240
timestamp 1604681595
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__D
timestamp 1604681595
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_
timestamp 1604681595
transform 1 0 26680 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1604681595
transform 1 0 26496 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__D
timestamp 1604681595
transform 1 0 26128 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1604681595
transform 1 0 25760 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_264
timestamp 1604681595
transform 1 0 25392 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_270
timestamp 1604681595
transform 1 0 25944 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_274
timestamp 1604681595
transform 1 0 26312 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604681595
transform 1 0 29164 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__D
timestamp 1604681595
transform 1 0 28704 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_297
timestamp 1604681595
transform 1 0 28428 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_302
timestamp 1604681595
transform 1 0 28888 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 29716 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 29532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_306
timestamp 1604681595
transform 1 0 29256 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 32292 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 32108 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 31740 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_330
timestamp 1604681595
transform 1 0 31464 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_335
timestamp 1604681595
transform 1 0 31924 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604681595
transform 1 0 34776 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 34224 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 35236 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 34592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_358
timestamp 1604681595
transform 1 0 34040 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_362
timestamp 1604681595
transform 1 0 34408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_367
timestamp 1604681595
transform 1 0 34868 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 35420 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_21_392
timestamp 1604681595
transform 1 0 37168 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 38824 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 37352 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_396
timestamp 1604681595
transform 1 0 37536 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_404
timestamp 1604681595
transform 1 0 38272 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1604681595
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1604681595
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1604681595
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1604681595
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_80
timestamp 1604681595
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_105
timestamp 1604681595
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_117
timestamp 1604681595
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_129
timestamp 1604681595
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1604681595
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1604681595
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1604681595
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1604681595
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__CLK
timestamp 1604681595
transform 1 0 21068 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_202
timestamp 1604681595
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_219
timestamp 1604681595
transform 1 0 21252 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_231
timestamp 1604681595
transform 1 0 22356 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604681595
transform 1 0 23460 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__CLK
timestamp 1604681595
transform 1 0 24472 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_252
timestamp 1604681595
transform 1 0 24288 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_256
timestamp 1604681595
transform 1 0 24656 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_268
timestamp 1604681595
transform 1 0 25760 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_274
timestamp 1604681595
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_
timestamp 1604681595
transform 1 0 28704 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1604681595
transform 1 0 27508 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_285
timestamp 1604681595
transform 1 0 27324 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_289
timestamp 1604681595
transform 1 0 27692 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_297
timestamp 1604681595
transform 1 0 28428 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_319
timestamp 1604681595
transform 1 0 30452 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_337
timestamp 1604681595
transform 1 0 32108 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_331
timestamp 1604681595
transform 1 0 31556 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 31832 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604681595
transform 1 0 32016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1604681595
transform 1 0 32200 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_345
timestamp 1604681595
transform 1 0 32844 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_341
timestamp 1604681595
transform 1 0 32476 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 32660 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 33028 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 33212 0 -1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_22_370
timestamp 1604681595
transform 1 0 35144 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 35880 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 35420 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_375
timestamp 1604681595
transform 1 0 35604 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_387
timestamp 1604681595
transform 1 0 36708 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 38824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604681595
transform 1 0 37628 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_395
timestamp 1604681595
transform 1 0 37444 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_398
timestamp 1604681595
transform 1 0 37720 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_406
timestamp 1604681595
transform 1 0 38456 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1604681595
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1604681595
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1604681595
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1604681595
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1604681595
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1604681595
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1604681595
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_110
timestamp 1604681595
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1604681595
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1604681595
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_159
timestamp 1604681595
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_171
timestamp 1604681595
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_196
timestamp 1604681595
transform 1 0 19136 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_
timestamp 1604681595
transform 1 0 21068 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__D
timestamp 1604681595
transform 1 0 20884 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__D
timestamp 1604681595
transform 1 0 20516 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__CLK
timestamp 1604681595
transform 1 0 20148 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_204
timestamp 1604681595
transform 1 0 19872 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_209
timestamp 1604681595
transform 1 0 20332 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_213
timestamp 1604681595
transform 1 0 20700 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_236
timestamp 1604681595
transform 1 0 22816 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_245
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_257
timestamp 1604681595
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604681595
transform 1 0 26588 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 26404 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 26036 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_269
timestamp 1604681595
transform 1 0 25852 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_273
timestamp 1604681595
transform 1 0 26220 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1604681595
transform 1 0 29164 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1604681595
transform 1 0 27600 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1604681595
transform 1 0 27968 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 28980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_286
timestamp 1604681595
transform 1 0 27416 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_290
timestamp 1604681595
transform 1 0 27784 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_294
timestamp 1604681595
transform 1 0 28152 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_302
timestamp 1604681595
transform 1 0 28888 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 31004 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604681595
transform 1 0 29808 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1604681595
transform 1 0 30452 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
timestamp 1604681595
transform 1 0 29624 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 30820 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_306
timestamp 1604681595
transform 1 0 29256 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_317
timestamp 1604681595
transform 1 0 30268 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_321
timestamp 1604681595
transform 1 0 30636 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 32292 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 32108 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 31740 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_329
timestamp 1604681595
transform 1 0 31372 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_335
timestamp 1604681595
transform 1 0 31924 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1604681595
transform 1 0 34776 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 35236 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 34592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_358
timestamp 1604681595
transform 1 0 34040 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_367
timestamp 1604681595
transform 1 0 34868 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 35420 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_23_392
timestamp 1604681595
transform 1 0 37168 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 38824 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_404
timestamp 1604681595
transform 1 0 38272 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1604681595
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1604681595
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1604681595
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1604681595
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1604681595
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1604681595
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1604681595
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1604681595
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1604681595
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1604681595
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1604681595
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1604681595
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_202
timestamp 1604681595
transform 1 0 19688 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_210
timestamp 1604681595
transform 1 0 20424 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_234
timestamp 1604681595
transform 1 0 22632 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_246
timestamp 1604681595
transform 1 0 23736 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_258
timestamp 1604681595
transform 1 0 24840 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 26680 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25484 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 27048 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_264
timestamp 1604681595
transform 1 0 25392 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_267
timestamp 1604681595
transform 1 0 25668 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_276
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_280
timestamp 1604681595
transform 1 0 26864 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604681595
transform 1 0 27324 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_24_284
timestamp 1604681595
transform 1 0 27232 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_294
timestamp 1604681595
transform 1 0 28152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 29716 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 30268 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_306
timestamp 1604681595
transform 1 0 29256 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_310
timestamp 1604681595
transform 1 0 29624 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_315
timestamp 1604681595
transform 1 0 30084 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_319
timestamp 1604681595
transform 1 0 30452 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 32384 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1604681595
transform 1 0 32016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_331
timestamp 1604681595
transform 1 0 31556 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_335
timestamp 1604681595
transform 1 0 31924 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_337
timestamp 1604681595
transform 1 0 32108 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_349
timestamp 1604681595
transform 1 0 33212 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_361
timestamp 1604681595
transform 1 0 34316 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 35420 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 35972 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_377
timestamp 1604681595
transform 1 0 35788 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_381
timestamp 1604681595
transform 1 0 36156 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_393
timestamp 1604681595
transform 1 0 37260 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 38824 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1604681595
transform 1 0 37628 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_398
timestamp 1604681595
transform 1 0 37720 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_406
timestamp 1604681595
transform 1 0 38456 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1604681595
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1604681595
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1604681595
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1604681595
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1604681595
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1604681595
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1604681595
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1604681595
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1604681595
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_147
timestamp 1604681595
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_159
timestamp 1604681595
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_171
timestamp 1604681595
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_184
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_192
timestamp 1604681595
transform 1 0 18768 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_195
timestamp 1604681595
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_
timestamp 1604681595
transform 1 0 20700 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 19228 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__D
timestamp 1604681595
transform 1 0 20516 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 19596 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__D
timestamp 1604681595
transform 1 0 20148 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_199
timestamp 1604681595
transform 1 0 19412 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_203
timestamp 1604681595
transform 1 0 19780 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_209
timestamp 1604681595
transform 1 0 20332 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__CLK
timestamp 1604681595
transform 1 0 22632 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_232
timestamp 1604681595
transform 1 0 22448 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_236
timestamp 1604681595
transform 1 0 22816 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23920 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24840 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 24288 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_245
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_250
timestamp 1604681595
transform 1 0 24104 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_254
timestamp 1604681595
transform 1 0 24472 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_260
timestamp 1604681595
transform 1 0 25024 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 25484 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 25300 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 27968 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1604681595
transform 1 0 29164 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 28520 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 27416 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_284
timestamp 1604681595
transform 1 0 27232 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_288
timestamp 1604681595
transform 1 0 27600 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_296
timestamp 1604681595
transform 1 0 28336 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_300
timestamp 1604681595
transform 1 0 28704 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_304
timestamp 1604681595
transform 1 0 29072 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 29256 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 29808 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 30176 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 30544 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_310
timestamp 1604681595
transform 1 0 29624 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_314
timestamp 1604681595
transform 1 0 29992 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_318
timestamp 1604681595
transform 1 0 30360 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_322
timestamp 1604681595
transform 1 0 30728 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_5.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 32384 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_334
timestamp 1604681595
transform 1 0 31832 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_342
timestamp 1604681595
transform 1 0 32568 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1604681595
transform 1 0 34776 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_354
timestamp 1604681595
transform 1 0 33672 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_367
timestamp 1604681595
transform 1 0 34868 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1604681595
transform 1 0 35420 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_376
timestamp 1604681595
transform 1 0 35696 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_388
timestamp 1604681595
transform 1 0 36800 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 38824 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_400
timestamp 1604681595
transform 1 0 37904 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_406
timestamp 1604681595
transform 1 0 38456 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1604681595
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1604681595
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1604681595
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1604681595
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1604681595
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1604681595
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1604681595
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1604681595
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1604681595
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1604681595
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1604681595
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1604681595
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1604681595
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1604681595
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1604681595
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_110
timestamp 1604681595
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1604681595
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_135
timestamp 1604681595
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_147
timestamp 1604681595
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1604681595
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_159
timestamp 1604681595
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_171
timestamp 1604681595
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604681595
transform 1 0 18952 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 18768 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 18952 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1604681595
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_190
timestamp 1604681595
transform 1 0 18584 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_196
timestamp 1604681595
transform 1 0 19136 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_203
timestamp 1604681595
transform 1 0 19780 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_206
timestamp 1604681595
transform 1 0 20056 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604681595
transform 1 0 19228 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_26_213
timestamp 1604681595
transform 1 0 20700 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_210
timestamp 1604681595
transform 1 0 20424 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__CLK
timestamp 1604681595
transform 1 0 20516 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__D
timestamp 1604681595
transform 1 0 20332 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_
timestamp 1604681595
transform 1 0 20516 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 22448 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_234
timestamp 1604681595
transform 1 0 22632 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_230
timestamp 1604681595
transform 1 0 22264 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_234
timestamp 1604681595
transform 1 0 22632 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_238
timestamp 1604681595
transform 1 0 23000 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_249
timestamp 1604681595
transform 1 0 24012 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_247
timestamp 1604681595
transform 1 0 23828 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_242
timestamp 1604681595
transform 1 0 23368 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
timestamp 1604681595
transform 1 0 23644 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
timestamp 1604681595
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_254
timestamp 1604681595
transform 1 0 24472 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 24288 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 24656 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 24840 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23920 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 26772 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 27140 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 25852 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_267
timestamp 1604681595
transform 1 0 25668 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_271
timestamp 1604681595
transform 1 0 26036 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_277
timestamp 1604681595
transform 1 0 26588 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1604681595
transform 1 0 26956 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_293
timestamp 1604681595
transform 1 0 28060 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_289
timestamp 1604681595
transform 1 0 27692 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_285
timestamp 1604681595
transform 1 0 27324 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 27876 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1604681595
transform 1 0 27416 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_297
timestamp 1604681595
transform 1 0 28428 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 28980 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 28244 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1604681595
transform 1 0 29164 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_295
timestamp 1604681595
transform 1 0 28244 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_310
timestamp 1604681595
transform 1 0 29624 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_306
timestamp 1604681595
transform 1 0 29256 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_307
timestamp 1604681595
transform 1 0 29348 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 29440 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 29992 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 29900 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_26_326
timestamp 1604681595
transform 1 0 31096 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_322
timestamp 1604681595
transform 1 0 30728 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 30912 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 30176 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_27_335
timestamp 1604681595
transform 1 0 31924 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_334
timestamp 1604681595
transform 1 0 31832 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 32108 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1604681595
transform 1 0 32016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_347
timestamp 1604681595
transform 1 0 33028 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_343
timestamp 1604681595
transform 1 0 32660 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_339
timestamp 1604681595
transform 1 0 32292 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 32844 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 32476 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_349
timestamp 1604681595
transform 1 0 33212 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_337
timestamp 1604681595
transform 1 0 32108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_360
timestamp 1604681595
transform 1 0 34224 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_355
timestamp 1604681595
transform 1 0 33764 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 33580 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 34040 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_371
timestamp 1604681595
transform 1 0 35236 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_367
timestamp 1604681595
transform 1 0 34868 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_364
timestamp 1604681595
transform 1 0 34592 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 35052 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 34408 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1604681595
transform 1 0 34776 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_361
timestamp 1604681595
transform 1 0 34316 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 35420 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 35420 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_375
timestamp 1604681595
transform 1 0 35604 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_387
timestamp 1604681595
transform 1 0 36708 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_392
timestamp 1604681595
transform 1 0 37168 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 38824 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 38824 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1604681595
transform 1 0 37628 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_395
timestamp 1604681595
transform 1 0 37444 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_398
timestamp 1604681595
transform 1 0 37720 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_406
timestamp 1604681595
transform 1 0 38456 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_404
timestamp 1604681595
transform 1 0 38272 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1604681595
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1604681595
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1604681595
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1604681595
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1604681595
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1604681595
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1604681595
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_129
timestamp 1604681595
transform 1 0 12972 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__CLK
timestamp 1604681595
transform 1 0 13984 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp 1604681595
transform 1 0 13708 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_142
timestamp 1604681595
transform 1 0 14168 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_150
timestamp 1604681595
transform 1 0 14904 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__CLK
timestamp 1604681595
transform 1 0 15456 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_154
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_158
timestamp 1604681595
transform 1 0 15640 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_170
timestamp 1604681595
transform 1 0 16744 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 18400 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 18952 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__CLK
timestamp 1604681595
transform 1 0 18032 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_182
timestamp 1604681595
transform 1 0 17848 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_186
timestamp 1604681595
transform 1 0 18216 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_190
timestamp 1604681595
transform 1 0 18584 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_196
timestamp 1604681595
transform 1 0 19136 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__D
timestamp 1604681595
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 19780 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 20148 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__CLK
timestamp 1604681595
transform 1 0 21068 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_202
timestamp 1604681595
transform 1 0 19688 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_205
timestamp 1604681595
transform 1 0 19964 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_209
timestamp 1604681595
transform 1 0 20332 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604681595
transform 1 0 21804 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 21620 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_219
timestamp 1604681595
transform 1 0 21252 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_234
timestamp 1604681595
transform 1 0 22632 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24840 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604681595
transform 1 0 23368 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 24656 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 24288 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23920 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_246
timestamp 1604681595
transform 1 0 23736 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1604681595
transform 1 0 24104 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_254
timestamp 1604681595
transform 1 0 24472 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 25852 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_267
timestamp 1604681595
transform 1 0 25668 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_271
timestamp 1604681595
transform 1 0 26036 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 27784 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 28152 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 29072 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_285
timestamp 1604681595
transform 1 0 27324 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_289
timestamp 1604681595
transform 1 0 27692 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_292
timestamp 1604681595
transform 1 0 27968 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_296
timestamp 1604681595
transform 1 0 28336 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 29256 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 31188 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_325
timestamp 1604681595
transform 1 0 31004 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 32108 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1604681595
transform 1 0 32016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 33212 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_329
timestamp 1604681595
transform 1 0 31372 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_335
timestamp 1604681595
transform 1 0 31924 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_346
timestamp 1604681595
transform 1 0 32936 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 34408 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 33580 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 33948 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_351
timestamp 1604681595
transform 1 0 33396 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_355
timestamp 1604681595
transform 1 0 33764 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_359
timestamp 1604681595
transform 1 0 34132 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_371
timestamp 1604681595
transform 1 0 35236 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _50_
timestamp 1604681595
transform 1 0 35972 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 35420 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 35788 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_375
timestamp 1604681595
transform 1 0 35604 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_382
timestamp 1604681595
transform 1 0 36248 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 38824 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1604681595
transform 1 0 37628 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_394
timestamp 1604681595
transform 1 0 37352 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_398
timestamp 1604681595
transform 1 0 37720 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_406
timestamp 1604681595
transform 1 0 38456 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1604681595
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1604681595
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1604681595
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1604681595
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1604681595
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_86
timestamp 1604681595
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_98
timestamp 1604681595
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_110
timestamp 1604681595
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_
timestamp 1604681595
transform 1 0 13984 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__D
timestamp 1604681595
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_135
timestamp 1604681595
transform 1 0 13524 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__D
timestamp 1604681595
transform 1 0 15916 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__CLK
timestamp 1604681595
transform 1 0 16284 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_159
timestamp 1604681595
transform 1 0 15732 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_163
timestamp 1604681595
transform 1 0 16100 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_167
timestamp 1604681595
transform 1 0 16468 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__D
timestamp 1604681595
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_179
timestamp 1604681595
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604681595
transform 1 0 19780 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_
timestamp 1604681595
transform 1 0 20608 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 22540 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 22908 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_231
timestamp 1604681595
transform 1 0 22356 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_235
timestamp 1604681595
transform 1 0 22724 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_239
timestamp 1604681595
transform 1 0 23092 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604681595
transform 1 0 24380 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 24196 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23828 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
timestamp 1604681595
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_245
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_249
timestamp 1604681595
transform 1 0 24012 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_262
timestamp 1604681595
transform 1 0 25208 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 25944 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 25392 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 25760 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_266
timestamp 1604681595
transform 1 0 25576 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 27784 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1604681595
transform 1 0 29164 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 28336 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 28704 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_294
timestamp 1604681595
transform 1 0 28152 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_298
timestamp 1604681595
transform 1 0 28520 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_302
timestamp 1604681595
transform 1 0 28888 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1604681595
transform 1 0 29532 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 30544 0 1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 30360 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 29992 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_306
timestamp 1604681595
transform 1 0 29256 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_312
timestamp 1604681595
transform 1 0 29808 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_316
timestamp 1604681595
transform 1 0 30176 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 33212 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 33028 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 32660 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_341
timestamp 1604681595
transform 1 0 32476 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_345
timestamp 1604681595
transform 1 0 32844 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 35052 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1604681595
transform 1 0 34776 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 34224 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 34592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_358
timestamp 1604681595
transform 1 0 34040 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_362
timestamp 1604681595
transform 1 0 34408 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_367
timestamp 1604681595
transform 1 0 34868 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_388
timestamp 1604681595
transform 1 0 36800 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 38824 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_400
timestamp 1604681595
transform 1 0 37904 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_406
timestamp 1604681595
transform 1 0 38456 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1604681595
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1604681595
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1604681595
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1604681595
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1604681595
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1604681595
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1604681595
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_117
timestamp 1604681595
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_129
timestamp 1604681595
transform 1 0 12972 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 13524 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_137
timestamp 1604681595
transform 1 0 13708 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 1604681595
transform 1 0 14812 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_173
timestamp 1604681595
transform 1 0 17020 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk
timestamp 1604681595
transform 1 0 18400 0 -1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__D
timestamp 1604681595
transform 1 0 18032 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__CLK
timestamp 1604681595
transform 1 0 17664 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_179
timestamp 1604681595
transform 1 0 17572 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_182
timestamp 1604681595
transform 1 0 17848 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_186
timestamp 1604681595
transform 1 0 18216 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 20424 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_208
timestamp 1604681595
transform 1 0 20240 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1604681595
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604681595
transform 1 0 21896 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__D
timestamp 1604681595
transform 1 0 21344 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 21712 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1604681595
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_222
timestamp 1604681595
transform 1 0 21528 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_235
timestamp 1604681595
transform 1 0 22724 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604681595
transform 1 0 24840 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604681595
transform 1 0 23736 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 24564 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_243
timestamp 1604681595
transform 1 0 23460 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_250
timestamp 1604681595
transform 1 0 24104 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_254
timestamp 1604681595
transform 1 0 24472 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_257
timestamp 1604681595
transform 1 0 24748 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 26864 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0__f_clk_A
timestamp 1604681595
transform 1 0 25944 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_267
timestamp 1604681595
transform 1 0 25668 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_272
timestamp 1604681595
transform 1 0 26128 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 27968 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 27416 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 27784 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 28980 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_284
timestamp 1604681595
transform 1 0 27232 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_288
timestamp 1604681595
transform 1 0 27600 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_301
timestamp 1604681595
transform 1 0 28796 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_305
timestamp 1604681595
transform 1 0 29164 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 29532 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 29348 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1604681595
transform 1 0 32108 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1604681595
transform 1 0 32016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 32568 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 31464 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_328
timestamp 1604681595
transform 1 0 31280 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_332
timestamp 1604681595
transform 1 0 31648 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_340
timestamp 1604681595
transform 1 0 32384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_344
timestamp 1604681595
transform 1 0 32752 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 33580 0 -1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 33396 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_350
timestamp 1604681595
transform 1 0 33304 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _49_
timestamp 1604681595
transform 1 0 36248 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 35696 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 36064 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_374
timestamp 1604681595
transform 1 0 35512 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_378
timestamp 1604681595
transform 1 0 35880 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_385
timestamp 1604681595
transform 1 0 36524 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 38824 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1604681595
transform 1 0 37628 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_398
timestamp 1604681595
transform 1 0 37720 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_406
timestamp 1604681595
transform 1 0 38456 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 1564 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_7
timestamp 1604681595
transform 1 0 1748 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_11
timestamp 1604681595
transform 1 0 2116 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_23
timestamp 1604681595
transform 1 0 3220 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_35
timestamp 1604681595
transform 1 0 4324 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_47
timestamp 1604681595
transform 1 0 5428 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1604681595
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1604681595
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1604681595
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__CLK
timestamp 1604681595
transform 1 0 12880 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1604681595
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_127
timestamp 1604681595
transform 1 0 12788 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_130
timestamp 1604681595
transform 1 0 13064 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_
timestamp 1604681595
transform 1 0 13432 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__D
timestamp 1604681595
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604681595
transform 1 0 15916 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1604681595
transform 1 0 15732 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__D
timestamp 1604681595
transform 1 0 15364 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1604681595
transform 1 0 16928 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_153
timestamp 1604681595
transform 1 0 15180 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_157
timestamp 1604681595
transform 1 0 15548 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_170
timestamp 1604681595
transform 1 0 16744 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_174
timestamp 1604681595
transform 1 0 17112 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1604681595
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1604681595
transform 1 0 17296 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_178
timestamp 1604681595
transform 1 0 17480 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_
timestamp 1604681595
transform 1 0 20976 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1604681595
transform 1 0 19964 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__D
timestamp 1604681595
transform 1 0 20792 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__CLK
timestamp 1604681595
transform 1 0 20424 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_203
timestamp 1604681595
transform 1 0 19780 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_207
timestamp 1604681595
transform 1 0 20148 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_212
timestamp 1604681595
transform 1 0 20608 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__CLK
timestamp 1604681595
transform 1 0 22908 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_235
timestamp 1604681595
transform 1 0 22724 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_239
timestamp 1604681595
transform 1 0 23092 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604681595
transform 1 0 24564 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 24380 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 24012 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_245
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_251
timestamp 1604681595
transform 1 0 24196 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 27048 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 26496 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 26864 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 25576 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 25944 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_264
timestamp 1604681595
transform 1 0 25392 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_268
timestamp 1604681595
transform 1 0 25760 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_272
timestamp 1604681595
transform 1 0 26128 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1604681595
transform 1 0 26680 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1604681595
transform 1 0 29164 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 28980 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 28060 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 28612 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_291
timestamp 1604681595
transform 1 0 27876 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_295
timestamp 1604681595
transform 1 0 28244 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_301
timestamp 1604681595
transform 1 0 28796 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 29624 0 1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 29440 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_306
timestamp 1604681595
transform 1 0 29256 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 32292 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 32108 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 31740 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_331
timestamp 1604681595
transform 1 0 31556 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_335
timestamp 1604681595
transform 1 0 31924 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_348
timestamp 1604681595
transform 1 0 33120 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_359
timestamp 1604681595
transform 1 0 34132 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_355
timestamp 1604681595
transform 1 0 33764 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_352
timestamp 1604681595
transform 1 0 33488 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 33948 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 33580 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_367
timestamp 1604681595
transform 1 0 34868 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_363
timestamp 1604681595
transform 1 0 34500 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 34592 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1604681595
transform 1 0 34776 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 35052 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 36984 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_388
timestamp 1604681595
transform 1 0 36800 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_392
timestamp 1604681595
transform 1 0 37168 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 38824 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_404
timestamp 1604681595
transform 1 0 38272 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_22
timestamp 1604681595
transform 1 0 3128 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_30
timestamp 1604681595
transform 1 0 3864 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1604681595
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1604681595
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1604681595
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1604681595
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1604681595
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__D
timestamp 1604681595
transform 1 0 13156 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__CLK
timestamp 1604681595
transform 1 0 12696 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_117
timestamp 1604681595
transform 1 0 11868 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_125
timestamp 1604681595
transform 1 0 12604 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_128
timestamp 1604681595
transform 1 0 12880 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_prog_clk
timestamp 1604681595
transform 1 0 13524 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__CLK
timestamp 1604681595
transform 1 0 13984 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_133
timestamp 1604681595
transform 1 0 13340 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1604681595
transform 1 0 13800 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_142
timestamp 1604681595
transform 1 0 14168 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_150
timestamp 1604681595
transform 1 0 14904 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_
timestamp 1604681595
transform 1 0 15916 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 15640 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_154
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_160
timestamp 1604681595
transform 1 0 15824 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604681595
transform 1 0 18400 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1604681595
transform 1 0 17848 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1604681595
transform 1 0 18216 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_180
timestamp 1604681595
transform 1 0 17664 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_184
timestamp 1604681595
transform 1 0 18032 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__CLK
timestamp 1604681595
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_197
timestamp 1604681595
transform 1 0 19228 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_209
timestamp 1604681595
transform 1 0 20332 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_213
timestamp 1604681595
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_
timestamp 1604681595
transform 1 0 21344 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_32_239
timestamp 1604681595
transform 1 0 23092 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1604681595
transform 1 0 23828 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604681595
transform 1 0 24840 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1604681595
transform 1 0 24288 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1604681595
transform 1 0 24656 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 23644 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 23276 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_243
timestamp 1604681595
transform 1 0 23460 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1604681595
transform 1 0 24104 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_254
timestamp 1604681595
transform 1 0 24472 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 27048 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 26220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1604681595
transform 1 0 25852 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_267
timestamp 1604681595
transform 1 0 25668 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_271
timestamp 1604681595
transform 1 0 26036 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_280
timestamp 1604681595
transform 1 0 26864 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 27876 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 27416 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_284
timestamp 1604681595
transform 1 0 27232 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_288
timestamp 1604681595
transform 1 0 27600 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 30360 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 29808 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 30176 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_310
timestamp 1604681595
transform 1 0 29624 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_314
timestamp 1604681595
transform 1 0 29992 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_327
timestamp 1604681595
transform 1 0 31188 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1604681595
transform 1 0 32016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 32292 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 31372 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 33212 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_331
timestamp 1604681595
transform 1 0 31556 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_335
timestamp 1604681595
transform 1 0 31924 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_337
timestamp 1604681595
transform 1 0 32108 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_341
timestamp 1604681595
transform 1 0 32476 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 33580 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 35144 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 34592 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 34960 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_351
timestamp 1604681595
transform 1 0 33396 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_362
timestamp 1604681595
transform 1 0 34408 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_366
timestamp 1604681595
transform 1 0 34776 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 36156 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_379
timestamp 1604681595
transform 1 0 35972 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_383
timestamp 1604681595
transform 1 0 36340 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 38824 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1604681595
transform 1 0 37628 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_395
timestamp 1604681595
transform 1 0 37444 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_398
timestamp 1604681595
transform 1 0 37720 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_406
timestamp 1604681595
transform 1 0 38456 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1604681595
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604681595
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1604681595
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1604681595
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1604681595
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_51
timestamp 1604681595
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1604681595
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1604681595
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_74
timestamp 1604681595
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_86
timestamp 1604681595
transform 1 0 9016 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1604681595
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1604681595
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 9476 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 9936 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_90
timestamp 1604681595
transform 1 0 9384 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_94
timestamp 1604681595
transform 1 0 9752 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_98
timestamp 1604681595
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1604681595
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_117
timestamp 1604681595
transform 1 0 11868 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_119
timestamp 1604681595
transform 1 0 12052 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_115
timestamp 1604681595
transform 1 0 11684 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1604681595
transform 1 0 11224 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 11868 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 11408 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_125
timestamp 1604681595
transform 1 0 12604 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_128
timestamp 1604681595
transform 1 0 12880 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_123
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__D
timestamp 1604681595
transform 1 0 12696 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_
timestamp 1604681595
transform 1 0 13156 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_
timestamp 1604681595
transform 1 0 12696 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 15088 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 14628 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_150
timestamp 1604681595
transform 1 0 14904 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_145
timestamp 1604681595
transform 1 0 14444 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_149
timestamp 1604681595
transform 1 0 14812 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_154
timestamp 1604681595
transform 1 0 15272 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 15456 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604681595
transform 1 0 15640 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_172
timestamp 1604681595
transform 1 0 16928 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_168
timestamp 1604681595
transform 1 0 16560 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_163
timestamp 1604681595
transform 1 0 16100 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_171
timestamp 1604681595
transform 1 0 16836 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_167
timestamp 1604681595
transform 1 0 16468 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 16744 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 16376 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 16652 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 17112 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1604681595
transform 1 0 17020 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_176
timestamp 1604681595
transform 1 0 17296 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_179
timestamp 1604681595
transform 1 0 17572 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_175
timestamp 1604681595
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__CLK
timestamp 1604681595
transform 1 0 17480 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1604681595
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__D
timestamp 1604681595
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604681595
transform 1 0 17664 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_34_193
timestamp 1604681595
transform 1 0 18860 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_189
timestamp 1604681595
transform 1 0 18492 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 18676 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_33_207
timestamp 1604681595
transform 1 0 20148 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_203
timestamp 1604681595
transform 1 0 19780 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
timestamp 1604681595
transform 1 0 19964 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604681595
transform 1 0 19228 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_215
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_213
timestamp 1604681595
transform 1 0 20700 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_216
timestamp 1604681595
transform 1 0 20976 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_213
timestamp 1604681595
transform 1 0 20700 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__CLK
timestamp 1604681595
transform 1 0 21068 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1604681595
transform 1 0 20792 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__D
timestamp 1604681595
transform 1 0 21160 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_201
timestamp 1604681595
transform 1 0 19596 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_219
timestamp 1604681595
transform 1 0 21252 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_220
timestamp 1604681595
transform 1 0 21344 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1604681595
transform 1 0 21528 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1604681595
transform 1 0 21528 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604681595
transform 1 0 21712 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_33_240
timestamp 1604681595
transform 1 0 23184 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_237
timestamp 1604681595
transform 1 0 22908 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_233
timestamp 1604681595
transform 1 0 22540 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 23000 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_
timestamp 1604681595
transform 1 0 21712 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604681595
transform 1 0 24472 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1604681595
transform 1 0 24196 0 -1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__D
timestamp 1604681595
transform 1 0 23920 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1604681595
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_243
timestamp 1604681595
transform 1 0 23460 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_247
timestamp 1604681595
transform 1 0 23828 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_250
timestamp 1604681595
transform 1 0 24104 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_271
timestamp 1604681595
transform 1 0 26036 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_269
timestamp 1604681595
transform 1 0 25852 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_263
timestamp 1604681595
transform 1 0 25300 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 26036 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 25484 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_273
timestamp 1604681595
transform 1 0 26220 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 26220 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 26496 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 26680 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_34_289
timestamp 1604681595
transform 1 0 27692 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_285
timestamp 1604681595
transform 1 0 27324 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 27508 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_297
timestamp 1604681595
transform 1 0 28428 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_301
timestamp 1604681595
transform 1 0 28796 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_297
timestamp 1604681595
transform 1 0 28428 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 28612 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 28060 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_305
timestamp 1604681595
transform 1 0 29164 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 28980 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1604681595
transform 1 0 29164 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_316
timestamp 1604681595
transform 1 0 30176 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_312
timestamp 1604681595
transform 1 0 29808 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_306
timestamp 1604681595
transform 1 0 29256 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 29256 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 29992 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 29440 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1604681595
transform 1 0 29532 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_317
timestamp 1604681595
transform 1 0 30268 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 30544 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 30360 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_322
timestamp 1604681595
transform 1 0 30728 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 30544 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 33212 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1604681595
transform 1 0 32016 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 33028 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 33212 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_339
timestamp 1604681595
transform 1 0 32292 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_334
timestamp 1604681595
transform 1 0 31832 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_337
timestamp 1604681595
transform 1 0 32108 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_351
timestamp 1604681595
transform 1 0 33396 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_358
timestamp 1604681595
transform 1 0 34040 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 33764 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 34224 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_367
timestamp 1604681595
transform 1 0 34868 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_362
timestamp 1604681595
transform 1 0 34408 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 34592 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1604681595
transform 1 0 34776 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 34960 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 33948 0 -1 21216
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _48_
timestamp 1604681595
transform 1 0 36616 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 36064 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_387
timestamp 1604681595
transform 1 0 36708 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_378
timestamp 1604681595
transform 1 0 35880 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_382
timestamp 1604681595
transform 1 0 36248 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_389
timestamp 1604681595
transform 1 0 36892 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 38824 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 38824 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1604681595
transform 1 0 37628 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_399
timestamp 1604681595
transform 1 0 37812 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_398
timestamp 1604681595
transform 1 0 37720 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_406
timestamp 1604681595
transform 1 0 38456 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604681595
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1604681595
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1604681595
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1604681595
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_51
timestamp 1604681595
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_59
timestamp 1604681595
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_62
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1604681595
transform 1 0 8556 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 9016 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_74
timestamp 1604681595
transform 1 0 7912 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_80
timestamp 1604681595
transform 1 0 8464 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_84
timestamp 1604681595
transform 1 0 8832 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_88
timestamp 1604681595
transform 1 0 9200 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_100
timestamp 1604681595
transform 1 0 10304 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1604681595
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__D
timestamp 1604681595
transform 1 0 13064 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 12696 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_112
timestamp 1604681595
transform 1 0 11408 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_123
timestamp 1604681595
transform 1 0 12420 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_128
timestamp 1604681595
transform 1 0 12880 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_
timestamp 1604681595
transform 1 0 13248 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_35_151
timestamp 1604681595
transform 1 0 14996 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604681595
transform 1 0 16376 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 15180 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 15548 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 15916 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_155
timestamp 1604681595
transform 1 0 15364 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_159
timestamp 1604681595
transform 1 0 15732 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_163
timestamp 1604681595
transform 1 0 16100 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_
timestamp 1604681595
transform 1 0 18584 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1604681595
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__D
timestamp 1604681595
transform 1 0 18400 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
timestamp 1604681595
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__CLK
timestamp 1604681595
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_175
timestamp 1604681595
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_179
timestamp 1604681595
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_184
timestamp 1604681595
transform 1 0 18032 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_
timestamp 1604681595
transform 1 0 21068 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__D
timestamp 1604681595
transform 1 0 20884 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_209
timestamp 1604681595
transform 1 0 20332 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1604681595
transform 1 0 23000 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_236
timestamp 1604681595
transform 1 0 22816 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_240
timestamp 1604681595
transform 1 0 23184 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_
timestamp 1604681595
transform 1 0 23644 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1604681595
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__D
timestamp 1604681595
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 26128 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 26680 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 25944 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__CLK
timestamp 1604681595
transform 1 0 25576 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 27048 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_264
timestamp 1604681595
transform 1 0 25392 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_268
timestamp 1604681595
transform 1 0 25760 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_276
timestamp 1604681595
transform 1 0 26496 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_280
timestamp 1604681595
transform 1 0 26864 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 27232 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1604681595
transform 1 0 29164 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 27784 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_288
timestamp 1604681595
transform 1 0 27600 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_292
timestamp 1604681595
transform 1 0 27968 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_304
timestamp 1604681595
transform 1 0 29072 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 29716 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 29532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_306
timestamp 1604681595
transform 1 0 29256 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_330
timestamp 1604681595
transform 1 0 31464 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_342
timestamp 1604681595
transform 1 0 32568 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 34868 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1604681595
transform 1 0 34776 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 34592 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 34224 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 33856 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_354
timestamp 1604681595
transform 1 0 33672 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_358
timestamp 1604681595
transform 1 0 34040 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_362
timestamp 1604681595
transform 1 0 34408 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_386
timestamp 1604681595
transform 1 0 36616 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 38824 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_398
timestamp 1604681595
transform 1 0 37720 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_406
timestamp 1604681595
transform 1 0 38456 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1604681595
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1604681595
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1604681595
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1604681595
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1604681595
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1604681595
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_56
timestamp 1604681595
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_68
timestamp 1604681595
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_80
timestamp 1604681595
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1604681595
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_93
timestamp 1604681595
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_105
timestamp 1604681595
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_prog_clk
timestamp 1604681595
transform 1 0 12972 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__CLK
timestamp 1604681595
transform 1 0 12788 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_117
timestamp 1604681595
transform 1 0 11868 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_125
timestamp 1604681595
transform 1 0 12604 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604681595
transform 1 0 13616 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
timestamp 1604681595
transform 1 0 14996 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 13432 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_132
timestamp 1604681595
transform 1 0 13248 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_145
timestamp 1604681595
transform 1 0 14444 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_149
timestamp 1604681595
transform 1 0 14812 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604681595
transform 1 0 16836 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1604681595
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 16376 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_163
timestamp 1604681595
transform 1 0 16100 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_168
timestamp 1604681595
transform 1 0 16560 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 18584 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 17388 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 18032 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 19136 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_175
timestamp 1604681595
transform 1 0 17204 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_179
timestamp 1604681595
transform 1 0 17572 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_183
timestamp 1604681595
transform 1 0 17940 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_186
timestamp 1604681595
transform 1 0 18216 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1604681595
transform 1 0 18952 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1604681595
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 19504 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 19872 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_198
timestamp 1604681595
transform 1 0 19320 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_202
timestamp 1604681595
transform 1 0 19688 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_206
timestamp 1604681595
transform 1 0 20056 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_215
timestamp 1604681595
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604681595
transform 1 0 22356 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1604681595
transform 1 0 22172 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_227
timestamp 1604681595
transform 1 0 21988 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_240
timestamp 1604681595
transform 1 0 23184 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_
timestamp 1604681595
transform 1 0 23920 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__CLK
timestamp 1604681595
transform 1 0 23644 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_244
timestamp 1604681595
transform 1 0 23552 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_247
timestamp 1604681595
transform 1 0 23828 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 26496 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1604681595
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_267
timestamp 1604681595
transform 1 0 25668 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_295
timestamp 1604681595
transform 1 0 28244 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 29532 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 29900 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_307
timestamp 1604681595
transform 1 0 29348 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_311
timestamp 1604681595
transform 1 0 29716 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_315
timestamp 1604681595
transform 1 0 30084 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_327
timestamp 1604681595
transform 1 0 31188 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1604681595
transform 1 0 32016 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_335
timestamp 1604681595
transform 1 0 31924 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_337
timestamp 1604681595
transform 1 0 32108 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_349
timestamp 1604681595
transform 1 0 33212 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 34592 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 33672 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 34408 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 34040 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_353
timestamp 1604681595
transform 1 0 33580 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_356
timestamp 1604681595
transform 1 0 33856 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_360
timestamp 1604681595
transform 1 0 34224 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_383
timestamp 1604681595
transform 1 0 36340 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 38824 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1604681595
transform 1 0 37628 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_395
timestamp 1604681595
transform 1 0 37444 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_398
timestamp 1604681595
transform 1 0 37720 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_406
timestamp 1604681595
transform 1 0 38456 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1604681595
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1604681595
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1604681595
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1604681595
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1604681595
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_51
timestamp 1604681595
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_59
timestamp 1604681595
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_62
timestamp 1604681595
transform 1 0 6808 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_prog_clk
timestamp 1604681595
transform 1 0 7544 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_73
timestamp 1604681595
transform 1 0 7820 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_77
timestamp 1604681595
transform 1 0 8188 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 10396 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_89
timestamp 1604681595
transform 1 0 9292 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_103
timestamp 1604681595
transform 1 0 10580 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1604681595
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 12880 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_115
timestamp 1604681595
transform 1 0 11684 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_121
timestamp 1604681595
transform 1 0 12236 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_123
timestamp 1604681595
transform 1 0 12420 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_127
timestamp 1604681595
transform 1 0 12788 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_130
timestamp 1604681595
transform 1 0 13064 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_
timestamp 1604681595
transform 1 0 13800 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__D
timestamp 1604681595
transform 1 0 13616 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 13248 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_134
timestamp 1604681595
transform 1 0 13432 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604681595
transform 1 0 16376 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 16192 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 15824 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_157
timestamp 1604681595
transform 1 0 15548 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_162
timestamp 1604681595
transform 1 0 16008 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_179
timestamp 1604681595
transform 1 0 17572 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_175
timestamp 1604681595
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1604681595
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 18032 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_192
timestamp 1604681595
transform 1 0 18768 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_188
timestamp 1604681595
transform 1 0 18400 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 18584 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 18952 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 19136 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_37_215
timestamp 1604681595
transform 1 0 20884 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1604681595
transform 1 0 22356 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_227
timestamp 1604681595
transform 1 0 21988 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_233
timestamp 1604681595
transform 1 0 22540 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_
timestamp 1604681595
transform 1 0 25116 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1604681595
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__D
timestamp 1604681595
transform 1 0 24932 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_241
timestamp 1604681595
transform 1 0 23276 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_245
timestamp 1604681595
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_257
timestamp 1604681595
transform 1 0 24748 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1604681595
transform 1 0 27048 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_280
timestamp 1604681595
transform 1 0 26864 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1604681595
transform 1 0 29164 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
timestamp 1604681595
transform 1 0 27416 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 28980 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 28612 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_284
timestamp 1604681595
transform 1 0 27232 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_288
timestamp 1604681595
transform 1 0 27600 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_296
timestamp 1604681595
transform 1 0 28336 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_301
timestamp 1604681595
transform 1 0 28796 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 29624 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 29440 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_306
timestamp 1604681595
transform 1 0 29256 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_prog_clk
timestamp 1604681595
transform 1 0 32108 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 32568 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_prog_clk_A
timestamp 1604681595
transform 1 0 32936 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_329
timestamp 1604681595
transform 1 0 31372 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_340
timestamp 1604681595
transform 1 0 32384 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_344
timestamp 1604681595
transform 1 0 32752 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_348
timestamp 1604681595
transform 1 0 33120 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_358
timestamp 1604681595
transform 1 0 34040 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_353
timestamp 1604681595
transform 1 0 33580 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 33396 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 33672 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_367
timestamp 1604681595
transform 1 0 34868 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_365
timestamp 1604681595
transform 1 0 34684 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_362
timestamp 1604681595
transform 1 0 34408 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 34500 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1604681595
transform 1 0 34776 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 35052 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 36064 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 36432 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 36800 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_378
timestamp 1604681595
transform 1 0 35880 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_382
timestamp 1604681595
transform 1 0 36248 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_386
timestamp 1604681595
transform 1 0 36616 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_390
timestamp 1604681595
transform 1 0 36984 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 38824 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_402
timestamp 1604681595
transform 1 0 38088 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_406
timestamp 1604681595
transform 1 0 38456 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1604681595
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1604681595
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1604681595
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1604681595
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1604681595
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__CLK
timestamp 1604681595
transform 1 0 7084 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_44
timestamp 1604681595
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_56
timestamp 1604681595
transform 1 0 6256 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_64
timestamp 1604681595
transform 1 0 6992 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__CLK
timestamp 1604681595
transform 1 0 7636 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_67
timestamp 1604681595
transform 1 0 7268 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_73
timestamp 1604681595
transform 1 0 7820 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_85
timestamp 1604681595
transform 1 0 8924 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_97
timestamp 1604681595
transform 1 0 10028 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_93
timestamp 1604681595
transform 1 0 9660 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_91
timestamp 1604681595
transform 1 0 9476 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 10120 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1604681595
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_104
timestamp 1604681595
transform 1 0 10672 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_100
timestamp 1604681595
transform 1 0 10304 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 10856 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_prog_clk
timestamp 1604681595
transform 1 0 10396 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_108
timestamp 1604681595
transform 1 0 11040 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_120
timestamp 1604681595
transform 1 0 12144 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604681595
transform 1 0 13616 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 13432 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_132
timestamp 1604681595
transform 1 0 13248 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_145
timestamp 1604681595
transform 1 0 14444 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16376 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604681595
transform 1 0 15272 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1604681595
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 15824 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 16192 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_158
timestamp 1604681595
transform 1 0 15640 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_162
timestamp 1604681595
transform 1 0 16008 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 18032 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 19044 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 18584 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_175
timestamp 1604681595
transform 1 0 17204 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_183
timestamp 1604681595
transform 1 0 17940 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_188
timestamp 1604681595
transform 1 0 18400 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_192
timestamp 1604681595
transform 1 0 18768 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1604681595
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 21068 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_215
timestamp 1604681595
transform 1 0 20884 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1__f_clk_A
timestamp 1604681595
transform 1 0 21436 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_219
timestamp 1604681595
transform 1 0 21252 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_223
timestamp 1604681595
transform 1 0 21620 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_235
timestamp 1604681595
transform 1 0 22724 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__CLK
timestamp 1604681595
transform 1 0 25116 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_247
timestamp 1604681595
transform 1 0 23828 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_259
timestamp 1604681595
transform 1 0 24932 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  ltile_clb_0.ltile_clb_m_default__fle_6.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604681595
transform 1 0 26496 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1604681595
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_263
timestamp 1604681595
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_281
timestamp 1604681595
transform 1 0 26956 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_293
timestamp 1604681595
transform 1 0 28060 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_305
timestamp 1604681595
transform 1 0 29164 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 29532 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 29348 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 32108 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1604681595
transform 1 0 32016 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_328
timestamp 1604681595
transform 1 0 31280 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_341
timestamp 1604681595
transform 1 0 32476 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_349
timestamp 1604681595
transform 1 0 33212 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 33396 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 34500 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 34316 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 33948 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_355
timestamp 1604681595
transform 1 0 33764 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_359
timestamp 1604681595
transform 1 0 34132 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1604681595
transform 1 0 36064 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 35512 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 35880 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 36524 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_372
timestamp 1604681595
transform 1 0 35328 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_376
timestamp 1604681595
transform 1 0 35696 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_383
timestamp 1604681595
transform 1 0 36340 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_387
timestamp 1604681595
transform 1 0 36708 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 38824 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1604681595
transform 1 0 37628 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_395
timestamp 1604681595
transform 1 0 37444 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_398
timestamp 1604681595
transform 1 0 37720 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_406
timestamp 1604681595
transform 1 0 38456 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1604681595
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1604681595
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1604681595
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1604681595
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1604681595
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1604681595
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1604681595
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1604681595
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1604681595
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_51
timestamp 1604681595
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_63
timestamp 1604681595
transform 1 0 6900 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_60
timestamp 1604681595
transform 1 0 6624 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_56
timestamp 1604681595
transform 1 0 6256 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_62
timestamp 1604681595
transform 1 0 6808 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_59
timestamp 1604681595
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__D
timestamp 1604681595
transform 1 0 6716 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__D
timestamp 1604681595
transform 1 0 7084 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1604681595
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_44
timestamp 1604681595
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_
timestamp 1604681595
transform 1 0 7084 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_
timestamp 1604681595
transform 1 0 7636 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__D
timestamp 1604681595
transform 1 0 7452 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_67
timestamp 1604681595
transform 1 0 7268 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_84
timestamp 1604681595
transform 1 0 8832 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_93
timestamp 1604681595
transform 1 0 9660 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_96
timestamp 1604681595
transform 1 0 9936 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_90
timestamp 1604681595
transform 1 0 9384 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__D
timestamp 1604681595
transform 1 0 9752 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1604681595
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604681595
transform 1 0 10120 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_39_107
timestamp 1604681595
transform 1 0 10948 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 11132 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_
timestamp 1604681595
transform 1 0 9752 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_40_117
timestamp 1604681595
transform 1 0 11868 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_113
timestamp 1604681595
transform 1 0 11500 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_115
timestamp 1604681595
transform 1 0 11684 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_111
timestamp 1604681595
transform 1 0 11316 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 11684 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__CLK
timestamp 1604681595
transform 1 0 11500 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_121
timestamp 1604681595
transform 1 0 12236 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 12420 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1604681595
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_125
timestamp 1604681595
transform 1 0 12604 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_123
timestamp 1604681595
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_
timestamp 1604681595
transform 1 0 14536 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__D
timestamp 1604681595
transform 1 0 14352 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__CLK
timestamp 1604681595
transform 1 0 14536 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_135
timestamp 1604681595
transform 1 0 13524 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_143
timestamp 1604681595
transform 1 0 14260 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_137
timestamp 1604681595
transform 1 0 13708 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_145
timestamp 1604681595
transform 1 0 14444 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_148
timestamp 1604681595
transform 1 0 14720 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15456 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 17020 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1604681595
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 16468 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 17020 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_165
timestamp 1604681595
transform 1 0 16284 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_169
timestamp 1604681595
transform 1 0 16652 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_154
timestamp 1604681595
transform 1 0 15272 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_165
timestamp 1604681595
transform 1 0 16284 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_177
timestamp 1604681595
transform 1 0 17388 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_39_184
timestamp 1604681595
transform 1 0 18032 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_175
timestamp 1604681595
transform 1 0 17204 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 17940 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1604681595
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_189
timestamp 1604681595
transform 1 0 18492 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_185
timestamp 1604681595
transform 1 0 18124 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_192
timestamp 1604681595
transform 1 0 18768 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
timestamp 1604681595
transform 1 0 18308 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1604681595
transform 1 0 18952 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604681595
transform 1 0 18308 0 1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604681595
transform 1 0 18584 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19136 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_207
timestamp 1604681595
transform 1 0 20148 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_203
timestamp 1604681595
transform 1 0 19780 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_199
timestamp 1604681595
transform 1 0 19412 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_205
timestamp 1604681595
transform 1 0 19964 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19964 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19596 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_211
timestamp 1604681595
transform 1 0 20516 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_210
timestamp 1604681595
transform 1 0 20424 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20332 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20240 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1604681595
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1604681595
transform 1 0 20792 0 1 23392
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 21896 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_234
timestamp 1604681595
transform 1 0 22632 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_224
timestamp 1604681595
transform 1 0 21712 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_228
timestamp 1604681595
transform 1 0 22080 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_240
timestamp 1604681595
transform 1 0 23184 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1604681595
transform 1 0 24656 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1604681595
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 25116 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_242
timestamp 1604681595
transform 1 0 23368 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_245
timestamp 1604681595
transform 1 0 23644 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_257
timestamp 1604681595
transform 1 0 24748 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_252
timestamp 1604681595
transform 1 0 24288 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_259
timestamp 1604681595
transform 1 0 24932 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_271
timestamp 1604681595
transform 1 0 26036 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_267
timestamp 1604681595
transform 1 0 25668 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_263
timestamp 1604681595
transform 1 0 25300 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 25484 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_prog_clk_A
timestamp 1604681595
transform 1 0 26128 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_274
timestamp 1604681595
transform 1 0 26312 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1604681595
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_276
timestamp 1604681595
transform 1 0 26496 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1604681595
transform 1 0 26956 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_269
timestamp 1604681595
transform 1 0 25852 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1604681595
transform 1 0 29164 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 28980 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 28612 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_293
timestamp 1604681595
transform 1 0 28060 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_301
timestamp 1604681595
transform 1 0 28796 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_288
timestamp 1604681595
transform 1 0 27600 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_300
timestamp 1604681595
transform 1 0 28704 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 29716 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 29532 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 29532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__CLK
timestamp 1604681595
transform 1 0 29348 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_306
timestamp 1604681595
transform 1 0 29256 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_40_306
timestamp 1604681595
transform 1 0 29256 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
timestamp 1604681595
transform 1 0 31648 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 31464 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_330
timestamp 1604681595
transform 1 0 31464 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_328
timestamp 1604681595
transform 1 0 31280 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_332
timestamp 1604681595
transform 1 0 31648 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1604681595
transform 1 0 32016 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 32016 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 31832 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1604681595
transform 1 0 31832 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604681595
transform 1 0 32108 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_346
timestamp 1604681595
transform 1 0 32936 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_346
timestamp 1604681595
transform 1 0 32936 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_342
timestamp 1604681595
transform 1 0 32568 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 32752 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604681595
transform 1 0 32200 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 33120 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 33120 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_360
timestamp 1604681595
transform 1 0 34224 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_356
timestamp 1604681595
transform 1 0 33856 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_350
timestamp 1604681595
transform 1 0 33304 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_358
timestamp 1604681595
transform 1 0 34040 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_350
timestamp 1604681595
transform 1 0 33304 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 34040 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 33488 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
timestamp 1604681595
transform 1 0 33672 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 33672 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_365
timestamp 1604681595
transform 1 0 34684 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_362
timestamp 1604681595
transform 1 0 34408 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 34500 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1604681595
transform 1 0 34776 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 34500 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 34868 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 36064 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 36800 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 35512 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 35880 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_386
timestamp 1604681595
transform 1 0 36616 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_390
timestamp 1604681595
transform 1 0 36984 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_372
timestamp 1604681595
transform 1 0 35328 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_376
timestamp 1604681595
transform 1 0 35696 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_384
timestamp 1604681595
transform 1 0 36432 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 38824 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 38824 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1604681595
transform 1 0 37628 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_402
timestamp 1604681595
transform 1 0 38088 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_406
timestamp 1604681595
transform 1 0 38456 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_396
timestamp 1604681595
transform 1 0 37536 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_398
timestamp 1604681595
transform 1 0 37720 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_406
timestamp 1604681595
transform 1 0 38456 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1604681595
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1604681595
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1604681595
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1604681595
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_
timestamp 1604681595
transform 1 0 6900 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1604681595
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__D
timestamp 1604681595
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__CLK
timestamp 1604681595
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__CLK
timestamp 1604681595
transform 1 0 5796 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_53
timestamp 1604681595
transform 1 0 5980 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1604681595
transform 1 0 6348 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_62
timestamp 1604681595
transform 1 0 6808 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 8924 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_82
timestamp 1604681595
transform 1 0 8648 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_87
timestamp 1604681595
transform 1 0 9108 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_
timestamp 1604681595
transform 1 0 9844 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 9660 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 9292 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_91
timestamp 1604681595
transform 1 0 9476 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 12420 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1604681595
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_114
timestamp 1604681595
transform 1 0 11592 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_118
timestamp 1604681595
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 15088 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 14720 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 14352 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_142
timestamp 1604681595
transform 1 0 14168 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_146
timestamp 1604681595
transform 1 0 14536 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_150
timestamp 1604681595
transform 1 0 14904 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 15272 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_41_173
timestamp 1604681595
transform 1 0 17020 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_177
timestamp 1604681595
transform 1 0 17388 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 17204 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_184
timestamp 1604681595
transform 1 0 18032 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1604681595
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_188
timestamp 1604681595
transform 1 0 18400 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18216 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_192
timestamp 1604681595
transform 1 0 18768 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 18584 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 18952 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 20056 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 19872 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 19504 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_198
timestamp 1604681595
transform 1 0 19320 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_202
timestamp 1604681595
transform 1 0 19688 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 21988 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 22356 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1604681595
transform 1 0 21804 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_229
timestamp 1604681595
transform 1 0 22172 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_233
timestamp 1604681595
transform 1 0 22540 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_249
timestamp 1604681595
transform 1 0 24012 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_245
timestamp 1604681595
transform 1 0 23644 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_241
timestamp 1604681595
transform 1 0 23276 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23828 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 24196 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1604681595
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_257
timestamp 1604681595
transform 1 0 24748 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_253
timestamp 1604681595
transform 1 0 24380 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 24564 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 25024 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_41_279
timestamp 1604681595
transform 1 0 26772 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_283
timestamp 1604681595
transform 1 0 27140 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1604681595
transform 1 0 29164 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 28980 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 27232 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_286
timestamp 1604681595
transform 1 0 27416 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_298
timestamp 1604681595
transform 1 0 28520 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_302
timestamp 1604681595
transform 1 0 28888 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_
timestamp 1604681595
transform 1 0 29624 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__D
timestamp 1604681595
transform 1 0 29440 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_306
timestamp 1604681595
transform 1 0 29256 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604681595
transform 1 0 32108 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 31924 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 31556 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 33120 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_329
timestamp 1604681595
transform 1 0 31372 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_333
timestamp 1604681595
transform 1 0 31740 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_346
timestamp 1604681595
transform 1 0 32936 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_358
timestamp 1604681595
transform 1 0 34040 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_350
timestamp 1604681595
transform 1 0 33304 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 33488 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 34224 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604681595
transform 1 0 33672 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_367
timestamp 1604681595
transform 1 0 34868 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_362
timestamp 1604681595
transform 1 0 34408 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 34592 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1604681595
transform 1 0 34776 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 35052 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 36984 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_388
timestamp 1604681595
transform 1 0 36800 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_392
timestamp 1604681595
transform 1 0 37168 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 38824 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_404
timestamp 1604681595
transform 1 0 38272 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 1564 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1604681595
transform 1 0 1380 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_7
timestamp 1604681595
transform 1 0 1748 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_19
timestamp 1604681595
transform 1 0 2852 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1604681595
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1604681595
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_
timestamp 1604681595
transform 1 0 6716 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 6440 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1604681595
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_56
timestamp 1604681595
transform 1 0 6256 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_60
timestamp 1604681595
transform 1 0 6624 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 8648 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_80
timestamp 1604681595
transform 1 0 8464 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_84
timestamp 1604681595
transform 1 0 8832 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10028 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1604681595
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__D
timestamp 1604681595
transform 1 0 9844 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 9292 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_88
timestamp 1604681595
transform 1 0 9200 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_91
timestamp 1604681595
transform 1 0 9476 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_93
timestamp 1604681595
transform 1 0 9660 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_106
timestamp 1604681595
transform 1 0 10856 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 11592 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1604681595
transform 1 0 14536 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13524 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_133
timestamp 1604681595
transform 1 0 13340 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_137
timestamp 1604681595
transform 1 0 13708 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_145
timestamp 1604681595
transform 1 0 14444 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_149
timestamp 1604681595
transform 1 0 14812 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 15456 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1604681595
transform 1 0 15180 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_154
timestamp 1604681595
transform 1 0 15272 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604681595
transform 1 0 17940 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_42_175
timestamp 1604681595
transform 1 0 17204 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1604681595
transform 1 0 18768 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_196
timestamp 1604681595
transform 1 0 19136 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _59_
timestamp 1604681595
transform 1 0 19596 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 20884 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1604681595
transform 1 0 20792 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19228 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 20608 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20056 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_199
timestamp 1604681595
transform 1 0 19412 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_204
timestamp 1604681595
transform 1 0 19872 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_208
timestamp 1604681595
transform 1 0 20240 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_234
timestamp 1604681595
transform 1 0 22632 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 24564 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 24380 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 24012 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_246
timestamp 1604681595
transform 1 0 23736 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_251
timestamp 1604681595
transform 1 0 24196 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1604681595
transform 1 0 26404 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_prog_clk
timestamp 1604681595
transform 1 0 26128 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 27048 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 26680 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_264
timestamp 1604681595
transform 1 0 25392 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_276
timestamp 1604681595
transform 1 0 26496 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_280
timestamp 1604681595
transform 1 0 26864 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 27232 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 27692 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 28888 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_287
timestamp 1604681595
transform 1 0 27508 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_291
timestamp 1604681595
transform 1 0 27876 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_299
timestamp 1604681595
transform 1 0 28612 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_304
timestamp 1604681595
transform 1 0 29072 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604681595
transform 1 0 30176 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 29992 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 29624 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 31188 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__CLK
timestamp 1604681595
transform 1 0 29256 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_308
timestamp 1604681595
transform 1 0 29440 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_312
timestamp 1604681595
transform 1 0 29808 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_325
timestamp 1604681595
transform 1 0 31004 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604681595
transform 1 0 32108 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1604681595
transform 1 0 32016 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 31740 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 33120 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 31556 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_329
timestamp 1604681595
transform 1 0 31372 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_346
timestamp 1604681595
transform 1 0 32936 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604681595
transform 1 0 33764 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__D
timestamp 1604681595
transform 1 0 35144 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 33488 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 34776 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_350
timestamp 1604681595
transform 1 0 33304 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_354
timestamp 1604681595
transform 1 0 33672 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_364
timestamp 1604681595
transform 1 0 34592 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_368
timestamp 1604681595
transform 1 0 34960 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604681595
transform 1 0 35328 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_42_381
timestamp 1604681595
transform 1 0 36156 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_393
timestamp 1604681595
transform 1 0 37260 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 38824 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1604681595
transform 1 0 37628 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_398
timestamp 1604681595
transform 1 0 37720 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_406
timestamp 1604681595
transform 1 0 38456 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1604681595
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 1564 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 2116 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 2484 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1604681595
transform 1 0 1380 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_7
timestamp 1604681595
transform 1 0 1748 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_13
timestamp 1604681595
transform 1 0 2300 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_17
timestamp 1604681595
transform 1 0 2668 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_29
timestamp 1604681595
transform 1 0 3772 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_41
timestamp 1604681595
transform 1 0 4876 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_
timestamp 1604681595
transform 1 0 6808 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1604681595
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 6440 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__D
timestamp 1604681595
transform 1 0 6072 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 5704 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_49
timestamp 1604681595
transform 1 0 5612 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_52
timestamp 1604681595
transform 1 0 5888 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_56
timestamp 1604681595
transform 1 0 6256 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_60
timestamp 1604681595
transform 1 0 6624 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 8740 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 9108 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_81
timestamp 1604681595
transform 1 0 8556 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_85
timestamp 1604681595
transform 1 0 8924 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9292 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10304 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10856 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_98
timestamp 1604681595
transform 1 0 10120 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_102
timestamp 1604681595
transform 1 0 10488 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_108
timestamp 1604681595
transform 1 0 11040 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1604681595
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 12144 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11224 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11592 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_112
timestamp 1604681595
transform 1 0 11408 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_116
timestamp 1604681595
transform 1 0 11776 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14352 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15088 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14720 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_142
timestamp 1604681595
transform 1 0 14168 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_146
timestamp 1604681595
transform 1 0 14536 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_150
timestamp 1604681595
transform 1 0 14904 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15640 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 15456 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16652 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 17020 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_154
timestamp 1604681595
transform 1 0 15272 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_167
timestamp 1604681595
transform 1 0 16468 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_171
timestamp 1604681595
transform 1 0 16836 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1604681595
transform 1 0 17940 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 18216 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 19044 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18676 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_175
timestamp 1604681595
transform 1 0 17204 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_184
timestamp 1604681595
transform 1 0 18032 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_188
timestamp 1604681595
transform 1 0 18400 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_193
timestamp 1604681595
transform 1 0 18860 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 20792 0 1 25568
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19228 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 20608 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 20240 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_206
timestamp 1604681595
transform 1 0 20056 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_210
timestamp 1604681595
transform 1 0 20424 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 22908 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_235
timestamp 1604681595
transform 1 0 22724 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_239
timestamp 1604681595
transform 1 0 23092 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 24380 0 1 25568
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1604681595
transform 1 0 23552 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 24196 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23828 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 23368 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_245
timestamp 1604681595
transform 1 0 23644 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_249
timestamp 1604681595
transform 1 0 24012 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 27048 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 26496 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 26864 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_274
timestamp 1604681595
transform 1 0 26312 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_278
timestamp 1604681595
transform 1 0 26680 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1604681595
transform 1 0 29164 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 28888 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 28060 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
timestamp 1604681595
transform 1 0 28704 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_291
timestamp 1604681595
transform 1 0 27876 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_295
timestamp 1604681595
transform 1 0 28244 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_299
timestamp 1604681595
transform 1 0 28612 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_
timestamp 1604681595
transform 1 0 29716 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__D
timestamp 1604681595
transform 1 0 29532 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_306
timestamp 1604681595
transform 1 0 29256 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604681595
transform 1 0 33028 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_prog_clk
timestamp 1604681595
transform 1 0 32200 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 31648 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 32016 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 32844 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_330
timestamp 1604681595
transform 1 0 31464 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_334
timestamp 1604681595
transform 1 0 31832 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_341
timestamp 1604681595
transform 1 0 32476 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1604681595
transform 1 0 34776 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 34040 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
timestamp 1604681595
transform 1 0 35236 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__CLK
timestamp 1604681595
transform 1 0 34592 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_356
timestamp 1604681595
transform 1 0 33856 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_360
timestamp 1604681595
transform 1 0 34224 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_367
timestamp 1604681595
transform 1 0 34868 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 36616 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604681595
transform 1 0 35420 0 1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1604681595
transform 1 0 36064 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 37168 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_378
timestamp 1604681595
transform 1 0 35880 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_382
timestamp 1604681595
transform 1 0 36248 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_390
timestamp 1604681595
transform 1 0 36984 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1604681595
transform -1 0 38824 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_394
timestamp 1604681595
transform 1 0 37352 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_406
timestamp 1604681595
transform 1 0 38456 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 1472 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1604681595
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_3
timestamp 1604681595
transform 1 0 1380 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1604681595
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__D
timestamp 1604681595
transform 1 0 4232 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 4600 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_23
timestamp 1604681595
transform 1 0 3220 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_32
timestamp 1604681595
transform 1 0 4048 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_36
timestamp 1604681595
transform 1 0 4416 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_40
timestamp 1604681595
transform 1 0 4784 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604681595
transform 1 0 6440 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_44_52
timestamp 1604681595
transform 1 0 5888 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604681595
transform 1 0 8004 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__CLK
timestamp 1604681595
transform 1 0 7452 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_67
timestamp 1604681595
transform 1 0 7268 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_71
timestamp 1604681595
transform 1 0 7636 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_84
timestamp 1604681595
transform 1 0 8832 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1604681595
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 9292 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_88
timestamp 1604681595
transform 1 0 9200 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_91
timestamp 1604681595
transform 1 0 9476 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_93
timestamp 1604681595
transform 1 0 9660 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_105
timestamp 1604681595
transform 1 0 10764 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_109
timestamp 1604681595
transform 1 0 11132 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12788 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11224 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12604 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 12236 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_119
timestamp 1604681595
transform 1 0 12052 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_123
timestamp 1604681595
transform 1 0 12420 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_136
timestamp 1604681595
transform 1 0 13616 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_148
timestamp 1604681595
transform 1 0 14720 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_152
timestamp 1604681595
transform 1 0 15088 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15548 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1604681595
transform 1 0 15180 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_154
timestamp 1604681595
transform 1 0 15272 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 18032 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19044 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_176
timestamp 1604681595
transform 1 0 17296 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_188
timestamp 1604681595
transform 1 0 18400 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_194
timestamp 1604681595
transform 1 0 18952 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 20884 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1604681595
transform 1 0 20792 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 20608 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 20240 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_206
timestamp 1604681595
transform 1 0 20056 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_210
timestamp 1604681595
transform 1 0 20424 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_234
timestamp 1604681595
transform 1 0 22632 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24656 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 24380 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24012 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_246
timestamp 1604681595
transform 1 0 23736 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_251
timestamp 1604681595
transform 1 0 24196 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_255
timestamp 1604681595
transform 1 0 24564 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 26496 0 -1 26656
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1604681595
transform 1 0 26404 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 25668 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 26220 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_265
timestamp 1604681595
transform 1 0 25484 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_269
timestamp 1604681595
transform 1 0 25852 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604681595
transform 1 0 29164 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_297
timestamp 1604681595
transform 1 0 28428 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604681595
transform 1 0 30268 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 30084 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__CLK
timestamp 1604681595
transform 1 0 29716 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_309
timestamp 1604681595
transform 1 0 29532 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_313
timestamp 1604681595
transform 1 0 29900 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_326
timestamp 1604681595
transform 1 0 31096 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604681595
transform 1 0 32108 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1604681595
transform 1 0 32016 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 31832 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1604681595
transform 1 0 33120 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 31464 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_332
timestamp 1604681595
transform 1 0 31648 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_346
timestamp 1604681595
transform 1 0 32936 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 34040 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_
timestamp 1604681595
transform 1 0 35144 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 34868 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_prog_clk_A
timestamp 1604681595
transform 1 0 33488 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_350
timestamp 1604681595
transform 1 0 33304 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_354
timestamp 1604681595
transform 1 0 33672 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_362
timestamp 1604681595
transform 1 0 34408 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_366
timestamp 1604681595
transform 1 0 34776 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_369
timestamp 1604681595
transform 1 0 35052 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1604681595
transform 1 0 37076 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_389
timestamp 1604681595
transform 1 0 36892 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_393
timestamp 1604681595
transform 1 0 37260 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1604681595
transform -1 0 38824 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1604681595
transform 1 0 37628 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_398
timestamp 1604681595
transform 1 0 37720 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_406
timestamp 1604681595
transform 1 0 38456 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1840 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1604681595
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 1656 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_3
timestamp 1604681595
transform 1 0 1380 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4324 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4140 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_27
timestamp 1604681595
transform 1 0 3588 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_31
timestamp 1604681595
transform 1 0 3956 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_52
timestamp 1604681595
transform 1 0 5888 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_48
timestamp 1604681595
transform 1 0 5520 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_44
timestamp 1604681595
transform 1 0 5152 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__CLK
timestamp 1604681595
transform 1 0 5704 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 5336 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_62
timestamp 1604681595
transform 1 0 6808 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_57
timestamp 1604681595
transform 1 0 6348 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__CLK
timestamp 1604681595
transform 1 0 6164 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__D
timestamp 1604681595
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1604681595
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_
timestamp 1604681595
transform 1 0 6900 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 8832 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_82
timestamp 1604681595
transform 1 0 8648 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_86
timestamp 1604681595
transform 1 0 9016 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_94
timestamp 1604681595
transform 1 0 9752 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_90
timestamp 1604681595
transform 1 0 9384 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 9568 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 9200 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604681595
transform 1 0 10028 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_105
timestamp 1604681595
transform 1 0 10764 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_101
timestamp 1604681595
transform 1 0 10396 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
timestamp 1604681595
transform 1 0 10580 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 10948 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_109
timestamp 1604681595
transform 1 0 11132 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1604681595
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_121
timestamp 1604681595
transform 1 0 12236 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_123
timestamp 1604681595
transform 1 0 12420 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_131
timestamp 1604681595
transform 1 0 13156 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 13432 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 13248 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 15548 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 15916 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_153
timestamp 1604681595
transform 1 0 15180 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_159
timestamp 1604681595
transform 1 0 15732 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_163
timestamp 1604681595
transform 1 0 16100 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 18032 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1604681595
transform 1 0 17940 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 18584 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_175
timestamp 1604681595
transform 1 0 17204 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_188
timestamp 1604681595
transform 1 0 18400 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_192
timestamp 1604681595
transform 1 0 18768 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_196
timestamp 1604681595
transform 1 0 19136 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _60_
timestamp 1604681595
transform 1 0 20148 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21160 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20976 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19228 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_199
timestamp 1604681595
transform 1 0 19412 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_210
timestamp 1604681595
transform 1 0 20424 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_214
timestamp 1604681595
transform 1 0 20792 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 22172 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 22540 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_227
timestamp 1604681595
transform 1 0 21988 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_231
timestamp 1604681595
transform 1 0 22356 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_235
timestamp 1604681595
transform 1 0 22724 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_249
timestamp 1604681595
transform 1 0 24012 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_245
timestamp 1604681595
transform 1 0 23644 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_243
timestamp 1604681595
transform 1 0 23460 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 24104 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1604681595
transform 1 0 23552 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_260
timestamp 1604681595
transform 1 0 25024 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_256
timestamp 1604681595
transform 1 0 24656 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_252
timestamp 1604681595
transform 1 0 24288 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 24472 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 24840 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 25208 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 27140 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1604681595
transform 1 0 26956 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1604681595
transform 1 0 27692 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1604681595
transform 1 0 29164 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__D
timestamp 1604681595
transform 1 0 28980 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 27508 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_285
timestamp 1604681595
transform 1 0 27324 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_292
timestamp 1604681595
transform 1 0 27968 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_300
timestamp 1604681595
transform 1 0 28704 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_
timestamp 1604681595
transform 1 0 29808 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__D
timestamp 1604681595
transform 1 0 29624 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_306
timestamp 1604681595
transform 1 0 29256 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604681595
transform 1 0 32292 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1604681595
transform 1 0 32108 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1604681595
transform 1 0 31740 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_331
timestamp 1604681595
transform 1 0 31556 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_335
timestamp 1604681595
transform 1 0 31924 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_348
timestamp 1604681595
transform 1 0 33120 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604681595
transform 1 0 34868 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1604681595
transform 1 0 34776 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 34040 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 33304 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 33672 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 34592 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_352
timestamp 1604681595
transform 1 0 33488 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_356
timestamp 1604681595
transform 1 0 33856 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_360
timestamp 1604681595
transform 1 0 34224 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604681595
transform 1 0 36432 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__D
timestamp 1604681595
transform 1 0 35880 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1604681595
transform 1 0 36248 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_376
timestamp 1604681595
transform 1 0 35696 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_380
timestamp 1604681595
transform 1 0 36064 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_393
timestamp 1604681595
transform 1 0 37260 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1604681595
transform -1 0 38824 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1604681595
transform 1 0 37444 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__CLK
timestamp 1604681595
transform 1 0 37812 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_397
timestamp 1604681595
transform 1 0 37628 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_401
timestamp 1604681595
transform 1 0 37996 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_9
timestamp 1604681595
transform 1 0 1932 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_3
timestamp 1604681595
transform 1 0 1380 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_10
timestamp 1604681595
transform 1 0 2024 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_7
timestamp 1604681595
transform 1 0 1748 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_3
timestamp 1604681595
transform 1 0 1380 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 1748 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 1840 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1604681595
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1604681595
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_20
timestamp 1604681595
transform 1 0 2944 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 2116 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2116 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 2300 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_47_32
timestamp 1604681595
transform 1 0 4048 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_28
timestamp 1604681595
transform 1 0 3680 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_24
timestamp 1604681595
transform 1 0 3312 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3128 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1604681595
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_36
timestamp 1604681595
transform 1 0 4416 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 4600 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__D
timestamp 1604681595
transform 1 0 4232 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4784 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_
timestamp 1604681595
transform 1 0 4048 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_47_53
timestamp 1604681595
transform 1 0 5980 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_49
timestamp 1604681595
transform 1 0 5612 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 5796 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_62
timestamp 1604681595
transform 1 0 6808 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_57
timestamp 1604681595
transform 1 0 6348 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_63
timestamp 1604681595
transform 1 0 6900 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__CLK
timestamp 1604681595
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__D
timestamp 1604681595
transform 1 0 7084 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 6164 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1604681595
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_51
timestamp 1604681595
transform 1 0 5796 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_66
timestamp 1604681595
transform 1 0 7176 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_71
timestamp 1604681595
transform 1 0 7636 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_67
timestamp 1604681595
transform 1 0 7268 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1604681595
transform 1 0 7820 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1604681595
transform 1 0 7452 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1604681595
transform 1 0 7268 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604681595
transform 1 0 8004 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604681595
transform 1 0 7452 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_47_78
timestamp 1604681595
transform 1 0 8280 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_84
timestamp 1604681595
transform 1 0 8832 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604681595
transform 1 0 9016 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_98
timestamp 1604681595
transform 1 0 10120 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_94
timestamp 1604681595
transform 1 0 9752 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_90
timestamp 1604681595
transform 1 0 9384 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
timestamp 1604681595
transform 1 0 9936 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
timestamp 1604681595
transform 1 0 9568 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1604681595
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_106
timestamp 1604681595
transform 1 0 10856 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_105
timestamp 1604681595
transform 1 0 10764 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 11040 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 10948 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_93
timestamp 1604681595
transform 1 0 9660 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_118
timestamp 1604681595
transform 1 0 11960 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_114
timestamp 1604681595
transform 1 0 11592 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_110
timestamp 1604681595
transform 1 0 11224 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11408 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_131
timestamp 1604681595
transform 1 0 13156 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_127
timestamp 1604681595
transform 1 0 12788 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_131
timestamp 1604681595
transform 1 0 13156 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_123
timestamp 1604681595
transform 1 0 12420 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 12972 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1604681595
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 12420 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_111
timestamp 1604681595
transform 1 0 11316 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_139
timestamp 1604681595
transform 1 0 13892 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_135
timestamp 1604681595
transform 1 0 13524 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 13432 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 13340 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 13708 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_147
timestamp 1604681595
transform 1 0 14628 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_143
timestamp 1604681595
transform 1 0 14260 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_152
timestamp 1604681595
transform 1 0 15088 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_148
timestamp 1604681595
transform 1 0 14720 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _55_
timestamp 1604681595
transform 1 0 14352 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_136
timestamp 1604681595
transform 1 0 13616 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15548 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1604681595
transform 1 0 15180 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15364 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15732 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16100 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_154
timestamp 1604681595
transform 1 0 15272 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_157
timestamp 1604681595
transform 1 0 15548 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_161
timestamp 1604681595
transform 1 0 15916 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_165
timestamp 1604681595
transform 1 0 16284 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_184
timestamp 1604681595
transform 1 0 18032 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_177
timestamp 1604681595
transform 1 0 17388 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1604681595
transform 1 0 17940 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_190
timestamp 1604681595
transform 1 0 18584 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_195
timestamp 1604681595
transform 1 0 19044 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_191
timestamp 1604681595
transform 1 0 18676 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_188
timestamp 1604681595
transform 1 0 18400 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 18492 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18860 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 18400 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 18768 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_176
timestamp 1604681595
transform 1 0 17296 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 18952 0 1 27744
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_46_206
timestamp 1604681595
transform 1 0 20056 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_199
timestamp 1604681595
transform 1 0 19412 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19596 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19228 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _61_
timestamp 1604681595
transform 1 0 19780 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_215
timestamp 1604681595
transform 1 0 20884 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_215
timestamp 1604681595
transform 1 0 20884 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21068 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1604681595
transform 1 0 20792 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 21068 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21620 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21436 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 22632 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_236
timestamp 1604681595
transform 1 0 22816 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_219
timestamp 1604681595
transform 1 0 21252 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_232
timestamp 1604681595
transform 1 0 22448 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_236
timestamp 1604681595
transform 1 0 22816 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_240
timestamp 1604681595
transform 1 0 23184 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_245
timestamp 1604681595
transform 1 0 23644 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_248
timestamp 1604681595
transform 1 0 23920 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23368 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 24012 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1604681595
transform 1 0 23552 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_251
timestamp 1604681595
transform 1 0 24196 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_257
timestamp 1604681595
transform 1 0 24748 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1604681595
transform 1 0 24380 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24196 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 24564 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 24380 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 24840 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24564 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_47_268
timestamp 1604681595
transform 1 0 25760 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_264
timestamp 1604681595
transform 1 0 25392 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_271
timestamp 1604681595
transform 1 0 26036 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_267
timestamp 1604681595
transform 1 0 25668 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25852 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 25944 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 25576 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 26220 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1604681595
transform 1 0 26404 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 26496 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 26128 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1604681595
transform 1 0 29164 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 28060 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_295
timestamp 1604681595
transform 1 0 28244 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_291
timestamp 1604681595
transform 1 0 27876 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_295
timestamp 1604681595
transform 1 0 28244 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_303
timestamp 1604681595
transform 1 0 28980 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_
timestamp 1604681595
transform 1 0 29532 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_
timestamp 1604681595
transform 1 0 30176 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__D
timestamp 1604681595
transform 1 0 29992 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 29624 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__CLK
timestamp 1604681595
transform 1 0 29348 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_306
timestamp 1604681595
transform 1 0 29256 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_312
timestamp 1604681595
transform 1 0 29808 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_335
timestamp 1604681595
transform 1 0 31924 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_328
timestamp 1604681595
transform 1 0 31280 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 31832 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__D
timestamp 1604681595
transform 1 0 32108 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1604681595
transform 1 0 32016 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604681595
transform 1 0 32108 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_47_345
timestamp 1604681595
transform 1 0 32844 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_339
timestamp 1604681595
transform 1 0 32292 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_346
timestamp 1604681595
transform 1 0 32936 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1604681595
transform 1 0 32660 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1604681595
transform 1 0 33028 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1604681595
transform 1 0 33212 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604681595
transform 1 0 33212 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_47_358
timestamp 1604681595
transform 1 0 34040 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_357
timestamp 1604681595
transform 1 0 33948 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_351
timestamp 1604681595
transform 1 0 33396 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__CLK
timestamp 1604681595
transform 1 0 34224 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 34040 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_367
timestamp 1604681595
transform 1 0 34868 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_362
timestamp 1604681595
transform 1 0 34408 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_366
timestamp 1604681595
transform 1 0 34776 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_362
timestamp 1604681595
transform 1 0 34408 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 34592 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__D
timestamp 1604681595
transform 1 0 34960 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__D
timestamp 1604681595
transform 1 0 34592 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1604681595
transform 1 0 34776 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_
timestamp 1604681595
transform 1 0 35144 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_
timestamp 1604681595
transform 1 0 34960 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_46_389
timestamp 1604681595
transform 1 0 36892 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_387
timestamp 1604681595
transform 1 0 36708 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1604681595
transform -1 0 38824 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1604681595
transform -1 0 38824 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1604681595
transform 1 0 37628 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_398
timestamp 1604681595
transform 1 0 37720 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_406
timestamp 1604681595
transform 1 0 38456 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_399
timestamp 1604681595
transform 1 0 37812 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1604681595
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2208 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 1840 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_3
timestamp 1604681595
transform 1 0 1380 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_7
timestamp 1604681595
transform 1 0 1748 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_10
timestamp 1604681595
transform 1 0 2024 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_
timestamp 1604681595
transform 1 0 4048 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1604681595
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_23
timestamp 1604681595
transform 1 0 3220 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_
timestamp 1604681595
transform 1 0 7084 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_48_51
timestamp 1604681595
transform 1 0 5796 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_63
timestamp 1604681595
transform 1 0 6900 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_84
timestamp 1604681595
transform 1 0 8832 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604681595
transform 1 0 11040 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604681595
transform 1 0 9660 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1604681595
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 10396 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 10764 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_97
timestamp 1604681595
transform 1 0 10028 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_103
timestamp 1604681595
transform 1 0 10580 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_107
timestamp 1604681595
transform 1 0 10948 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 12604 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_117
timestamp 1604681595
transform 1 0 11868 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_129
timestamp 1604681595
transform 1 0 12972 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 13708 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 13432 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14260 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_133
timestamp 1604681595
transform 1 0 13340 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_136
timestamp 1604681595
transform 1 0 13616 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1604681595
transform 1 0 14076 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_145
timestamp 1604681595
transform 1 0 14444 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15364 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1604681595
transform 1 0 15180 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16376 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_154
timestamp 1604681595
transform 1 0 15272 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_164
timestamp 1604681595
transform 1 0 16192 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_168
timestamp 1604681595
transform 1 0 16560 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _62_
timestamp 1604681595
transform 1 0 18216 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 18952 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_180
timestamp 1604681595
transform 1 0 17664 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_189
timestamp 1604681595
transform 1 0 18492 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_193
timestamp 1604681595
transform 1 0 18860 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_196
timestamp 1604681595
transform 1 0 19136 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 20884 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1604681595
transform 1 0 20792 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 20240 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_206
timestamp 1604681595
transform 1 0 20056 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_210
timestamp 1604681595
transform 1 0 20424 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_234
timestamp 1604681595
transform 1 0 22632 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 24840 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 24656 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 23920 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 24288 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_246
timestamp 1604681595
transform 1 0 23736 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1604681595
transform 1 0 24104 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_254
timestamp 1604681595
transform 1 0 24472 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 26496 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1604681595
transform 1 0 26404 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25852 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 26220 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_267
timestamp 1604681595
transform 1 0 25668 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_271
timestamp 1604681595
transform 1 0 26036 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_295
timestamp 1604681595
transform 1 0 28244 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604681595
transform 1 0 30452 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 30268 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__CLK
timestamp 1604681595
transform 1 0 29900 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_307
timestamp 1604681595
transform 1 0 29348 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_48_315
timestamp 1604681595
transform 1 0 30084 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_
timestamp 1604681595
transform 1 0 32108 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1604681595
transform 1 0 32016 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__CLK
timestamp 1604681595
transform 1 0 31832 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_328
timestamp 1604681595
transform 1 0 31280 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_
timestamp 1604681595
transform 1 0 34592 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__CLK
timestamp 1604681595
transform 1 0 34408 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_356
timestamp 1604681595
transform 1 0 33856 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_48_383
timestamp 1604681595
transform 1 0 36340 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1604681595
transform -1 0 38824 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1604681595
transform 1 0 37628 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_395
timestamp 1604681595
transform 1 0 37444 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_398
timestamp 1604681595
transform 1 0 37720 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_406
timestamp 1604681595
transform 1 0 38456 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1604681595
transform 1 0 1380 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1604681595
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_7
timestamp 1604681595
transform 1 0 1748 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__D
timestamp 1604681595
transform 1 0 1564 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_11
timestamp 1604681595
transform 1 0 2116 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__D
timestamp 1604681595
transform 1 0 1932 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_15
timestamp 1604681595
transform 1 0 2484 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__CLK
timestamp 1604681595
transform 1 0 2300 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_19
timestamp 1604681595
transform 1 0 2852 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__CLK
timestamp 1604681595
transform 1 0 2668 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 3128 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_
timestamp 1604681595
transform 1 0 4232 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__D
timestamp 1604681595
transform 1 0 4048 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 3680 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_26
timestamp 1604681595
transform 1 0 3496 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_30
timestamp 1604681595
transform 1 0 3864 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1604681595
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__D
timestamp 1604681595
transform 1 0 6164 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 6992 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_53
timestamp 1604681595
transform 1 0 5980 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_57
timestamp 1604681595
transform 1 0 6348 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_62
timestamp 1604681595
transform 1 0 6808 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_
timestamp 1604681595
transform 1 0 7912 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__D
timestamp 1604681595
transform 1 0 7728 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 7360 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_66
timestamp 1604681595
transform 1 0 7176 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_70
timestamp 1604681595
transform 1 0 7544 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604681595
transform 1 0 10396 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__D
timestamp 1604681595
transform 1 0 9844 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 10212 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_93
timestamp 1604681595
transform 1 0 9660 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_97
timestamp 1604681595
transform 1 0 10028 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_114
timestamp 1604681595
transform 1 0 11592 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_110
timestamp 1604681595
transform 1 0 11224 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__CLK
timestamp 1604681595
transform 1 0 11408 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12144 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1604681595
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_127
timestamp 1604681595
transform 1 0 12788 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_123
timestamp 1604681595
transform 1 0 12420 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 12604 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12972 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_131
timestamp 1604681595
transform 1 0 13156 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 13432 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15916 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15732 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15364 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 16928 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_153
timestamp 1604681595
transform 1 0 15180 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_157
timestamp 1604681595
transform 1 0 15548 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_170
timestamp 1604681595
transform 1 0 16744 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_174
timestamp 1604681595
transform 1 0 17112 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_178
timestamp 1604681595
transform 1 0 17480 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 17296 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_184
timestamp 1604681595
transform 1 0 18032 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_182
timestamp 1604681595
transform 1 0 17848 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1604681595
transform 1 0 17940 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18400 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_194
timestamp 1604681595
transform 1 0 18952 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_190
timestamp 1604681595
transform 1 0 18584 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 18768 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 19136 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 19596 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_49_198
timestamp 1604681595
transform 1 0 19320 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_220
timestamp 1604681595
transform 1 0 21344 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_232
timestamp 1604681595
transform 1 0 22448 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_240
timestamp 1604681595
transform 1 0 23184 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 23920 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 25024 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1604681595
transform 1 0 23552 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 24656 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 23368 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_245
timestamp 1604681595
transform 1 0 23644 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_252
timestamp 1604681595
transform 1 0 24288 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_258
timestamp 1604681595
transform 1 0 24840 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_279
timestamp 1604681595
transform 1 0 26772 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _63_
timestamp 1604681595
transform 1 0 27508 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1604681595
transform 1 0 29164 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_prog_clk_A
timestamp 1604681595
transform 1 0 27968 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_290
timestamp 1604681595
transform 1 0 27784 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_294
timestamp 1604681595
transform 1 0 28152 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_302
timestamp 1604681595
transform 1 0 28888 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__D
timestamp 1604681595
transform 1 0 31096 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 30452 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_306
timestamp 1604681595
transform 1 0 29256 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_318
timestamp 1604681595
transform 1 0 30360 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_321
timestamp 1604681595
transform 1 0 30636 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_325
timestamp 1604681595
transform 1 0 31004 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_
timestamp 1604681595
transform 1 0 31280 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__D
timestamp 1604681595
transform 1 0 33212 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_347
timestamp 1604681595
transform 1 0 33028 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_
timestamp 1604681595
transform 1 0 34868 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1604681595
transform 1 0 34776 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1604681595
transform 1 0 34592 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__CLK
timestamp 1604681595
transform 1 0 33580 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__CLK
timestamp 1604681595
transform 1 0 34224 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_351
timestamp 1604681595
transform 1 0 33396 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_355
timestamp 1604681595
transform 1 0 33764 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_359
timestamp 1604681595
transform 1 0 34132 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_362
timestamp 1604681595
transform 1 0 34408 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_386
timestamp 1604681595
transform 1 0 36616 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1604681595
transform -1 0 38824 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_398
timestamp 1604681595
transform 1 0 37720 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_406
timestamp 1604681595
transform 1 0 38456 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_
timestamp 1604681595
transform 1 0 1380 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1604681595
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_
timestamp 1604681595
transform 1 0 4692 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1604681595
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 4416 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__CLK
timestamp 1604681595
transform 1 0 3312 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_22
timestamp 1604681595
transform 1 0 3128 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_26
timestamp 1604681595
transform 1 0 3496 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_32
timestamp 1604681595
transform 1 0 4048 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_38
timestamp 1604681595
transform 1 0 4600 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__CLK
timestamp 1604681595
transform 1 0 7084 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_58
timestamp 1604681595
transform 1 0 6440 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_64
timestamp 1604681595
transform 1 0 6992 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604681595
transform 1 0 8004 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1604681595
transform 1 0 7820 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 7452 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_67
timestamp 1604681595
transform 1 0 7268 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_71
timestamp 1604681595
transform 1 0 7636 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_84
timestamp 1604681595
transform 1 0 8832 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_
timestamp 1604681595
transform 1 0 9660 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1604681595
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_88
timestamp 1604681595
transform 1 0 9200 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12144 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_50_112
timestamp 1604681595
transform 1 0 11408 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 14996 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 14168 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14628 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_139
timestamp 1604681595
transform 1 0 13892 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_144
timestamp 1604681595
transform 1 0 14352 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_149
timestamp 1604681595
transform 1 0 14812 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15640 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1604681595
transform 1 0 15180 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15456 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_154
timestamp 1604681595
transform 1 0 15272 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _58_
timestamp 1604681595
transform 1 0 18124 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19136 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 17572 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 17940 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18584 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_177
timestamp 1604681595
transform 1 0 17388 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_181
timestamp 1604681595
transform 1 0 17756 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_188
timestamp 1604681595
transform 1 0 18400 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_192
timestamp 1604681595
transform 1 0 18768 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1604681595
transform 1 0 20792 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 20148 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 21068 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_205
timestamp 1604681595
transform 1 0 19964 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_209
timestamp 1604681595
transform 1 0 20332 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_213
timestamp 1604681595
transform 1 0 20700 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_215
timestamp 1604681595
transform 1 0 20884 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 21436 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_219
timestamp 1604681595
transform 1 0 21252 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_223
timestamp 1604681595
transform 1 0 21620 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_235
timestamp 1604681595
transform 1 0 22724 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 23552 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 24656 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24472 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 24104 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_243
timestamp 1604681595
transform 1 0 23460 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_248
timestamp 1604681595
transform 1 0 23920 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_252
timestamp 1604681595
transform 1 0 24288 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1604681595
transform 1 0 26496 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1604681595
transform 1 0 26404 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 25668 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_265
timestamp 1604681595
transform 1 0 25484 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_269
timestamp 1604681595
transform 1 0 25852 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_279
timestamp 1604681595
transform 1 0 26772 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_prog_clk
timestamp 1604681595
transform 1 0 27508 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_290
timestamp 1604681595
transform 1 0 27784 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_302
timestamp 1604681595
transform 1 0 28888 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_314
timestamp 1604681595
transform 1 0 29992 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_326
timestamp 1604681595
transform 1 0 31096 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_
timestamp 1604681595
transform 1 0 32200 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1604681595
transform 1 0 32016 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__CLK
timestamp 1604681595
transform 1 0 31280 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_330
timestamp 1604681595
transform 1 0 31464 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_337
timestamp 1604681595
transform 1 0 32108 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_7.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__D
timestamp 1604681595
transform 1 0 34868 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_357
timestamp 1604681595
transform 1 0 33948 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_365
timestamp 1604681595
transform 1 0 34684 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_369
timestamp 1604681595
transform 1 0 35052 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604681595
transform 1 0 35420 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1604681595
transform 1 0 35788 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_389
timestamp 1604681595
transform 1 0 36892 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1604681595
transform -1 0 38824 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1604681595
transform 1 0 37628 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_398
timestamp 1604681595
transform 1 0 37720 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_406
timestamp 1604681595
transform 1 0 38456 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_
timestamp 1604681595
transform 1 0 1380 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1604681595
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604681595
transform 1 0 4600 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 4416 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 4048 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 3680 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3312 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_22
timestamp 1604681595
transform 1 0 3128 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_26
timestamp 1604681595
transform 1 0 3496 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_30
timestamp 1604681595
transform 1 0 3864 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_34
timestamp 1604681595
transform 1 0 4232 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604681595
transform 1 0 6808 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1604681595
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
timestamp 1604681595
transform 1 0 5980 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 5612 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_47
timestamp 1604681595
transform 1 0 5428 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_51
timestamp 1604681595
transform 1 0 5796 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_55
timestamp 1604681595
transform 1 0 6164 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_
timestamp 1604681595
transform 1 0 8556 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
timestamp 1604681595
transform 1 0 7360 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1604681595
transform 1 0 8004 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__D
timestamp 1604681595
transform 1 0 8372 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_66
timestamp 1604681595
transform 1 0 7176 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_70
timestamp 1604681595
transform 1 0 7544 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_74
timestamp 1604681595
transform 1 0 7912 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_77
timestamp 1604681595
transform 1 0 8188 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__D
timestamp 1604681595
transform 1 0 10488 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__CLK
timestamp 1604681595
transform 1 0 10856 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_100
timestamp 1604681595
transform 1 0 10304 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_104
timestamp 1604681595
transform 1 0 10672 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_108
timestamp 1604681595
transform 1 0 11040 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 11224 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1604681595
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 11776 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_114
timestamp 1604681595
transform 1 0 11592 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_118
timestamp 1604681595
transform 1 0 11960 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_132
timestamp 1604681595
transform 1 0 13248 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13432 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_140
timestamp 1604681595
transform 1 0 13984 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_136
timestamp 1604681595
transform 1 0 13616 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13800 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 14168 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_150
timestamp 1604681595
transform 1 0 14904 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_146
timestamp 1604681595
transform 1 0 14536 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 14720 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 15088 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 15272 0 1 29920
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1604681595
transform 1 0 17940 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 17388 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19044 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_175
timestamp 1604681595
transform 1 0 17204 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_179
timestamp 1604681595
transform 1 0 17572 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_193
timestamp 1604681595
transform 1 0 18860 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 20148 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 19964 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_197
timestamp 1604681595
transform 1 0 19228 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_226
timestamp 1604681595
transform 1 0 21896 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_238
timestamp 1604681595
transform 1 0 23000 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 24656 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1604681595
transform 1 0 23552 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 24472 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 24104 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 23368 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_245
timestamp 1604681595
transform 1 0 23644 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_249
timestamp 1604681595
transform 1 0 24012 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_252
timestamp 1604681595
transform 1 0 24288 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 26588 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_275
timestamp 1604681595
transform 1 0 26404 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_279
timestamp 1604681595
transform 1 0 26772 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1604681595
transform 1 0 29164 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__D
timestamp 1604681595
transform 1 0 28336 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__CLK
timestamp 1604681595
transform 1 0 28704 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_291
timestamp 1604681595
transform 1 0 27876 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_295
timestamp 1604681595
transform 1 0 28244 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_298
timestamp 1604681595
transform 1 0 28520 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_302
timestamp 1604681595
transform 1 0 28888 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_306
timestamp 1604681595
transform 1 0 29256 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_318
timestamp 1604681595
transform 1 0 30360 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_330
timestamp 1604681595
transform 1 0 31464 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_342
timestamp 1604681595
transform 1 0 32568 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1604681595
transform 1 0 34776 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1604681595
transform 1 0 35236 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_354
timestamp 1604681595
transform 1 0 33672 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_367
timestamp 1604681595
transform 1 0 34868 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604681595
transform 1 0 35420 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1604681595
transform 1 0 35972 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_377
timestamp 1604681595
transform 1 0 35788 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_381
timestamp 1604681595
transform 1 0 36156 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1604681595
transform 1 0 37260 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1604681595
transform -1 0 38824 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1604681595
transform 1 0 38364 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_
timestamp 1604681595
transform 1 0 1472 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_
timestamp 1604681595
transform 1 0 2208 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1604681595
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1604681595
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__D
timestamp 1604681595
transform 1 0 2024 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__D
timestamp 1604681595
transform 1 0 1564 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_3
timestamp 1604681595
transform 1 0 1380 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1604681595
transform 1 0 1380 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_7
timestamp 1604681595
transform 1 0 1748 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_31
timestamp 1604681595
transform 1 0 3956 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_23
timestamp 1604681595
transform 1 0 3220 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1604681595
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_35
timestamp 1604681595
transform 1 0 4324 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_32
timestamp 1604681595
transform 1 0 4048 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1604681595
transform 1 0 4232 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1604681595
transform 1 0 4508 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1604681595
transform 1 0 4140 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604681595
transform 1 0 4692 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4416 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_53_53
timestamp 1604681595
transform 1 0 5980 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_48
timestamp 1604681595
transform 1 0 5520 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_49
timestamp 1604681595
transform 1 0 5612 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_45
timestamp 1604681595
transform 1 0 5244 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 5428 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 5796 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604681595
transform 1 0 5980 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_62
timestamp 1604681595
transform 1 0 6808 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_57
timestamp 1604681595
transform 1 0 6348 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1604681595
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_57
timestamp 1604681595
transform 1 0 6348 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_70
timestamp 1604681595
transform 1 0 7544 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_69
timestamp 1604681595
transform 1 0 7452 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1604681595
transform 1 0 7820 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604681595
transform 1 0 8004 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 7728 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_84
timestamp 1604681595
transform 1 0 8832 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_80
timestamp 1604681595
transform 1 0 8464 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_76
timestamp 1604681595
transform 1 0 8096 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_84
timestamp 1604681595
transform 1 0 8832 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 8648 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 8280 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1604681595
transform 1 0 9108 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_98
timestamp 1604681595
transform 1 0 10120 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_97
timestamp 1604681595
transform 1 0 10028 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_93
timestamp 1604681595
transform 1 0 9660 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_91
timestamp 1604681595
transform 1 0 9476 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_88
timestamp 1604681595
transform 1 0 9200 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 9844 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1604681595
transform 1 0 9292 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1604681595
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604681595
transform 1 0 9292 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_52_101
timestamp 1604681595
transform 1 0 10396 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1604681595
transform 1 0 10304 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_102
timestamp 1604681595
transform 1 0 10488 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_
timestamp 1604681595
transform 1 0 10488 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_53_114
timestamp 1604681595
transform 1 0 11592 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_128
timestamp 1604681595
transform 1 0 12880 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_125
timestamp 1604681595
transform 1 0 12604 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_121
timestamp 1604681595
transform 1 0 12236 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 12788 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 12420 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
timestamp 1604681595
transform 1 0 12144 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1604681595
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 31008
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1604681595
transform 1 0 13064 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12972 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_53_132
timestamp 1604681595
transform 1 0 13248 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_138
timestamp 1604681595
transform 1 0 13800 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 13616 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_144
timestamp 1604681595
transform 1 0 14352 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_140
timestamp 1604681595
transform 1 0 13984 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_146
timestamp 1604681595
transform 1 0 14536 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14720 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 14168 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_150
timestamp 1604681595
transform 1 0 14904 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_149
timestamp 1604681595
transform 1 0 14812 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 15088 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 17112 0 -1 31008
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15272 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15548 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1604681595
transform 1 0 15180 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 16928 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_154
timestamp 1604681595
transform 1 0 15272 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_166
timestamp 1604681595
transform 1 0 16376 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_173
timestamp 1604681595
transform 1 0 17020 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1604681595
transform 1 0 17940 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17572 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18216 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 17204 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_195
timestamp 1604681595
transform 1 0 19044 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_177
timestamp 1604681595
transform 1 0 17388 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_181
timestamp 1604681595
transform 1 0 17756 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_184
timestamp 1604681595
transform 1 0 18032 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_188
timestamp 1604681595
transform 1 0 18400 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_200
timestamp 1604681595
transform 1 0 19504 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 20148 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_214
timestamp 1604681595
transform 1 0 20792 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_210
timestamp 1604681595
transform 1 0 20424 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_213
timestamp 1604681595
transform 1 0 20700 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_209
timestamp 1604681595
transform 1 0 20332 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20240 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 20608 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20976 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1604681595
transform 1 0 20792 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21160 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 20884 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 22172 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 22540 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_234
timestamp 1604681595
transform 1 0 22632 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_227
timestamp 1604681595
transform 1 0 21988 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_231
timestamp 1604681595
transform 1 0 22356 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_235
timestamp 1604681595
transform 1 0 22724 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 23552 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1604681595
transform 1 0 23552 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 23368 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_242
timestamp 1604681595
transform 1 0 23368 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_241
timestamp 1604681595
transform 1 0 23276 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_245
timestamp 1604681595
transform 1 0 23644 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_248
timestamp 1604681595
transform 1 0 23920 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_249
timestamp 1604681595
transform 1 0 24012 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 24104 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 24104 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_252
timestamp 1604681595
transform 1 0 24288 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_252
timestamp 1604681595
transform 1 0 24288 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 24472 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 24472 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24656 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 24656 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_52_269
timestamp 1604681595
transform 1 0 25852 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_52_265
timestamp 1604681595
transform 1 0 25484 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 25668 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_279
timestamp 1604681595
transform 1 0 26772 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_275
timestamp 1604681595
transform 1 0 26404 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1604681595
transform 1 0 26588 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1604681595
transform 1 0 26404 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 26496 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_283
timestamp 1604681595
transform 1 0 27140 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_280
timestamp 1604681595
transform 1 0 26864 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
timestamp 1604681595
transform 1 0 26956 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_294
timestamp 1604681595
transform 1 0 28152 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_290
timestamp 1604681595
transform 1 0 27784 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1604681595
transform 1 0 27968 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1604681595
transform 1 0 27600 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1604681595
transform 1 0 27416 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604681595
transform 1 0 27600 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_53_301
timestamp 1604681595
transform 1 0 28796 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_297
timestamp 1604681595
transform 1 0 28428 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__CLK
timestamp 1604681595
transform 1 0 28980 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__D
timestamp 1604681595
transform 1 0 28612 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1604681595
transform 1 0 29164 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_
timestamp 1604681595
transform 1 0 28336 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_52_315
timestamp 1604681595
transform 1 0 30084 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_327
timestamp 1604681595
transform 1 0 31188 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_306
timestamp 1604681595
transform 1 0 29256 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_318
timestamp 1604681595
transform 1 0 30360 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1604681595
transform 1 0 32016 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_335
timestamp 1604681595
transform 1 0 31924 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_337
timestamp 1604681595
transform 1 0 32108 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_349
timestamp 1604681595
transform 1 0 33212 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_330
timestamp 1604681595
transform 1 0 31464 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_342
timestamp 1604681595
transform 1 0 32568 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1604681595
transform 1 0 34776 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_361
timestamp 1604681595
transform 1 0 34316 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_354
timestamp 1604681595
transform 1 0 33672 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_367
timestamp 1604681595
transform 1 0 34868 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604681595
transform 1 0 35420 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1604681595
transform 1 0 35420 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1604681595
transform 1 0 35788 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_389
timestamp 1604681595
transform 1 0 36892 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_375
timestamp 1604681595
transform 1 0 35604 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_387
timestamp 1604681595
transform 1 0 36708 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1604681595
transform -1 0 38824 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1604681595
transform -1 0 38824 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1604681595
transform 1 0 37628 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_398
timestamp 1604681595
transform 1 0 37720 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_406
timestamp 1604681595
transform 1 0 38456 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_399
timestamp 1604681595
transform 1 0 37812 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604681595
transform 1 0 1932 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1604681595
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 1748 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__CLK
timestamp 1604681595
transform 1 0 2944 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_3
timestamp 1604681595
transform 1 0 1380 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_18
timestamp 1604681595
transform 1 0 2760 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604681595
transform 1 0 4048 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1604681595
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 5060 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_22
timestamp 1604681595
transform 1 0 3128 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_30
timestamp 1604681595
transform 1 0 3864 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_41
timestamp 1604681595
transform 1 0 4876 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604681595
transform 1 0 5796 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 5428 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 6808 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_45
timestamp 1604681595
transform 1 0 5244 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_49
timestamp 1604681595
transform 1 0 5612 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_60
timestamp 1604681595
transform 1 0 6624 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_64
timestamp 1604681595
transform 1 0 6992 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 7820 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_prog_clk
timestamp 1604681595
transform 1 0 9016 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
timestamp 1604681595
transform 1 0 8372 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_72
timestamp 1604681595
transform 1 0 7728 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_77
timestamp 1604681595
transform 1 0 8188 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_81
timestamp 1604681595
transform 1 0 8556 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_85
timestamp 1604681595
transform 1 0 8924 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1604681595
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9844 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 10672 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_89
timestamp 1604681595
transform 1 0 9292 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_93
timestamp 1604681595
transform 1 0 9660 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_97
timestamp 1604681595
transform 1 0 10028 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_103
timestamp 1604681595
transform 1 0 10580 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_106
timestamp 1604681595
transform 1 0 10856 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_118
timestamp 1604681595
transform 1 0 11960 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_130
timestamp 1604681595
transform 1 0 13064 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _54_
timestamp 1604681595
transform 1 0 14076 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 14536 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14904 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_138
timestamp 1604681595
transform 1 0 13800 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_144
timestamp 1604681595
transform 1 0 14352 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_148
timestamp 1604681595
transform 1 0 14720 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_152
timestamp 1604681595
transform 1 0 15088 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_154
timestamp 1604681595
transform 1 0 15272 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCD
timestamp 1604681595
transform 1 0 15456 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1604681595
transform 1 0 15180 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_158
timestamp 1604681595
transform 1 0 15640 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 15824 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_prog_clk
timestamp 1604681595
transform 1 0 16008 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_165
timestamp 1604681595
transform 1 0 16284 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 16468 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_169
timestamp 1604681595
transform 1 0 16652 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 17020 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 17572 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 18584 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 17388 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 18952 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_175
timestamp 1604681595
transform 1 0 17204 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_188
timestamp 1604681595
transform 1 0 18400 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_192
timestamp 1604681595
transform 1 0 18768 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_196
timestamp 1604681595
transform 1 0 19136 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 20976 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1604681595
transform 1 0 20792 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 20608 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_208
timestamp 1604681595
transform 1 0 20240 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_215
timestamp 1604681595
transform 1 0 20884 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 22908 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_235
timestamp 1604681595
transform 1 0 22724 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_239
timestamp 1604681595
transform 1 0 23092 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604681595
transform 1 0 24656 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 23460 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23276 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 24012 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 24472 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_247
timestamp 1604681595
transform 1 0 23828 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_251
timestamp 1604681595
transform 1 0 24196 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604681595
transform 1 0 26496 0 -1 32096
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1604681595
transform 1 0 26404 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 26036 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 25668 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 27140 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_265
timestamp 1604681595
transform 1 0 25484 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_269
timestamp 1604681595
transform 1 0 25852 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_273
timestamp 1604681595
transform 1 0 26220 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_281
timestamp 1604681595
transform 1 0 26956 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_
timestamp 1604681595
transform 1 0 28152 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1604681595
transform 1 0 27600 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__CLK
timestamp 1604681595
transform 1 0 27968 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_285
timestamp 1604681595
transform 1 0 27324 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_290
timestamp 1604681595
transform 1 0 27784 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__CLK
timestamp 1604681595
transform 1 0 30084 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_313
timestamp 1604681595
transform 1 0 29900 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_317
timestamp 1604681595
transform 1 0 30268 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1604681595
transform 1 0 32016 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_329
timestamp 1604681595
transform 1 0 31372 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_335
timestamp 1604681595
transform 1 0 31924 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_337
timestamp 1604681595
transform 1 0 32108 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_349
timestamp 1604681595
transform 1 0 33212 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_361
timestamp 1604681595
transform 1 0 34316 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604681595
transform 1 0 35420 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1604681595
transform 1 0 35788 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_389
timestamp 1604681595
transform 1 0 36892 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1604681595
transform -1 0 38824 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1604681595
transform 1 0 37628 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_398
timestamp 1604681595
transform 1 0 37720 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_406
timestamp 1604681595
transform 1 0 38456 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1604681595
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__D
timestamp 1604681595
transform 1 0 2944 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 1932 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 2300 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_3
timestamp 1604681595
transform 1 0 1380 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_11
timestamp 1604681595
transform 1 0 2116 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_15
timestamp 1604681595
transform 1 0 2484 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_19
timestamp 1604681595
transform 1 0 2852 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_
timestamp 1604681595
transform 1 0 3128 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__D
timestamp 1604681595
transform 1 0 5060 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_41
timestamp 1604681595
transform 1 0 4876 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_45
timestamp 1604681595
transform 1 0 5244 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__CLK
timestamp 1604681595
transform 1 0 5428 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_53
timestamp 1604681595
transform 1 0 5980 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604681595
transform 1 0 5612 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_57
timestamp 1604681595
transform 1 0 6348 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
timestamp 1604681595
transform 1 0 6164 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_62
timestamp 1604681595
transform 1 0 6808 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1604681595
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 6992 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1604681595
transform 1 0 7728 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 7544 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 9108 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 8740 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_66
timestamp 1604681595
transform 1 0 7176 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_81
timestamp 1604681595
transform 1 0 8556 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_85
timestamp 1604681595
transform 1 0 8924 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 9292 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 10672 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9844 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10212 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_93
timestamp 1604681595
transform 1 0 9660 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_97
timestamp 1604681595
transform 1 0 10028 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_101
timestamp 1604681595
transform 1 0 10396 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_107
timestamp 1604681595
transform 1 0 10948 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_112
timestamp 1604681595
transform 1 0 11408 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11224 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_116
timestamp 1604681595
transform 1 0 11776 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11592 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_120
timestamp 1604681595
transform 1 0 12144 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11960 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_123
timestamp 1604681595
transform 1 0 12420 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1604681595
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_128
timestamp 1604681595
transform 1 0 12880 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 12696 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13064 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 14352 0 1 32096
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1604681595
transform 1 0 14168 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13800 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_132
timestamp 1604681595
transform 1 0 13248 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_136
timestamp 1604681595
transform 1 0 13616 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_140
timestamp 1604681595
transform 1 0 13984 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_prog_clk
timestamp 1604681595
transform 1 0 17020 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 16468 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 16836 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_165
timestamp 1604681595
transform 1 0 16284 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1604681595
transform 1 0 16652 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18032 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1604681595
transform 1 0 17940 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 17756 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_176
timestamp 1604681595
transform 1 0 17296 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_180
timestamp 1604681595
transform 1 0 17664 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 20976 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 20792 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 20424 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 20056 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_203
timestamp 1604681595
transform 1 0 19780 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_208
timestamp 1604681595
transform 1 0 20240 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_212
timestamp 1604681595
transform 1 0 20608 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 22908 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_235
timestamp 1604681595
transform 1 0 22724 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_239
timestamp 1604681595
transform 1 0 23092 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1604681595
transform 1 0 23552 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 23368 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 24840 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 25208 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_254
timestamp 1604681595
transform 1 0 24472 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_260
timestamp 1604681595
transform 1 0 25024 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604681595
transform 1 0 26036 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 27048 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 25852 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_264
timestamp 1604681595
transform 1 0 25392 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_268
timestamp 1604681595
transform 1 0 25760 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_280
timestamp 1604681595
transform 1 0 26864 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604681595
transform 1 0 27600 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1604681595
transform 1 0 29164 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__D
timestamp 1604681595
transform 1 0 28980 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1604681595
transform 1 0 27416 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__D
timestamp 1604681595
transform 1 0 28612 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_284
timestamp 1604681595
transform 1 0 27232 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_297
timestamp 1604681595
transform 1 0 28428 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_301
timestamp 1604681595
transform 1 0 28796 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_
timestamp 1604681595
transform 1 0 29256 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_55_325
timestamp 1604681595
transform 1 0 31004 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_337
timestamp 1604681595
transform 1 0 32108 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_349
timestamp 1604681595
transform 1 0 33212 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1604681595
transform 1 0 34776 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_361
timestamp 1604681595
transform 1 0 34316 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_365
timestamp 1604681595
transform 1 0 34684 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_367
timestamp 1604681595
transform 1 0 34868 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_379
timestamp 1604681595
transform 1 0 35972 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_391
timestamp 1604681595
transform 1 0 37076 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1604681595
transform -1 0 38824 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_403
timestamp 1604681595
transform 1 0 38180 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1604681595
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1604681595
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_15
timestamp 1604681595
transform 1 0 2484 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_21
timestamp 1604681595
transform 1 0 3036 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_
timestamp 1604681595
transform 1 0 4048 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1604681595
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__CLK
timestamp 1604681595
transform 1 0 3128 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_24
timestamp 1604681595
transform 1 0 3312 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_30
timestamp 1604681595
transform 1 0 3864 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604681595
transform 1 0 6532 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__CLK
timestamp 1604681595
transform 1 0 5980 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_51
timestamp 1604681595
transform 1 0 5796 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_55
timestamp 1604681595
transform 1 0 6164 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1604681595
transform 1 0 8096 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8648 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 7728 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9016 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_68
timestamp 1604681595
transform 1 0 7360 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_74
timestamp 1604681595
transform 1 0 7912 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_80
timestamp 1604681595
transform 1 0 8464 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_84
timestamp 1604681595
transform 1 0 8832 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1604681595
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 9384 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_88
timestamp 1604681595
transform 1 0 9200 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_102
timestamp 1604681595
transform 1 0 10488 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11224 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 12788 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_119
timestamp 1604681595
transform 1 0 12052 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_130
timestamp 1604681595
transform 1 0 13064 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13432 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_default_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__D
timestamp 1604681595
transform 1 0 14444 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 13248 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_143
timestamp 1604681595
transform 1 0 14260 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_147
timestamp 1604681595
transform 1 0 14628 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_default_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1604681595
transform 1 0 15272 0 -1 33184
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1604681595
transform 1 0 15180 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 17940 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 17756 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 17388 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_175
timestamp 1604681595
transform 1 0 17204 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_179
timestamp 1604681595
transform 1 0 17572 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1604681595
transform 1 0 20792 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__D
timestamp 1604681595
transform 1 0 21068 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_202
timestamp 1604681595
transform 1 0 19688 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_210
timestamp 1604681595
transform 1 0 20424 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_215
timestamp 1604681595
transform 1 0 20884 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1604681595
transform 1 0 21344 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1604681595
transform 1 0 22908 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 22724 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_219
timestamp 1604681595
transform 1 0 21252 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_229
timestamp 1604681595
transform 1 0 22172 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1604681595
transform 1 0 24840 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 23920 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 24288 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 24656 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_246
timestamp 1604681595
transform 1 0 23736 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1604681595
transform 1 0 24104 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_254
timestamp 1604681595
transform 1 0 24472 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1604681595
transform 1 0 26496 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1604681595
transform 1 0 26404 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 25852 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 26220 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_267
timestamp 1604681595
transform 1 0 25668 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_271
timestamp 1604681595
transform 1 0 26036 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_
timestamp 1604681595
transform 1 0 28336 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1604681595
transform 1 0 27600 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
timestamp 1604681595
transform 1 0 27968 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_285
timestamp 1604681595
transform 1 0 27324 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_290
timestamp 1604681595
transform 1 0 27784 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_294
timestamp 1604681595
transform 1 0 28152 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_315
timestamp 1604681595
transform 1 0 30084 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_327
timestamp 1604681595
transform 1 0 31188 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1604681595
transform 1 0 32016 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_335
timestamp 1604681595
transform 1 0 31924 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_337
timestamp 1604681595
transform 1 0 32108 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_349
timestamp 1604681595
transform 1 0 33212 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_361
timestamp 1604681595
transform 1 0 34316 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_373
timestamp 1604681595
transform 1 0 35420 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_385
timestamp 1604681595
transform 1 0 36524 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1604681595
transform -1 0 38824 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1604681595
transform 1 0 37628 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_398
timestamp 1604681595
transform 1 0 37720 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_406
timestamp 1604681595
transform 1 0 38456 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1604681595
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1604681595
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_15
timestamp 1604681595
transform 1 0 2484 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_
timestamp 1604681595
transform 1 0 4232 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1604681595
transform 1 0 4048 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__D
timestamp 1604681595
transform 1 0 3680 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__CLK
timestamp 1604681595
transform 1 0 3312 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_23
timestamp 1604681595
transform 1 0 3220 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_26
timestamp 1604681595
transform 1 0 3496 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_30
timestamp 1604681595
transform 1 0 3864 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1604681595
transform 1 0 6808 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1604681595
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__D
timestamp 1604681595
transform 1 0 6164 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1604681595
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_53
timestamp 1604681595
transform 1 0 5980 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_57
timestamp 1604681595
transform 1 0 6348 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 8740 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_prog_clk
timestamp 1604681595
transform 1 0 8464 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8004 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_71
timestamp 1604681595
transform 1 0 7636 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_57_77
timestamp 1604681595
transform 1 0 8188 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 10672 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11040 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_102
timestamp 1604681595
transform 1 0 10488 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_106
timestamp 1604681595
transform 1 0 10856 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _52_
timestamp 1604681595
transform 1 0 11224 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 12972 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1604681595
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 12144 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 12788 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11776 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_113
timestamp 1604681595
transform 1 0 11500 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_118
timestamp 1604681595
transform 1 0 11960 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_123
timestamp 1604681595
transform 1 0 12420 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 14904 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_148
timestamp 1604681595
transform 1 0 14720 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_152
timestamp 1604681595
transform 1 0 15088 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15456 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15272 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 18032 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1604681595
transform 1 0 17940 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17388 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 17756 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_175
timestamp 1604681595
transform 1 0 17204 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_179
timestamp 1604681595
transform 1 0 17572 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_
timestamp 1604681595
transform 1 0 20700 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__D
timestamp 1604681595
transform 1 0 20516 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__CLK
timestamp 1604681595
transform 1 0 20148 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_203
timestamp 1604681595
transform 1 0 19780 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_209
timestamp 1604681595
transform 1 0 20332 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 23000 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 22632 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_232
timestamp 1604681595
transform 1 0 22448 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_236
timestamp 1604681595
transform 1 0 22816 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_240
timestamp 1604681595
transform 1 0 23184 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1604681595
transform 1 0 23552 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 23368 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 24656 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_254
timestamp 1604681595
transform 1 0 24472 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_258
timestamp 1604681595
transform 1 0 24840 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_262
timestamp 1604681595
transform 1 0 25208 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1604681595
transform 1 0 25852 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
timestamp 1604681595
transform 1 0 26864 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 25668 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
timestamp 1604681595
transform 1 0 25300 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_265
timestamp 1604681595
transform 1 0 25484 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_278
timestamp 1604681595
transform 1 0 26680 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_282
timestamp 1604681595
transform 1 0 27048 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1604681595
transform 1 0 27416 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1604681595
transform 1 0 29164 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
timestamp 1604681595
transform 1 0 27232 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__D
timestamp 1604681595
transform 1 0 28428 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__CLK
timestamp 1604681595
transform 1 0 28796 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_295
timestamp 1604681595
transform 1 0 28244 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_299
timestamp 1604681595
transform 1 0 28612 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_303
timestamp 1604681595
transform 1 0 28980 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_306
timestamp 1604681595
transform 1 0 29256 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_318
timestamp 1604681595
transform 1 0 30360 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_330
timestamp 1604681595
transform 1 0 31464 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_342
timestamp 1604681595
transform 1 0 32568 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1604681595
transform 1 0 34776 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1604681595
transform 1 0 35236 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_354
timestamp 1604681595
transform 1 0 33672 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_367
timestamp 1604681595
transform 1 0 34868 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1604681595
transform 1 0 35420 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1604681595
transform 1 0 35972 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_377
timestamp 1604681595
transform 1 0 35788 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_381
timestamp 1604681595
transform 1 0 36156 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1604681595
transform 1 0 37260 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1604681595
transform -1 0 38824 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1604681595
transform 1 0 38364 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1604681595
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1604681595
transform 1 0 1564 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_3
timestamp 1604681595
transform 1 0 1380 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_7
timestamp 1604681595
transform 1 0 1748 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_19
timestamp 1604681595
transform 1 0 2852 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1604681595
transform 1 0 4048 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1604681595
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 4600 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 4968 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_36
timestamp 1604681595
transform 1 0 4416 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_40
timestamp 1604681595
transform 1 0 4784 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_
timestamp 1604681595
transform 1 0 5244 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_58_44
timestamp 1604681595
transform 1 0 5152 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_64
timestamp 1604681595
transform 1 0 6992 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1604681595
transform 1 0 7176 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
timestamp 1604681595
transform 1 0 7544 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 9016 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_68
timestamp 1604681595
transform 1 0 7360 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_72
timestamp 1604681595
transform 1 0 7728 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_84
timestamp 1604681595
transform 1 0 8832 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9660 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1604681595
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_88
timestamp 1604681595
transform 1 0 9200 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 12144 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11592 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_112
timestamp 1604681595
transform 1 0 11408 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_116
timestamp 1604681595
transform 1 0 11776 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 14628 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14076 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 14444 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_139
timestamp 1604681595
transform 1 0 13892 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_143
timestamp 1604681595
transform 1 0 14260 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_150
timestamp 1604681595
transform 1 0 14904 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15824 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1604681595
transform 1 0 15180 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15456 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 16836 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_154
timestamp 1604681595
transform 1 0 15272 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_158
timestamp 1604681595
transform 1 0 15640 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_169
timestamp 1604681595
transform 1 0 16652 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_173
timestamp 1604681595
transform 1 0 17020 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 17388 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 17204 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_196
timestamp 1604681595
transform 1 0 19136 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_
timestamp 1604681595
transform 1 0 20884 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1604681595
transform 1 0 20792 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_208
timestamp 1604681595
transform 1 0 20240 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__CLK
timestamp 1604681595
transform 1 0 22816 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_234
timestamp 1604681595
transform 1 0 22632 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_238
timestamp 1604681595
transform 1 0 23000 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1604681595
transform 1 0 23368 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 24380 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_251
timestamp 1604681595
transform 1 0 24196 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_255
timestamp 1604681595
transform 1 0 24564 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1604681595
transform 1 0 25300 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1604681595
transform 1 0 26496 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1604681595
transform 1 0 26404 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
timestamp 1604681595
transform 1 0 27048 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 25852 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_267
timestamp 1604681595
transform 1 0 25668 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_271
timestamp 1604681595
transform 1 0 26036 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_280
timestamp 1604681595
transform 1 0 26864 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_
timestamp 1604681595
transform 1 0 27876 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__D
timestamp 1604681595
transform 1 0 27416 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_284
timestamp 1604681595
transform 1 0 27232 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_288
timestamp 1604681595
transform 1 0 27600 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_310
timestamp 1604681595
transform 1 0 29624 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_322
timestamp 1604681595
transform 1 0 30728 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1604681595
transform 1 0 32016 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_334
timestamp 1604681595
transform 1 0 31832 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_337
timestamp 1604681595
transform 1 0 32108 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_349
timestamp 1604681595
transform 1 0 33212 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_361
timestamp 1604681595
transform 1 0 34316 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604681595
transform 1 0 35420 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1604681595
transform 1 0 35788 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_389
timestamp 1604681595
transform 1 0 36892 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1604681595
transform -1 0 38824 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1604681595
transform 1 0 37628 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_398
timestamp 1604681595
transform 1 0 37720 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_406
timestamp 1604681595
transform 1 0 38456 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_7
timestamp 1604681595
transform 1 0 1748 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1604681595
transform 1 0 1932 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1604681595
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1604681595
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1604681595
transform 1 0 1380 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1604681595
transform 1 0 1380 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_19
timestamp 1604681595
transform 1 0 2852 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_11
timestamp 1604681595
transform 1 0 2116 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1604681595
transform 1 0 3036 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1604681595
transform 1 0 2484 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_19
timestamp 1604681595
transform 1 0 2852 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_7
timestamp 1604681595
transform 1 0 1748 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_30
timestamp 1604681595
transform 1 0 3864 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_27
timestamp 1604681595
transform 1 0 3588 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_23
timestamp 1604681595
transform 1 0 3220 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
timestamp 1604681595
transform 1 0 3680 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1604681595
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_36
timestamp 1604681595
transform 1 0 4416 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_32
timestamp 1604681595
transform 1 0 4048 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1604681595
transform 1 0 4232 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1604681595
transform 1 0 4048 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4600 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1604681595
transform 1 0 4232 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_59_43
timestamp 1604681595
transform 1 0 5060 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_47
timestamp 1604681595
transform 1 0 5428 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 5244 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_59
timestamp 1604681595
transform 1 0 6532 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_57
timestamp 1604681595
transform 1 0 6348 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__D
timestamp 1604681595
transform 1 0 6164 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 6532 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1604681595
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 6808 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_47
timestamp 1604681595
transform 1 0 5428 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_
timestamp 1604681595
transform 1 0 6808 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1604681595
transform 1 0 8096 0 -1 35360
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1604681595
transform 1 0 8740 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
timestamp 1604681595
transform 1 0 9108 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__CLK
timestamp 1604681595
transform 1 0 7360 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_81
timestamp 1604681595
transform 1 0 8556 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_85
timestamp 1604681595
transform 1 0 8924 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_66
timestamp 1604681595
transform 1 0 7176 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_70
timestamp 1604681595
transform 1 0 7544 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_60_81
timestamp 1604681595
transform 1 0 8556 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_96
timestamp 1604681595
transform 1 0 9936 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_89
timestamp 1604681595
transform 1 0 9292 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_89
timestamp 1604681595
transform 1 0 9292 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 10120 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9568 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1604681595
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _51_
timestamp 1604681595
transform 1 0 9660 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_60_100
timestamp 1604681595
transform 1 0 10304 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10856 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9752 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_60_115
timestamp 1604681595
transform 1 0 11684 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_117
timestamp 1604681595
transform 1 0 11868 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_113
timestamp 1604681595
transform 1 0 11500 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 12052 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12052 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11684 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_125
timestamp 1604681595
transform 1 0 12604 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_121
timestamp 1604681595
transform 1 0 12236 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_121
timestamp 1604681595
transform 1 0 12236 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12972 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12420 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1604681595
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13156 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_60_140
timestamp 1604681595
transform 1 0 13984 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_152
timestamp 1604681595
transform 1 0 15088 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_148
timestamp 1604681595
transform 1 0 14720 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_146
timestamp 1604681595
transform 1 0 14536 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_142
timestamp 1604681595
transform 1 0 14168 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14536 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 14904 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14720 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14352 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 14904 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 16836 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1604681595
transform 1 0 15180 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_2.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 16836 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_169
timestamp 1604681595
transform 1 0 16652 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_173
timestamp 1604681595
transform 1 0 17020 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_163
timestamp 1604681595
transform 1 0 16100 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_175
timestamp 1604681595
transform 1 0 17204 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_179
timestamp 1604681595
transform 1 0 17572 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17388 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1604681595
transform 1 0 17940 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _57_
timestamp 1604681595
transform 1 0 17940 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_186
timestamp 1604681595
transform 1 0 18216 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18400 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_190
timestamp 1604681595
transform 1 0 18584 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_193
timestamp 1604681595
transform 1 0 18860 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 19964 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_215
timestamp 1604681595
transform 1 0 20884 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_213
timestamp 1604681595
transform 1 0 20700 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_209
timestamp 1604681595
transform 1 0 20332 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__CLK
timestamp 1604681595
transform 1 0 21068 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__D
timestamp 1604681595
transform 1 0 20884 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 20516 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1604681595
transform 1 0 20792 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_202
timestamp 1604681595
transform 1 0 19688 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_
timestamp 1604681595
transform 1 0 21068 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1604681595
transform 1 0 21252 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_
timestamp 1604681595
transform 1 0 22356 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__D
timestamp 1604681595
transform 1 0 23000 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
timestamp 1604681595
transform 1 0 21804 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_236
timestamp 1604681595
transform 1 0 22816 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_240
timestamp 1604681595
transform 1 0 23184 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_223
timestamp 1604681595
transform 1 0 21620 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_227
timestamp 1604681595
transform 1 0 21988 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_
timestamp 1604681595
transform 1 0 24196 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1604681595
transform 1 0 23552 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__D
timestamp 1604681595
transform 1 0 24012 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__CLK
timestamp 1604681595
transform 1 0 24288 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_245
timestamp 1604681595
transform 1 0 23644 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1604681595
transform 1 0 24104 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_254
timestamp 1604681595
transform 1 0 24472 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_269
timestamp 1604681595
transform 1 0 25852 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_266
timestamp 1604681595
transform 1 0 25576 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_270
timestamp 1604681595
transform 1 0 25944 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__CLK
timestamp 1604681595
transform 1 0 25668 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_280
timestamp 1604681595
transform 1 0 26864 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_276
timestamp 1604681595
transform 1 0 26496 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__CLK
timestamp 1604681595
transform 1 0 26680 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__D
timestamp 1604681595
transform 1 0 26496 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1604681595
transform 1 0 26404 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_
timestamp 1604681595
transform 1 0 26680 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_
timestamp 1604681595
transform 1 0 27416 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1604681595
transform 1 0 29164 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__CLK
timestamp 1604681595
transform 1 0 28612 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_297
timestamp 1604681595
transform 1 0 28428 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_301
timestamp 1604681595
transform 1 0 28796 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_305
timestamp 1604681595
transform 1 0 29164 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_306
timestamp 1604681595
transform 1 0 29256 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_318
timestamp 1604681595
transform 1 0 30360 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_317
timestamp 1604681595
transform 1 0 30268 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1604681595
transform 1 0 32016 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_330
timestamp 1604681595
transform 1 0 31464 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_342
timestamp 1604681595
transform 1 0 32568 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_329
timestamp 1604681595
transform 1 0 31372 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_335
timestamp 1604681595
transform 1 0 31924 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_337
timestamp 1604681595
transform 1 0 32108 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_349
timestamp 1604681595
transform 1 0 33212 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1604681595
transform 1 0 34776 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1604681595
transform 1 0 35236 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_354
timestamp 1604681595
transform 1 0 33672 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_367
timestamp 1604681595
transform 1 0 34868 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_361
timestamp 1604681595
transform 1 0 34316 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_369
timestamp 1604681595
transform 1 0 35052 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_381
timestamp 1604681595
transform 1 0 36156 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_377
timestamp 1604681595
transform 1 0 35788 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1604681595
transform 1 0 35972 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604681595
transform 1 0 35420 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604681595
transform 1 0 35328 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_388
timestamp 1604681595
transform 1 0 36800 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_389
timestamp 1604681595
transform 1 0 36892 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1604681595
transform 1 0 37076 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1604681595
transform 1 0 36524 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_376
timestamp 1604681595
transform 1 0 35696 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1604681595
transform 1 0 37260 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1604681595
transform -1 0 38824 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1604681595
transform -1 0 38824 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1604681595
transform 1 0 37628 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1604681595
transform 1 0 38364 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_396
timestamp 1604681595
transform 1 0 37536 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_398
timestamp 1604681595
transform 1 0 37720 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_406
timestamp 1604681595
transform 1 0 38456 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1604681595
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1604681595
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1604681595
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1604681595
transform 1 0 4324 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__80__A
timestamp 1604681595
transform 1 0 4876 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_27
timestamp 1604681595
transform 1 0 3588 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_39
timestamp 1604681595
transform 1 0 4692 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_43
timestamp 1604681595
transform 1 0 5060 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 6808 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 5612 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1604681595
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 6164 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__81__A
timestamp 1604681595
transform 1 0 5428 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__82__A
timestamp 1604681595
transform 1 0 6532 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_53
timestamp 1604681595
transform 1 0 5980 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_57
timestamp 1604681595
transform 1 0 6348 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1604681595
transform 1 0 7912 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 7360 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__83__A
timestamp 1604681595
transform 1 0 8464 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_66
timestamp 1604681595
transform 1 0 7176 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_70
timestamp 1604681595
transform 1 0 7544 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_78
timestamp 1604681595
transform 1 0 8280 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_82
timestamp 1604681595
transform 1 0 8648 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_94
timestamp 1604681595
transform 1 0 9752 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_106
timestamp 1604681595
transform 1 0 10856 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _53_
timestamp 1604681595
transform 1 0 13064 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1604681595
transform 1 0 11224 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1604681595
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_1.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1604681595
transform 1 0 11776 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_114
timestamp 1604681595
transform 1 0 11592 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_118
timestamp 1604681595
transform 1 0 11960 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_123
timestamp 1604681595
transform 1 0 12420 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_129
timestamp 1604681595
transform 1 0 12972 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14076 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13892 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13524 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_133
timestamp 1604681595
transform 1 0 13340 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_137
timestamp 1604681595
transform 1 0 13708 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_150
timestamp 1604681595
transform 1 0 14904 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _56_
timestamp 1604681595
transform 1 0 16744 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 15272 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_156
timestamp 1604681595
transform 1 0 15456 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_168
timestamp 1604681595
transform 1 0 16560 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_173
timestamp 1604681595
transform 1 0 17020 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1604681595
transform 1 0 17940 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_181
timestamp 1604681595
transform 1 0 17756 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_184
timestamp 1604681595
transform 1 0 18032 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_196
timestamp 1604681595
transform 1 0 19136 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 21160 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 20792 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_208
timestamp 1604681595
transform 1 0 20240 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_61_216
timestamp 1604681595
transform 1 0 20976 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1604681595
transform 1 0 21344 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1604681595
transform 1 0 22356 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_229
timestamp 1604681595
transform 1 0 22172 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_233
timestamp 1604681595
transform 1 0 22540 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1604681595
transform 1 0 23644 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1604681595
transform 1 0 23552 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
timestamp 1604681595
transform 1 0 24196 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_241
timestamp 1604681595
transform 1 0 23276 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_249
timestamp 1604681595
transform 1 0 24012 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_253
timestamp 1604681595
transform 1 0 24380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_
timestamp 1604681595
transform 1 0 25668 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__D
timestamp 1604681595
transform 1 0 25484 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1604681595
transform 1 0 29164 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_286
timestamp 1604681595
transform 1 0 27416 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_298
timestamp 1604681595
transform 1 0 28520 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_304
timestamp 1604681595
transform 1 0 29072 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_306
timestamp 1604681595
transform 1 0 29256 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_318
timestamp 1604681595
transform 1 0 30360 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_330
timestamp 1604681595
transform 1 0 31464 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_342
timestamp 1604681595
transform 1 0 32568 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1604681595
transform 1 0 34776 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_354
timestamp 1604681595
transform 1 0 33672 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_367
timestamp 1604681595
transform 1 0 34868 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1604681595
transform 1 0 35420 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1604681595
transform 1 0 35972 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_377
timestamp 1604681595
transform 1 0 35788 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_381
timestamp 1604681595
transform 1 0 36156 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1604681595
transform 1 0 37260 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1604681595
transform -1 0 38824 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1604681595
transform 1 0 38364 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1604681595
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1604681595
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1604681595
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1604681595
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_27
timestamp 1604681595
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_32
timestamp 1604681595
transform 1 0 4048 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1604681595
transform 1 0 5428 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1604681595
transform 1 0 6624 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_44
timestamp 1604681595
transform 1 0 5152 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_51
timestamp 1604681595
transform 1 0 5796 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_59
timestamp 1604681595
transform 1 0 6532 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_64
timestamp 1604681595
transform 1 0 6992 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_76
timestamp 1604681595
transform 1 0 8096 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1604681595
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_88
timestamp 1604681595
transform 1 0 9200 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_93
timestamp 1604681595
transform 1 0 9660 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_105
timestamp 1604681595
transform 1 0 10764 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_117
timestamp 1604681595
transform 1 0 11868 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_129
timestamp 1604681595
transform 1 0 12972 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_0.ltile_clb_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14076 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_143
timestamp 1604681595
transform 1 0 14260 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_151
timestamp 1604681595
transform 1 0 14996 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1604681595
transform 1 0 15180 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_154
timestamp 1604681595
transform 1 0 15272 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_166
timestamp 1604681595
transform 1 0 16376 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_178
timestamp 1604681595
transform 1 0 17480 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_190
timestamp 1604681595
transform 1 0 18584 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1604681595
transform 1 0 20792 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_202
timestamp 1604681595
transform 1 0 19688 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_215
timestamp 1604681595
transform 1 0 20884 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1604681595
transform 1 0 22356 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_0.ltile_clb_m_default__fle_3.ltile_clb_fabric_0.ltile_clb_m_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 21344 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_219
timestamp 1604681595
transform 1 0 21252 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_222
timestamp 1604681595
transform 1 0 21528 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_230
timestamp 1604681595
transform 1 0 22264 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_235
timestamp 1604681595
transform 1 0 22724 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_247
timestamp 1604681595
transform 1 0 23828 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_259
timestamp 1604681595
transform 1 0 24932 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1604681595
transform 1 0 26404 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_271
timestamp 1604681595
transform 1 0 26036 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_276
timestamp 1604681595
transform 1 0 26496 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_288
timestamp 1604681595
transform 1 0 27600 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_300
timestamp 1604681595
transform 1 0 28704 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_312
timestamp 1604681595
transform 1 0 29808 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_324
timestamp 1604681595
transform 1 0 30912 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1604681595
transform 1 0 32016 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_337
timestamp 1604681595
transform 1 0 32108 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_349
timestamp 1604681595
transform 1 0 33212 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_361
timestamp 1604681595
transform 1 0 34316 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_373
timestamp 1604681595
transform 1 0 35420 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_385
timestamp 1604681595
transform 1 0 36524 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1604681595
transform -1 0 38824 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1604681595
transform 1 0 37628 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_398
timestamp 1604681595
transform 1 0 37720 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_406
timestamp 1604681595
transform 1 0 38456 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1604681595
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1604681595
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1604681595
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1604681595
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1604681595
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1604681595
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_51
timestamp 1604681595
transform 1 0 5796 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_59
timestamp 1604681595
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_62
timestamp 1604681595
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_74
timestamp 1604681595
transform 1 0 7912 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_86
timestamp 1604681595
transform 1 0 9016 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_98
timestamp 1604681595
transform 1 0 10120 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1604681595
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_110
timestamp 1604681595
transform 1 0 11224 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_123
timestamp 1604681595
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_135
timestamp 1604681595
transform 1 0 13524 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_147
timestamp 1604681595
transform 1 0 14628 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_159
timestamp 1604681595
transform 1 0 15732 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_171
timestamp 1604681595
transform 1 0 16836 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1604681595
transform 1 0 17940 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_184
timestamp 1604681595
transform 1 0 18032 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_196
timestamp 1604681595
transform 1 0 19136 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_208
timestamp 1604681595
transform 1 0 20240 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_220
timestamp 1604681595
transform 1 0 21344 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_232
timestamp 1604681595
transform 1 0 22448 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1604681595
transform 1 0 23552 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_245
timestamp 1604681595
transform 1 0 23644 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_257
timestamp 1604681595
transform 1 0 24748 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_269
timestamp 1604681595
transform 1 0 25852 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1604681595
transform 1 0 26956 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1604681595
transform 1 0 29164 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1604681595
transform 1 0 28060 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_306
timestamp 1604681595
transform 1 0 29256 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_318
timestamp 1604681595
transform 1 0 30360 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_330
timestamp 1604681595
transform 1 0 31464 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_342
timestamp 1604681595
transform 1 0 32568 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1604681595
transform 1 0 34776 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_354
timestamp 1604681595
transform 1 0 33672 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_367
timestamp 1604681595
transform 1 0 34868 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_379
timestamp 1604681595
transform 1 0 35972 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_391
timestamp 1604681595
transform 1 0 37076 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1604681595
transform -1 0 38824 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_403
timestamp 1604681595
transform 1 0 38180 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1604681595
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1604681595
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1604681595
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1604681595
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_27
timestamp 1604681595
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_32
timestamp 1604681595
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1604681595
transform 1 0 6808 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_44
timestamp 1604681595
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_56
timestamp 1604681595
transform 1 0 6256 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_63
timestamp 1604681595
transform 1 0 6900 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_75
timestamp 1604681595
transform 1 0 8004 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_87
timestamp 1604681595
transform 1 0 9108 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1604681595
transform 1 0 9660 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_94
timestamp 1604681595
transform 1 0 9752 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_106
timestamp 1604681595
transform 1 0 10856 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1604681595
transform 1 0 12512 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_118
timestamp 1604681595
transform 1 0 11960 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_125
timestamp 1604681595
transform 1 0 12604 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_137
timestamp 1604681595
transform 1 0 13708 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_149
timestamp 1604681595
transform 1 0 14812 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1604681595
transform 1 0 15364 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_156
timestamp 1604681595
transform 1 0 15456 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_168
timestamp 1604681595
transform 1 0 16560 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1604681595
transform 1 0 18216 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_180
timestamp 1604681595
transform 1 0 17664 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_187
timestamp 1604681595
transform 1 0 18308 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1604681595
transform 1 0 21068 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_199
timestamp 1604681595
transform 1 0 19412 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_211
timestamp 1604681595
transform 1 0 20516 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_218
timestamp 1604681595
transform 1 0 21160 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_230
timestamp 1604681595
transform 1 0 22264 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1604681595
transform 1 0 23920 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_242
timestamp 1604681595
transform 1 0 23368 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_249
timestamp 1604681595
transform 1 0 24012 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_261
timestamp 1604681595
transform 1 0 25116 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1604681595
transform 1 0 26772 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_273
timestamp 1604681595
transform 1 0 26220 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_280
timestamp 1604681595
transform 1 0 26864 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_292
timestamp 1604681595
transform 1 0 27968 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_304
timestamp 1604681595
transform 1 0 29072 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1604681595
transform 1 0 29624 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_311
timestamp 1604681595
transform 1 0 29716 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_323
timestamp 1604681595
transform 1 0 30820 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1604681595
transform 1 0 32476 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_335
timestamp 1604681595
transform 1 0 31924 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_342
timestamp 1604681595
transform 1 0 32568 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_354
timestamp 1604681595
transform 1 0 33672 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_366
timestamp 1604681595
transform 1 0 34776 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1604681595
transform 1 0 35328 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_373
timestamp 1604681595
transform 1 0 35420 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_385
timestamp 1604681595
transform 1 0 36524 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1604681595
transform -1 0 38824 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1604681595
transform 1 0 38180 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_397
timestamp 1604681595
transform 1 0 37628 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_64_404
timestamp 1604681595
transform 1 0 38272 0 -1 37536
box -38 -48 314 592
<< labels >>
rlabel metal2 s 30010 0 30066 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 38290 39520 38346 40000 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 36634 0 36690 480 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 39394 39520 39450 40000 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal2 s 16670 0 16726 480 6 Test_en
port 4 nsew default input
rlabel metal2 s 3330 0 3386 480 6 bottom_width_0_height_0__pin_50_
port 5 nsew default tristate
rlabel metal2 s 9954 0 10010 480 6 bottom_width_0_height_0__pin_51_
port 6 nsew default tristate
rlabel metal3 s 0 20000 480 20120 6 ccff_head
port 7 nsew default input
rlabel metal3 s 39520 10208 40000 10328 6 ccff_tail
port 8 nsew default tristate
rlabel metal2 s 23294 0 23350 480 6 clk
port 9 nsew default input
rlabel metal3 s 0 33328 480 33448 6 left_width_0_height_0__pin_52_
port 10 nsew default input
rlabel metal3 s 0 6672 480 6792 6 prog_clk
port 11 nsew default input
rlabel metal3 s 39520 11432 40000 11552 6 right_width_0_height_0__pin_16_
port 12 nsew default input
rlabel metal3 s 39520 12656 40000 12776 6 right_width_0_height_0__pin_17_
port 13 nsew default input
rlabel metal3 s 39520 13880 40000 14000 6 right_width_0_height_0__pin_18_
port 14 nsew default input
rlabel metal3 s 39520 14968 40000 15088 6 right_width_0_height_0__pin_19_
port 15 nsew default input
rlabel metal3 s 39520 16192 40000 16312 6 right_width_0_height_0__pin_20_
port 16 nsew default input
rlabel metal3 s 39520 17416 40000 17536 6 right_width_0_height_0__pin_21_
port 17 nsew default input
rlabel metal3 s 39520 18640 40000 18760 6 right_width_0_height_0__pin_22_
port 18 nsew default input
rlabel metal3 s 39520 19864 40000 19984 6 right_width_0_height_0__pin_23_
port 19 nsew default input
rlabel metal3 s 39520 21088 40000 21208 6 right_width_0_height_0__pin_24_
port 20 nsew default input
rlabel metal3 s 39520 22312 40000 22432 6 right_width_0_height_0__pin_25_
port 21 nsew default input
rlabel metal3 s 39520 23536 40000 23656 6 right_width_0_height_0__pin_26_
port 22 nsew default input
rlabel metal3 s 39520 24760 40000 24880 6 right_width_0_height_0__pin_27_
port 23 nsew default input
rlabel metal3 s 39520 25984 40000 26104 6 right_width_0_height_0__pin_28_
port 24 nsew default input
rlabel metal3 s 39520 27208 40000 27328 6 right_width_0_height_0__pin_29_
port 25 nsew default input
rlabel metal3 s 39520 28296 40000 28416 6 right_width_0_height_0__pin_30_
port 26 nsew default input
rlabel metal3 s 39520 29520 40000 29640 6 right_width_0_height_0__pin_31_
port 27 nsew default input
rlabel metal3 s 39520 552 40000 672 6 right_width_0_height_0__pin_42_lower
port 28 nsew default tristate
rlabel metal3 s 39520 30744 40000 30864 6 right_width_0_height_0__pin_42_upper
port 29 nsew default tristate
rlabel metal3 s 39520 1640 40000 1760 6 right_width_0_height_0__pin_43_lower
port 30 nsew default tristate
rlabel metal3 s 39520 31968 40000 32088 6 right_width_0_height_0__pin_43_upper
port 31 nsew default tristate
rlabel metal3 s 39520 2864 40000 2984 6 right_width_0_height_0__pin_44_lower
port 32 nsew default tristate
rlabel metal3 s 39520 33192 40000 33312 6 right_width_0_height_0__pin_44_upper
port 33 nsew default tristate
rlabel metal3 s 39520 4088 40000 4208 6 right_width_0_height_0__pin_45_lower
port 34 nsew default tristate
rlabel metal3 s 39520 34416 40000 34536 6 right_width_0_height_0__pin_45_upper
port 35 nsew default tristate
rlabel metal3 s 39520 5312 40000 5432 6 right_width_0_height_0__pin_46_lower
port 36 nsew default tristate
rlabel metal3 s 39520 35640 40000 35760 6 right_width_0_height_0__pin_46_upper
port 37 nsew default tristate
rlabel metal3 s 39520 6536 40000 6656 6 right_width_0_height_0__pin_47_lower
port 38 nsew default tristate
rlabel metal3 s 39520 36864 40000 36984 6 right_width_0_height_0__pin_47_upper
port 39 nsew default tristate
rlabel metal3 s 39520 7760 40000 7880 6 right_width_0_height_0__pin_48_lower
port 40 nsew default tristate
rlabel metal3 s 39520 38088 40000 38208 6 right_width_0_height_0__pin_48_upper
port 41 nsew default tristate
rlabel metal3 s 39520 8984 40000 9104 6 right_width_0_height_0__pin_49_lower
port 42 nsew default tristate
rlabel metal3 s 39520 39312 40000 39432 6 right_width_0_height_0__pin_49_upper
port 43 nsew default tristate
rlabel metal2 s 9402 39520 9458 40000 6 top_width_0_height_0__pin_0_
port 44 nsew default input
rlabel metal2 s 20534 39520 20590 40000 6 top_width_0_height_0__pin_10_
port 45 nsew default input
rlabel metal2 s 21638 39520 21694 40000 6 top_width_0_height_0__pin_11_
port 46 nsew default input
rlabel metal2 s 22742 39520 22798 40000 6 top_width_0_height_0__pin_12_
port 47 nsew default input
rlabel metal2 s 23846 39520 23902 40000 6 top_width_0_height_0__pin_13_
port 48 nsew default input
rlabel metal2 s 24950 39520 25006 40000 6 top_width_0_height_0__pin_14_
port 49 nsew default input
rlabel metal2 s 26054 39520 26110 40000 6 top_width_0_height_0__pin_15_
port 50 nsew default input
rlabel metal2 s 10506 39520 10562 40000 6 top_width_0_height_0__pin_1_
port 51 nsew default input
rlabel metal2 s 11610 39520 11666 40000 6 top_width_0_height_0__pin_2_
port 52 nsew default input
rlabel metal2 s 27250 39520 27306 40000 6 top_width_0_height_0__pin_32_
port 53 nsew default input
rlabel metal2 s 28354 39520 28410 40000 6 top_width_0_height_0__pin_33_
port 54 nsew default input
rlabel metal2 s 29458 39520 29514 40000 6 top_width_0_height_0__pin_34_lower
port 55 nsew default tristate
rlabel metal2 s 570 39520 626 40000 6 top_width_0_height_0__pin_34_upper
port 56 nsew default tristate
rlabel metal2 s 30562 39520 30618 40000 6 top_width_0_height_0__pin_35_lower
port 57 nsew default tristate
rlabel metal2 s 1674 39520 1730 40000 6 top_width_0_height_0__pin_35_upper
port 58 nsew default tristate
rlabel metal2 s 31666 39520 31722 40000 6 top_width_0_height_0__pin_36_lower
port 59 nsew default tristate
rlabel metal2 s 2778 39520 2834 40000 6 top_width_0_height_0__pin_36_upper
port 60 nsew default tristate
rlabel metal2 s 32770 39520 32826 40000 6 top_width_0_height_0__pin_37_lower
port 61 nsew default tristate
rlabel metal2 s 3882 39520 3938 40000 6 top_width_0_height_0__pin_37_upper
port 62 nsew default tristate
rlabel metal2 s 33874 39520 33930 40000 6 top_width_0_height_0__pin_38_lower
port 63 nsew default tristate
rlabel metal2 s 4986 39520 5042 40000 6 top_width_0_height_0__pin_38_upper
port 64 nsew default tristate
rlabel metal2 s 34978 39520 35034 40000 6 top_width_0_height_0__pin_39_lower
port 65 nsew default tristate
rlabel metal2 s 6090 39520 6146 40000 6 top_width_0_height_0__pin_39_upper
port 66 nsew default tristate
rlabel metal2 s 12714 39520 12770 40000 6 top_width_0_height_0__pin_3_
port 67 nsew default input
rlabel metal2 s 36082 39520 36138 40000 6 top_width_0_height_0__pin_40_lower
port 68 nsew default tristate
rlabel metal2 s 7194 39520 7250 40000 6 top_width_0_height_0__pin_40_upper
port 69 nsew default tristate
rlabel metal2 s 37186 39520 37242 40000 6 top_width_0_height_0__pin_41_lower
port 70 nsew default tristate
rlabel metal2 s 8298 39520 8354 40000 6 top_width_0_height_0__pin_41_upper
port 71 nsew default tristate
rlabel metal2 s 13910 39520 13966 40000 6 top_width_0_height_0__pin_4_
port 72 nsew default input
rlabel metal2 s 15014 39520 15070 40000 6 top_width_0_height_0__pin_5_
port 73 nsew default input
rlabel metal2 s 16118 39520 16174 40000 6 top_width_0_height_0__pin_6_
port 74 nsew default input
rlabel metal2 s 17222 39520 17278 40000 6 top_width_0_height_0__pin_7_
port 75 nsew default input
rlabel metal2 s 18326 39520 18382 40000 6 top_width_0_height_0__pin_8_
port 76 nsew default input
rlabel metal2 s 19430 39520 19486 40000 6 top_width_0_height_0__pin_9_
port 77 nsew default input
rlabel metal4 s 4208 2128 4528 37584 6 VPWR
port 78 nsew default input
rlabel metal4 s 19568 2128 19888 37584 6 VGND
port 79 nsew default input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
