magic
tech sky130A
magscale 1 2
timestamp 1605199094
<< locali >>
rect 5549 18751 5583 18921
rect 18061 17187 18095 17289
rect 4169 15351 4203 15657
rect 16037 15419 16071 15657
rect 6561 11611 6595 11781
rect 12265 7259 12299 7429
rect 6929 6103 6963 6341
rect 3433 5015 3467 5253
rect 13277 1411 13311 1921
<< viali >>
rect 7113 20553 7147 20587
rect 8217 20553 8251 20587
rect 17325 20553 17359 20587
rect 20177 20553 20211 20587
rect 5365 20485 5399 20519
rect 10977 20485 11011 20519
rect 11621 20417 11655 20451
rect 13553 20417 13587 20451
rect 13737 20417 13771 20451
rect 15945 20417 15979 20451
rect 16129 20417 16163 20451
rect 18889 20417 18923 20451
rect 1777 20349 1811 20383
rect 2881 20349 2915 20383
rect 4077 20349 4111 20383
rect 5181 20349 5215 20383
rect 6929 20349 6963 20383
rect 8033 20349 8067 20383
rect 9873 20349 9907 20383
rect 17141 20349 17175 20383
rect 18705 20349 18739 20383
rect 19993 20349 20027 20383
rect 13461 20281 13495 20315
rect 1961 20213 1995 20247
rect 3065 20213 3099 20247
rect 4261 20213 4295 20247
rect 10057 20213 10091 20247
rect 11345 20213 11379 20247
rect 11437 20213 11471 20247
rect 13093 20213 13127 20247
rect 15485 20213 15519 20247
rect 15853 20213 15887 20247
rect 18337 20213 18371 20247
rect 18797 20213 18831 20247
rect 8125 20009 8159 20043
rect 17969 20009 18003 20043
rect 19073 20009 19107 20043
rect 19533 20009 19567 20043
rect 1777 19873 1811 19907
rect 2881 19873 2915 19907
rect 4077 19873 4111 19907
rect 5549 19873 5583 19907
rect 7012 19873 7046 19907
rect 9945 19873 9979 19907
rect 12532 19873 12566 19907
rect 15557 19873 15591 19907
rect 17877 19873 17911 19907
rect 19441 19873 19475 19907
rect 5641 19805 5675 19839
rect 5825 19805 5859 19839
rect 6745 19805 6779 19839
rect 9689 19805 9723 19839
rect 12265 19805 12299 19839
rect 15301 19805 15335 19839
rect 18153 19805 18187 19839
rect 19625 19805 19659 19839
rect 1961 19669 1995 19703
rect 3065 19669 3099 19703
rect 4261 19669 4295 19703
rect 5181 19669 5215 19703
rect 11069 19669 11103 19703
rect 13645 19669 13679 19703
rect 16681 19669 16715 19703
rect 17509 19669 17543 19703
rect 6837 19465 6871 19499
rect 19625 19465 19659 19499
rect 5089 19329 5123 19363
rect 7389 19329 7423 19363
rect 9321 19329 9355 19363
rect 10793 19329 10827 19363
rect 16405 19329 16439 19363
rect 18613 19329 18647 19363
rect 20177 19329 20211 19363
rect 1777 19261 1811 19295
rect 2881 19261 2915 19295
rect 4813 19261 4847 19295
rect 9045 19261 9079 19295
rect 12541 19261 12575 19295
rect 13645 19261 13679 19295
rect 16221 19261 16255 19295
rect 7297 19193 7331 19227
rect 10609 19193 10643 19227
rect 13912 19193 13946 19227
rect 16313 19193 16347 19227
rect 18429 19193 18463 19227
rect 18521 19193 18555 19227
rect 20085 19193 20119 19227
rect 1961 19125 1995 19159
rect 3065 19125 3099 19159
rect 7205 19125 7239 19159
rect 8677 19125 8711 19159
rect 9137 19125 9171 19159
rect 10241 19125 10275 19159
rect 10701 19125 10735 19159
rect 12725 19125 12759 19159
rect 15025 19125 15059 19159
rect 15853 19125 15887 19159
rect 18061 19125 18095 19159
rect 19993 19125 20027 19159
rect 5549 18921 5583 18955
rect 7021 18921 7055 18955
rect 8309 18921 8343 18955
rect 11069 18921 11103 18955
rect 13277 18921 13311 18955
rect 15301 18921 15335 18955
rect 15669 18921 15703 18955
rect 19901 18921 19935 18955
rect 1777 18785 1811 18819
rect 2881 18785 2915 18819
rect 4077 18785 4111 18819
rect 5908 18853 5942 18887
rect 18521 18853 18555 18887
rect 8217 18785 8251 18819
rect 9956 18785 9990 18819
rect 12164 18785 12198 18819
rect 14105 18785 14139 18819
rect 15761 18785 15795 18819
rect 16957 18785 16991 18819
rect 18429 18785 18463 18819
rect 19717 18785 19751 18819
rect 5549 18717 5583 18751
rect 5641 18717 5675 18751
rect 8401 18717 8435 18751
rect 9689 18717 9723 18751
rect 11897 18717 11931 18751
rect 15853 18717 15887 18751
rect 18705 18717 18739 18751
rect 1961 18649 1995 18683
rect 14289 18649 14323 18683
rect 3065 18581 3099 18615
rect 4261 18581 4295 18615
rect 7849 18581 7883 18615
rect 17141 18581 17175 18615
rect 18061 18581 18095 18615
rect 6837 18377 6871 18411
rect 15945 18309 15979 18343
rect 18061 18309 18095 18343
rect 5733 18241 5767 18275
rect 7389 18241 7423 18275
rect 11161 18241 11195 18275
rect 13001 18241 13035 18275
rect 14933 18241 14967 18275
rect 16497 18241 16531 18275
rect 18613 18241 18647 18275
rect 20177 18241 20211 18275
rect 1593 18173 1627 18207
rect 2697 18173 2731 18207
rect 5457 18173 5491 18207
rect 7297 18173 7331 18207
rect 8401 18173 8435 18207
rect 10977 18173 11011 18207
rect 2964 18105 2998 18139
rect 8668 18105 8702 18139
rect 11069 18105 11103 18139
rect 12817 18105 12851 18139
rect 12909 18105 12943 18139
rect 14749 18105 14783 18139
rect 16313 18105 16347 18139
rect 19993 18105 20027 18139
rect 20085 18105 20119 18139
rect 1777 18037 1811 18071
rect 4077 18037 4111 18071
rect 7205 18037 7239 18071
rect 9781 18037 9815 18071
rect 10609 18037 10643 18071
rect 12449 18037 12483 18071
rect 14381 18037 14415 18071
rect 14841 18037 14875 18071
rect 16405 18037 16439 18071
rect 18429 18037 18463 18071
rect 18521 18037 18555 18071
rect 19625 18037 19659 18071
rect 7113 17833 7147 17867
rect 10517 17833 10551 17867
rect 12541 17833 12575 17867
rect 15577 17833 15611 17867
rect 2329 17765 2363 17799
rect 5150 17765 5184 17799
rect 7481 17765 7515 17799
rect 12449 17765 12483 17799
rect 19349 17765 19383 17799
rect 2053 17697 2087 17731
rect 10885 17697 10919 17731
rect 10977 17697 11011 17731
rect 14013 17697 14047 17731
rect 15393 17697 15427 17731
rect 16764 17697 16798 17731
rect 19441 17697 19475 17731
rect 4905 17629 4939 17663
rect 7573 17629 7607 17663
rect 7757 17629 7791 17663
rect 11069 17629 11103 17663
rect 12725 17629 12759 17663
rect 14105 17629 14139 17663
rect 14289 17629 14323 17663
rect 16497 17629 16531 17663
rect 19533 17629 19567 17663
rect 18981 17561 19015 17595
rect 6285 17493 6319 17527
rect 12081 17493 12115 17527
rect 13645 17493 13679 17527
rect 17877 17493 17911 17527
rect 8401 17289 8435 17323
rect 15485 17289 15519 17323
rect 18061 17289 18095 17323
rect 19533 17289 19567 17323
rect 10517 17221 10551 17255
rect 7389 17153 7423 17187
rect 9045 17153 9079 17187
rect 11161 17153 11195 17187
rect 12633 17153 12667 17187
rect 14289 17153 14323 17187
rect 17049 17153 17083 17187
rect 18061 17153 18095 17187
rect 18153 17153 18187 17187
rect 1961 17085 1995 17119
rect 3525 17085 3559 17119
rect 3792 17085 3826 17119
rect 5733 17085 5767 17119
rect 12449 17085 12483 17119
rect 14105 17085 14139 17119
rect 15301 17085 15335 17119
rect 20361 17085 20395 17119
rect 2237 17017 2271 17051
rect 7205 17017 7239 17051
rect 8861 17017 8895 17051
rect 10977 17017 11011 17051
rect 18409 17017 18443 17051
rect 20637 17017 20671 17051
rect 4905 16949 4939 16983
rect 6837 16949 6871 16983
rect 7297 16949 7331 16983
rect 8769 16949 8803 16983
rect 10885 16949 10919 16983
rect 13737 16949 13771 16983
rect 14197 16949 14231 16983
rect 16405 16949 16439 16983
rect 16773 16949 16807 16983
rect 16865 16949 16899 16983
rect 2421 16745 2455 16779
rect 4169 16745 4203 16779
rect 8033 16745 8067 16779
rect 8493 16745 8527 16779
rect 9873 16745 9907 16779
rect 13185 16745 13219 16779
rect 13645 16745 13679 16779
rect 14105 16745 14139 16779
rect 15577 16745 15611 16779
rect 16037 16745 16071 16779
rect 18797 16745 18831 16779
rect 19901 16745 19935 16779
rect 1409 16677 1443 16711
rect 4537 16677 4571 16711
rect 15945 16677 15979 16711
rect 17662 16677 17696 16711
rect 2789 16609 2823 16643
rect 4629 16609 4663 16643
rect 5733 16609 5767 16643
rect 6000 16609 6034 16643
rect 8401 16609 8435 16643
rect 9689 16609 9723 16643
rect 10977 16609 11011 16643
rect 11244 16609 11278 16643
rect 13369 16609 13403 16643
rect 14013 16609 14047 16643
rect 19717 16609 19751 16643
rect 2881 16541 2915 16575
rect 3065 16541 3099 16575
rect 4721 16541 4755 16575
rect 8677 16541 8711 16575
rect 14289 16541 14323 16575
rect 16221 16541 16255 16575
rect 17417 16541 17451 16575
rect 7113 16405 7147 16439
rect 12357 16405 12391 16439
rect 3065 16201 3099 16235
rect 4629 16201 4663 16235
rect 6837 16201 6871 16235
rect 9781 16201 9815 16235
rect 16497 16201 16531 16235
rect 20729 16201 20763 16235
rect 14289 16133 14323 16167
rect 1961 16065 1995 16099
rect 2145 16065 2179 16099
rect 3709 16065 3743 16099
rect 5181 16065 5215 16099
rect 7389 16065 7423 16099
rect 11437 16065 11471 16099
rect 1869 15997 1903 16031
rect 3433 15997 3467 16031
rect 3525 15997 3559 16031
rect 8401 15997 8435 16031
rect 8657 15997 8691 16031
rect 12909 15997 12943 16031
rect 13176 15997 13210 16031
rect 15117 15997 15151 16031
rect 18153 15997 18187 16031
rect 19257 15997 19291 16031
rect 20545 15997 20579 16031
rect 4997 15929 5031 15963
rect 7205 15929 7239 15963
rect 11253 15929 11287 15963
rect 15362 15929 15396 15963
rect 19533 15929 19567 15963
rect 1501 15861 1535 15895
rect 5089 15861 5123 15895
rect 7297 15861 7331 15895
rect 10793 15861 10827 15895
rect 11161 15861 11195 15895
rect 18337 15861 18371 15895
rect 1409 15657 1443 15691
rect 2421 15657 2455 15691
rect 4169 15657 4203 15691
rect 6469 15657 6503 15691
rect 6929 15657 6963 15691
rect 8033 15657 8067 15691
rect 8493 15657 8527 15691
rect 9689 15657 9723 15691
rect 10057 15657 10091 15691
rect 11897 15657 11931 15691
rect 11989 15657 12023 15691
rect 13093 15657 13127 15691
rect 16037 15657 16071 15691
rect 16497 15657 16531 15691
rect 16589 15657 16623 15691
rect 17693 15657 17727 15691
rect 19901 15657 19935 15691
rect 2789 15521 2823 15555
rect 2881 15521 2915 15555
rect 2973 15453 3007 15487
rect 4261 15521 4295 15555
rect 4528 15521 4562 15555
rect 6837 15521 6871 15555
rect 8401 15521 8435 15555
rect 10149 15521 10183 15555
rect 13461 15521 13495 15555
rect 13553 15521 13587 15555
rect 7021 15453 7055 15487
rect 8677 15453 8711 15487
rect 10241 15453 10275 15487
rect 12173 15453 12207 15487
rect 13737 15453 13771 15487
rect 18061 15521 18095 15555
rect 19717 15521 19751 15555
rect 16681 15453 16715 15487
rect 18153 15453 18187 15487
rect 18245 15453 18279 15487
rect 5641 15385 5675 15419
rect 11529 15385 11563 15419
rect 16037 15385 16071 15419
rect 4169 15317 4203 15351
rect 16129 15317 16163 15351
rect 10425 15113 10459 15147
rect 11437 15113 11471 15147
rect 20729 15113 20763 15147
rect 1961 15045 1995 15079
rect 2513 14977 2547 15011
rect 9045 14977 9079 15011
rect 19441 14977 19475 15011
rect 3525 14909 3559 14943
rect 6837 14909 6871 14943
rect 11253 14909 11287 14943
rect 13093 14909 13127 14943
rect 15301 14909 15335 14943
rect 19349 14909 19383 14943
rect 20545 14909 20579 14943
rect 2329 14841 2363 14875
rect 3792 14841 3826 14875
rect 7104 14841 7138 14875
rect 9290 14841 9324 14875
rect 13338 14841 13372 14875
rect 15546 14841 15580 14875
rect 2421 14773 2455 14807
rect 4905 14773 4939 14807
rect 5733 14773 5767 14807
rect 8217 14773 8251 14807
rect 14473 14773 14507 14807
rect 16681 14773 16715 14807
rect 18889 14773 18923 14807
rect 19257 14773 19291 14807
rect 2789 14569 2823 14603
rect 7205 14569 7239 14603
rect 8033 14569 8067 14603
rect 9873 14569 9907 14603
rect 12449 14569 12483 14603
rect 13737 14569 13771 14603
rect 1409 14501 1443 14535
rect 8401 14501 8435 14535
rect 13645 14501 13679 14535
rect 15568 14501 15602 14535
rect 19809 14501 19843 14535
rect 2881 14433 2915 14467
rect 4445 14433 4479 14467
rect 6092 14433 6126 14467
rect 9689 14433 9723 14467
rect 11336 14433 11370 14467
rect 15025 14433 15059 14467
rect 15301 14433 15335 14467
rect 18429 14433 18463 14467
rect 19543 14433 19577 14467
rect 3065 14365 3099 14399
rect 4537 14365 4571 14399
rect 4629 14365 4663 14399
rect 5825 14365 5859 14399
rect 8493 14365 8527 14399
rect 8585 14365 8619 14399
rect 11069 14365 11103 14399
rect 13921 14365 13955 14399
rect 14841 14297 14875 14331
rect 2421 14229 2455 14263
rect 4077 14229 4111 14263
rect 13277 14229 13311 14263
rect 16681 14229 16715 14263
rect 18613 14229 18647 14263
rect 1685 14025 1719 14059
rect 4813 14025 4847 14059
rect 18245 14025 18279 14059
rect 11529 13957 11563 13991
rect 14013 13957 14047 13991
rect 2605 13889 2639 13923
rect 5365 13889 5399 13923
rect 7481 13889 7515 13923
rect 8953 13889 8987 13923
rect 10149 13889 10183 13923
rect 13001 13889 13035 13923
rect 14565 13889 14599 13923
rect 16405 13889 16439 13923
rect 16497 13889 16531 13923
rect 18705 13889 18739 13923
rect 18797 13889 18831 13923
rect 1501 13821 1535 13855
rect 2872 13821 2906 13855
rect 5273 13821 5307 13855
rect 6561 13821 6595 13855
rect 14473 13821 14507 13855
rect 16313 13821 16347 13855
rect 20545 13821 20579 13855
rect 8769 13753 8803 13787
rect 10416 13753 10450 13787
rect 14381 13753 14415 13787
rect 18613 13753 18647 13787
rect 3985 13685 4019 13719
rect 5181 13685 5215 13719
rect 6377 13685 6411 13719
rect 6837 13685 6871 13719
rect 7205 13685 7239 13719
rect 7297 13685 7331 13719
rect 8401 13685 8435 13719
rect 8861 13685 8895 13719
rect 12449 13685 12483 13719
rect 12817 13685 12851 13719
rect 12909 13685 12943 13719
rect 15945 13685 15979 13719
rect 20729 13685 20763 13719
rect 2881 13481 2915 13515
rect 5917 13481 5951 13515
rect 7113 13481 7147 13515
rect 7481 13481 7515 13515
rect 8677 13481 8711 13515
rect 9689 13481 9723 13515
rect 11253 13481 11287 13515
rect 12265 13481 12299 13515
rect 15301 13481 15335 13515
rect 15761 13481 15795 13515
rect 10057 13413 10091 13447
rect 12633 13413 12667 13447
rect 14197 13413 14231 13447
rect 19349 13413 19383 13447
rect 2789 13345 2823 13379
rect 4077 13345 4111 13379
rect 6009 13345 6043 13379
rect 8861 13345 8895 13379
rect 10149 13345 10183 13379
rect 13921 13345 13955 13379
rect 15669 13345 15703 13379
rect 17693 13345 17727 13379
rect 19257 13345 19291 13379
rect 1409 13277 1443 13311
rect 3065 13277 3099 13311
rect 4261 13277 4295 13311
rect 6193 13277 6227 13311
rect 7573 13277 7607 13311
rect 7665 13277 7699 13311
rect 10241 13277 10275 13311
rect 12725 13277 12759 13311
rect 12817 13277 12851 13311
rect 15853 13277 15887 13311
rect 17785 13277 17819 13311
rect 17969 13277 18003 13311
rect 19441 13277 19475 13311
rect 2421 13209 2455 13243
rect 5549 13209 5583 13243
rect 17325 13141 17359 13175
rect 18889 13141 18923 13175
rect 2329 12937 2363 12971
rect 4077 12937 4111 12971
rect 4997 12937 5031 12971
rect 6837 12937 6871 12971
rect 8401 12937 8435 12971
rect 9229 12937 9263 12971
rect 10793 12937 10827 12971
rect 12449 12937 12483 12971
rect 14013 12937 14047 12971
rect 15945 12937 15979 12971
rect 14381 12869 14415 12903
rect 2973 12801 3007 12835
rect 5641 12801 5675 12835
rect 7481 12801 7515 12835
rect 9781 12801 9815 12835
rect 11437 12801 11471 12835
rect 12909 12801 12943 12835
rect 13001 12801 13035 12835
rect 14933 12801 14967 12835
rect 16497 12801 16531 12835
rect 18797 12801 18831 12835
rect 3893 12733 3927 12767
rect 8585 12733 8619 12767
rect 14197 12733 14231 12767
rect 14841 12733 14875 12767
rect 16313 12733 16347 12767
rect 2789 12665 2823 12699
rect 9689 12665 9723 12699
rect 11253 12665 11287 12699
rect 12817 12665 12851 12699
rect 14749 12665 14783 12699
rect 16405 12665 16439 12699
rect 19064 12665 19098 12699
rect 2697 12597 2731 12631
rect 5365 12597 5399 12631
rect 5457 12597 5491 12631
rect 7205 12597 7239 12631
rect 7297 12597 7331 12631
rect 9597 12597 9631 12631
rect 11161 12597 11195 12631
rect 20177 12597 20211 12631
rect 2697 12393 2731 12427
rect 5457 12393 5491 12427
rect 7205 12393 7239 12427
rect 12265 12393 12299 12427
rect 13829 12393 13863 12427
rect 15669 12393 15703 12427
rect 19901 12393 19935 12427
rect 10057 12325 10091 12359
rect 13921 12325 13955 12359
rect 15761 12325 15795 12359
rect 2605 12257 2639 12291
rect 4077 12257 4111 12291
rect 8493 12257 8527 12291
rect 17141 12257 17175 12291
rect 17397 12257 17431 12291
rect 19717 12257 19751 12291
rect 2881 12189 2915 12223
rect 5549 12189 5583 12223
rect 5641 12189 5675 12223
rect 7297 12189 7331 12223
rect 7389 12189 7423 12223
rect 10149 12189 10183 12223
rect 10333 12189 10367 12223
rect 12357 12189 12391 12223
rect 12449 12189 12483 12223
rect 14013 12189 14047 12223
rect 15945 12189 15979 12223
rect 2237 12121 2271 12155
rect 6837 12121 6871 12155
rect 9689 12121 9723 12155
rect 13461 12121 13495 12155
rect 5089 12053 5123 12087
rect 8677 12053 8711 12087
rect 11897 12053 11931 12087
rect 15301 12053 15335 12087
rect 18521 12053 18555 12087
rect 3433 11849 3467 11883
rect 4997 11849 5031 11883
rect 7389 11849 7423 11883
rect 12081 11849 12115 11883
rect 14381 11849 14415 11883
rect 16405 11849 16439 11883
rect 19073 11849 19107 11883
rect 1869 11781 1903 11815
rect 6561 11781 6595 11815
rect 11069 11781 11103 11815
rect 2329 11713 2363 11747
rect 2513 11713 2547 11747
rect 4077 11713 4111 11747
rect 5549 11713 5583 11747
rect 7941 11713 7975 11747
rect 9689 11713 9723 11747
rect 13001 11713 13035 11747
rect 17049 11713 17083 11747
rect 18061 11713 18095 11747
rect 19625 11713 19659 11747
rect 20637 11713 20671 11747
rect 9956 11645 9990 11679
rect 12265 11645 12299 11679
rect 15301 11645 15335 11679
rect 19533 11645 19567 11679
rect 2237 11577 2271 11611
rect 3893 11577 3927 11611
rect 5457 11577 5491 11611
rect 6561 11577 6595 11611
rect 13268 11577 13302 11611
rect 16865 11577 16899 11611
rect 3801 11509 3835 11543
rect 5365 11509 5399 11543
rect 7757 11509 7791 11543
rect 7849 11509 7883 11543
rect 15485 11509 15519 11543
rect 16773 11509 16807 11543
rect 19441 11509 19475 11543
rect 2421 11305 2455 11339
rect 2789 11305 2823 11339
rect 8769 11305 8803 11339
rect 13645 11305 13679 11339
rect 14105 11305 14139 11339
rect 16957 11305 16991 11339
rect 18245 11305 18279 11339
rect 2881 11237 2915 11271
rect 4353 11237 4387 11271
rect 7634 11237 7668 11271
rect 10425 11237 10459 11271
rect 12532 11237 12566 11271
rect 19809 11237 19843 11271
rect 4077 11169 4111 11203
rect 5733 11169 5767 11203
rect 7389 11169 7423 11203
rect 15844 11169 15878 11203
rect 18153 11169 18187 11203
rect 19533 11169 19567 11203
rect 1409 11101 1443 11135
rect 2973 11101 3007 11135
rect 5825 11101 5859 11135
rect 6009 11101 6043 11135
rect 12265 11101 12299 11135
rect 14197 11101 14231 11135
rect 14289 11101 14323 11135
rect 15577 11101 15611 11135
rect 18337 11101 18371 11135
rect 5365 11033 5399 11067
rect 11713 11033 11747 11067
rect 13737 10965 13771 10999
rect 17785 10965 17819 10999
rect 5181 10761 5215 10795
rect 8217 10761 8251 10795
rect 13277 10761 13311 10795
rect 18521 10761 18555 10795
rect 4261 10693 4295 10727
rect 14841 10693 14875 10727
rect 5825 10625 5859 10659
rect 10057 10625 10091 10659
rect 13737 10625 13771 10659
rect 13921 10625 13955 10659
rect 15301 10625 15335 10659
rect 15393 10625 15427 10659
rect 16865 10625 16899 10659
rect 17049 10625 17083 10659
rect 1603 10557 1637 10591
rect 2881 10557 2915 10591
rect 3148 10557 3182 10591
rect 5549 10557 5583 10591
rect 6837 10557 6871 10591
rect 9229 10557 9263 10591
rect 10333 10557 10367 10591
rect 11253 10557 11287 10591
rect 16773 10557 16807 10591
rect 18337 10557 18371 10591
rect 19441 10557 19475 10591
rect 1869 10489 1903 10523
rect 7104 10489 7138 10523
rect 9965 10489 9999 10523
rect 15209 10489 15243 10523
rect 19686 10489 19720 10523
rect 5641 10421 5675 10455
rect 9045 10421 9079 10455
rect 9505 10421 9539 10455
rect 9873 10421 9907 10455
rect 10517 10421 10551 10455
rect 11437 10421 11471 10455
rect 13645 10421 13679 10455
rect 16405 10421 16439 10455
rect 20821 10421 20855 10455
rect 2513 10217 2547 10251
rect 6745 10217 6779 10251
rect 8493 10217 8527 10251
rect 12081 10217 12115 10251
rect 15853 10217 15887 10251
rect 18337 10217 18371 10251
rect 19717 10217 19751 10251
rect 7113 10149 7147 10183
rect 14013 10149 14047 10183
rect 2421 10081 2455 10115
rect 4537 10081 4571 10115
rect 4804 10081 4838 10115
rect 8309 10081 8343 10115
rect 9689 10081 9723 10115
rect 9956 10081 9990 10115
rect 12449 10081 12483 10115
rect 14105 10081 14139 10115
rect 15761 10081 15795 10115
rect 16957 10081 16991 10115
rect 17224 10081 17258 10115
rect 19625 10081 19659 10115
rect 2697 10013 2731 10047
rect 7205 10013 7239 10047
rect 7297 10013 7331 10047
rect 12541 10013 12575 10047
rect 12725 10013 12759 10047
rect 14197 10013 14231 10047
rect 16037 10013 16071 10047
rect 19901 10013 19935 10047
rect 5917 9945 5951 9979
rect 13645 9945 13679 9979
rect 2053 9877 2087 9911
rect 11069 9877 11103 9911
rect 15393 9877 15427 9911
rect 19257 9877 19291 9911
rect 6837 9673 6871 9707
rect 5181 9605 5215 9639
rect 9781 9605 9815 9639
rect 13829 9605 13863 9639
rect 2513 9537 2547 9571
rect 4169 9537 4203 9571
rect 5733 9537 5767 9571
rect 7389 9537 7423 9571
rect 10241 9537 10275 9571
rect 10425 9537 10459 9571
rect 15301 9537 15335 9571
rect 15485 9537 15519 9571
rect 16957 9537 16991 9571
rect 2237 9469 2271 9503
rect 4077 9469 4111 9503
rect 5549 9469 5583 9503
rect 8677 9469 8711 9503
rect 12449 9469 12483 9503
rect 12716 9469 12750 9503
rect 16773 9469 16807 9503
rect 18061 9469 18095 9503
rect 19257 9469 19291 9503
rect 19524 9469 19558 9503
rect 7297 9401 7331 9435
rect 10149 9401 10183 9435
rect 16865 9401 16899 9435
rect 1869 9333 1903 9367
rect 2329 9333 2363 9367
rect 3617 9333 3651 9367
rect 3985 9333 4019 9367
rect 5641 9333 5675 9367
rect 7205 9333 7239 9367
rect 8861 9333 8895 9367
rect 11345 9333 11379 9367
rect 14841 9333 14875 9367
rect 15209 9333 15243 9367
rect 16405 9333 16439 9367
rect 18245 9333 18279 9367
rect 20637 9333 20671 9367
rect 3157 9129 3191 9163
rect 14381 9129 14415 9163
rect 15485 9129 15519 9163
rect 17785 9129 17819 9163
rect 4322 9061 4356 9095
rect 7205 9061 7239 9095
rect 10784 9061 10818 9095
rect 2044 8993 2078 9027
rect 6653 8993 6687 9027
rect 7113 8993 7147 9027
rect 8493 8993 8527 9027
rect 12909 8993 12943 9027
rect 13268 8993 13302 9027
rect 15301 8993 15335 9027
rect 16405 8993 16439 9027
rect 16672 8993 16706 9027
rect 18981 8993 19015 9027
rect 1777 8925 1811 8959
rect 4077 8925 4111 8959
rect 7297 8925 7331 8959
rect 10517 8925 10551 8959
rect 13001 8925 13035 8959
rect 19073 8925 19107 8959
rect 19165 8925 19199 8959
rect 6745 8857 6779 8891
rect 5457 8789 5491 8823
rect 6469 8789 6503 8823
rect 8677 8789 8711 8823
rect 11897 8789 11931 8823
rect 12725 8789 12759 8823
rect 18613 8789 18647 8823
rect 2145 8585 2179 8619
rect 6009 8585 6043 8619
rect 10609 8585 10643 8619
rect 12449 8585 12483 8619
rect 16405 8585 16439 8619
rect 18061 8585 18095 8619
rect 7021 8517 7055 8551
rect 12081 8517 12115 8551
rect 15577 8517 15611 8551
rect 2789 8449 2823 8483
rect 4905 8449 4939 8483
rect 5089 8449 5123 8483
rect 7481 8449 7515 8483
rect 7665 8449 7699 8483
rect 13001 8449 13035 8483
rect 14197 8449 14231 8483
rect 17049 8449 17083 8483
rect 18705 8449 18739 8483
rect 20545 8449 20579 8483
rect 20637 8449 20671 8483
rect 2513 8381 2547 8415
rect 4813 8381 4847 8415
rect 6193 8381 6227 8415
rect 9229 8381 9263 8415
rect 12265 8381 12299 8415
rect 12817 8381 12851 8415
rect 14464 8381 14498 8415
rect 16773 8381 16807 8415
rect 2605 8313 2639 8347
rect 7389 8313 7423 8347
rect 9496 8313 9530 8347
rect 12909 8313 12943 8347
rect 16865 8313 16899 8347
rect 20453 8313 20487 8347
rect 4445 8245 4479 8279
rect 18429 8245 18463 8279
rect 18521 8245 18555 8279
rect 20085 8245 20119 8279
rect 1869 8041 1903 8075
rect 2145 8041 2179 8075
rect 6193 8041 6227 8075
rect 7113 8041 7147 8075
rect 7573 8041 7607 8075
rect 9689 8041 9723 8075
rect 17509 8041 17543 8075
rect 19349 8041 19383 8075
rect 5080 7973 5114 8007
rect 11796 7973 11830 8007
rect 15546 7973 15580 8007
rect 18236 7973 18270 8007
rect 2513 7905 2547 7939
rect 4813 7905 4847 7939
rect 7481 7905 7515 7939
rect 8861 7905 8895 7939
rect 10057 7905 10091 7939
rect 13921 7905 13955 7939
rect 15301 7905 15335 7939
rect 17693 7905 17727 7939
rect 17969 7905 18003 7939
rect 2605 7837 2639 7871
rect 2789 7837 2823 7871
rect 7665 7837 7699 7871
rect 10149 7837 10183 7871
rect 10333 7837 10367 7871
rect 11529 7837 11563 7871
rect 14105 7837 14139 7871
rect 8677 7701 8711 7735
rect 12909 7701 12943 7735
rect 16681 7701 16715 7735
rect 1409 7497 1443 7531
rect 2421 7497 2455 7531
rect 4813 7497 4847 7531
rect 9781 7497 9815 7531
rect 10609 7497 10643 7531
rect 14013 7497 14047 7531
rect 20821 7497 20855 7531
rect 3985 7429 4019 7463
rect 12265 7429 12299 7463
rect 12449 7429 12483 7463
rect 1961 7361 1995 7395
rect 5365 7361 5399 7395
rect 7389 7361 7423 7395
rect 11161 7361 11195 7395
rect 1869 7293 1903 7327
rect 2237 7293 2271 7327
rect 2605 7293 2639 7327
rect 5181 7293 5215 7327
rect 8401 7293 8435 7327
rect 11069 7293 11103 7327
rect 12909 7361 12943 7395
rect 13093 7361 13127 7395
rect 14565 7361 14599 7395
rect 15761 7361 15795 7395
rect 18153 7361 18187 7395
rect 19441 7361 19475 7395
rect 19708 7293 19742 7327
rect 1777 7225 1811 7259
rect 2872 7225 2906 7259
rect 7297 7225 7331 7259
rect 8646 7225 8680 7259
rect 12265 7225 12299 7259
rect 14473 7225 14507 7259
rect 16028 7225 16062 7259
rect 5273 7157 5307 7191
rect 6837 7157 6871 7191
rect 7205 7157 7239 7191
rect 10977 7157 11011 7191
rect 12817 7157 12851 7191
rect 14381 7157 14415 7191
rect 17141 7157 17175 7191
rect 2329 6953 2363 6987
rect 2789 6953 2823 6987
rect 8217 6953 8251 6987
rect 12449 6953 12483 6987
rect 14013 6953 14047 6987
rect 14105 6953 14139 6987
rect 5089 6885 5123 6919
rect 2881 6817 2915 6851
rect 5181 6817 5215 6851
rect 6653 6817 6687 6851
rect 10057 6817 10091 6851
rect 12357 6817 12391 6851
rect 16109 6817 16143 6851
rect 19533 6817 19567 6851
rect 2973 6749 3007 6783
rect 5365 6749 5399 6783
rect 6745 6749 6779 6783
rect 6929 6749 6963 6783
rect 8309 6749 8343 6783
rect 8401 6749 8435 6783
rect 10149 6749 10183 6783
rect 10333 6749 10367 6783
rect 12633 6749 12667 6783
rect 14289 6749 14323 6783
rect 15853 6749 15887 6783
rect 18153 6749 18187 6783
rect 19625 6749 19659 6783
rect 19717 6749 19751 6783
rect 4721 6681 4755 6715
rect 9689 6681 9723 6715
rect 11989 6681 12023 6715
rect 2421 6613 2455 6647
rect 6285 6613 6319 6647
rect 7849 6613 7883 6647
rect 13645 6613 13679 6647
rect 17233 6613 17267 6647
rect 19165 6613 19199 6647
rect 5917 6409 5951 6443
rect 8401 6409 8435 6443
rect 10793 6409 10827 6443
rect 13829 6409 13863 6443
rect 18061 6409 18095 6443
rect 2605 6341 2639 6375
rect 6929 6341 6963 6375
rect 2053 6273 2087 6307
rect 2237 6273 2271 6307
rect 4537 6273 4571 6307
rect 2421 6205 2455 6239
rect 3433 6205 3467 6239
rect 4804 6137 4838 6171
rect 15577 6273 15611 6307
rect 16957 6273 16991 6307
rect 18613 6273 18647 6307
rect 19625 6273 19659 6307
rect 7021 6205 7055 6239
rect 7288 6205 7322 6239
rect 9413 6205 9447 6239
rect 12449 6205 12483 6239
rect 15393 6205 15427 6239
rect 18429 6205 18463 6239
rect 18521 6205 18555 6239
rect 9680 6137 9714 6171
rect 12716 6137 12750 6171
rect 15301 6137 15335 6171
rect 1593 6069 1627 6103
rect 1961 6069 1995 6103
rect 3617 6069 3651 6103
rect 6929 6069 6963 6103
rect 14933 6069 14967 6103
rect 20637 6069 20671 6103
rect 1409 5865 1443 5899
rect 4077 5865 4111 5899
rect 8033 5865 8067 5899
rect 10057 5865 10091 5899
rect 10425 5865 10459 5899
rect 14197 5865 14231 5899
rect 15669 5865 15703 5899
rect 15761 5865 15795 5899
rect 18613 5865 18647 5899
rect 7941 5797 7975 5831
rect 19717 5797 19751 5831
rect 1777 5729 1811 5763
rect 2789 5729 2823 5763
rect 5632 5729 5666 5763
rect 12256 5729 12290 5763
rect 17233 5729 17267 5763
rect 17500 5729 17534 5763
rect 19441 5729 19475 5763
rect 1869 5661 1903 5695
rect 2053 5661 2087 5695
rect 2881 5661 2915 5695
rect 2973 5661 3007 5695
rect 5365 5661 5399 5695
rect 8217 5661 8251 5695
rect 10517 5661 10551 5695
rect 10701 5661 10735 5695
rect 11989 5661 12023 5695
rect 15853 5661 15887 5695
rect 2329 5593 2363 5627
rect 2421 5525 2455 5559
rect 6745 5525 6779 5559
rect 7573 5525 7607 5559
rect 13369 5525 13403 5559
rect 15301 5525 15335 5559
rect 14381 5321 14415 5355
rect 20821 5321 20855 5355
rect 3433 5253 3467 5287
rect 9873 5253 9907 5287
rect 1676 5117 1710 5151
rect 4169 5185 4203 5219
rect 4353 5185 4387 5219
rect 5641 5185 5675 5219
rect 6837 5185 6871 5219
rect 8861 5185 8895 5219
rect 10333 5185 10367 5219
rect 10517 5185 10551 5219
rect 12725 5185 12759 5219
rect 16957 5185 16991 5219
rect 18429 5185 18463 5219
rect 8033 5117 8067 5151
rect 12541 5117 12575 5151
rect 14197 5117 14231 5151
rect 15301 5117 15335 5151
rect 19441 5117 19475 5151
rect 19708 5117 19742 5151
rect 3617 5049 3651 5083
rect 4077 5049 4111 5083
rect 5549 5049 5583 5083
rect 16773 5049 16807 5083
rect 2789 4981 2823 5015
rect 3433 4981 3467 5015
rect 3709 4981 3743 5015
rect 5089 4981 5123 5015
rect 5457 4981 5491 5015
rect 10241 4981 10275 5015
rect 15485 4981 15519 5015
rect 16405 4981 16439 5015
rect 16865 4981 16899 5015
rect 2789 4777 2823 4811
rect 2881 4777 2915 4811
rect 4537 4777 4571 4811
rect 4905 4777 4939 4811
rect 5733 4777 5767 4811
rect 14105 4777 14139 4811
rect 16037 4777 16071 4811
rect 19625 4777 19659 4811
rect 19809 4777 19843 4811
rect 3249 4709 3283 4743
rect 3341 4709 3375 4743
rect 12992 4709 13026 4743
rect 17846 4709 17880 4743
rect 1676 4641 1710 4675
rect 4445 4641 4479 4675
rect 5273 4641 5307 4675
rect 7389 4641 7423 4675
rect 7656 4641 7690 4675
rect 10057 4641 10091 4675
rect 11437 4641 11471 4675
rect 12725 4641 12759 4675
rect 16405 4641 16439 4675
rect 16497 4641 16531 4675
rect 3433 4573 3467 4607
rect 4721 4573 4755 4607
rect 5365 4573 5399 4607
rect 5457 4573 5491 4607
rect 10149 4573 10183 4607
rect 10241 4573 10275 4607
rect 11713 4573 11747 4607
rect 16681 4573 16715 4607
rect 17601 4573 17635 4607
rect 4077 4505 4111 4539
rect 8769 4505 8803 4539
rect 3893 4437 3927 4471
rect 9689 4437 9723 4471
rect 18981 4437 19015 4471
rect 2881 4165 2915 4199
rect 4353 4165 4387 4199
rect 18521 4165 18555 4199
rect 5733 4097 5767 4131
rect 11161 4097 11195 4131
rect 13921 4097 13955 4131
rect 14105 4097 14139 4131
rect 15209 4097 15243 4131
rect 19073 4097 19107 4131
rect 1501 4029 1535 4063
rect 2973 4029 3007 4063
rect 4445 4029 4479 4063
rect 7481 4029 7515 4063
rect 9505 4029 9539 4063
rect 10977 4029 11011 4063
rect 15025 4029 15059 4063
rect 18889 4029 18923 4063
rect 20545 4029 20579 4063
rect 1768 3961 1802 3995
rect 3240 3961 3274 3995
rect 4721 3961 4755 3995
rect 5549 3961 5583 3995
rect 7757 3961 7791 3995
rect 18981 3961 19015 3995
rect 5181 3893 5215 3927
rect 5641 3893 5675 3927
rect 9689 3893 9723 3927
rect 10609 3893 10643 3927
rect 11069 3893 11103 3927
rect 12449 3893 12483 3927
rect 13461 3893 13495 3927
rect 13829 3893 13863 3927
rect 16313 3893 16347 3927
rect 20729 3893 20763 3927
rect 2973 3689 3007 3723
rect 3065 3689 3099 3723
rect 6009 3689 6043 3723
rect 6653 3689 6687 3723
rect 7021 3689 7055 3723
rect 8585 3689 8619 3723
rect 12265 3689 12299 3723
rect 13553 3689 13587 3723
rect 13921 3689 13955 3723
rect 1860 3621 1894 3655
rect 7113 3621 7147 3655
rect 10609 3621 10643 3655
rect 14013 3621 14047 3655
rect 18880 3621 18914 3655
rect 1593 3553 1627 3587
rect 3433 3553 3467 3587
rect 3525 3553 3559 3587
rect 4344 3553 4378 3587
rect 5917 3553 5951 3587
rect 10701 3553 10735 3587
rect 12173 3553 12207 3587
rect 15669 3553 15703 3587
rect 15761 3553 15795 3587
rect 17141 3553 17175 3587
rect 3617 3485 3651 3519
rect 6101 3485 6135 3519
rect 7205 3485 7239 3519
rect 10885 3485 10919 3519
rect 12449 3485 12483 3519
rect 14105 3485 14139 3519
rect 15945 3485 15979 3519
rect 17325 3485 17359 3519
rect 18613 3485 18647 3519
rect 10241 3417 10275 3451
rect 11805 3417 11839 3451
rect 5457 3349 5491 3383
rect 5549 3349 5583 3383
rect 15301 3349 15335 3383
rect 19993 3349 20027 3383
rect 2881 3145 2915 3179
rect 6837 3145 6871 3179
rect 10701 3145 10735 3179
rect 12817 3145 12851 3179
rect 14381 3145 14415 3179
rect 2789 3077 2823 3111
rect 5181 3077 5215 3111
rect 5273 3077 5307 3111
rect 19625 3077 19659 3111
rect 3525 3009 3559 3043
rect 5825 3009 5859 3043
rect 6377 3009 6411 3043
rect 7297 3009 7331 3043
rect 7481 3009 7515 3043
rect 13369 3009 13403 3043
rect 15025 3009 15059 3043
rect 16129 3009 16163 3043
rect 18245 3009 18279 3043
rect 1409 2941 1443 2975
rect 3801 2941 3835 2975
rect 4057 2941 4091 2975
rect 5733 2941 5767 2975
rect 6101 2941 6135 2975
rect 7849 2941 7883 2975
rect 9321 2941 9355 2975
rect 9588 2941 9622 2975
rect 14749 2941 14783 2975
rect 15945 2941 15979 2975
rect 18061 2941 18095 2975
rect 19441 2941 19475 2975
rect 20545 2941 20579 2975
rect 1676 2873 1710 2907
rect 3249 2873 3283 2907
rect 7205 2873 7239 2907
rect 7757 2873 7791 2907
rect 8125 2873 8159 2907
rect 13185 2873 13219 2907
rect 14841 2873 14875 2907
rect 3341 2805 3375 2839
rect 5641 2805 5675 2839
rect 13277 2805 13311 2839
rect 20729 2805 20763 2839
rect 2881 2601 2915 2635
rect 3249 2601 3283 2635
rect 3341 2601 3375 2635
rect 5549 2601 5583 2635
rect 5917 2601 5951 2635
rect 6929 2601 6963 2635
rect 7389 2601 7423 2635
rect 8769 2601 8803 2635
rect 10149 2601 10183 2635
rect 10241 2601 10275 2635
rect 12633 2601 12667 2635
rect 20177 2601 20211 2635
rect 4344 2533 4378 2567
rect 7297 2533 7331 2567
rect 13093 2533 13127 2567
rect 15761 2533 15795 2567
rect 1409 2465 1443 2499
rect 1676 2465 1710 2499
rect 6009 2465 6043 2499
rect 6377 2465 6411 2499
rect 8125 2465 8159 2499
rect 8585 2465 8619 2499
rect 11437 2465 11471 2499
rect 13001 2465 13035 2499
rect 14197 2465 14231 2499
rect 15485 2465 15519 2499
rect 16865 2465 16899 2499
rect 18705 2465 18739 2499
rect 19993 2465 20027 2499
rect 3525 2397 3559 2431
rect 6193 2397 6227 2431
rect 7481 2397 7515 2431
rect 8217 2397 8251 2431
rect 8309 2397 8343 2431
rect 10425 2397 10459 2431
rect 13277 2397 13311 2431
rect 17049 2397 17083 2431
rect 18889 2397 18923 2431
rect 7757 2329 7791 2363
rect 9781 2329 9815 2363
rect 11621 2329 11655 2363
rect 2789 2261 2823 2295
rect 5457 2261 5491 2295
rect 6561 2261 6595 2295
rect 14381 2261 14415 2295
rect 13277 1921 13311 1955
rect 13277 1377 13311 1411
<< metal1 >>
rect 3510 21292 3516 21344
rect 3568 21332 3574 21344
rect 9306 21332 9312 21344
rect 3568 21304 9312 21332
rect 3568 21292 3574 21304
rect 9306 21292 9312 21304
rect 9364 21292 9370 21344
rect 3142 21088 3148 21140
rect 3200 21128 3206 21140
rect 7650 21128 7656 21140
rect 3200 21100 7656 21128
rect 3200 21088 3206 21100
rect 7650 21088 7656 21100
rect 7708 21088 7714 21140
rect 4062 20816 4068 20868
rect 4120 20856 4126 20868
rect 8202 20856 8208 20868
rect 4120 20828 8208 20856
rect 4120 20816 4126 20828
rect 8202 20816 8208 20828
rect 8260 20816 8266 20868
rect 1104 20698 21896 20720
rect 1104 20646 4447 20698
rect 4499 20646 4511 20698
rect 4563 20646 4575 20698
rect 4627 20646 4639 20698
rect 4691 20646 11378 20698
rect 11430 20646 11442 20698
rect 11494 20646 11506 20698
rect 11558 20646 11570 20698
rect 11622 20646 18308 20698
rect 18360 20646 18372 20698
rect 18424 20646 18436 20698
rect 18488 20646 18500 20698
rect 18552 20646 21896 20698
rect 1104 20624 21896 20646
rect 3970 20544 3976 20596
rect 4028 20584 4034 20596
rect 7101 20587 7159 20593
rect 7101 20584 7113 20587
rect 4028 20556 7113 20584
rect 4028 20544 4034 20556
rect 7101 20553 7113 20556
rect 7147 20553 7159 20587
rect 8202 20584 8208 20596
rect 8163 20556 8208 20584
rect 7101 20547 7159 20553
rect 8202 20544 8208 20556
rect 8260 20544 8266 20596
rect 17313 20587 17371 20593
rect 17313 20553 17325 20587
rect 17359 20584 17371 20587
rect 18046 20584 18052 20596
rect 17359 20556 18052 20584
rect 17359 20553 17371 20556
rect 17313 20547 17371 20553
rect 18046 20544 18052 20556
rect 18104 20544 18110 20596
rect 20162 20584 20168 20596
rect 20123 20556 20168 20584
rect 20162 20544 20168 20556
rect 20220 20544 20226 20596
rect 4062 20476 4068 20528
rect 4120 20516 4126 20528
rect 5353 20519 5411 20525
rect 5353 20516 5365 20519
rect 4120 20488 5365 20516
rect 4120 20476 4126 20488
rect 5353 20485 5365 20488
rect 5399 20485 5411 20519
rect 5353 20479 5411 20485
rect 10965 20519 11023 20525
rect 10965 20485 10977 20519
rect 11011 20516 11023 20519
rect 11011 20488 13584 20516
rect 11011 20485 11023 20488
rect 10965 20479 11023 20485
rect 8202 20448 8208 20460
rect 1780 20420 8208 20448
rect 1780 20389 1808 20420
rect 8202 20408 8208 20420
rect 8260 20408 8266 20460
rect 11609 20451 11667 20457
rect 11609 20417 11621 20451
rect 11655 20448 11667 20451
rect 12526 20448 12532 20460
rect 11655 20420 12532 20448
rect 11655 20417 11667 20420
rect 11609 20411 11667 20417
rect 12526 20408 12532 20420
rect 12584 20408 12590 20460
rect 13556 20457 13584 20488
rect 13630 20476 13636 20528
rect 13688 20516 13694 20528
rect 18138 20516 18144 20528
rect 13688 20488 18144 20516
rect 13688 20476 13694 20488
rect 13541 20451 13599 20457
rect 13541 20417 13553 20451
rect 13587 20417 13599 20451
rect 13541 20411 13599 20417
rect 13725 20451 13783 20457
rect 13725 20417 13737 20451
rect 13771 20448 13783 20451
rect 13906 20448 13912 20460
rect 13771 20420 13912 20448
rect 13771 20417 13783 20420
rect 13725 20411 13783 20417
rect 13906 20408 13912 20420
rect 13964 20408 13970 20460
rect 13998 20408 14004 20460
rect 14056 20448 14062 20460
rect 16132 20457 16160 20488
rect 18138 20476 18144 20488
rect 18196 20476 18202 20528
rect 18230 20476 18236 20528
rect 18288 20516 18294 20528
rect 18288 20488 20024 20516
rect 18288 20476 18294 20488
rect 15933 20451 15991 20457
rect 15933 20448 15945 20451
rect 14056 20420 15945 20448
rect 14056 20408 14062 20420
rect 15933 20417 15945 20420
rect 15979 20417 15991 20451
rect 15933 20411 15991 20417
rect 16117 20451 16175 20457
rect 16117 20417 16129 20451
rect 16163 20417 16175 20451
rect 18874 20448 18880 20460
rect 16117 20411 16175 20417
rect 16224 20420 18276 20448
rect 1765 20383 1823 20389
rect 1765 20349 1777 20383
rect 1811 20349 1823 20383
rect 1765 20343 1823 20349
rect 2869 20383 2927 20389
rect 2869 20349 2881 20383
rect 2915 20380 2927 20383
rect 3786 20380 3792 20392
rect 2915 20352 3792 20380
rect 2915 20349 2927 20352
rect 2869 20343 2927 20349
rect 3786 20340 3792 20352
rect 3844 20340 3850 20392
rect 4065 20383 4123 20389
rect 4065 20349 4077 20383
rect 4111 20349 4123 20383
rect 5166 20380 5172 20392
rect 5127 20352 5172 20380
rect 4065 20343 4123 20349
rect 4080 20312 4108 20343
rect 5166 20340 5172 20352
rect 5224 20340 5230 20392
rect 6917 20383 6975 20389
rect 6917 20349 6929 20383
rect 6963 20380 6975 20383
rect 7190 20380 7196 20392
rect 6963 20352 7196 20380
rect 6963 20349 6975 20352
rect 6917 20343 6975 20349
rect 7190 20340 7196 20352
rect 7248 20340 7254 20392
rect 7558 20340 7564 20392
rect 7616 20380 7622 20392
rect 8021 20383 8079 20389
rect 8021 20380 8033 20383
rect 7616 20352 8033 20380
rect 7616 20340 7622 20352
rect 8021 20349 8033 20352
rect 8067 20349 8079 20383
rect 8021 20343 8079 20349
rect 9861 20383 9919 20389
rect 9861 20349 9873 20383
rect 9907 20380 9919 20383
rect 12618 20380 12624 20392
rect 9907 20352 12624 20380
rect 9907 20349 9919 20352
rect 9861 20343 9919 20349
rect 12618 20340 12624 20352
rect 12676 20340 12682 20392
rect 16224 20380 16252 20420
rect 13372 20352 16252 20380
rect 17129 20383 17187 20389
rect 5442 20312 5448 20324
rect 4080 20284 5448 20312
rect 5442 20272 5448 20284
rect 5500 20272 5506 20324
rect 12158 20272 12164 20324
rect 12216 20312 12222 20324
rect 13372 20312 13400 20352
rect 17129 20349 17141 20383
rect 17175 20380 17187 20383
rect 17218 20380 17224 20392
rect 17175 20352 17224 20380
rect 17175 20349 17187 20352
rect 17129 20343 17187 20349
rect 17218 20340 17224 20352
rect 17276 20340 17282 20392
rect 18248 20380 18276 20420
rect 18432 20420 18880 20448
rect 18432 20380 18460 20420
rect 18874 20408 18880 20420
rect 18932 20408 18938 20460
rect 18248 20352 18460 20380
rect 18693 20383 18751 20389
rect 18693 20349 18705 20383
rect 18739 20380 18751 20383
rect 18782 20380 18788 20392
rect 18739 20352 18788 20380
rect 18739 20349 18751 20352
rect 18693 20343 18751 20349
rect 18782 20340 18788 20352
rect 18840 20340 18846 20392
rect 19996 20389 20024 20488
rect 19981 20383 20039 20389
rect 19981 20349 19993 20383
rect 20027 20349 20039 20383
rect 19981 20343 20039 20349
rect 12216 20284 13400 20312
rect 13449 20315 13507 20321
rect 12216 20272 12222 20284
rect 13449 20281 13461 20315
rect 13495 20312 13507 20315
rect 13495 20284 15516 20312
rect 13495 20281 13507 20284
rect 13449 20275 13507 20281
rect 1946 20244 1952 20256
rect 1907 20216 1952 20244
rect 1946 20204 1952 20216
rect 2004 20204 2010 20256
rect 2866 20204 2872 20256
rect 2924 20244 2930 20256
rect 3053 20247 3111 20253
rect 3053 20244 3065 20247
rect 2924 20216 3065 20244
rect 2924 20204 2930 20216
rect 3053 20213 3065 20216
rect 3099 20213 3111 20247
rect 3053 20207 3111 20213
rect 3326 20204 3332 20256
rect 3384 20244 3390 20256
rect 4249 20247 4307 20253
rect 4249 20244 4261 20247
rect 3384 20216 4261 20244
rect 3384 20204 3390 20216
rect 4249 20213 4261 20216
rect 4295 20213 4307 20247
rect 10042 20244 10048 20256
rect 10003 20216 10048 20244
rect 4249 20207 4307 20213
rect 10042 20204 10048 20216
rect 10100 20204 10106 20256
rect 11330 20244 11336 20256
rect 11291 20216 11336 20244
rect 11330 20204 11336 20216
rect 11388 20204 11394 20256
rect 11425 20247 11483 20253
rect 11425 20213 11437 20247
rect 11471 20244 11483 20247
rect 12434 20244 12440 20256
rect 11471 20216 12440 20244
rect 11471 20213 11483 20216
rect 11425 20207 11483 20213
rect 12434 20204 12440 20216
rect 12492 20204 12498 20256
rect 13081 20247 13139 20253
rect 13081 20213 13093 20247
rect 13127 20244 13139 20247
rect 15194 20244 15200 20256
rect 13127 20216 15200 20244
rect 13127 20213 13139 20216
rect 13081 20207 13139 20213
rect 15194 20204 15200 20216
rect 15252 20204 15258 20256
rect 15488 20253 15516 20284
rect 18046 20272 18052 20324
rect 18104 20312 18110 20324
rect 18104 20284 18828 20312
rect 18104 20272 18110 20284
rect 15473 20247 15531 20253
rect 15473 20213 15485 20247
rect 15519 20213 15531 20247
rect 15838 20244 15844 20256
rect 15799 20216 15844 20244
rect 15473 20207 15531 20213
rect 15838 20204 15844 20216
rect 15896 20204 15902 20256
rect 18325 20247 18383 20253
rect 18325 20213 18337 20247
rect 18371 20244 18383 20247
rect 18598 20244 18604 20256
rect 18371 20216 18604 20244
rect 18371 20213 18383 20216
rect 18325 20207 18383 20213
rect 18598 20204 18604 20216
rect 18656 20204 18662 20256
rect 18800 20253 18828 20284
rect 18785 20247 18843 20253
rect 18785 20213 18797 20247
rect 18831 20213 18843 20247
rect 18785 20207 18843 20213
rect 1104 20154 21896 20176
rect 1104 20102 7912 20154
rect 7964 20102 7976 20154
rect 8028 20102 8040 20154
rect 8092 20102 8104 20154
rect 8156 20102 14843 20154
rect 14895 20102 14907 20154
rect 14959 20102 14971 20154
rect 15023 20102 15035 20154
rect 15087 20102 21896 20154
rect 1104 20080 21896 20102
rect 8113 20043 8171 20049
rect 8113 20009 8125 20043
rect 8159 20040 8171 20043
rect 8159 20012 9996 20040
rect 8159 20009 8171 20012
rect 8113 20003 8171 20009
rect 8128 19972 8156 20003
rect 5828 19944 8156 19972
rect 9968 19972 9996 20012
rect 10042 20000 10048 20052
rect 10100 20040 10106 20052
rect 17862 20040 17868 20052
rect 10100 20012 17868 20040
rect 10100 20000 10106 20012
rect 17862 20000 17868 20012
rect 17920 20000 17926 20052
rect 17957 20043 18015 20049
rect 17957 20009 17969 20043
rect 18003 20040 18015 20043
rect 19061 20043 19119 20049
rect 19061 20040 19073 20043
rect 18003 20012 19073 20040
rect 18003 20009 18015 20012
rect 17957 20003 18015 20009
rect 19061 20009 19073 20012
rect 19107 20009 19119 20043
rect 19061 20003 19119 20009
rect 19150 20000 19156 20052
rect 19208 20040 19214 20052
rect 19521 20043 19579 20049
rect 19521 20040 19533 20043
rect 19208 20012 19533 20040
rect 19208 20000 19214 20012
rect 19521 20009 19533 20012
rect 19567 20009 19579 20043
rect 19521 20003 19579 20009
rect 14366 19972 14372 19984
rect 9968 19944 14372 19972
rect 1762 19904 1768 19916
rect 1723 19876 1768 19904
rect 1762 19864 1768 19876
rect 1820 19864 1826 19916
rect 2869 19907 2927 19913
rect 2869 19873 2881 19907
rect 2915 19873 2927 19907
rect 2869 19867 2927 19873
rect 2884 19768 2912 19867
rect 3234 19864 3240 19916
rect 3292 19904 3298 19916
rect 4065 19907 4123 19913
rect 4065 19904 4077 19907
rect 3292 19876 4077 19904
rect 3292 19864 3298 19876
rect 4065 19873 4077 19876
rect 4111 19873 4123 19907
rect 5534 19904 5540 19916
rect 5495 19876 5540 19904
rect 4065 19867 4123 19873
rect 5534 19864 5540 19876
rect 5592 19864 5598 19916
rect 5626 19836 5632 19848
rect 5587 19808 5632 19836
rect 5626 19796 5632 19808
rect 5684 19796 5690 19848
rect 5828 19845 5856 19944
rect 14366 19932 14372 19944
rect 14424 19932 14430 19984
rect 15654 19932 15660 19984
rect 15712 19972 15718 19984
rect 18230 19972 18236 19984
rect 15712 19944 18236 19972
rect 15712 19932 15718 19944
rect 18230 19932 18236 19944
rect 18288 19932 18294 19984
rect 7000 19907 7058 19913
rect 7000 19873 7012 19907
rect 7046 19904 7058 19907
rect 7374 19904 7380 19916
rect 7046 19876 7380 19904
rect 7046 19873 7058 19876
rect 7000 19867 7058 19873
rect 7374 19864 7380 19876
rect 7432 19864 7438 19916
rect 8570 19864 8576 19916
rect 8628 19904 8634 19916
rect 12526 19913 12532 19916
rect 9933 19907 9991 19913
rect 9933 19904 9945 19907
rect 8628 19876 9945 19904
rect 8628 19864 8634 19876
rect 9933 19873 9945 19876
rect 9979 19873 9991 19907
rect 12520 19904 12532 19913
rect 12439 19876 12532 19904
rect 9933 19867 9991 19873
rect 12520 19867 12532 19876
rect 12584 19904 12590 19916
rect 13630 19904 13636 19916
rect 12584 19876 13636 19904
rect 12526 19864 12532 19867
rect 12584 19864 12590 19876
rect 13630 19864 13636 19876
rect 13688 19864 13694 19916
rect 15378 19864 15384 19916
rect 15436 19904 15442 19916
rect 15545 19907 15603 19913
rect 15545 19904 15557 19907
rect 15436 19876 15557 19904
rect 15436 19864 15442 19876
rect 15545 19873 15557 19876
rect 15591 19873 15603 19907
rect 15545 19867 15603 19873
rect 17865 19907 17923 19913
rect 17865 19873 17877 19907
rect 17911 19904 17923 19907
rect 19334 19904 19340 19916
rect 17911 19876 19340 19904
rect 17911 19873 17923 19876
rect 17865 19867 17923 19873
rect 19334 19864 19340 19876
rect 19392 19864 19398 19916
rect 19429 19907 19487 19913
rect 19429 19873 19441 19907
rect 19475 19904 19487 19907
rect 20070 19904 20076 19916
rect 19475 19876 20076 19904
rect 19475 19873 19487 19876
rect 19429 19867 19487 19873
rect 20070 19864 20076 19876
rect 20128 19864 20134 19916
rect 5813 19839 5871 19845
rect 5813 19805 5825 19839
rect 5859 19805 5871 19839
rect 6730 19836 6736 19848
rect 6691 19808 6736 19836
rect 5813 19799 5871 19805
rect 6730 19796 6736 19808
rect 6788 19796 6794 19848
rect 9674 19836 9680 19848
rect 9635 19808 9680 19836
rect 9674 19796 9680 19808
rect 9732 19796 9738 19848
rect 11882 19796 11888 19848
rect 11940 19836 11946 19848
rect 12253 19839 12311 19845
rect 12253 19836 12265 19839
rect 11940 19808 12265 19836
rect 11940 19796 11946 19808
rect 12253 19805 12265 19808
rect 12299 19805 12311 19839
rect 12253 19799 12311 19805
rect 15289 19839 15347 19845
rect 15289 19805 15301 19839
rect 15335 19805 15347 19839
rect 18138 19836 18144 19848
rect 18099 19808 18144 19836
rect 15289 19799 15347 19805
rect 5718 19768 5724 19780
rect 2884 19740 5724 19768
rect 5718 19728 5724 19740
rect 5776 19728 5782 19780
rect 11330 19728 11336 19780
rect 11388 19768 11394 19780
rect 11974 19768 11980 19780
rect 11388 19740 11980 19768
rect 11388 19728 11394 19740
rect 11974 19728 11980 19740
rect 12032 19728 12038 19780
rect 1949 19703 2007 19709
rect 1949 19669 1961 19703
rect 1995 19700 2007 19703
rect 2774 19700 2780 19712
rect 1995 19672 2780 19700
rect 1995 19669 2007 19672
rect 1949 19663 2007 19669
rect 2774 19660 2780 19672
rect 2832 19660 2838 19712
rect 3050 19700 3056 19712
rect 3011 19672 3056 19700
rect 3050 19660 3056 19672
rect 3108 19660 3114 19712
rect 4154 19660 4160 19712
rect 4212 19700 4218 19712
rect 4249 19703 4307 19709
rect 4249 19700 4261 19703
rect 4212 19672 4261 19700
rect 4212 19660 4218 19672
rect 4249 19669 4261 19672
rect 4295 19669 4307 19703
rect 4249 19663 4307 19669
rect 4798 19660 4804 19712
rect 4856 19700 4862 19712
rect 5169 19703 5227 19709
rect 5169 19700 5181 19703
rect 4856 19672 5181 19700
rect 4856 19660 4862 19672
rect 5169 19669 5181 19672
rect 5215 19669 5227 19703
rect 5169 19663 5227 19669
rect 11057 19703 11115 19709
rect 11057 19669 11069 19703
rect 11103 19700 11115 19703
rect 12158 19700 12164 19712
rect 11103 19672 12164 19700
rect 11103 19669 11115 19672
rect 11057 19663 11115 19669
rect 12158 19660 12164 19672
rect 12216 19660 12222 19712
rect 13633 19703 13691 19709
rect 13633 19669 13645 19703
rect 13679 19700 13691 19703
rect 13906 19700 13912 19712
rect 13679 19672 13912 19700
rect 13679 19669 13691 19672
rect 13633 19663 13691 19669
rect 13906 19660 13912 19672
rect 13964 19660 13970 19712
rect 15304 19700 15332 19799
rect 18138 19796 18144 19808
rect 18196 19796 18202 19848
rect 18874 19796 18880 19848
rect 18932 19836 18938 19848
rect 19613 19839 19671 19845
rect 19613 19836 19625 19839
rect 18932 19808 19625 19836
rect 18932 19796 18938 19808
rect 19613 19805 19625 19808
rect 19659 19836 19671 19839
rect 20162 19836 20168 19848
rect 19659 19808 20168 19836
rect 19659 19805 19671 19808
rect 19613 19799 19671 19805
rect 20162 19796 20168 19808
rect 20220 19796 20226 19848
rect 16390 19700 16396 19712
rect 15304 19672 16396 19700
rect 16390 19660 16396 19672
rect 16448 19660 16454 19712
rect 16666 19700 16672 19712
rect 16627 19672 16672 19700
rect 16666 19660 16672 19672
rect 16724 19660 16730 19712
rect 16758 19660 16764 19712
rect 16816 19700 16822 19712
rect 17497 19703 17555 19709
rect 17497 19700 17509 19703
rect 16816 19672 17509 19700
rect 16816 19660 16822 19672
rect 17497 19669 17509 19672
rect 17543 19669 17555 19703
rect 17497 19663 17555 19669
rect 1104 19610 21896 19632
rect 1104 19558 4447 19610
rect 4499 19558 4511 19610
rect 4563 19558 4575 19610
rect 4627 19558 4639 19610
rect 4691 19558 11378 19610
rect 11430 19558 11442 19610
rect 11494 19558 11506 19610
rect 11558 19558 11570 19610
rect 11622 19558 18308 19610
rect 18360 19558 18372 19610
rect 18424 19558 18436 19610
rect 18488 19558 18500 19610
rect 18552 19558 21896 19610
rect 1104 19536 21896 19558
rect 5534 19456 5540 19508
rect 5592 19496 5598 19508
rect 6825 19499 6883 19505
rect 6825 19496 6837 19499
rect 5592 19468 6837 19496
rect 5592 19456 5598 19468
rect 6825 19465 6837 19468
rect 6871 19465 6883 19499
rect 6825 19459 6883 19465
rect 19334 19456 19340 19508
rect 19392 19496 19398 19508
rect 19613 19499 19671 19505
rect 19613 19496 19625 19499
rect 19392 19468 19625 19496
rect 19392 19456 19398 19468
rect 19613 19465 19625 19468
rect 19659 19465 19671 19499
rect 19613 19459 19671 19465
rect 5077 19363 5135 19369
rect 5077 19329 5089 19363
rect 5123 19360 5135 19363
rect 5166 19360 5172 19372
rect 5123 19332 5172 19360
rect 5123 19329 5135 19332
rect 5077 19323 5135 19329
rect 5166 19320 5172 19332
rect 5224 19320 5230 19372
rect 5810 19360 5816 19372
rect 5368 19332 5816 19360
rect 1765 19295 1823 19301
rect 1765 19261 1777 19295
rect 1811 19292 1823 19295
rect 2682 19292 2688 19304
rect 1811 19264 2688 19292
rect 1811 19261 1823 19264
rect 1765 19255 1823 19261
rect 2682 19252 2688 19264
rect 2740 19252 2746 19304
rect 2869 19295 2927 19301
rect 2869 19261 2881 19295
rect 2915 19292 2927 19295
rect 4798 19292 4804 19304
rect 2915 19264 4660 19292
rect 4759 19264 4804 19292
rect 2915 19261 2927 19264
rect 2869 19255 2927 19261
rect 3510 19224 3516 19236
rect 1964 19196 3516 19224
rect 1964 19165 1992 19196
rect 3510 19184 3516 19196
rect 3568 19184 3574 19236
rect 4632 19224 4660 19264
rect 4798 19252 4804 19264
rect 4856 19252 4862 19304
rect 5368 19224 5396 19332
rect 5810 19320 5816 19332
rect 5868 19320 5874 19372
rect 7374 19360 7380 19372
rect 7335 19332 7380 19360
rect 7374 19320 7380 19332
rect 7432 19320 7438 19372
rect 9309 19363 9367 19369
rect 9309 19329 9321 19363
rect 9355 19360 9367 19363
rect 10778 19360 10784 19372
rect 9355 19332 10784 19360
rect 9355 19329 9367 19332
rect 9309 19323 9367 19329
rect 10778 19320 10784 19332
rect 10836 19320 10842 19372
rect 15378 19320 15384 19372
rect 15436 19360 15442 19372
rect 16393 19363 16451 19369
rect 16393 19360 16405 19363
rect 15436 19332 16405 19360
rect 15436 19320 15442 19332
rect 16393 19329 16405 19332
rect 16439 19329 16451 19363
rect 16393 19323 16451 19329
rect 18138 19320 18144 19372
rect 18196 19360 18202 19372
rect 18601 19363 18659 19369
rect 18601 19360 18613 19363
rect 18196 19332 18613 19360
rect 18196 19320 18202 19332
rect 18601 19329 18613 19332
rect 18647 19329 18659 19363
rect 20162 19360 20168 19372
rect 20123 19332 20168 19360
rect 18601 19323 18659 19329
rect 20162 19320 20168 19332
rect 20220 19320 20226 19372
rect 4632 19196 5396 19224
rect 5460 19264 7420 19292
rect 1949 19159 2007 19165
rect 1949 19125 1961 19159
rect 1995 19125 2007 19159
rect 1949 19119 2007 19125
rect 2958 19116 2964 19168
rect 3016 19156 3022 19168
rect 3053 19159 3111 19165
rect 3053 19156 3065 19159
rect 3016 19128 3065 19156
rect 3016 19116 3022 19128
rect 3053 19125 3065 19128
rect 3099 19125 3111 19159
rect 3053 19119 3111 19125
rect 3142 19116 3148 19168
rect 3200 19156 3206 19168
rect 5460 19156 5488 19264
rect 7098 19184 7104 19236
rect 7156 19224 7162 19236
rect 7285 19227 7343 19233
rect 7285 19224 7297 19227
rect 7156 19196 7297 19224
rect 7156 19184 7162 19196
rect 7285 19193 7297 19196
rect 7331 19193 7343 19227
rect 7392 19224 7420 19264
rect 8846 19252 8852 19304
rect 8904 19292 8910 19304
rect 9033 19295 9091 19301
rect 9033 19292 9045 19295
rect 8904 19264 9045 19292
rect 8904 19252 8910 19264
rect 9033 19261 9045 19264
rect 9079 19261 9091 19295
rect 9033 19255 9091 19261
rect 12529 19295 12587 19301
rect 12529 19261 12541 19295
rect 12575 19292 12587 19295
rect 12802 19292 12808 19304
rect 12575 19264 12808 19292
rect 12575 19261 12587 19264
rect 12529 19255 12587 19261
rect 12802 19252 12808 19264
rect 12860 19252 12866 19304
rect 13633 19295 13691 19301
rect 13633 19261 13645 19295
rect 13679 19261 13691 19295
rect 13633 19255 13691 19261
rect 8570 19224 8576 19236
rect 7392 19196 8576 19224
rect 7285 19187 7343 19193
rect 8570 19184 8576 19196
rect 8628 19184 8634 19236
rect 10410 19224 10416 19236
rect 8680 19196 10416 19224
rect 3200 19128 5488 19156
rect 3200 19116 3206 19128
rect 5534 19116 5540 19168
rect 5592 19156 5598 19168
rect 8680 19165 8708 19196
rect 10410 19184 10416 19196
rect 10468 19184 10474 19236
rect 10594 19224 10600 19236
rect 10555 19196 10600 19224
rect 10594 19184 10600 19196
rect 10652 19184 10658 19236
rect 11882 19184 11888 19236
rect 11940 19224 11946 19236
rect 13648 19224 13676 19255
rect 15194 19252 15200 19304
rect 15252 19292 15258 19304
rect 16209 19295 16267 19301
rect 16209 19292 16221 19295
rect 15252 19264 16221 19292
rect 15252 19252 15258 19264
rect 16209 19261 16221 19264
rect 16255 19261 16267 19295
rect 16209 19255 16267 19261
rect 13906 19233 13912 19236
rect 13900 19224 13912 19233
rect 11940 19196 13676 19224
rect 13867 19196 13912 19224
rect 11940 19184 11946 19196
rect 13900 19187 13912 19196
rect 13906 19184 13912 19187
rect 13964 19184 13970 19236
rect 15286 19184 15292 19236
rect 15344 19224 15350 19236
rect 16301 19227 16359 19233
rect 16301 19224 16313 19227
rect 15344 19196 16313 19224
rect 15344 19184 15350 19196
rect 16301 19193 16313 19196
rect 16347 19193 16359 19227
rect 16301 19187 16359 19193
rect 17126 19184 17132 19236
rect 17184 19224 17190 19236
rect 18417 19227 18475 19233
rect 18417 19224 18429 19227
rect 17184 19196 18429 19224
rect 17184 19184 17190 19196
rect 18417 19193 18429 19196
rect 18463 19193 18475 19227
rect 18417 19187 18475 19193
rect 18509 19227 18567 19233
rect 18509 19193 18521 19227
rect 18555 19224 18567 19227
rect 18598 19224 18604 19236
rect 18555 19196 18604 19224
rect 18555 19193 18567 19196
rect 18509 19187 18567 19193
rect 18598 19184 18604 19196
rect 18656 19184 18662 19236
rect 18966 19184 18972 19236
rect 19024 19224 19030 19236
rect 20073 19227 20131 19233
rect 20073 19224 20085 19227
rect 19024 19196 20085 19224
rect 19024 19184 19030 19196
rect 20073 19193 20085 19196
rect 20119 19193 20131 19227
rect 20073 19187 20131 19193
rect 7193 19159 7251 19165
rect 7193 19156 7205 19159
rect 5592 19128 7205 19156
rect 5592 19116 5598 19128
rect 7193 19125 7205 19128
rect 7239 19125 7251 19159
rect 7193 19119 7251 19125
rect 8665 19159 8723 19165
rect 8665 19125 8677 19159
rect 8711 19125 8723 19159
rect 8665 19119 8723 19125
rect 8754 19116 8760 19168
rect 8812 19156 8818 19168
rect 9125 19159 9183 19165
rect 9125 19156 9137 19159
rect 8812 19128 9137 19156
rect 8812 19116 8818 19128
rect 9125 19125 9137 19128
rect 9171 19125 9183 19159
rect 10226 19156 10232 19168
rect 10187 19128 10232 19156
rect 9125 19119 9183 19125
rect 10226 19116 10232 19128
rect 10284 19116 10290 19168
rect 10686 19156 10692 19168
rect 10647 19128 10692 19156
rect 10686 19116 10692 19128
rect 10744 19116 10750 19168
rect 12710 19156 12716 19168
rect 12671 19128 12716 19156
rect 12710 19116 12716 19128
rect 12768 19116 12774 19168
rect 15013 19159 15071 19165
rect 15013 19125 15025 19159
rect 15059 19156 15071 19159
rect 15378 19156 15384 19168
rect 15059 19128 15384 19156
rect 15059 19125 15071 19128
rect 15013 19119 15071 19125
rect 15378 19116 15384 19128
rect 15436 19116 15442 19168
rect 15746 19116 15752 19168
rect 15804 19156 15810 19168
rect 15841 19159 15899 19165
rect 15841 19156 15853 19159
rect 15804 19128 15853 19156
rect 15804 19116 15810 19128
rect 15841 19125 15853 19128
rect 15887 19125 15899 19159
rect 18046 19156 18052 19168
rect 18007 19128 18052 19156
rect 15841 19119 15899 19125
rect 18046 19116 18052 19128
rect 18104 19116 18110 19168
rect 19058 19116 19064 19168
rect 19116 19156 19122 19168
rect 19981 19159 20039 19165
rect 19981 19156 19993 19159
rect 19116 19128 19993 19156
rect 19116 19116 19122 19128
rect 19981 19125 19993 19128
rect 20027 19125 20039 19159
rect 19981 19119 20039 19125
rect 1104 19066 21896 19088
rect 1104 19014 7912 19066
rect 7964 19014 7976 19066
rect 8028 19014 8040 19066
rect 8092 19014 8104 19066
rect 8156 19014 14843 19066
rect 14895 19014 14907 19066
rect 14959 19014 14971 19066
rect 15023 19014 15035 19066
rect 15087 19014 21896 19066
rect 1104 18992 21896 19014
rect 2682 18912 2688 18964
rect 2740 18952 2746 18964
rect 5166 18952 5172 18964
rect 2740 18924 5172 18952
rect 2740 18912 2746 18924
rect 5166 18912 5172 18924
rect 5224 18912 5230 18964
rect 5537 18955 5595 18961
rect 5537 18921 5549 18955
rect 5583 18952 5595 18955
rect 6730 18952 6736 18964
rect 5583 18924 6736 18952
rect 5583 18921 5595 18924
rect 5537 18915 5595 18921
rect 6730 18912 6736 18924
rect 6788 18912 6794 18964
rect 7009 18955 7067 18961
rect 7009 18921 7021 18955
rect 7055 18952 7067 18955
rect 7374 18952 7380 18964
rect 7055 18924 7380 18952
rect 7055 18921 7067 18924
rect 7009 18915 7067 18921
rect 7374 18912 7380 18924
rect 7432 18912 7438 18964
rect 8202 18912 8208 18964
rect 8260 18952 8266 18964
rect 8297 18955 8355 18961
rect 8297 18952 8309 18955
rect 8260 18924 8309 18952
rect 8260 18912 8266 18924
rect 8297 18921 8309 18924
rect 8343 18921 8355 18955
rect 8297 18915 8355 18921
rect 8570 18912 8576 18964
rect 8628 18952 8634 18964
rect 10134 18952 10140 18964
rect 8628 18924 10140 18952
rect 8628 18912 8634 18924
rect 10134 18912 10140 18924
rect 10192 18912 10198 18964
rect 11057 18955 11115 18961
rect 11057 18921 11069 18955
rect 11103 18921 11115 18955
rect 11057 18915 11115 18921
rect 13265 18955 13323 18961
rect 13265 18921 13277 18955
rect 13311 18952 13323 18955
rect 13630 18952 13636 18964
rect 13311 18924 13636 18952
rect 13311 18921 13323 18924
rect 13265 18915 13323 18921
rect 5896 18887 5954 18893
rect 2884 18856 5856 18884
rect 2884 18825 2912 18856
rect 1765 18819 1823 18825
rect 1765 18785 1777 18819
rect 1811 18785 1823 18819
rect 1765 18779 1823 18785
rect 2869 18819 2927 18825
rect 2869 18785 2881 18819
rect 2915 18785 2927 18819
rect 4062 18816 4068 18828
rect 4023 18788 4068 18816
rect 2869 18779 2927 18785
rect 1780 18748 1808 18779
rect 4062 18776 4068 18788
rect 4120 18776 4126 18828
rect 5828 18816 5856 18856
rect 5896 18853 5908 18887
rect 5942 18884 5954 18887
rect 7742 18884 7748 18896
rect 5942 18856 7748 18884
rect 5942 18853 5954 18856
rect 5896 18847 5954 18853
rect 7742 18844 7748 18856
rect 7800 18884 7806 18896
rect 11072 18884 11100 18915
rect 13630 18912 13636 18924
rect 13688 18912 13694 18964
rect 15286 18952 15292 18964
rect 15247 18924 15292 18952
rect 15286 18912 15292 18924
rect 15344 18912 15350 18964
rect 15657 18955 15715 18961
rect 15657 18921 15669 18955
rect 15703 18952 15715 18955
rect 18046 18952 18052 18964
rect 15703 18924 18052 18952
rect 15703 18921 15715 18924
rect 15657 18915 15715 18921
rect 18046 18912 18052 18924
rect 18104 18912 18110 18964
rect 19242 18912 19248 18964
rect 19300 18952 19306 18964
rect 19889 18955 19947 18961
rect 19889 18952 19901 18955
rect 19300 18924 19901 18952
rect 19300 18912 19306 18924
rect 19889 18921 19901 18924
rect 19935 18921 19947 18955
rect 19889 18915 19947 18921
rect 11146 18884 11152 18896
rect 7800 18856 11152 18884
rect 7800 18844 7806 18856
rect 6730 18816 6736 18828
rect 5828 18788 6736 18816
rect 6730 18776 6736 18788
rect 6788 18776 6794 18828
rect 7466 18776 7472 18828
rect 7524 18816 7530 18828
rect 8205 18819 8263 18825
rect 8205 18816 8217 18819
rect 7524 18788 8217 18816
rect 7524 18776 7530 18788
rect 8205 18785 8217 18788
rect 8251 18785 8263 18819
rect 8205 18779 8263 18785
rect 3694 18748 3700 18760
rect 1780 18720 3700 18748
rect 3694 18708 3700 18720
rect 3752 18708 3758 18760
rect 4798 18708 4804 18760
rect 4856 18748 4862 18760
rect 8404 18757 8432 18856
rect 11146 18844 11152 18856
rect 11204 18844 11210 18896
rect 12066 18884 12072 18896
rect 11992 18856 12072 18884
rect 9950 18825 9956 18828
rect 9944 18816 9956 18825
rect 9911 18788 9956 18816
rect 9944 18779 9956 18788
rect 9950 18776 9956 18779
rect 10008 18776 10014 18828
rect 5537 18751 5595 18757
rect 5537 18748 5549 18751
rect 4856 18720 5549 18748
rect 4856 18708 4862 18720
rect 5537 18717 5549 18720
rect 5583 18748 5595 18751
rect 5629 18751 5687 18757
rect 5629 18748 5641 18751
rect 5583 18720 5641 18748
rect 5583 18717 5595 18720
rect 5537 18711 5595 18717
rect 5629 18717 5641 18720
rect 5675 18717 5687 18751
rect 5629 18711 5687 18717
rect 8389 18751 8447 18757
rect 8389 18717 8401 18751
rect 8435 18717 8447 18751
rect 8389 18711 8447 18717
rect 9674 18708 9680 18760
rect 9732 18748 9738 18760
rect 11882 18748 11888 18760
rect 9732 18720 9777 18748
rect 11795 18720 11888 18748
rect 9732 18708 9738 18720
rect 11882 18708 11888 18720
rect 11940 18748 11946 18760
rect 11992 18748 12020 18856
rect 12066 18844 12072 18856
rect 12124 18844 12130 18896
rect 12342 18844 12348 18896
rect 12400 18884 12406 18896
rect 17126 18884 17132 18896
rect 12400 18856 17132 18884
rect 12400 18844 12406 18856
rect 17126 18844 17132 18856
rect 17184 18844 17190 18896
rect 17310 18844 17316 18896
rect 17368 18884 17374 18896
rect 18509 18887 18567 18893
rect 18509 18884 18521 18887
rect 17368 18856 18521 18884
rect 17368 18844 17374 18856
rect 18509 18853 18521 18856
rect 18555 18884 18567 18887
rect 18966 18884 18972 18896
rect 18555 18856 18972 18884
rect 18555 18853 18567 18856
rect 18509 18847 18567 18853
rect 18966 18844 18972 18856
rect 19024 18844 19030 18896
rect 12158 18825 12164 18828
rect 12152 18816 12164 18825
rect 12119 18788 12164 18816
rect 12152 18779 12164 18788
rect 12158 18776 12164 18779
rect 12216 18776 12222 18828
rect 13998 18776 14004 18828
rect 14056 18816 14062 18828
rect 14093 18819 14151 18825
rect 14093 18816 14105 18819
rect 14056 18788 14105 18816
rect 14056 18776 14062 18788
rect 14093 18785 14105 18788
rect 14139 18785 14151 18819
rect 14093 18779 14151 18785
rect 15749 18819 15807 18825
rect 15749 18785 15761 18819
rect 15795 18816 15807 18819
rect 16758 18816 16764 18828
rect 15795 18788 16764 18816
rect 15795 18785 15807 18788
rect 15749 18779 15807 18785
rect 16758 18776 16764 18788
rect 16816 18776 16822 18828
rect 16850 18776 16856 18828
rect 16908 18816 16914 18828
rect 16945 18819 17003 18825
rect 16945 18816 16957 18819
rect 16908 18788 16957 18816
rect 16908 18776 16914 18788
rect 16945 18785 16957 18788
rect 16991 18785 17003 18819
rect 16945 18779 17003 18785
rect 17034 18776 17040 18828
rect 17092 18816 17098 18828
rect 18417 18819 18475 18825
rect 18417 18816 18429 18819
rect 17092 18788 18429 18816
rect 17092 18776 17098 18788
rect 18417 18785 18429 18788
rect 18463 18785 18475 18819
rect 18417 18779 18475 18785
rect 19426 18776 19432 18828
rect 19484 18816 19490 18828
rect 19705 18819 19763 18825
rect 19705 18816 19717 18819
rect 19484 18788 19717 18816
rect 19484 18776 19490 18788
rect 19705 18785 19717 18788
rect 19751 18785 19763 18819
rect 19705 18779 19763 18785
rect 11940 18720 12020 18748
rect 11940 18708 11946 18720
rect 13906 18708 13912 18760
rect 13964 18748 13970 18760
rect 15841 18751 15899 18757
rect 15841 18748 15853 18751
rect 13964 18720 15853 18748
rect 13964 18708 13970 18720
rect 15841 18717 15853 18720
rect 15887 18717 15899 18751
rect 15841 18711 15899 18717
rect 18693 18751 18751 18757
rect 18693 18717 18705 18751
rect 18739 18748 18751 18751
rect 19334 18748 19340 18760
rect 18739 18720 19340 18748
rect 18739 18717 18751 18720
rect 18693 18711 18751 18717
rect 19334 18708 19340 18720
rect 19392 18708 19398 18760
rect 1026 18640 1032 18692
rect 1084 18680 1090 18692
rect 1949 18683 2007 18689
rect 1949 18680 1961 18683
rect 1084 18652 1961 18680
rect 1084 18640 1090 18652
rect 1949 18649 1961 18652
rect 1995 18649 2007 18683
rect 1949 18643 2007 18649
rect 14277 18683 14335 18689
rect 14277 18649 14289 18683
rect 14323 18680 14335 18683
rect 17770 18680 17776 18692
rect 14323 18652 17776 18680
rect 14323 18649 14335 18652
rect 14277 18643 14335 18649
rect 17770 18640 17776 18652
rect 17828 18640 17834 18692
rect 18138 18640 18144 18692
rect 18196 18680 18202 18692
rect 19978 18680 19984 18692
rect 18196 18652 19984 18680
rect 18196 18640 18202 18652
rect 19978 18640 19984 18652
rect 20036 18640 20042 18692
rect 3053 18615 3111 18621
rect 3053 18581 3065 18615
rect 3099 18612 3111 18615
rect 3326 18612 3332 18624
rect 3099 18584 3332 18612
rect 3099 18581 3111 18584
rect 3053 18575 3111 18581
rect 3326 18572 3332 18584
rect 3384 18572 3390 18624
rect 4154 18572 4160 18624
rect 4212 18612 4218 18624
rect 4249 18615 4307 18621
rect 4249 18612 4261 18615
rect 4212 18584 4261 18612
rect 4212 18572 4218 18584
rect 4249 18581 4261 18584
rect 4295 18581 4307 18615
rect 4249 18575 4307 18581
rect 7282 18572 7288 18624
rect 7340 18612 7346 18624
rect 7837 18615 7895 18621
rect 7837 18612 7849 18615
rect 7340 18584 7849 18612
rect 7340 18572 7346 18584
rect 7837 18581 7849 18584
rect 7883 18581 7895 18615
rect 7837 18575 7895 18581
rect 8202 18572 8208 18624
rect 8260 18612 8266 18624
rect 12894 18612 12900 18624
rect 8260 18584 12900 18612
rect 8260 18572 8266 18584
rect 12894 18572 12900 18584
rect 12952 18572 12958 18624
rect 17129 18615 17187 18621
rect 17129 18581 17141 18615
rect 17175 18612 17187 18615
rect 17862 18612 17868 18624
rect 17175 18584 17868 18612
rect 17175 18581 17187 18584
rect 17129 18575 17187 18581
rect 17862 18572 17868 18584
rect 17920 18572 17926 18624
rect 18046 18612 18052 18624
rect 18007 18584 18052 18612
rect 18046 18572 18052 18584
rect 18104 18572 18110 18624
rect 1104 18522 21896 18544
rect 1104 18470 4447 18522
rect 4499 18470 4511 18522
rect 4563 18470 4575 18522
rect 4627 18470 4639 18522
rect 4691 18470 11378 18522
rect 11430 18470 11442 18522
rect 11494 18470 11506 18522
rect 11558 18470 11570 18522
rect 11622 18470 18308 18522
rect 18360 18470 18372 18522
rect 18424 18470 18436 18522
rect 18488 18470 18500 18522
rect 18552 18470 21896 18522
rect 1104 18448 21896 18470
rect 5626 18368 5632 18420
rect 5684 18408 5690 18420
rect 6825 18411 6883 18417
rect 6825 18408 6837 18411
rect 5684 18380 6837 18408
rect 5684 18368 5690 18380
rect 6825 18377 6837 18380
rect 6871 18377 6883 18411
rect 6825 18371 6883 18377
rect 7466 18368 7472 18420
rect 7524 18408 7530 18420
rect 7524 18380 12664 18408
rect 7524 18368 7530 18380
rect 4062 18300 4068 18352
rect 4120 18340 4126 18352
rect 6914 18340 6920 18352
rect 4120 18312 6920 18340
rect 4120 18300 4126 18312
rect 6914 18300 6920 18312
rect 6972 18300 6978 18352
rect 12636 18340 12664 18380
rect 12710 18368 12716 18420
rect 12768 18408 12774 18420
rect 18598 18408 18604 18420
rect 12768 18380 18604 18408
rect 12768 18368 12774 18380
rect 18598 18368 18604 18380
rect 18656 18368 18662 18420
rect 12636 18312 13124 18340
rect 5718 18272 5724 18284
rect 5679 18244 5724 18272
rect 5718 18232 5724 18244
rect 5776 18232 5782 18284
rect 7374 18272 7380 18284
rect 7335 18244 7380 18272
rect 7374 18232 7380 18244
rect 7432 18232 7438 18284
rect 11146 18272 11152 18284
rect 11107 18244 11152 18272
rect 11146 18232 11152 18244
rect 11204 18232 11210 18284
rect 12989 18275 13047 18281
rect 12989 18241 13001 18275
rect 13035 18241 13047 18275
rect 12989 18235 13047 18241
rect 1581 18207 1639 18213
rect 1581 18173 1593 18207
rect 1627 18173 1639 18207
rect 1581 18167 1639 18173
rect 2685 18207 2743 18213
rect 2685 18173 2697 18207
rect 2731 18204 2743 18207
rect 4798 18204 4804 18216
rect 2731 18176 4804 18204
rect 2731 18173 2743 18176
rect 2685 18167 2743 18173
rect 1596 18136 1624 18167
rect 4798 18164 4804 18176
rect 4856 18164 4862 18216
rect 5445 18207 5503 18213
rect 5445 18173 5457 18207
rect 5491 18204 5503 18207
rect 6822 18204 6828 18216
rect 5491 18176 6828 18204
rect 5491 18173 5503 18176
rect 5445 18167 5503 18173
rect 6822 18164 6828 18176
rect 6880 18164 6886 18216
rect 7282 18204 7288 18216
rect 7243 18176 7288 18204
rect 7282 18164 7288 18176
rect 7340 18164 7346 18216
rect 8386 18204 8392 18216
rect 8299 18176 8392 18204
rect 8386 18164 8392 18176
rect 8444 18204 8450 18216
rect 9674 18204 9680 18216
rect 8444 18176 9680 18204
rect 8444 18164 8450 18176
rect 9674 18164 9680 18176
rect 9732 18164 9738 18216
rect 10226 18164 10232 18216
rect 10284 18204 10290 18216
rect 10965 18207 11023 18213
rect 10284 18176 10916 18204
rect 10284 18164 10290 18176
rect 2952 18139 3010 18145
rect 1596 18108 2912 18136
rect 1765 18071 1823 18077
rect 1765 18037 1777 18071
rect 1811 18068 1823 18071
rect 2774 18068 2780 18080
rect 1811 18040 2780 18068
rect 1811 18037 1823 18040
rect 1765 18031 1823 18037
rect 2774 18028 2780 18040
rect 2832 18028 2838 18080
rect 2884 18068 2912 18108
rect 2952 18105 2964 18139
rect 2998 18136 3010 18139
rect 3602 18136 3608 18148
rect 2998 18108 3608 18136
rect 2998 18105 3010 18108
rect 2952 18099 3010 18105
rect 3602 18096 3608 18108
rect 3660 18096 3666 18148
rect 8662 18145 8668 18148
rect 8656 18099 8668 18145
rect 8720 18136 8726 18148
rect 10888 18136 10916 18176
rect 10965 18173 10977 18207
rect 11011 18204 11023 18207
rect 12434 18204 12440 18216
rect 11011 18176 12440 18204
rect 11011 18173 11023 18176
rect 10965 18167 11023 18173
rect 12434 18164 12440 18176
rect 12492 18164 12498 18216
rect 12710 18164 12716 18216
rect 12768 18204 12774 18216
rect 13004 18204 13032 18235
rect 12768 18176 13032 18204
rect 13096 18204 13124 18312
rect 13814 18300 13820 18352
rect 13872 18340 13878 18352
rect 15933 18343 15991 18349
rect 15933 18340 15945 18343
rect 13872 18312 15945 18340
rect 13872 18300 13878 18312
rect 15933 18309 15945 18312
rect 15979 18309 15991 18343
rect 18046 18340 18052 18352
rect 15933 18303 15991 18309
rect 16132 18312 17908 18340
rect 18007 18312 18052 18340
rect 14550 18232 14556 18284
rect 14608 18272 14614 18284
rect 14921 18275 14979 18281
rect 14921 18272 14933 18275
rect 14608 18244 14933 18272
rect 14608 18232 14614 18244
rect 14921 18241 14933 18244
rect 14967 18272 14979 18275
rect 16132 18272 16160 18312
rect 14967 18244 16160 18272
rect 14967 18241 14979 18244
rect 14921 18235 14979 18241
rect 16206 18232 16212 18284
rect 16264 18272 16270 18284
rect 16485 18275 16543 18281
rect 16485 18272 16497 18275
rect 16264 18244 16497 18272
rect 16264 18232 16270 18244
rect 16485 18241 16497 18244
rect 16531 18241 16543 18275
rect 17880 18272 17908 18312
rect 18046 18300 18052 18312
rect 18104 18300 18110 18352
rect 18601 18275 18659 18281
rect 18601 18272 18613 18275
rect 17880 18244 18613 18272
rect 16485 18235 16543 18241
rect 18601 18241 18613 18244
rect 18647 18272 18659 18275
rect 19334 18272 19340 18284
rect 18647 18244 19340 18272
rect 18647 18241 18659 18244
rect 18601 18235 18659 18241
rect 19334 18232 19340 18244
rect 19392 18272 19398 18284
rect 20165 18275 20223 18281
rect 20165 18272 20177 18275
rect 19392 18244 20177 18272
rect 19392 18232 19398 18244
rect 20165 18241 20177 18244
rect 20211 18241 20223 18275
rect 20165 18235 20223 18241
rect 18782 18204 18788 18216
rect 13096 18176 18788 18204
rect 12768 18164 12774 18176
rect 18782 18164 18788 18176
rect 18840 18164 18846 18216
rect 11057 18139 11115 18145
rect 11057 18136 11069 18139
rect 8720 18108 8756 18136
rect 8864 18108 10640 18136
rect 10888 18108 11069 18136
rect 8662 18096 8668 18099
rect 8720 18096 8726 18108
rect 3878 18068 3884 18080
rect 2884 18040 3884 18068
rect 3878 18028 3884 18040
rect 3936 18028 3942 18080
rect 4062 18068 4068 18080
rect 4023 18040 4068 18068
rect 4062 18028 4068 18040
rect 4120 18028 4126 18080
rect 7193 18071 7251 18077
rect 7193 18037 7205 18071
rect 7239 18068 7251 18071
rect 8864 18068 8892 18108
rect 9766 18068 9772 18080
rect 7239 18040 8892 18068
rect 9727 18040 9772 18068
rect 7239 18037 7251 18040
rect 7193 18031 7251 18037
rect 9766 18028 9772 18040
rect 9824 18028 9830 18080
rect 10612 18077 10640 18108
rect 11057 18105 11069 18108
rect 11103 18105 11115 18139
rect 11057 18099 11115 18105
rect 10597 18071 10655 18077
rect 10597 18037 10609 18071
rect 10643 18037 10655 18071
rect 11072 18068 11100 18099
rect 11146 18096 11152 18148
rect 11204 18136 11210 18148
rect 12805 18139 12863 18145
rect 12805 18136 12817 18139
rect 11204 18108 12817 18136
rect 11204 18096 11210 18108
rect 12805 18105 12817 18108
rect 12851 18105 12863 18139
rect 12805 18099 12863 18105
rect 12897 18139 12955 18145
rect 12897 18105 12909 18139
rect 12943 18136 12955 18139
rect 12986 18136 12992 18148
rect 12943 18108 12992 18136
rect 12943 18105 12955 18108
rect 12897 18099 12955 18105
rect 12986 18096 12992 18108
rect 13044 18096 13050 18148
rect 13906 18096 13912 18148
rect 13964 18136 13970 18148
rect 14737 18139 14795 18145
rect 14737 18136 14749 18139
rect 13964 18108 14749 18136
rect 13964 18096 13970 18108
rect 14737 18105 14749 18108
rect 14783 18105 14795 18139
rect 14737 18099 14795 18105
rect 16301 18139 16359 18145
rect 16301 18105 16313 18139
rect 16347 18136 16359 18139
rect 16347 18108 16528 18136
rect 16347 18105 16359 18108
rect 16301 18099 16359 18105
rect 12342 18068 12348 18080
rect 11072 18040 12348 18068
rect 10597 18031 10655 18037
rect 12342 18028 12348 18040
rect 12400 18028 12406 18080
rect 12437 18071 12495 18077
rect 12437 18037 12449 18071
rect 12483 18068 12495 18071
rect 13262 18068 13268 18080
rect 12483 18040 13268 18068
rect 12483 18037 12495 18040
rect 12437 18031 12495 18037
rect 13262 18028 13268 18040
rect 13320 18028 13326 18080
rect 14366 18068 14372 18080
rect 14327 18040 14372 18068
rect 14366 18028 14372 18040
rect 14424 18028 14430 18080
rect 14829 18071 14887 18077
rect 14829 18037 14841 18071
rect 14875 18068 14887 18071
rect 15930 18068 15936 18080
rect 14875 18040 15936 18068
rect 14875 18037 14887 18040
rect 14829 18031 14887 18037
rect 15930 18028 15936 18040
rect 15988 18028 15994 18080
rect 16114 18028 16120 18080
rect 16172 18068 16178 18080
rect 16393 18071 16451 18077
rect 16393 18068 16405 18071
rect 16172 18040 16405 18068
rect 16172 18028 16178 18040
rect 16393 18037 16405 18040
rect 16439 18037 16451 18071
rect 16500 18068 16528 18108
rect 16574 18096 16580 18148
rect 16632 18136 16638 18148
rect 18230 18136 18236 18148
rect 16632 18108 18236 18136
rect 16632 18096 16638 18108
rect 18230 18096 18236 18108
rect 18288 18096 18294 18148
rect 19978 18136 19984 18148
rect 19939 18108 19984 18136
rect 19978 18096 19984 18108
rect 20036 18096 20042 18148
rect 20073 18139 20131 18145
rect 20073 18105 20085 18139
rect 20119 18136 20131 18139
rect 20162 18136 20168 18148
rect 20119 18108 20168 18136
rect 20119 18105 20131 18108
rect 20073 18099 20131 18105
rect 20162 18096 20168 18108
rect 20220 18136 20226 18148
rect 20438 18136 20444 18148
rect 20220 18108 20444 18136
rect 20220 18096 20226 18108
rect 20438 18096 20444 18108
rect 20496 18096 20502 18148
rect 16758 18068 16764 18080
rect 16500 18040 16764 18068
rect 16393 18031 16451 18037
rect 16758 18028 16764 18040
rect 16816 18068 16822 18080
rect 17034 18068 17040 18080
rect 16816 18040 17040 18068
rect 16816 18028 16822 18040
rect 17034 18028 17040 18040
rect 17092 18028 17098 18080
rect 17586 18028 17592 18080
rect 17644 18068 17650 18080
rect 18417 18071 18475 18077
rect 18417 18068 18429 18071
rect 17644 18040 18429 18068
rect 17644 18028 17650 18040
rect 18417 18037 18429 18040
rect 18463 18037 18475 18071
rect 18417 18031 18475 18037
rect 18506 18028 18512 18080
rect 18564 18068 18570 18080
rect 19058 18068 19064 18080
rect 18564 18040 19064 18068
rect 18564 18028 18570 18040
rect 19058 18028 19064 18040
rect 19116 18028 19122 18080
rect 19242 18028 19248 18080
rect 19300 18068 19306 18080
rect 19613 18071 19671 18077
rect 19613 18068 19625 18071
rect 19300 18040 19625 18068
rect 19300 18028 19306 18040
rect 19613 18037 19625 18040
rect 19659 18037 19671 18071
rect 19613 18031 19671 18037
rect 1104 17978 21896 18000
rect 1104 17926 7912 17978
rect 7964 17926 7976 17978
rect 8028 17926 8040 17978
rect 8092 17926 8104 17978
rect 8156 17926 14843 17978
rect 14895 17926 14907 17978
rect 14959 17926 14971 17978
rect 15023 17926 15035 17978
rect 15087 17926 21896 17978
rect 1104 17904 21896 17926
rect 3142 17824 3148 17876
rect 3200 17864 3206 17876
rect 7098 17864 7104 17876
rect 3200 17836 5304 17864
rect 7059 17836 7104 17864
rect 3200 17824 3206 17836
rect 1762 17756 1768 17808
rect 1820 17796 1826 17808
rect 2317 17799 2375 17805
rect 2317 17796 2329 17799
rect 1820 17768 2329 17796
rect 1820 17756 1826 17768
rect 2317 17765 2329 17768
rect 2363 17765 2375 17799
rect 2317 17759 2375 17765
rect 4890 17756 4896 17808
rect 4948 17796 4954 17808
rect 5138 17799 5196 17805
rect 5138 17796 5150 17799
rect 4948 17768 5150 17796
rect 4948 17756 4954 17768
rect 5138 17765 5150 17768
rect 5184 17765 5196 17799
rect 5276 17796 5304 17836
rect 7098 17824 7104 17836
rect 7156 17824 7162 17876
rect 10505 17867 10563 17873
rect 10505 17833 10517 17867
rect 10551 17864 10563 17867
rect 11146 17864 11152 17876
rect 10551 17836 11152 17864
rect 10551 17833 10563 17836
rect 10505 17827 10563 17833
rect 11146 17824 11152 17836
rect 11204 17824 11210 17876
rect 12529 17867 12587 17873
rect 12529 17833 12541 17867
rect 12575 17864 12587 17867
rect 13814 17864 13820 17876
rect 12575 17836 13820 17864
rect 12575 17833 12587 17836
rect 12529 17827 12587 17833
rect 13814 17824 13820 17836
rect 13872 17824 13878 17876
rect 15565 17867 15623 17873
rect 15565 17833 15577 17867
rect 15611 17864 15623 17867
rect 18690 17864 18696 17876
rect 15611 17836 18696 17864
rect 15611 17833 15623 17836
rect 15565 17827 15623 17833
rect 18690 17824 18696 17836
rect 18748 17824 18754 17876
rect 7469 17799 7527 17805
rect 7469 17796 7481 17799
rect 5276 17768 7481 17796
rect 5138 17759 5196 17765
rect 7469 17765 7481 17768
rect 7515 17765 7527 17799
rect 7469 17759 7527 17765
rect 10410 17756 10416 17808
rect 10468 17796 10474 17808
rect 12437 17799 12495 17805
rect 12437 17796 12449 17799
rect 10468 17768 12449 17796
rect 10468 17756 10474 17768
rect 12437 17765 12449 17768
rect 12483 17765 12495 17799
rect 15838 17796 15844 17808
rect 12437 17759 12495 17765
rect 12544 17768 15844 17796
rect 2041 17731 2099 17737
rect 2041 17697 2053 17731
rect 2087 17728 2099 17731
rect 6638 17728 6644 17740
rect 2087 17700 6644 17728
rect 2087 17697 2099 17700
rect 2041 17691 2099 17697
rect 6638 17688 6644 17700
rect 6696 17688 6702 17740
rect 10870 17728 10876 17740
rect 10831 17700 10876 17728
rect 10870 17688 10876 17700
rect 10928 17688 10934 17740
rect 10962 17688 10968 17740
rect 11020 17728 11026 17740
rect 11020 17700 11065 17728
rect 11020 17688 11026 17700
rect 4798 17620 4804 17672
rect 4856 17660 4862 17672
rect 4893 17663 4951 17669
rect 4893 17660 4905 17663
rect 4856 17632 4905 17660
rect 4856 17620 4862 17632
rect 4893 17629 4905 17632
rect 4939 17629 4951 17663
rect 4893 17623 4951 17629
rect 6086 17620 6092 17672
rect 6144 17660 6150 17672
rect 7561 17663 7619 17669
rect 7561 17660 7573 17663
rect 6144 17632 7573 17660
rect 6144 17620 6150 17632
rect 7561 17629 7573 17632
rect 7607 17629 7619 17663
rect 7742 17660 7748 17672
rect 7703 17632 7748 17660
rect 7561 17623 7619 17629
rect 7742 17620 7748 17632
rect 7800 17620 7806 17672
rect 10778 17620 10784 17672
rect 10836 17660 10842 17672
rect 11057 17663 11115 17669
rect 11057 17660 11069 17663
rect 10836 17632 11069 17660
rect 10836 17620 10842 17632
rect 11057 17629 11069 17632
rect 11103 17629 11115 17663
rect 11057 17623 11115 17629
rect 11698 17620 11704 17672
rect 11756 17660 11762 17672
rect 12544 17660 12572 17768
rect 15838 17756 15844 17768
rect 15896 17756 15902 17808
rect 16850 17756 16856 17808
rect 16908 17796 16914 17808
rect 19337 17799 19395 17805
rect 19337 17796 19349 17799
rect 16908 17768 19349 17796
rect 16908 17756 16914 17768
rect 19337 17765 19349 17768
rect 19383 17765 19395 17799
rect 19337 17759 19395 17765
rect 13170 17688 13176 17740
rect 13228 17728 13234 17740
rect 14001 17731 14059 17737
rect 14001 17728 14013 17731
rect 13228 17700 14013 17728
rect 13228 17688 13234 17700
rect 14001 17697 14013 17700
rect 14047 17697 14059 17731
rect 15378 17728 15384 17740
rect 15339 17700 15384 17728
rect 14001 17691 14059 17697
rect 15378 17688 15384 17700
rect 15436 17688 15442 17740
rect 16752 17731 16810 17737
rect 16752 17697 16764 17731
rect 16798 17728 16810 17731
rect 17034 17728 17040 17740
rect 16798 17700 17040 17728
rect 16798 17697 16810 17700
rect 16752 17691 16810 17697
rect 17034 17688 17040 17700
rect 17092 17688 17098 17740
rect 19429 17731 19487 17737
rect 19429 17697 19441 17731
rect 19475 17728 19487 17731
rect 19794 17728 19800 17740
rect 19475 17700 19800 17728
rect 19475 17697 19487 17700
rect 19429 17691 19487 17697
rect 19794 17688 19800 17700
rect 19852 17688 19858 17740
rect 12710 17660 12716 17672
rect 11756 17632 12572 17660
rect 12671 17632 12716 17660
rect 11756 17620 11762 17632
rect 12710 17620 12716 17632
rect 12768 17620 12774 17672
rect 14090 17660 14096 17672
rect 14051 17632 14096 17660
rect 14090 17620 14096 17632
rect 14148 17620 14154 17672
rect 14277 17663 14335 17669
rect 14277 17629 14289 17663
rect 14323 17660 14335 17663
rect 14550 17660 14556 17672
rect 14323 17632 14556 17660
rect 14323 17629 14335 17632
rect 14277 17623 14335 17629
rect 14550 17620 14556 17632
rect 14608 17620 14614 17672
rect 16482 17660 16488 17672
rect 16443 17632 16488 17660
rect 16482 17620 16488 17632
rect 16540 17620 16546 17672
rect 19334 17620 19340 17672
rect 19392 17660 19398 17672
rect 19521 17663 19579 17669
rect 19521 17660 19533 17663
rect 19392 17632 19533 17660
rect 19392 17620 19398 17632
rect 19521 17629 19533 17632
rect 19567 17629 19579 17663
rect 19521 17623 19579 17629
rect 6196 17564 16528 17592
rect 1762 17484 1768 17536
rect 1820 17524 1826 17536
rect 6196 17524 6224 17564
rect 1820 17496 6224 17524
rect 6273 17527 6331 17533
rect 1820 17484 1826 17496
rect 6273 17493 6285 17527
rect 6319 17524 6331 17527
rect 6362 17524 6368 17536
rect 6319 17496 6368 17524
rect 6319 17493 6331 17496
rect 6273 17487 6331 17493
rect 6362 17484 6368 17496
rect 6420 17484 6426 17536
rect 9122 17484 9128 17536
rect 9180 17524 9186 17536
rect 11882 17524 11888 17536
rect 9180 17496 11888 17524
rect 9180 17484 9186 17496
rect 11882 17484 11888 17496
rect 11940 17484 11946 17536
rect 12069 17527 12127 17533
rect 12069 17493 12081 17527
rect 12115 17524 12127 17527
rect 12986 17524 12992 17536
rect 12115 17496 12992 17524
rect 12115 17493 12127 17496
rect 12069 17487 12127 17493
rect 12986 17484 12992 17496
rect 13044 17484 13050 17536
rect 13633 17527 13691 17533
rect 13633 17493 13645 17527
rect 13679 17524 13691 17527
rect 14734 17524 14740 17536
rect 13679 17496 14740 17524
rect 13679 17493 13691 17496
rect 13633 17487 13691 17493
rect 14734 17484 14740 17496
rect 14792 17484 14798 17536
rect 16500 17524 16528 17564
rect 17494 17552 17500 17604
rect 17552 17592 17558 17604
rect 18969 17595 19027 17601
rect 18969 17592 18981 17595
rect 17552 17564 18981 17592
rect 17552 17552 17558 17564
rect 18969 17561 18981 17564
rect 19015 17561 19027 17595
rect 18969 17555 19027 17561
rect 17402 17524 17408 17536
rect 16500 17496 17408 17524
rect 17402 17484 17408 17496
rect 17460 17484 17466 17536
rect 17862 17524 17868 17536
rect 17823 17496 17868 17524
rect 17862 17484 17868 17496
rect 17920 17484 17926 17536
rect 1104 17434 21896 17456
rect 1104 17382 4447 17434
rect 4499 17382 4511 17434
rect 4563 17382 4575 17434
rect 4627 17382 4639 17434
rect 4691 17382 11378 17434
rect 11430 17382 11442 17434
rect 11494 17382 11506 17434
rect 11558 17382 11570 17434
rect 11622 17382 18308 17434
rect 18360 17382 18372 17434
rect 18424 17382 18436 17434
rect 18488 17382 18500 17434
rect 18552 17382 21896 17434
rect 1104 17360 21896 17382
rect 6822 17280 6828 17332
rect 6880 17320 6886 17332
rect 8389 17323 8447 17329
rect 8389 17320 8401 17323
rect 6880 17292 8401 17320
rect 6880 17280 6886 17292
rect 8389 17289 8401 17292
rect 8435 17289 8447 17323
rect 11790 17320 11796 17332
rect 8389 17283 8447 17289
rect 8496 17292 11796 17320
rect 7190 17212 7196 17264
rect 7248 17252 7254 17264
rect 8496 17252 8524 17292
rect 11790 17280 11796 17292
rect 11848 17280 11854 17332
rect 11882 17280 11888 17332
rect 11940 17320 11946 17332
rect 14090 17320 14096 17332
rect 11940 17292 14096 17320
rect 11940 17280 11946 17292
rect 14090 17280 14096 17292
rect 14148 17280 14154 17332
rect 15473 17323 15531 17329
rect 15473 17289 15485 17323
rect 15519 17320 15531 17323
rect 16574 17320 16580 17332
rect 15519 17292 16580 17320
rect 15519 17289 15531 17292
rect 15473 17283 15531 17289
rect 16574 17280 16580 17292
rect 16632 17280 16638 17332
rect 18049 17323 18107 17329
rect 18049 17289 18061 17323
rect 18095 17320 18107 17323
rect 19521 17323 19579 17329
rect 19521 17320 19533 17323
rect 18095 17292 19533 17320
rect 18095 17289 18107 17292
rect 18049 17283 18107 17289
rect 19521 17289 19533 17292
rect 19567 17289 19579 17323
rect 19521 17283 19579 17289
rect 9858 17252 9864 17264
rect 7248 17224 8524 17252
rect 8588 17224 9864 17252
rect 7248 17212 7254 17224
rect 5994 17144 6000 17196
rect 6052 17184 6058 17196
rect 7377 17187 7435 17193
rect 7377 17184 7389 17187
rect 6052 17156 7389 17184
rect 6052 17144 6058 17156
rect 7377 17153 7389 17156
rect 7423 17153 7435 17187
rect 7377 17147 7435 17153
rect 7650 17144 7656 17196
rect 7708 17184 7714 17196
rect 8588 17184 8616 17224
rect 9858 17212 9864 17224
rect 9916 17212 9922 17264
rect 10505 17255 10563 17261
rect 10505 17221 10517 17255
rect 10551 17252 10563 17255
rect 10551 17224 13299 17252
rect 10551 17221 10563 17224
rect 10505 17215 10563 17221
rect 7708 17156 8616 17184
rect 9033 17187 9091 17193
rect 7708 17144 7714 17156
rect 9033 17153 9045 17187
rect 9079 17184 9091 17187
rect 9766 17184 9772 17196
rect 9079 17156 9772 17184
rect 9079 17153 9091 17156
rect 9033 17147 9091 17153
rect 9766 17144 9772 17156
rect 9824 17144 9830 17196
rect 11149 17187 11207 17193
rect 11149 17153 11161 17187
rect 11195 17184 11207 17187
rect 11238 17184 11244 17196
rect 11195 17156 11244 17184
rect 11195 17153 11207 17156
rect 11149 17147 11207 17153
rect 11238 17144 11244 17156
rect 11296 17144 11302 17196
rect 12618 17184 12624 17196
rect 12579 17156 12624 17184
rect 12618 17144 12624 17156
rect 12676 17144 12682 17196
rect 13170 17184 13176 17196
rect 13096 17156 13176 17184
rect 1949 17119 2007 17125
rect 1949 17085 1961 17119
rect 1995 17116 2007 17119
rect 3050 17116 3056 17128
rect 1995 17088 3056 17116
rect 1995 17085 2007 17088
rect 1949 17079 2007 17085
rect 3050 17076 3056 17088
rect 3108 17076 3114 17128
rect 3513 17119 3571 17125
rect 3513 17085 3525 17119
rect 3559 17085 3571 17119
rect 3513 17079 3571 17085
rect 3780 17119 3838 17125
rect 3780 17085 3792 17119
rect 3826 17116 3838 17119
rect 4062 17116 4068 17128
rect 3826 17088 4068 17116
rect 3826 17085 3838 17088
rect 3780 17079 3838 17085
rect 1486 17008 1492 17060
rect 1544 17048 1550 17060
rect 2225 17051 2283 17057
rect 2225 17048 2237 17051
rect 1544 17020 2237 17048
rect 1544 17008 1550 17020
rect 2225 17017 2237 17020
rect 2271 17017 2283 17051
rect 3528 17048 3556 17079
rect 4062 17076 4068 17088
rect 4120 17076 4126 17128
rect 5721 17119 5779 17125
rect 5721 17085 5733 17119
rect 5767 17116 5779 17119
rect 11698 17116 11704 17128
rect 5767 17088 11704 17116
rect 5767 17085 5779 17088
rect 5721 17079 5779 17085
rect 11698 17076 11704 17088
rect 11756 17076 11762 17128
rect 12437 17119 12495 17125
rect 12437 17085 12449 17119
rect 12483 17116 12495 17119
rect 12526 17116 12532 17128
rect 12483 17088 12532 17116
rect 12483 17085 12495 17088
rect 12437 17079 12495 17085
rect 12526 17076 12532 17088
rect 12584 17076 12590 17128
rect 4798 17048 4804 17060
rect 3528 17020 4804 17048
rect 2225 17011 2283 17017
rect 4798 17008 4804 17020
rect 4856 17048 4862 17060
rect 5350 17048 5356 17060
rect 4856 17020 5356 17048
rect 4856 17008 4862 17020
rect 5350 17008 5356 17020
rect 5408 17008 5414 17060
rect 6454 17008 6460 17060
rect 6512 17048 6518 17060
rect 6730 17048 6736 17060
rect 6512 17020 6736 17048
rect 6512 17008 6518 17020
rect 6730 17008 6736 17020
rect 6788 17048 6794 17060
rect 7190 17048 7196 17060
rect 6788 17020 6960 17048
rect 7151 17020 7196 17048
rect 6788 17008 6794 17020
rect 4890 16980 4896 16992
rect 4851 16952 4896 16980
rect 4890 16940 4896 16952
rect 4948 16940 4954 16992
rect 6822 16980 6828 16992
rect 6783 16952 6828 16980
rect 6822 16940 6828 16952
rect 6880 16940 6886 16992
rect 6932 16980 6960 17020
rect 7190 17008 7196 17020
rect 7248 17008 7254 17060
rect 8202 17008 8208 17060
rect 8260 17048 8266 17060
rect 8849 17051 8907 17057
rect 8849 17048 8861 17051
rect 8260 17020 8861 17048
rect 8260 17008 8266 17020
rect 8849 17017 8861 17020
rect 8895 17017 8907 17051
rect 8849 17011 8907 17017
rect 9030 17008 9036 17060
rect 9088 17048 9094 17060
rect 10965 17051 11023 17057
rect 10965 17048 10977 17051
rect 9088 17020 10977 17048
rect 9088 17008 9094 17020
rect 10965 17017 10977 17020
rect 11011 17017 11023 17051
rect 13096 17048 13124 17156
rect 13170 17144 13176 17156
rect 13228 17144 13234 17196
rect 13271 17116 13299 17224
rect 16482 17212 16488 17264
rect 16540 17252 16546 17264
rect 17126 17252 17132 17264
rect 16540 17224 17132 17252
rect 16540 17212 16546 17224
rect 17126 17212 17132 17224
rect 17184 17252 17190 17264
rect 17184 17224 18184 17252
rect 17184 17212 17190 17224
rect 14274 17184 14280 17196
rect 14235 17156 14280 17184
rect 14274 17144 14280 17156
rect 14332 17144 14338 17196
rect 17034 17184 17040 17196
rect 16947 17156 17040 17184
rect 17034 17144 17040 17156
rect 17092 17184 17098 17196
rect 18156 17193 18184 17224
rect 18049 17187 18107 17193
rect 18049 17184 18061 17187
rect 17092 17156 18061 17184
rect 17092 17144 17098 17156
rect 18049 17153 18061 17156
rect 18095 17153 18107 17187
rect 18049 17147 18107 17153
rect 18141 17187 18199 17193
rect 18141 17153 18153 17187
rect 18187 17153 18199 17187
rect 18141 17147 18199 17153
rect 14093 17119 14151 17125
rect 14093 17116 14105 17119
rect 13271 17088 14105 17116
rect 14093 17085 14105 17088
rect 14139 17085 14151 17119
rect 14093 17079 14151 17085
rect 15289 17119 15347 17125
rect 15289 17085 15301 17119
rect 15335 17116 15347 17119
rect 17862 17116 17868 17128
rect 15335 17088 17868 17116
rect 15335 17085 15347 17088
rect 15289 17079 15347 17085
rect 17862 17076 17868 17088
rect 17920 17076 17926 17128
rect 20349 17119 20407 17125
rect 20349 17116 20361 17119
rect 18248 17088 20361 17116
rect 10965 17011 11023 17017
rect 11716 17020 13124 17048
rect 11716 16992 11744 17020
rect 14458 17008 14464 17060
rect 14516 17048 14522 17060
rect 18248 17048 18276 17088
rect 20349 17085 20361 17088
rect 20395 17085 20407 17119
rect 20349 17079 20407 17085
rect 14516 17020 18276 17048
rect 18397 17051 18455 17057
rect 14516 17008 14522 17020
rect 18397 17017 18409 17051
rect 18443 17017 18455 17051
rect 18397 17011 18455 17017
rect 7285 16983 7343 16989
rect 7285 16980 7297 16983
rect 6932 16952 7297 16980
rect 7285 16949 7297 16952
rect 7331 16949 7343 16983
rect 7285 16943 7343 16949
rect 8294 16940 8300 16992
rect 8352 16980 8358 16992
rect 8757 16983 8815 16989
rect 8757 16980 8769 16983
rect 8352 16952 8769 16980
rect 8352 16940 8358 16952
rect 8757 16949 8769 16952
rect 8803 16949 8815 16983
rect 8757 16943 8815 16949
rect 8938 16940 8944 16992
rect 8996 16980 9002 16992
rect 10873 16983 10931 16989
rect 10873 16980 10885 16983
rect 8996 16952 10885 16980
rect 8996 16940 9002 16952
rect 10873 16949 10885 16952
rect 10919 16949 10931 16983
rect 10873 16943 10931 16949
rect 11698 16940 11704 16992
rect 11756 16940 11762 16992
rect 13722 16980 13728 16992
rect 13683 16952 13728 16980
rect 13722 16940 13728 16952
rect 13780 16940 13786 16992
rect 14182 16940 14188 16992
rect 14240 16980 14246 16992
rect 14240 16952 14285 16980
rect 14240 16940 14246 16952
rect 16022 16940 16028 16992
rect 16080 16980 16086 16992
rect 16393 16983 16451 16989
rect 16393 16980 16405 16983
rect 16080 16952 16405 16980
rect 16080 16940 16086 16952
rect 16393 16949 16405 16952
rect 16439 16949 16451 16983
rect 16393 16943 16451 16949
rect 16574 16940 16580 16992
rect 16632 16980 16638 16992
rect 16761 16983 16819 16989
rect 16761 16980 16773 16983
rect 16632 16952 16773 16980
rect 16632 16940 16638 16952
rect 16761 16949 16773 16952
rect 16807 16949 16819 16983
rect 16761 16943 16819 16949
rect 16853 16983 16911 16989
rect 16853 16949 16865 16983
rect 16899 16980 16911 16983
rect 16942 16980 16948 16992
rect 16899 16952 16948 16980
rect 16899 16949 16911 16952
rect 16853 16943 16911 16949
rect 16942 16940 16948 16952
rect 17000 16940 17006 16992
rect 17402 16940 17408 16992
rect 17460 16980 17466 16992
rect 18401 16980 18429 17011
rect 19702 17008 19708 17060
rect 19760 17048 19766 17060
rect 20625 17051 20683 17057
rect 20625 17048 20637 17051
rect 19760 17020 20637 17048
rect 19760 17008 19766 17020
rect 20625 17017 20637 17020
rect 20671 17017 20683 17051
rect 20625 17011 20683 17017
rect 18598 16980 18604 16992
rect 17460 16952 18604 16980
rect 17460 16940 17466 16952
rect 18598 16940 18604 16952
rect 18656 16940 18662 16992
rect 1104 16890 21896 16912
rect 1104 16838 7912 16890
rect 7964 16838 7976 16890
rect 8028 16838 8040 16890
rect 8092 16838 8104 16890
rect 8156 16838 14843 16890
rect 14895 16838 14907 16890
rect 14959 16838 14971 16890
rect 15023 16838 15035 16890
rect 15087 16838 21896 16890
rect 1104 16816 21896 16838
rect 2409 16779 2467 16785
rect 2409 16745 2421 16779
rect 2455 16776 2467 16779
rect 3418 16776 3424 16788
rect 2455 16748 3424 16776
rect 2455 16745 2467 16748
rect 2409 16739 2467 16745
rect 3418 16736 3424 16748
rect 3476 16736 3482 16788
rect 4154 16776 4160 16788
rect 4115 16748 4160 16776
rect 4154 16736 4160 16748
rect 4212 16736 4218 16788
rect 5534 16776 5540 16788
rect 4448 16748 5540 16776
rect 1397 16711 1455 16717
rect 1397 16677 1409 16711
rect 1443 16708 1455 16711
rect 4448 16708 4476 16748
rect 5534 16736 5540 16748
rect 5592 16736 5598 16788
rect 8021 16779 8079 16785
rect 8021 16745 8033 16779
rect 8067 16776 8079 16779
rect 8202 16776 8208 16788
rect 8067 16748 8208 16776
rect 8067 16745 8079 16748
rect 8021 16739 8079 16745
rect 8202 16736 8208 16748
rect 8260 16736 8266 16788
rect 8481 16779 8539 16785
rect 8481 16745 8493 16779
rect 8527 16776 8539 16779
rect 9674 16776 9680 16788
rect 8527 16748 9680 16776
rect 8527 16745 8539 16748
rect 8481 16739 8539 16745
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 9858 16776 9864 16788
rect 9819 16748 9864 16776
rect 9858 16736 9864 16748
rect 9916 16736 9922 16788
rect 12066 16776 12072 16788
rect 10980 16748 12072 16776
rect 1443 16680 4476 16708
rect 4525 16711 4583 16717
rect 1443 16677 1455 16680
rect 1397 16671 1455 16677
rect 4525 16677 4537 16711
rect 4571 16708 4583 16711
rect 6730 16708 6736 16720
rect 4571 16680 6736 16708
rect 4571 16677 4583 16680
rect 4525 16671 4583 16677
rect 6730 16668 6736 16680
rect 6788 16668 6794 16720
rect 9030 16708 9036 16720
rect 6840 16680 9036 16708
rect 2777 16643 2835 16649
rect 2777 16609 2789 16643
rect 2823 16640 2835 16643
rect 4338 16640 4344 16652
rect 2823 16612 4344 16640
rect 2823 16609 2835 16612
rect 2777 16603 2835 16609
rect 4338 16600 4344 16612
rect 4396 16600 4402 16652
rect 4617 16643 4675 16649
rect 4617 16609 4629 16643
rect 4663 16640 4675 16643
rect 5534 16640 5540 16652
rect 4663 16612 5540 16640
rect 4663 16609 4675 16612
rect 4617 16603 4675 16609
rect 5534 16600 5540 16612
rect 5592 16600 5598 16652
rect 5994 16649 6000 16652
rect 5721 16643 5779 16649
rect 5721 16640 5733 16643
rect 5644 16612 5733 16640
rect 2406 16532 2412 16584
rect 2464 16572 2470 16584
rect 2869 16575 2927 16581
rect 2869 16572 2881 16575
rect 2464 16544 2881 16572
rect 2464 16532 2470 16544
rect 2869 16541 2881 16544
rect 2915 16541 2927 16575
rect 2869 16535 2927 16541
rect 3053 16575 3111 16581
rect 3053 16541 3065 16575
rect 3099 16541 3111 16575
rect 3053 16535 3111 16541
rect 4709 16575 4767 16581
rect 4709 16541 4721 16575
rect 4755 16541 4767 16575
rect 4709 16535 4767 16541
rect 2590 16464 2596 16516
rect 2648 16504 2654 16516
rect 2774 16504 2780 16516
rect 2648 16476 2780 16504
rect 2648 16464 2654 16476
rect 2774 16464 2780 16476
rect 2832 16464 2838 16516
rect 3068 16504 3096 16535
rect 4062 16504 4068 16516
rect 3068 16476 4068 16504
rect 4062 16464 4068 16476
rect 4120 16504 4126 16516
rect 4724 16504 4752 16535
rect 5350 16532 5356 16584
rect 5408 16572 5414 16584
rect 5644 16572 5672 16612
rect 5721 16609 5733 16612
rect 5767 16609 5779 16643
rect 5988 16640 6000 16649
rect 5955 16612 6000 16640
rect 5721 16603 5779 16609
rect 5988 16603 6000 16612
rect 5994 16600 6000 16603
rect 6052 16600 6058 16652
rect 6546 16600 6552 16652
rect 6604 16640 6610 16652
rect 6840 16640 6868 16680
rect 9030 16668 9036 16680
rect 9088 16668 9094 16720
rect 6604 16612 6868 16640
rect 8389 16643 8447 16649
rect 6604 16600 6610 16612
rect 8389 16609 8401 16643
rect 8435 16640 8447 16643
rect 9214 16640 9220 16652
rect 8435 16612 9220 16640
rect 8435 16609 8447 16612
rect 8389 16603 8447 16609
rect 9214 16600 9220 16612
rect 9272 16600 9278 16652
rect 9677 16643 9735 16649
rect 9677 16609 9689 16643
rect 9723 16640 9735 16643
rect 10042 16640 10048 16652
rect 9723 16612 10048 16640
rect 9723 16609 9735 16612
rect 9677 16603 9735 16609
rect 10042 16600 10048 16612
rect 10100 16600 10106 16652
rect 10980 16649 11008 16748
rect 12066 16736 12072 16748
rect 12124 16776 12130 16788
rect 12618 16776 12624 16788
rect 12124 16748 12624 16776
rect 12124 16736 12130 16748
rect 12618 16736 12624 16748
rect 12676 16776 12682 16788
rect 13173 16779 13231 16785
rect 13173 16776 13185 16779
rect 12676 16748 13185 16776
rect 12676 16736 12682 16748
rect 13173 16745 13185 16748
rect 13219 16745 13231 16779
rect 13354 16776 13360 16788
rect 13173 16739 13231 16745
rect 13280 16748 13360 16776
rect 12526 16668 12532 16720
rect 12584 16708 12590 16720
rect 13280 16708 13308 16748
rect 13354 16736 13360 16748
rect 13412 16736 13418 16788
rect 13633 16779 13691 16785
rect 13633 16745 13645 16779
rect 13679 16745 13691 16779
rect 13633 16739 13691 16745
rect 13538 16708 13544 16720
rect 12584 16680 13308 16708
rect 13372 16680 13544 16708
rect 12584 16668 12590 16680
rect 11238 16649 11244 16652
rect 10965 16643 11023 16649
rect 10965 16609 10977 16643
rect 11011 16609 11023 16643
rect 11232 16640 11244 16649
rect 11199 16612 11244 16640
rect 10965 16603 11023 16609
rect 11232 16603 11244 16612
rect 11238 16600 11244 16603
rect 11296 16600 11302 16652
rect 13372 16649 13400 16680
rect 13538 16668 13544 16680
rect 13596 16668 13602 16720
rect 13648 16708 13676 16739
rect 13722 16736 13728 16788
rect 13780 16776 13786 16788
rect 14093 16779 14151 16785
rect 14093 16776 14105 16779
rect 13780 16748 14105 16776
rect 13780 16736 13786 16748
rect 14093 16745 14105 16748
rect 14139 16745 14151 16779
rect 14093 16739 14151 16745
rect 14182 16736 14188 16788
rect 14240 16776 14246 16788
rect 15565 16779 15623 16785
rect 15565 16776 15577 16779
rect 14240 16748 15577 16776
rect 14240 16736 14246 16748
rect 15565 16745 15577 16748
rect 15611 16745 15623 16779
rect 16022 16776 16028 16788
rect 15983 16748 16028 16776
rect 15565 16739 15623 16745
rect 16022 16736 16028 16748
rect 16080 16736 16086 16788
rect 18598 16736 18604 16788
rect 18656 16776 18662 16788
rect 18785 16779 18843 16785
rect 18785 16776 18797 16779
rect 18656 16748 18797 16776
rect 18656 16736 18662 16748
rect 18785 16745 18797 16748
rect 18831 16745 18843 16779
rect 18785 16739 18843 16745
rect 19889 16779 19947 16785
rect 19889 16745 19901 16779
rect 19935 16776 19947 16779
rect 19978 16776 19984 16788
rect 19935 16748 19984 16776
rect 19935 16745 19947 16748
rect 19889 16739 19947 16745
rect 19978 16736 19984 16748
rect 20036 16736 20042 16788
rect 14458 16708 14464 16720
rect 13648 16680 14464 16708
rect 14458 16668 14464 16680
rect 14516 16668 14522 16720
rect 15930 16708 15936 16720
rect 15891 16680 15936 16708
rect 15930 16668 15936 16680
rect 15988 16668 15994 16720
rect 16574 16668 16580 16720
rect 16632 16708 16638 16720
rect 17310 16708 17316 16720
rect 16632 16680 17316 16708
rect 16632 16668 16638 16680
rect 17310 16668 17316 16680
rect 17368 16668 17374 16720
rect 17402 16668 17408 16720
rect 17460 16708 17466 16720
rect 17650 16711 17708 16717
rect 17650 16708 17662 16711
rect 17460 16680 17662 16708
rect 17460 16668 17466 16680
rect 17650 16677 17662 16680
rect 17696 16677 17708 16711
rect 17650 16671 17708 16677
rect 17862 16668 17868 16720
rect 17920 16708 17926 16720
rect 19610 16708 19616 16720
rect 17920 16680 19616 16708
rect 17920 16668 17926 16680
rect 19610 16668 19616 16680
rect 19668 16668 19674 16720
rect 13357 16643 13415 16649
rect 13357 16609 13369 16643
rect 13403 16609 13415 16643
rect 13357 16603 13415 16609
rect 13446 16600 13452 16652
rect 13504 16640 13510 16652
rect 14001 16643 14059 16649
rect 14001 16640 14013 16643
rect 13504 16612 14013 16640
rect 13504 16600 13510 16612
rect 14001 16609 14013 16612
rect 14047 16609 14059 16643
rect 14001 16603 14059 16609
rect 16942 16600 16948 16652
rect 17000 16640 17006 16652
rect 19150 16640 19156 16652
rect 17000 16612 19156 16640
rect 17000 16600 17006 16612
rect 19150 16600 19156 16612
rect 19208 16600 19214 16652
rect 19702 16640 19708 16652
rect 19663 16612 19708 16640
rect 19702 16600 19708 16612
rect 19760 16600 19766 16652
rect 8662 16572 8668 16584
rect 5408 16544 5672 16572
rect 8623 16544 8668 16572
rect 5408 16532 5414 16544
rect 8662 16532 8668 16544
rect 8720 16532 8726 16584
rect 14274 16572 14280 16584
rect 14235 16544 14280 16572
rect 14274 16532 14280 16544
rect 14332 16532 14338 16584
rect 16209 16575 16267 16581
rect 16209 16541 16221 16575
rect 16255 16572 16267 16575
rect 16255 16544 16344 16572
rect 16255 16541 16267 16544
rect 16209 16535 16267 16541
rect 4120 16476 4752 16504
rect 4120 16464 4126 16476
rect 9766 16464 9772 16516
rect 9824 16504 9830 16516
rect 10962 16504 10968 16516
rect 9824 16476 10968 16504
rect 9824 16464 9830 16476
rect 10962 16464 10968 16476
rect 11020 16464 11026 16516
rect 11900 16476 14044 16504
rect 1946 16396 1952 16448
rect 2004 16436 2010 16448
rect 6086 16436 6092 16448
rect 2004 16408 6092 16436
rect 2004 16396 2010 16408
rect 6086 16396 6092 16408
rect 6144 16396 6150 16448
rect 7006 16396 7012 16448
rect 7064 16436 7070 16448
rect 7101 16439 7159 16445
rect 7101 16436 7113 16439
rect 7064 16408 7113 16436
rect 7064 16396 7070 16408
rect 7101 16405 7113 16408
rect 7147 16405 7159 16439
rect 7101 16399 7159 16405
rect 10318 16396 10324 16448
rect 10376 16436 10382 16448
rect 10778 16436 10784 16448
rect 10376 16408 10784 16436
rect 10376 16396 10382 16408
rect 10778 16396 10784 16408
rect 10836 16436 10842 16448
rect 11900 16436 11928 16476
rect 10836 16408 11928 16436
rect 10836 16396 10842 16408
rect 12158 16396 12164 16448
rect 12216 16436 12222 16448
rect 12345 16439 12403 16445
rect 12345 16436 12357 16439
rect 12216 16408 12357 16436
rect 12216 16396 12222 16408
rect 12345 16405 12357 16408
rect 12391 16436 12403 16439
rect 13170 16436 13176 16448
rect 12391 16408 13176 16436
rect 12391 16405 12403 16408
rect 12345 16399 12403 16405
rect 13170 16396 13176 16408
rect 13228 16396 13234 16448
rect 14016 16436 14044 16476
rect 16206 16436 16212 16448
rect 14016 16408 16212 16436
rect 16206 16396 16212 16408
rect 16264 16396 16270 16448
rect 16316 16436 16344 16544
rect 17126 16532 17132 16584
rect 17184 16572 17190 16584
rect 17405 16575 17463 16581
rect 17405 16572 17417 16575
rect 17184 16544 17417 16572
rect 17184 16532 17190 16544
rect 17405 16541 17417 16544
rect 17451 16541 17463 16575
rect 17405 16535 17463 16541
rect 18782 16464 18788 16516
rect 18840 16504 18846 16516
rect 19242 16504 19248 16516
rect 18840 16476 19248 16504
rect 18840 16464 18846 16476
rect 19242 16464 19248 16476
rect 19300 16464 19306 16516
rect 16574 16436 16580 16448
rect 16316 16408 16580 16436
rect 16574 16396 16580 16408
rect 16632 16436 16638 16448
rect 17678 16436 17684 16448
rect 16632 16408 17684 16436
rect 16632 16396 16638 16408
rect 17678 16396 17684 16408
rect 17736 16396 17742 16448
rect 1104 16346 21896 16368
rect 1104 16294 4447 16346
rect 4499 16294 4511 16346
rect 4563 16294 4575 16346
rect 4627 16294 4639 16346
rect 4691 16294 11378 16346
rect 11430 16294 11442 16346
rect 11494 16294 11506 16346
rect 11558 16294 11570 16346
rect 11622 16294 18308 16346
rect 18360 16294 18372 16346
rect 18424 16294 18436 16346
rect 18488 16294 18500 16346
rect 18552 16294 21896 16346
rect 1104 16272 21896 16294
rect 3050 16232 3056 16244
rect 3011 16204 3056 16232
rect 3050 16192 3056 16204
rect 3108 16192 3114 16244
rect 4338 16192 4344 16244
rect 4396 16232 4402 16244
rect 4617 16235 4675 16241
rect 4617 16232 4629 16235
rect 4396 16204 4629 16232
rect 4396 16192 4402 16204
rect 4617 16201 4629 16204
rect 4663 16201 4675 16235
rect 4617 16195 4675 16201
rect 6730 16192 6736 16244
rect 6788 16232 6794 16244
rect 6825 16235 6883 16241
rect 6825 16232 6837 16235
rect 6788 16204 6837 16232
rect 6788 16192 6794 16204
rect 6825 16201 6837 16204
rect 6871 16201 6883 16235
rect 8570 16232 8576 16244
rect 6825 16195 6883 16201
rect 8404 16204 8576 16232
rect 3620 16136 5212 16164
rect 3620 16108 3648 16136
rect 1946 16096 1952 16108
rect 1907 16068 1952 16096
rect 1946 16056 1952 16068
rect 2004 16056 2010 16108
rect 2130 16096 2136 16108
rect 2091 16068 2136 16096
rect 2130 16056 2136 16068
rect 2188 16056 2194 16108
rect 2958 16056 2964 16108
rect 3016 16096 3022 16108
rect 3602 16096 3608 16108
rect 3016 16068 3608 16096
rect 3016 16056 3022 16068
rect 3602 16056 3608 16068
rect 3660 16056 3666 16108
rect 3697 16099 3755 16105
rect 3697 16065 3709 16099
rect 3743 16096 3755 16099
rect 4890 16096 4896 16108
rect 3743 16068 4896 16096
rect 3743 16065 3755 16068
rect 3697 16059 3755 16065
rect 4890 16056 4896 16068
rect 4948 16056 4954 16108
rect 5184 16105 5212 16136
rect 5169 16099 5227 16105
rect 5169 16065 5181 16099
rect 5215 16096 5227 16099
rect 7006 16096 7012 16108
rect 5215 16068 7012 16096
rect 5215 16065 5227 16068
rect 5169 16059 5227 16065
rect 7006 16056 7012 16068
rect 7064 16096 7070 16108
rect 7377 16099 7435 16105
rect 7377 16096 7389 16099
rect 7064 16068 7389 16096
rect 7064 16056 7070 16068
rect 7377 16065 7389 16068
rect 7423 16065 7435 16099
rect 8404 16096 8432 16204
rect 8570 16192 8576 16204
rect 8628 16192 8634 16244
rect 8662 16192 8668 16244
rect 8720 16232 8726 16244
rect 9769 16235 9827 16241
rect 9769 16232 9781 16235
rect 8720 16204 9781 16232
rect 8720 16192 8726 16204
rect 9769 16201 9781 16204
rect 9815 16201 9827 16235
rect 9769 16195 9827 16201
rect 10042 16192 10048 16244
rect 10100 16232 10106 16244
rect 10100 16204 16160 16232
rect 10100 16192 10106 16204
rect 14274 16164 14280 16176
rect 14187 16136 14280 16164
rect 14274 16124 14280 16136
rect 14332 16164 14338 16176
rect 16132 16164 16160 16204
rect 16206 16192 16212 16244
rect 16264 16232 16270 16244
rect 16485 16235 16543 16241
rect 16485 16232 16497 16235
rect 16264 16204 16497 16232
rect 16264 16192 16270 16204
rect 16485 16201 16497 16204
rect 16531 16201 16543 16235
rect 20714 16232 20720 16244
rect 20675 16204 20720 16232
rect 16485 16195 16543 16201
rect 20714 16192 20720 16204
rect 20772 16192 20778 16244
rect 17770 16164 17776 16176
rect 14332 16136 14780 16164
rect 16132 16136 17776 16164
rect 14332 16124 14338 16136
rect 11422 16096 11428 16108
rect 8404 16068 8524 16096
rect 11383 16068 11428 16096
rect 7377 16059 7435 16065
rect 1857 16031 1915 16037
rect 1857 15997 1869 16031
rect 1903 16028 1915 16031
rect 2590 16028 2596 16040
rect 1903 16000 2596 16028
rect 1903 15997 1915 16000
rect 1857 15991 1915 15997
rect 2590 15988 2596 16000
rect 2648 15988 2654 16040
rect 3418 16028 3424 16040
rect 3379 16000 3424 16028
rect 3418 15988 3424 16000
rect 3476 15988 3482 16040
rect 3513 16031 3571 16037
rect 3513 15997 3525 16031
rect 3559 16028 3571 16031
rect 4154 16028 4160 16040
rect 3559 16000 4160 16028
rect 3559 15997 3571 16000
rect 3513 15991 3571 15997
rect 4154 15988 4160 16000
rect 4212 15988 4218 16040
rect 8386 16028 8392 16040
rect 8347 16000 8392 16028
rect 8386 15988 8392 16000
rect 8444 15988 8450 16040
rect 8496 16028 8524 16068
rect 11422 16056 11428 16068
rect 11480 16056 11486 16108
rect 8645 16031 8703 16037
rect 8645 16028 8657 16031
rect 8496 16000 8657 16028
rect 8645 15997 8657 16000
rect 8691 15997 8703 16031
rect 11882 16028 11888 16040
rect 8645 15991 8703 15997
rect 10980 16000 11888 16028
rect 4985 15963 5043 15969
rect 4985 15960 4997 15963
rect 2976 15932 4997 15960
rect 1489 15895 1547 15901
rect 1489 15861 1501 15895
rect 1535 15892 1547 15895
rect 1946 15892 1952 15904
rect 1535 15864 1952 15892
rect 1535 15861 1547 15864
rect 1489 15855 1547 15861
rect 1946 15852 1952 15864
rect 2004 15852 2010 15904
rect 2038 15852 2044 15904
rect 2096 15892 2102 15904
rect 2976 15892 3004 15932
rect 4985 15929 4997 15932
rect 5031 15929 5043 15963
rect 4985 15923 5043 15929
rect 7193 15963 7251 15969
rect 7193 15929 7205 15963
rect 7239 15960 7251 15963
rect 10980 15960 11008 16000
rect 11882 15988 11888 16000
rect 11940 15988 11946 16040
rect 12618 15988 12624 16040
rect 12676 16028 12682 16040
rect 13170 16037 13176 16040
rect 12897 16031 12955 16037
rect 12897 16028 12909 16031
rect 12676 16000 12909 16028
rect 12676 15988 12682 16000
rect 12897 15997 12909 16000
rect 12943 15997 12955 16031
rect 13164 16028 13176 16037
rect 13083 16000 13176 16028
rect 12897 15991 12955 15997
rect 13164 15991 13176 16000
rect 13228 16028 13234 16040
rect 14182 16028 14188 16040
rect 13228 16000 14188 16028
rect 13170 15988 13176 15991
rect 13228 15988 13234 16000
rect 14182 15988 14188 16000
rect 14240 15988 14246 16040
rect 7239 15932 11008 15960
rect 7239 15929 7251 15932
rect 7193 15923 7251 15929
rect 11054 15920 11060 15972
rect 11112 15960 11118 15972
rect 11241 15963 11299 15969
rect 11241 15960 11253 15963
rect 11112 15932 11253 15960
rect 11112 15920 11118 15932
rect 11241 15929 11253 15932
rect 11287 15960 11299 15963
rect 11514 15960 11520 15972
rect 11287 15932 11520 15960
rect 11287 15929 11299 15932
rect 11241 15923 11299 15929
rect 11514 15920 11520 15932
rect 11572 15920 11578 15972
rect 11974 15920 11980 15972
rect 12032 15960 12038 15972
rect 14752 15960 14780 16136
rect 17770 16124 17776 16136
rect 17828 16124 17834 16176
rect 15105 16031 15163 16037
rect 15105 15997 15117 16031
rect 15151 16028 15163 16031
rect 15194 16028 15200 16040
rect 15151 16000 15200 16028
rect 15151 15997 15163 16000
rect 15105 15991 15163 15997
rect 15194 15988 15200 16000
rect 15252 15988 15258 16040
rect 18141 16031 18199 16037
rect 18141 16028 18153 16031
rect 15488 16000 18153 16028
rect 15350 15963 15408 15969
rect 15350 15960 15362 15963
rect 12032 15932 14688 15960
rect 14752 15932 15362 15960
rect 12032 15920 12038 15932
rect 2096 15864 3004 15892
rect 2096 15852 2102 15864
rect 3418 15852 3424 15904
rect 3476 15892 3482 15904
rect 5077 15895 5135 15901
rect 5077 15892 5089 15895
rect 3476 15864 5089 15892
rect 3476 15852 3482 15864
rect 5077 15861 5089 15864
rect 5123 15861 5135 15895
rect 5077 15855 5135 15861
rect 7285 15895 7343 15901
rect 7285 15861 7297 15895
rect 7331 15892 7343 15895
rect 8386 15892 8392 15904
rect 7331 15864 8392 15892
rect 7331 15861 7343 15864
rect 7285 15855 7343 15861
rect 8386 15852 8392 15864
rect 8444 15892 8450 15904
rect 8938 15892 8944 15904
rect 8444 15864 8944 15892
rect 8444 15852 8450 15864
rect 8938 15852 8944 15864
rect 8996 15852 9002 15904
rect 10778 15892 10784 15904
rect 10739 15864 10784 15892
rect 10778 15852 10784 15864
rect 10836 15852 10842 15904
rect 11146 15892 11152 15904
rect 11107 15864 11152 15892
rect 11146 15852 11152 15864
rect 11204 15852 11210 15904
rect 14660 15892 14688 15932
rect 15350 15929 15362 15932
rect 15396 15929 15408 15963
rect 15350 15923 15408 15929
rect 15488 15892 15516 16000
rect 18141 15997 18153 16000
rect 18187 15997 18199 16031
rect 18141 15991 18199 15997
rect 19245 16031 19303 16037
rect 19245 15997 19257 16031
rect 19291 15997 19303 16031
rect 19245 15991 19303 15997
rect 20533 16031 20591 16037
rect 20533 15997 20545 16031
rect 20579 15997 20591 16031
rect 20533 15991 20591 15997
rect 15562 15920 15568 15972
rect 15620 15960 15626 15972
rect 19260 15960 19288 15991
rect 15620 15932 19288 15960
rect 15620 15920 15626 15932
rect 19426 15920 19432 15972
rect 19484 15960 19490 15972
rect 19521 15963 19579 15969
rect 19521 15960 19533 15963
rect 19484 15932 19533 15960
rect 19484 15920 19490 15932
rect 19521 15929 19533 15932
rect 19567 15929 19579 15963
rect 19521 15923 19579 15929
rect 14660 15864 15516 15892
rect 18325 15895 18383 15901
rect 18325 15861 18337 15895
rect 18371 15892 18383 15895
rect 18598 15892 18604 15904
rect 18371 15864 18604 15892
rect 18371 15861 18383 15864
rect 18325 15855 18383 15861
rect 18598 15852 18604 15864
rect 18656 15852 18662 15904
rect 18874 15852 18880 15904
rect 18932 15892 18938 15904
rect 20548 15892 20576 15991
rect 18932 15864 20576 15892
rect 18932 15852 18938 15864
rect 1104 15802 21896 15824
rect 1104 15750 7912 15802
rect 7964 15750 7976 15802
rect 8028 15750 8040 15802
rect 8092 15750 8104 15802
rect 8156 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 15035 15802
rect 15087 15750 21896 15802
rect 1104 15728 21896 15750
rect 1397 15691 1455 15697
rect 1397 15657 1409 15691
rect 1443 15688 1455 15691
rect 2038 15688 2044 15700
rect 1443 15660 2044 15688
rect 1443 15657 1455 15660
rect 1397 15651 1455 15657
rect 2038 15648 2044 15660
rect 2096 15648 2102 15700
rect 2406 15688 2412 15700
rect 2367 15660 2412 15688
rect 2406 15648 2412 15660
rect 2464 15648 2470 15700
rect 4157 15691 4215 15697
rect 4157 15688 4169 15691
rect 2516 15660 4169 15688
rect 1394 15512 1400 15564
rect 1452 15552 1458 15564
rect 2516 15552 2544 15660
rect 4157 15657 4169 15660
rect 4203 15657 4215 15691
rect 5350 15688 5356 15700
rect 4157 15651 4215 15657
rect 4264 15660 5356 15688
rect 1452 15524 2544 15552
rect 1452 15512 1458 15524
rect 2590 15512 2596 15564
rect 2648 15552 2654 15564
rect 2777 15555 2835 15561
rect 2777 15552 2789 15555
rect 2648 15524 2789 15552
rect 2648 15512 2654 15524
rect 2777 15521 2789 15524
rect 2823 15521 2835 15555
rect 2777 15515 2835 15521
rect 2869 15555 2927 15561
rect 2869 15521 2881 15555
rect 2915 15552 2927 15555
rect 4154 15552 4160 15564
rect 2915 15524 4160 15552
rect 2915 15521 2927 15524
rect 2869 15515 2927 15521
rect 4154 15512 4160 15524
rect 4212 15512 4218 15564
rect 4264 15561 4292 15660
rect 5350 15648 5356 15660
rect 5408 15648 5414 15700
rect 5534 15648 5540 15700
rect 5592 15688 5598 15700
rect 6457 15691 6515 15697
rect 6457 15688 6469 15691
rect 5592 15660 6469 15688
rect 5592 15648 5598 15660
rect 6457 15657 6469 15660
rect 6503 15657 6515 15691
rect 6457 15651 6515 15657
rect 6822 15648 6828 15700
rect 6880 15688 6886 15700
rect 6917 15691 6975 15697
rect 6917 15688 6929 15691
rect 6880 15660 6929 15688
rect 6880 15648 6886 15660
rect 6917 15657 6929 15660
rect 6963 15657 6975 15691
rect 6917 15651 6975 15657
rect 8021 15691 8079 15697
rect 8021 15657 8033 15691
rect 8067 15688 8079 15691
rect 8294 15688 8300 15700
rect 8067 15660 8300 15688
rect 8067 15657 8079 15660
rect 8021 15651 8079 15657
rect 8294 15648 8300 15660
rect 8352 15648 8358 15700
rect 8481 15691 8539 15697
rect 8481 15657 8493 15691
rect 8527 15688 8539 15691
rect 9490 15688 9496 15700
rect 8527 15660 9496 15688
rect 8527 15657 8539 15660
rect 8481 15651 8539 15657
rect 9490 15648 9496 15660
rect 9548 15648 9554 15700
rect 9674 15688 9680 15700
rect 9635 15660 9680 15688
rect 9674 15648 9680 15660
rect 9732 15648 9738 15700
rect 10042 15688 10048 15700
rect 10003 15660 10048 15688
rect 10042 15648 10048 15660
rect 10100 15648 10106 15700
rect 10778 15648 10784 15700
rect 10836 15688 10842 15700
rect 11885 15691 11943 15697
rect 11885 15688 11897 15691
rect 10836 15660 11897 15688
rect 10836 15648 10842 15660
rect 11885 15657 11897 15660
rect 11931 15657 11943 15691
rect 11885 15651 11943 15657
rect 11977 15691 12035 15697
rect 11977 15657 11989 15691
rect 12023 15688 12035 15691
rect 13081 15691 13139 15697
rect 13081 15688 13093 15691
rect 12023 15660 13093 15688
rect 12023 15657 12035 15660
rect 11977 15651 12035 15657
rect 13081 15657 13093 15660
rect 13127 15657 13139 15691
rect 13081 15651 13139 15657
rect 15194 15648 15200 15700
rect 15252 15688 15258 15700
rect 15654 15688 15660 15700
rect 15252 15660 15660 15688
rect 15252 15648 15258 15660
rect 15654 15648 15660 15660
rect 15712 15648 15718 15700
rect 16025 15691 16083 15697
rect 16025 15657 16037 15691
rect 16071 15688 16083 15691
rect 16485 15691 16543 15697
rect 16485 15688 16497 15691
rect 16071 15660 16497 15688
rect 16071 15657 16083 15660
rect 16025 15651 16083 15657
rect 16485 15657 16497 15660
rect 16531 15657 16543 15691
rect 16485 15651 16543 15657
rect 16577 15691 16635 15697
rect 16577 15657 16589 15691
rect 16623 15688 16635 15691
rect 17494 15688 17500 15700
rect 16623 15660 17500 15688
rect 16623 15657 16635 15660
rect 16577 15651 16635 15657
rect 17494 15648 17500 15660
rect 17552 15648 17558 15700
rect 17681 15691 17739 15697
rect 17681 15657 17693 15691
rect 17727 15657 17739 15691
rect 19886 15688 19892 15700
rect 19847 15660 19892 15688
rect 17681 15651 17739 15657
rect 17696 15620 17724 15651
rect 19886 15648 19892 15660
rect 19944 15648 19950 15700
rect 4347 15592 17724 15620
rect 4249 15555 4307 15561
rect 4249 15521 4261 15555
rect 4295 15521 4307 15555
rect 4249 15515 4307 15521
rect 2958 15444 2964 15496
rect 3016 15484 3022 15496
rect 4347 15484 4375 15592
rect 4516 15555 4574 15561
rect 4516 15521 4528 15555
rect 4562 15552 4574 15555
rect 4890 15552 4896 15564
rect 4562 15524 4896 15552
rect 4562 15521 4574 15524
rect 4516 15515 4574 15521
rect 4890 15512 4896 15524
rect 4948 15512 4954 15564
rect 6178 15512 6184 15564
rect 6236 15552 6242 15564
rect 6546 15552 6552 15564
rect 6236 15524 6552 15552
rect 6236 15512 6242 15524
rect 6546 15512 6552 15524
rect 6604 15552 6610 15564
rect 6825 15555 6883 15561
rect 6825 15552 6837 15555
rect 6604 15524 6837 15552
rect 6604 15512 6610 15524
rect 6825 15521 6837 15524
rect 6871 15521 6883 15555
rect 6825 15515 6883 15521
rect 6914 15512 6920 15564
rect 6972 15552 6978 15564
rect 6972 15524 8248 15552
rect 6972 15512 6978 15524
rect 7006 15484 7012 15496
rect 3016 15456 3061 15484
rect 3252 15456 4375 15484
rect 6967 15456 7012 15484
rect 3016 15444 3022 15456
rect 1578 15308 1584 15360
rect 1636 15348 1642 15360
rect 3252 15348 3280 15456
rect 7006 15444 7012 15456
rect 7064 15444 7070 15496
rect 8220 15484 8248 15524
rect 8294 15512 8300 15564
rect 8352 15552 8358 15564
rect 8389 15555 8447 15561
rect 8389 15552 8401 15555
rect 8352 15524 8401 15552
rect 8352 15512 8358 15524
rect 8389 15521 8401 15524
rect 8435 15521 8447 15555
rect 10137 15555 10195 15561
rect 10137 15552 10149 15555
rect 8389 15515 8447 15521
rect 8588 15524 10149 15552
rect 8588 15484 8616 15524
rect 10137 15521 10149 15524
rect 10183 15552 10195 15555
rect 10183 15524 11376 15552
rect 10183 15521 10195 15524
rect 10137 15515 10195 15521
rect 8220 15456 8616 15484
rect 8662 15444 8668 15496
rect 8720 15484 8726 15496
rect 10229 15487 10287 15493
rect 8720 15456 8765 15484
rect 8720 15444 8726 15456
rect 10229 15453 10241 15487
rect 10275 15453 10287 15487
rect 11348 15484 11376 15524
rect 11422 15512 11428 15564
rect 11480 15552 11486 15564
rect 11480 15524 12480 15552
rect 11480 15512 11486 15524
rect 12066 15484 12072 15496
rect 11348 15456 12072 15484
rect 10229 15447 10287 15453
rect 5629 15419 5687 15425
rect 5629 15385 5641 15419
rect 5675 15416 5687 15419
rect 5994 15416 6000 15428
rect 5675 15388 6000 15416
rect 5675 15385 5687 15388
rect 5629 15379 5687 15385
rect 5994 15376 6000 15388
rect 6052 15376 6058 15428
rect 8570 15376 8576 15428
rect 8628 15416 8634 15428
rect 10244 15416 10272 15447
rect 12066 15444 12072 15456
rect 12124 15444 12130 15496
rect 12158 15444 12164 15496
rect 12216 15484 12222 15496
rect 12452 15484 12480 15524
rect 12526 15512 12532 15564
rect 12584 15552 12590 15564
rect 13449 15555 13507 15561
rect 13449 15552 13461 15555
rect 12584 15524 13461 15552
rect 12584 15512 12590 15524
rect 13449 15521 13461 15524
rect 13495 15521 13507 15555
rect 13449 15515 13507 15521
rect 13538 15512 13544 15564
rect 13596 15552 13602 15564
rect 18046 15552 18052 15564
rect 13596 15524 13641 15552
rect 18007 15524 18052 15552
rect 13596 15512 13602 15524
rect 18046 15512 18052 15524
rect 18104 15512 18110 15564
rect 19705 15555 19763 15561
rect 19705 15521 19717 15555
rect 19751 15552 19763 15555
rect 19794 15552 19800 15564
rect 19751 15524 19800 15552
rect 19751 15521 19763 15524
rect 19705 15515 19763 15521
rect 19794 15512 19800 15524
rect 19852 15512 19858 15564
rect 13725 15487 13783 15493
rect 13725 15484 13737 15487
rect 12216 15456 12261 15484
rect 12452 15456 13737 15484
rect 12216 15444 12222 15456
rect 13725 15453 13737 15456
rect 13771 15484 13783 15487
rect 16390 15484 16396 15496
rect 13771 15456 16396 15484
rect 13771 15453 13783 15456
rect 13725 15447 13783 15453
rect 16390 15444 16396 15456
rect 16448 15444 16454 15496
rect 16574 15444 16580 15496
rect 16632 15484 16638 15496
rect 16669 15487 16727 15493
rect 16669 15484 16681 15487
rect 16632 15456 16681 15484
rect 16632 15444 16638 15456
rect 16669 15453 16681 15456
rect 16715 15453 16727 15487
rect 18138 15484 18144 15496
rect 18099 15456 18144 15484
rect 16669 15447 16727 15453
rect 18138 15444 18144 15456
rect 18196 15444 18202 15496
rect 18233 15487 18291 15493
rect 18233 15453 18245 15487
rect 18279 15453 18291 15487
rect 18233 15447 18291 15453
rect 10410 15416 10416 15428
rect 8628 15388 10416 15416
rect 8628 15376 8634 15388
rect 10410 15376 10416 15388
rect 10468 15376 10474 15428
rect 11517 15419 11575 15425
rect 11517 15385 11529 15419
rect 11563 15416 11575 15419
rect 13446 15416 13452 15428
rect 11563 15388 13452 15416
rect 11563 15385 11575 15388
rect 11517 15379 11575 15385
rect 13446 15376 13452 15388
rect 13504 15376 13510 15428
rect 16025 15419 16083 15425
rect 16025 15385 16037 15419
rect 16071 15416 16083 15419
rect 16071 15388 17172 15416
rect 16071 15385 16083 15388
rect 16025 15379 16083 15385
rect 1636 15320 3280 15348
rect 4157 15351 4215 15357
rect 1636 15308 1642 15320
rect 4157 15317 4169 15351
rect 4203 15348 4215 15351
rect 15562 15348 15568 15360
rect 4203 15320 15568 15348
rect 4203 15317 4215 15320
rect 4157 15311 4215 15317
rect 15562 15308 15568 15320
rect 15620 15308 15626 15360
rect 15654 15308 15660 15360
rect 15712 15348 15718 15360
rect 16117 15351 16175 15357
rect 16117 15348 16129 15351
rect 15712 15320 16129 15348
rect 15712 15308 15718 15320
rect 16117 15317 16129 15320
rect 16163 15317 16175 15351
rect 17144 15348 17172 15388
rect 17402 15376 17408 15428
rect 17460 15416 17466 15428
rect 18248 15416 18276 15447
rect 17460 15388 18276 15416
rect 17460 15376 17466 15388
rect 18322 15376 18328 15428
rect 18380 15416 18386 15428
rect 19334 15416 19340 15428
rect 18380 15388 19340 15416
rect 18380 15376 18386 15388
rect 19334 15376 19340 15388
rect 19392 15376 19398 15428
rect 18046 15348 18052 15360
rect 17144 15320 18052 15348
rect 16117 15311 16175 15317
rect 18046 15308 18052 15320
rect 18104 15308 18110 15360
rect 1104 15258 21896 15280
rect 1104 15206 4447 15258
rect 4499 15206 4511 15258
rect 4563 15206 4575 15258
rect 4627 15206 4639 15258
rect 4691 15206 11378 15258
rect 11430 15206 11442 15258
rect 11494 15206 11506 15258
rect 11558 15206 11570 15258
rect 11622 15206 18308 15258
rect 18360 15206 18372 15258
rect 18424 15206 18436 15258
rect 18488 15206 18500 15258
rect 18552 15206 21896 15258
rect 1104 15184 21896 15206
rect 10410 15144 10416 15156
rect 10371 15116 10416 15144
rect 10410 15104 10416 15116
rect 10468 15104 10474 15156
rect 11425 15147 11483 15153
rect 11425 15113 11437 15147
rect 11471 15144 11483 15147
rect 12250 15144 12256 15156
rect 11471 15116 12256 15144
rect 11471 15113 11483 15116
rect 11425 15107 11483 15113
rect 12250 15104 12256 15116
rect 12308 15104 12314 15156
rect 18690 15144 18696 15156
rect 12360 15116 18696 15144
rect 1949 15079 2007 15085
rect 1949 15045 1961 15079
rect 1995 15076 2007 15079
rect 2866 15076 2872 15088
rect 1995 15048 2872 15076
rect 1995 15045 2007 15048
rect 1949 15039 2007 15045
rect 2866 15036 2872 15048
rect 2924 15036 2930 15088
rect 10502 15036 10508 15088
rect 10560 15076 10566 15088
rect 12360 15076 12388 15116
rect 18690 15104 18696 15116
rect 18748 15104 18754 15156
rect 20714 15144 20720 15156
rect 20675 15116 20720 15144
rect 20714 15104 20720 15116
rect 20772 15104 20778 15156
rect 10560 15048 12388 15076
rect 10560 15036 10566 15048
rect 12434 15036 12440 15088
rect 12492 15076 12498 15088
rect 13078 15076 13084 15088
rect 12492 15048 13084 15076
rect 12492 15036 12498 15048
rect 13078 15036 13084 15048
rect 13136 15036 13142 15088
rect 2130 14968 2136 15020
rect 2188 15008 2194 15020
rect 2501 15011 2559 15017
rect 2501 15008 2513 15011
rect 2188 14980 2513 15008
rect 2188 14968 2194 14980
rect 2501 14977 2513 14980
rect 2547 14977 2559 15011
rect 2501 14971 2559 14977
rect 8478 14968 8484 15020
rect 8536 15008 8542 15020
rect 9033 15011 9091 15017
rect 9033 15008 9045 15011
rect 8536 14980 9045 15008
rect 8536 14968 8542 14980
rect 9033 14977 9045 14980
rect 9079 14977 9091 15011
rect 9033 14971 9091 14977
rect 10134 14968 10140 15020
rect 10192 15008 10198 15020
rect 10410 15008 10416 15020
rect 10192 14980 10416 15008
rect 10192 14968 10198 14980
rect 10410 14968 10416 14980
rect 10468 14968 10474 15020
rect 19429 15011 19487 15017
rect 19429 15008 19441 15011
rect 17328 14980 19441 15008
rect 3326 14900 3332 14952
rect 3384 14940 3390 14952
rect 3513 14943 3571 14949
rect 3513 14940 3525 14943
rect 3384 14912 3525 14940
rect 3384 14900 3390 14912
rect 3513 14909 3525 14912
rect 3559 14940 3571 14943
rect 5350 14940 5356 14952
rect 3559 14912 5356 14940
rect 3559 14909 3571 14912
rect 3513 14903 3571 14909
rect 5350 14900 5356 14912
rect 5408 14900 5414 14952
rect 6825 14943 6883 14949
rect 6825 14909 6837 14943
rect 6871 14940 6883 14943
rect 8496 14940 8524 14968
rect 6871 14912 8524 14940
rect 6871 14909 6883 14912
rect 6825 14903 6883 14909
rect 10042 14900 10048 14952
rect 10100 14940 10106 14952
rect 10594 14940 10600 14952
rect 10100 14912 10600 14940
rect 10100 14900 10106 14912
rect 10594 14900 10600 14912
rect 10652 14940 10658 14952
rect 11241 14943 11299 14949
rect 11241 14940 11253 14943
rect 10652 14912 11253 14940
rect 10652 14900 10658 14912
rect 11241 14909 11253 14912
rect 11287 14909 11299 14943
rect 11241 14903 11299 14909
rect 13081 14943 13139 14949
rect 13081 14909 13093 14943
rect 13127 14940 13139 14943
rect 15286 14940 15292 14952
rect 13127 14912 15292 14940
rect 13127 14909 13139 14912
rect 13081 14903 13139 14909
rect 15286 14900 15292 14912
rect 15344 14900 15350 14952
rect 2222 14832 2228 14884
rect 2280 14872 2286 14884
rect 2317 14875 2375 14881
rect 2317 14872 2329 14875
rect 2280 14844 2329 14872
rect 2280 14832 2286 14844
rect 2317 14841 2329 14844
rect 2363 14872 2375 14875
rect 3780 14875 3838 14881
rect 2363 14844 3740 14872
rect 2363 14841 2375 14844
rect 2317 14835 2375 14841
rect 2409 14807 2467 14813
rect 2409 14773 2421 14807
rect 2455 14804 2467 14807
rect 3050 14804 3056 14816
rect 2455 14776 3056 14804
rect 2455 14773 2467 14776
rect 2409 14767 2467 14773
rect 3050 14764 3056 14776
rect 3108 14764 3114 14816
rect 3712 14804 3740 14844
rect 3780 14841 3792 14875
rect 3826 14872 3838 14875
rect 3970 14872 3976 14884
rect 3826 14844 3976 14872
rect 3826 14841 3838 14844
rect 3780 14835 3838 14841
rect 3970 14832 3976 14844
rect 4028 14832 4034 14884
rect 6914 14872 6920 14884
rect 4080 14844 6920 14872
rect 4080 14804 4108 14844
rect 6914 14832 6920 14844
rect 6972 14832 6978 14884
rect 7092 14875 7150 14881
rect 7092 14841 7104 14875
rect 7138 14872 7150 14875
rect 7190 14872 7196 14884
rect 7138 14844 7196 14872
rect 7138 14841 7150 14844
rect 7092 14835 7150 14841
rect 7190 14832 7196 14844
rect 7248 14832 7254 14884
rect 9278 14875 9336 14881
rect 9278 14872 9290 14875
rect 8220 14844 9290 14872
rect 8220 14816 8248 14844
rect 9278 14841 9290 14844
rect 9324 14841 9336 14875
rect 9278 14835 9336 14841
rect 12434 14832 12440 14884
rect 12492 14872 12498 14884
rect 13326 14875 13384 14881
rect 13326 14872 13338 14875
rect 12492 14844 13338 14872
rect 12492 14832 12498 14844
rect 13326 14841 13338 14844
rect 13372 14841 13384 14875
rect 14550 14872 14556 14884
rect 14463 14844 14556 14872
rect 13326 14835 13384 14841
rect 4890 14804 4896 14816
rect 3712 14776 4108 14804
rect 4851 14776 4896 14804
rect 4890 14764 4896 14776
rect 4948 14764 4954 14816
rect 5721 14807 5779 14813
rect 5721 14773 5733 14807
rect 5767 14804 5779 14807
rect 7742 14804 7748 14816
rect 5767 14776 7748 14804
rect 5767 14773 5779 14776
rect 5721 14767 5779 14773
rect 7742 14764 7748 14776
rect 7800 14764 7806 14816
rect 8202 14804 8208 14816
rect 8163 14776 8208 14804
rect 8202 14764 8208 14776
rect 8260 14764 8266 14816
rect 9950 14764 9956 14816
rect 10008 14804 10014 14816
rect 12526 14804 12532 14816
rect 10008 14776 12532 14804
rect 10008 14764 10014 14776
rect 12526 14764 12532 14776
rect 12584 14764 12590 14816
rect 14476 14813 14504 14844
rect 14550 14832 14556 14844
rect 14608 14872 14614 14884
rect 15534 14875 15592 14881
rect 15534 14872 15546 14875
rect 14608 14844 15546 14872
rect 14608 14832 14614 14844
rect 15534 14841 15546 14844
rect 15580 14872 15592 14875
rect 17328 14872 17356 14980
rect 19429 14977 19441 14980
rect 19475 14977 19487 15011
rect 19429 14971 19487 14977
rect 19242 14900 19248 14952
rect 19300 14940 19306 14952
rect 19337 14943 19395 14949
rect 19337 14940 19349 14943
rect 19300 14912 19349 14940
rect 19300 14900 19306 14912
rect 19337 14909 19349 14912
rect 19383 14909 19395 14943
rect 19337 14903 19395 14909
rect 20533 14943 20591 14949
rect 20533 14909 20545 14943
rect 20579 14909 20591 14943
rect 20533 14903 20591 14909
rect 15580 14844 17356 14872
rect 15580 14841 15592 14844
rect 15534 14835 15592 14841
rect 17494 14832 17500 14884
rect 17552 14872 17558 14884
rect 20548 14872 20576 14903
rect 17552 14844 20576 14872
rect 17552 14832 17558 14844
rect 14461 14807 14519 14813
rect 14461 14773 14473 14807
rect 14507 14773 14519 14807
rect 14461 14767 14519 14773
rect 16114 14764 16120 14816
rect 16172 14804 16178 14816
rect 16482 14804 16488 14816
rect 16172 14776 16488 14804
rect 16172 14764 16178 14776
rect 16482 14764 16488 14776
rect 16540 14804 16546 14816
rect 16669 14807 16727 14813
rect 16669 14804 16681 14807
rect 16540 14776 16681 14804
rect 16540 14764 16546 14776
rect 16669 14773 16681 14776
rect 16715 14773 16727 14807
rect 16669 14767 16727 14773
rect 18690 14764 18696 14816
rect 18748 14804 18754 14816
rect 18877 14807 18935 14813
rect 18877 14804 18889 14807
rect 18748 14776 18889 14804
rect 18748 14764 18754 14776
rect 18877 14773 18889 14776
rect 18923 14773 18935 14807
rect 19242 14804 19248 14816
rect 19203 14776 19248 14804
rect 18877 14767 18935 14773
rect 19242 14764 19248 14776
rect 19300 14764 19306 14816
rect 1104 14714 21896 14736
rect 1104 14662 7912 14714
rect 7964 14662 7976 14714
rect 8028 14662 8040 14714
rect 8092 14662 8104 14714
rect 8156 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 15035 14714
rect 15087 14662 21896 14714
rect 1104 14640 21896 14662
rect 2777 14603 2835 14609
rect 2777 14569 2789 14603
rect 2823 14600 2835 14603
rect 3418 14600 3424 14612
rect 2823 14572 3424 14600
rect 2823 14569 2835 14572
rect 2777 14563 2835 14569
rect 3418 14560 3424 14572
rect 3476 14560 3482 14612
rect 7190 14600 7196 14612
rect 4264 14572 4476 14600
rect 7151 14572 7196 14600
rect 1397 14535 1455 14541
rect 1397 14501 1409 14535
rect 1443 14532 1455 14535
rect 4264 14532 4292 14572
rect 1443 14504 4292 14532
rect 4448 14532 4476 14572
rect 7190 14560 7196 14572
rect 7248 14600 7254 14612
rect 7650 14600 7656 14612
rect 7248 14572 7656 14600
rect 7248 14560 7254 14572
rect 7650 14560 7656 14572
rect 7708 14560 7714 14612
rect 8021 14603 8079 14609
rect 8021 14569 8033 14603
rect 8067 14600 8079 14603
rect 8294 14600 8300 14612
rect 8067 14572 8300 14600
rect 8067 14569 8079 14572
rect 8021 14563 8079 14569
rect 8294 14560 8300 14572
rect 8352 14560 8358 14612
rect 9858 14600 9864 14612
rect 9819 14572 9864 14600
rect 9858 14560 9864 14572
rect 9916 14560 9922 14612
rect 12434 14600 12440 14612
rect 12395 14572 12440 14600
rect 12434 14560 12440 14572
rect 12492 14560 12498 14612
rect 13725 14603 13783 14609
rect 13725 14569 13737 14603
rect 13771 14600 13783 14603
rect 14642 14600 14648 14612
rect 13771 14572 14648 14600
rect 13771 14569 13783 14572
rect 13725 14563 13783 14569
rect 14642 14560 14648 14572
rect 14700 14600 14706 14612
rect 15378 14600 15384 14612
rect 14700 14572 15384 14600
rect 14700 14560 14706 14572
rect 15378 14560 15384 14572
rect 15436 14560 15442 14612
rect 16206 14560 16212 14612
rect 16264 14600 16270 14612
rect 19242 14600 19248 14612
rect 16264 14572 19248 14600
rect 16264 14560 16270 14572
rect 19242 14560 19248 14572
rect 19300 14560 19306 14612
rect 19610 14560 19616 14612
rect 19668 14560 19674 14612
rect 8389 14535 8447 14541
rect 8389 14532 8401 14535
rect 4448 14504 8401 14532
rect 1443 14501 1455 14504
rect 1397 14495 1455 14501
rect 8389 14501 8401 14504
rect 8435 14501 8447 14535
rect 13633 14535 13691 14541
rect 13633 14532 13645 14535
rect 8389 14495 8447 14501
rect 9048 14504 13645 14532
rect 2869 14467 2927 14473
rect 2869 14433 2881 14467
rect 2915 14464 2927 14467
rect 3142 14464 3148 14476
rect 2915 14436 3148 14464
rect 2915 14433 2927 14436
rect 2869 14427 2927 14433
rect 3142 14424 3148 14436
rect 3200 14464 3206 14476
rect 3510 14464 3516 14476
rect 3200 14436 3516 14464
rect 3200 14424 3206 14436
rect 3510 14424 3516 14436
rect 3568 14424 3574 14476
rect 4433 14467 4491 14473
rect 4433 14433 4445 14467
rect 4479 14464 4491 14467
rect 4798 14464 4804 14476
rect 4479 14436 4804 14464
rect 4479 14433 4491 14436
rect 4433 14427 4491 14433
rect 4798 14424 4804 14436
rect 4856 14424 4862 14476
rect 6080 14467 6138 14473
rect 6080 14433 6092 14467
rect 6126 14464 6138 14467
rect 6362 14464 6368 14476
rect 6126 14436 6368 14464
rect 6126 14433 6138 14436
rect 6080 14427 6138 14433
rect 6362 14424 6368 14436
rect 6420 14424 6426 14476
rect 7742 14424 7748 14476
rect 7800 14464 7806 14476
rect 9048 14464 9076 14504
rect 13633 14501 13645 14504
rect 13679 14501 13691 14535
rect 13633 14495 13691 14501
rect 15556 14535 15614 14541
rect 15556 14501 15568 14535
rect 15602 14532 15614 14535
rect 16666 14532 16672 14544
rect 15602 14504 16672 14532
rect 15602 14501 15614 14504
rect 15556 14495 15614 14501
rect 16666 14492 16672 14504
rect 16724 14492 16730 14544
rect 19426 14532 19432 14544
rect 18432 14504 19432 14532
rect 7800 14436 9076 14464
rect 7800 14424 7806 14436
rect 9306 14424 9312 14476
rect 9364 14464 9370 14476
rect 11330 14473 11336 14476
rect 9677 14467 9735 14473
rect 9677 14464 9689 14467
rect 9364 14436 9689 14464
rect 9364 14424 9370 14436
rect 9677 14433 9689 14436
rect 9723 14433 9735 14467
rect 11324 14464 11336 14473
rect 11291 14436 11336 14464
rect 9677 14427 9735 14433
rect 11324 14427 11336 14436
rect 11330 14424 11336 14427
rect 11388 14424 11394 14476
rect 13814 14424 13820 14476
rect 13872 14464 13878 14476
rect 15013 14467 15071 14473
rect 15013 14464 15025 14467
rect 13872 14436 15025 14464
rect 13872 14424 13878 14436
rect 15013 14433 15025 14436
rect 15059 14433 15071 14467
rect 15286 14464 15292 14476
rect 15199 14436 15292 14464
rect 15013 14427 15071 14433
rect 15286 14424 15292 14436
rect 15344 14464 15350 14476
rect 17126 14464 17132 14476
rect 15344 14436 17132 14464
rect 15344 14424 15350 14436
rect 17126 14424 17132 14436
rect 17184 14424 17190 14476
rect 18432 14473 18460 14504
rect 19426 14492 19432 14504
rect 19484 14492 19490 14544
rect 19628 14532 19656 14560
rect 19797 14535 19855 14541
rect 19797 14532 19809 14535
rect 19628 14504 19809 14532
rect 19797 14501 19809 14504
rect 19843 14501 19855 14535
rect 19797 14495 19855 14501
rect 18417 14467 18475 14473
rect 18417 14433 18429 14467
rect 18463 14433 18475 14467
rect 18417 14427 18475 14433
rect 19334 14424 19340 14476
rect 19392 14424 19398 14476
rect 19531 14467 19589 14473
rect 19531 14433 19543 14467
rect 19577 14464 19589 14467
rect 19577 14436 19656 14464
rect 19577 14433 19589 14436
rect 19531 14427 19589 14433
rect 2130 14356 2136 14408
rect 2188 14396 2194 14408
rect 3053 14399 3111 14405
rect 3053 14396 3065 14399
rect 2188 14368 3065 14396
rect 2188 14356 2194 14368
rect 3053 14365 3065 14368
rect 3099 14396 3111 14399
rect 3694 14396 3700 14408
rect 3099 14368 3700 14396
rect 3099 14365 3111 14368
rect 3053 14359 3111 14365
rect 3694 14356 3700 14368
rect 3752 14356 3758 14408
rect 4154 14356 4160 14408
rect 4212 14396 4218 14408
rect 4525 14399 4583 14405
rect 4525 14396 4537 14399
rect 4212 14368 4537 14396
rect 4212 14356 4218 14368
rect 4525 14365 4537 14368
rect 4571 14365 4583 14399
rect 4525 14359 4583 14365
rect 4617 14399 4675 14405
rect 4617 14365 4629 14399
rect 4663 14365 4675 14399
rect 4617 14359 4675 14365
rect 3970 14288 3976 14340
rect 4028 14328 4034 14340
rect 4632 14328 4660 14359
rect 5350 14356 5356 14408
rect 5408 14396 5414 14408
rect 5813 14399 5871 14405
rect 5813 14396 5825 14399
rect 5408 14368 5825 14396
rect 5408 14356 5414 14368
rect 5813 14365 5825 14368
rect 5859 14365 5871 14399
rect 5813 14359 5871 14365
rect 4028 14300 4660 14328
rect 4028 14288 4034 14300
rect 2406 14260 2412 14272
rect 2367 14232 2412 14260
rect 2406 14220 2412 14232
rect 2464 14220 2470 14272
rect 4062 14260 4068 14272
rect 4023 14232 4068 14260
rect 4062 14220 4068 14232
rect 4120 14220 4126 14272
rect 5828 14260 5856 14359
rect 6914 14356 6920 14408
rect 6972 14396 6978 14408
rect 8481 14399 8539 14405
rect 8481 14396 8493 14399
rect 6972 14368 8493 14396
rect 6972 14356 6978 14368
rect 8481 14365 8493 14368
rect 8527 14365 8539 14399
rect 8481 14359 8539 14365
rect 8570 14356 8576 14408
rect 8628 14396 8634 14408
rect 11057 14399 11115 14405
rect 8628 14368 8673 14396
rect 8628 14356 8634 14368
rect 11057 14365 11069 14399
rect 11103 14365 11115 14399
rect 11057 14359 11115 14365
rect 6546 14260 6552 14272
rect 5828 14232 6552 14260
rect 6546 14220 6552 14232
rect 6604 14220 6610 14272
rect 11072 14260 11100 14359
rect 12158 14356 12164 14408
rect 12216 14396 12222 14408
rect 12618 14396 12624 14408
rect 12216 14368 12624 14396
rect 12216 14356 12222 14368
rect 12618 14356 12624 14368
rect 12676 14356 12682 14408
rect 12894 14356 12900 14408
rect 12952 14396 12958 14408
rect 13262 14396 13268 14408
rect 12952 14368 13268 14396
rect 12952 14356 12958 14368
rect 13262 14356 13268 14368
rect 13320 14356 13326 14408
rect 13909 14399 13967 14405
rect 13909 14365 13921 14399
rect 13955 14396 13967 14399
rect 13955 14368 14044 14396
rect 13955 14365 13967 14368
rect 13909 14359 13967 14365
rect 12158 14260 12164 14272
rect 11072 14232 12164 14260
rect 12158 14220 12164 14232
rect 12216 14220 12222 14272
rect 12618 14220 12624 14272
rect 12676 14260 12682 14272
rect 13265 14263 13323 14269
rect 13265 14260 13277 14263
rect 12676 14232 13277 14260
rect 12676 14220 12682 14232
rect 13265 14229 13277 14232
rect 13311 14229 13323 14263
rect 13265 14223 13323 14229
rect 13446 14220 13452 14272
rect 13504 14260 13510 14272
rect 14016 14260 14044 14368
rect 14829 14331 14887 14337
rect 14829 14297 14841 14331
rect 14875 14328 14887 14331
rect 15304 14328 15332 14424
rect 19352 14396 19380 14424
rect 19426 14396 19432 14408
rect 19352 14368 19432 14396
rect 19426 14356 19432 14368
rect 19484 14356 19490 14408
rect 14875 14300 15332 14328
rect 14875 14297 14887 14300
rect 14829 14291 14887 14297
rect 19334 14288 19340 14340
rect 19392 14328 19398 14340
rect 19628 14328 19656 14436
rect 19392 14300 19656 14328
rect 19392 14288 19398 14300
rect 16022 14260 16028 14272
rect 13504 14232 16028 14260
rect 13504 14220 13510 14232
rect 16022 14220 16028 14232
rect 16080 14260 16086 14272
rect 16669 14263 16727 14269
rect 16669 14260 16681 14263
rect 16080 14232 16681 14260
rect 16080 14220 16086 14232
rect 16669 14229 16681 14232
rect 16715 14229 16727 14263
rect 18598 14260 18604 14272
rect 18559 14232 18604 14260
rect 16669 14223 16727 14229
rect 18598 14220 18604 14232
rect 18656 14220 18662 14272
rect 1104 14170 21896 14192
rect 1104 14118 4447 14170
rect 4499 14118 4511 14170
rect 4563 14118 4575 14170
rect 4627 14118 4639 14170
rect 4691 14118 11378 14170
rect 11430 14118 11442 14170
rect 11494 14118 11506 14170
rect 11558 14118 11570 14170
rect 11622 14118 18308 14170
rect 18360 14118 18372 14170
rect 18424 14118 18436 14170
rect 18488 14118 18500 14170
rect 18552 14118 21896 14170
rect 1104 14096 21896 14118
rect 1670 14056 1676 14068
rect 1631 14028 1676 14056
rect 1670 14016 1676 14028
rect 1728 14016 1734 14068
rect 3326 14056 3332 14068
rect 2608 14028 3332 14056
rect 2608 13929 2636 14028
rect 3326 14016 3332 14028
rect 3384 14016 3390 14068
rect 4798 14056 4804 14068
rect 4759 14028 4804 14056
rect 4798 14016 4804 14028
rect 4856 14016 4862 14068
rect 6362 14016 6368 14068
rect 6420 14056 6426 14068
rect 6420 14028 8800 14056
rect 6420 14016 6426 14028
rect 6270 13948 6276 14000
rect 6328 13988 6334 14000
rect 6328 13960 8340 13988
rect 6328 13948 6334 13960
rect 2593 13923 2651 13929
rect 2593 13889 2605 13923
rect 2639 13889 2651 13923
rect 5353 13923 5411 13929
rect 5353 13920 5365 13923
rect 2593 13883 2651 13889
rect 3712 13892 5365 13920
rect 1486 13852 1492 13864
rect 1447 13824 1492 13852
rect 1486 13812 1492 13824
rect 1544 13812 1550 13864
rect 2860 13855 2918 13861
rect 2860 13821 2872 13855
rect 2906 13852 2918 13855
rect 3712 13852 3740 13892
rect 5353 13889 5365 13892
rect 5399 13889 5411 13923
rect 5353 13883 5411 13889
rect 7469 13923 7527 13929
rect 7469 13889 7481 13923
rect 7515 13920 7527 13923
rect 8202 13920 8208 13932
rect 7515 13892 8208 13920
rect 7515 13889 7527 13892
rect 7469 13883 7527 13889
rect 8202 13880 8208 13892
rect 8260 13880 8266 13932
rect 5258 13852 5264 13864
rect 2906 13824 3740 13852
rect 5219 13824 5264 13852
rect 2906 13821 2918 13824
rect 2860 13815 2918 13821
rect 2976 13796 3004 13824
rect 5258 13812 5264 13824
rect 5316 13812 5322 13864
rect 6549 13855 6607 13861
rect 6549 13821 6561 13855
rect 6595 13852 6607 13855
rect 7742 13852 7748 13864
rect 6595 13824 7748 13852
rect 6595 13821 6607 13824
rect 6549 13815 6607 13821
rect 7742 13812 7748 13824
rect 7800 13812 7806 13864
rect 8312 13852 8340 13960
rect 8772 13920 8800 14028
rect 8938 14016 8944 14068
rect 8996 14056 9002 14068
rect 8996 14028 11376 14056
rect 8996 14016 9002 14028
rect 8941 13923 8999 13929
rect 8941 13920 8953 13923
rect 8772 13892 8953 13920
rect 8941 13889 8953 13892
rect 8987 13889 8999 13923
rect 8941 13883 8999 13889
rect 9398 13880 9404 13932
rect 9456 13920 9462 13932
rect 10137 13923 10195 13929
rect 10137 13920 10149 13923
rect 9456 13892 10149 13920
rect 9456 13880 9462 13892
rect 10137 13889 10149 13892
rect 10183 13889 10195 13923
rect 10137 13883 10195 13889
rect 11348 13852 11376 14028
rect 13722 14016 13728 14068
rect 13780 14056 13786 14068
rect 17494 14056 17500 14068
rect 13780 14028 17500 14056
rect 13780 14016 13786 14028
rect 17494 14016 17500 14028
rect 17552 14016 17558 14068
rect 18138 14016 18144 14068
rect 18196 14056 18202 14068
rect 18233 14059 18291 14065
rect 18233 14056 18245 14059
rect 18196 14028 18245 14056
rect 18196 14016 18202 14028
rect 18233 14025 18245 14028
rect 18279 14025 18291 14059
rect 18233 14019 18291 14025
rect 11514 13988 11520 14000
rect 11475 13960 11520 13988
rect 11514 13948 11520 13960
rect 11572 13948 11578 14000
rect 12894 13948 12900 14000
rect 12952 13988 12958 14000
rect 14001 13991 14059 13997
rect 14001 13988 14013 13991
rect 12952 13960 14013 13988
rect 12952 13948 12958 13960
rect 14001 13957 14013 13960
rect 14047 13957 14059 13991
rect 14001 13951 14059 13957
rect 16114 13948 16120 14000
rect 16172 13988 16178 14000
rect 16172 13960 18828 13988
rect 16172 13948 16178 13960
rect 12434 13880 12440 13932
rect 12492 13920 12498 13932
rect 12989 13923 13047 13929
rect 12989 13920 13001 13923
rect 12492 13892 13001 13920
rect 12492 13880 12498 13892
rect 12989 13889 13001 13892
rect 13035 13889 13047 13923
rect 14550 13920 14556 13932
rect 14511 13892 14556 13920
rect 12989 13883 13047 13889
rect 14550 13880 14556 13892
rect 14608 13880 14614 13932
rect 16206 13880 16212 13932
rect 16264 13920 16270 13932
rect 16393 13923 16451 13929
rect 16393 13920 16405 13923
rect 16264 13892 16405 13920
rect 16264 13880 16270 13892
rect 16393 13889 16405 13892
rect 16439 13889 16451 13923
rect 16393 13883 16451 13889
rect 16485 13923 16543 13929
rect 16485 13889 16497 13923
rect 16531 13920 16543 13923
rect 16666 13920 16672 13932
rect 16531 13892 16672 13920
rect 16531 13889 16543 13892
rect 16485 13883 16543 13889
rect 16666 13880 16672 13892
rect 16724 13880 16730 13932
rect 18690 13920 18696 13932
rect 18651 13892 18696 13920
rect 18690 13880 18696 13892
rect 18748 13880 18754 13932
rect 18800 13929 18828 13960
rect 18785 13923 18843 13929
rect 18785 13889 18797 13923
rect 18831 13889 18843 13923
rect 18785 13883 18843 13889
rect 13906 13852 13912 13864
rect 8312 13824 10364 13852
rect 11348 13824 13912 13852
rect 2958 13744 2964 13796
rect 3016 13744 3022 13796
rect 6914 13744 6920 13796
rect 6972 13784 6978 13796
rect 7558 13784 7564 13796
rect 6972 13756 7564 13784
rect 6972 13744 6978 13756
rect 7558 13744 7564 13756
rect 7616 13784 7622 13796
rect 8202 13784 8208 13796
rect 7616 13756 8208 13784
rect 7616 13744 7622 13756
rect 8202 13744 8208 13756
rect 8260 13744 8266 13796
rect 8754 13784 8760 13796
rect 8667 13756 8760 13784
rect 8754 13744 8760 13756
rect 8812 13784 8818 13796
rect 9122 13784 9128 13796
rect 8812 13756 9128 13784
rect 8812 13744 8818 13756
rect 9122 13744 9128 13756
rect 9180 13744 9186 13796
rect 3326 13676 3332 13728
rect 3384 13716 3390 13728
rect 3970 13716 3976 13728
rect 3384 13688 3976 13716
rect 3384 13676 3390 13688
rect 3970 13676 3976 13688
rect 4028 13676 4034 13728
rect 4982 13676 4988 13728
rect 5040 13716 5046 13728
rect 5169 13719 5227 13725
rect 5169 13716 5181 13719
rect 5040 13688 5181 13716
rect 5040 13676 5046 13688
rect 5169 13685 5181 13688
rect 5215 13685 5227 13719
rect 5169 13679 5227 13685
rect 6365 13719 6423 13725
rect 6365 13685 6377 13719
rect 6411 13716 6423 13719
rect 6546 13716 6552 13728
rect 6411 13688 6552 13716
rect 6411 13685 6423 13688
rect 6365 13679 6423 13685
rect 6546 13676 6552 13688
rect 6604 13676 6610 13728
rect 6638 13676 6644 13728
rect 6696 13716 6702 13728
rect 6825 13719 6883 13725
rect 6825 13716 6837 13719
rect 6696 13688 6837 13716
rect 6696 13676 6702 13688
rect 6825 13685 6837 13688
rect 6871 13685 6883 13719
rect 7190 13716 7196 13728
rect 7151 13688 7196 13716
rect 6825 13679 6883 13685
rect 7190 13676 7196 13688
rect 7248 13676 7254 13728
rect 7282 13676 7288 13728
rect 7340 13716 7346 13728
rect 8386 13716 8392 13728
rect 7340 13688 7385 13716
rect 8347 13688 8392 13716
rect 7340 13676 7346 13688
rect 8386 13676 8392 13688
rect 8444 13676 8450 13728
rect 8849 13719 8907 13725
rect 8849 13685 8861 13719
rect 8895 13716 8907 13719
rect 8938 13716 8944 13728
rect 8895 13688 8944 13716
rect 8895 13685 8907 13688
rect 8849 13679 8907 13685
rect 8938 13676 8944 13688
rect 8996 13676 9002 13728
rect 10336 13716 10364 13824
rect 13906 13812 13912 13824
rect 13964 13812 13970 13864
rect 14461 13855 14519 13861
rect 14461 13821 14473 13855
rect 14507 13852 14519 13855
rect 15286 13852 15292 13864
rect 14507 13824 15292 13852
rect 14507 13821 14519 13824
rect 14461 13815 14519 13821
rect 15286 13812 15292 13824
rect 15344 13812 15350 13864
rect 16301 13855 16359 13861
rect 16301 13852 16313 13855
rect 16224 13824 16313 13852
rect 16224 13796 16252 13824
rect 16301 13821 16313 13824
rect 16347 13852 16359 13855
rect 17954 13852 17960 13864
rect 16347 13824 17960 13852
rect 16347 13821 16359 13824
rect 16301 13815 16359 13821
rect 17954 13812 17960 13824
rect 18012 13812 18018 13864
rect 19242 13812 19248 13864
rect 19300 13852 19306 13864
rect 19978 13852 19984 13864
rect 19300 13824 19984 13852
rect 19300 13812 19306 13824
rect 19978 13812 19984 13824
rect 20036 13812 20042 13864
rect 20346 13812 20352 13864
rect 20404 13852 20410 13864
rect 20533 13855 20591 13861
rect 20533 13852 20545 13855
rect 20404 13824 20545 13852
rect 20404 13812 20410 13824
rect 20533 13821 20545 13824
rect 20579 13821 20591 13855
rect 20533 13815 20591 13821
rect 10404 13787 10462 13793
rect 10404 13753 10416 13787
rect 10450 13784 10462 13787
rect 10594 13784 10600 13796
rect 10450 13756 10600 13784
rect 10450 13753 10462 13756
rect 10404 13747 10462 13753
rect 10594 13744 10600 13756
rect 10652 13744 10658 13796
rect 10778 13744 10784 13796
rect 10836 13784 10842 13796
rect 14369 13787 14427 13793
rect 14369 13784 14381 13787
rect 10836 13756 14381 13784
rect 10836 13744 10842 13756
rect 14369 13753 14381 13756
rect 14415 13753 14427 13787
rect 14369 13747 14427 13753
rect 16206 13744 16212 13796
rect 16264 13744 16270 13796
rect 18601 13787 18659 13793
rect 18601 13753 18613 13787
rect 18647 13784 18659 13787
rect 18782 13784 18788 13796
rect 18647 13756 18788 13784
rect 18647 13753 18659 13756
rect 18601 13747 18659 13753
rect 18782 13744 18788 13756
rect 18840 13744 18846 13796
rect 12437 13719 12495 13725
rect 12437 13716 12449 13719
rect 10336 13688 12449 13716
rect 12437 13685 12449 13688
rect 12483 13685 12495 13719
rect 12802 13716 12808 13728
rect 12763 13688 12808 13716
rect 12437 13679 12495 13685
rect 12802 13676 12808 13688
rect 12860 13676 12866 13728
rect 12894 13676 12900 13728
rect 12952 13716 12958 13728
rect 15930 13716 15936 13728
rect 12952 13688 12997 13716
rect 15891 13688 15936 13716
rect 12952 13676 12958 13688
rect 15930 13676 15936 13688
rect 15988 13676 15994 13728
rect 20714 13716 20720 13728
rect 20675 13688 20720 13716
rect 20714 13676 20720 13688
rect 20772 13676 20778 13728
rect 1104 13626 21896 13648
rect 1104 13574 7912 13626
rect 7964 13574 7976 13626
rect 8028 13574 8040 13626
rect 8092 13574 8104 13626
rect 8156 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 15035 13626
rect 15087 13574 21896 13626
rect 1104 13552 21896 13574
rect 2869 13515 2927 13521
rect 2869 13481 2881 13515
rect 2915 13512 2927 13515
rect 4062 13512 4068 13524
rect 2915 13484 4068 13512
rect 2915 13481 2927 13484
rect 2869 13475 2927 13481
rect 4062 13472 4068 13484
rect 4120 13472 4126 13524
rect 5905 13515 5963 13521
rect 5905 13481 5917 13515
rect 5951 13512 5963 13515
rect 6914 13512 6920 13524
rect 5951 13484 6920 13512
rect 5951 13481 5963 13484
rect 5905 13475 5963 13481
rect 6914 13472 6920 13484
rect 6972 13472 6978 13524
rect 7101 13515 7159 13521
rect 7101 13481 7113 13515
rect 7147 13512 7159 13515
rect 7282 13512 7288 13524
rect 7147 13484 7288 13512
rect 7147 13481 7159 13484
rect 7101 13475 7159 13481
rect 7282 13472 7288 13484
rect 7340 13472 7346 13524
rect 7469 13515 7527 13521
rect 7469 13481 7481 13515
rect 7515 13512 7527 13515
rect 8386 13512 8392 13524
rect 7515 13484 8392 13512
rect 7515 13481 7527 13484
rect 7469 13475 7527 13481
rect 8386 13472 8392 13484
rect 8444 13472 8450 13524
rect 8478 13472 8484 13524
rect 8536 13512 8542 13524
rect 8662 13512 8668 13524
rect 8536 13484 8668 13512
rect 8536 13472 8542 13484
rect 8662 13472 8668 13484
rect 8720 13512 8726 13524
rect 9398 13512 9404 13524
rect 8720 13484 9404 13512
rect 8720 13472 8726 13484
rect 9398 13472 9404 13484
rect 9456 13472 9462 13524
rect 9490 13472 9496 13524
rect 9548 13512 9554 13524
rect 9677 13515 9735 13521
rect 9677 13512 9689 13515
rect 9548 13484 9689 13512
rect 9548 13472 9554 13484
rect 9677 13481 9689 13484
rect 9723 13481 9735 13515
rect 9677 13475 9735 13481
rect 11146 13472 11152 13524
rect 11204 13512 11210 13524
rect 11241 13515 11299 13521
rect 11241 13512 11253 13515
rect 11204 13484 11253 13512
rect 11204 13472 11210 13484
rect 11241 13481 11253 13484
rect 11287 13481 11299 13515
rect 11241 13475 11299 13481
rect 12253 13515 12311 13521
rect 12253 13481 12265 13515
rect 12299 13512 12311 13515
rect 12802 13512 12808 13524
rect 12299 13484 12808 13512
rect 12299 13481 12311 13484
rect 12253 13475 12311 13481
rect 12802 13472 12808 13484
rect 12860 13472 12866 13524
rect 12986 13472 12992 13524
rect 13044 13512 13050 13524
rect 13354 13512 13360 13524
rect 13044 13484 13360 13512
rect 13044 13472 13050 13484
rect 13354 13472 13360 13484
rect 13412 13472 13418 13524
rect 15286 13512 15292 13524
rect 15247 13484 15292 13512
rect 15286 13472 15292 13484
rect 15344 13472 15350 13524
rect 15749 13515 15807 13521
rect 15749 13481 15761 13515
rect 15795 13512 15807 13515
rect 15930 13512 15936 13524
rect 15795 13484 15936 13512
rect 15795 13481 15807 13484
rect 15749 13475 15807 13481
rect 15930 13472 15936 13484
rect 15988 13472 15994 13524
rect 19150 13512 19156 13524
rect 17788 13484 19156 13512
rect 4890 13444 4896 13456
rect 3068 13416 4896 13444
rect 2314 13336 2320 13388
rect 2372 13376 2378 13388
rect 2777 13379 2835 13385
rect 2777 13376 2789 13379
rect 2372 13348 2789 13376
rect 2372 13336 2378 13348
rect 2777 13345 2789 13348
rect 2823 13345 2835 13379
rect 2777 13339 2835 13345
rect 3068 13317 3096 13416
rect 4890 13404 4896 13416
rect 4948 13404 4954 13456
rect 5350 13404 5356 13456
rect 5408 13444 5414 13456
rect 10045 13447 10103 13453
rect 10045 13444 10057 13447
rect 5408 13416 10057 13444
rect 5408 13404 5414 13416
rect 10045 13413 10057 13416
rect 10091 13413 10103 13447
rect 12618 13444 12624 13456
rect 12579 13416 12624 13444
rect 10045 13407 10103 13413
rect 12618 13404 12624 13416
rect 12676 13404 12682 13456
rect 14185 13447 14243 13453
rect 14185 13413 14197 13447
rect 14231 13444 14243 13447
rect 17788 13444 17816 13484
rect 19150 13472 19156 13484
rect 19208 13472 19214 13524
rect 14231 13416 17816 13444
rect 14231 13413 14243 13416
rect 14185 13407 14243 13413
rect 17862 13404 17868 13456
rect 17920 13444 17926 13456
rect 19337 13447 19395 13453
rect 19337 13444 19349 13447
rect 17920 13416 19349 13444
rect 17920 13404 17926 13416
rect 19337 13413 19349 13416
rect 19383 13413 19395 13447
rect 19337 13407 19395 13413
rect 4065 13379 4123 13385
rect 4065 13376 4077 13379
rect 3436 13348 4077 13376
rect 1397 13311 1455 13317
rect 1397 13277 1409 13311
rect 1443 13277 1455 13311
rect 1397 13271 1455 13277
rect 3053 13311 3111 13317
rect 3053 13277 3065 13311
rect 3099 13277 3111 13311
rect 3053 13271 3111 13277
rect 1412 13172 1440 13271
rect 2409 13243 2467 13249
rect 2409 13209 2421 13243
rect 2455 13240 2467 13243
rect 3436 13240 3464 13348
rect 4065 13345 4077 13348
rect 4111 13345 4123 13379
rect 4065 13339 4123 13345
rect 5810 13336 5816 13388
rect 5868 13376 5874 13388
rect 5997 13379 6055 13385
rect 5997 13376 6009 13379
rect 5868 13348 6009 13376
rect 5868 13336 5874 13348
rect 5997 13345 6009 13348
rect 6043 13376 6055 13379
rect 6546 13376 6552 13388
rect 6043 13348 6552 13376
rect 6043 13345 6055 13348
rect 5997 13339 6055 13345
rect 6546 13336 6552 13348
rect 6604 13336 6610 13388
rect 7742 13336 7748 13388
rect 7800 13376 7806 13388
rect 8849 13379 8907 13385
rect 8849 13376 8861 13379
rect 7800 13348 8861 13376
rect 7800 13336 7806 13348
rect 8849 13345 8861 13348
rect 8895 13345 8907 13379
rect 8849 13339 8907 13345
rect 10137 13379 10195 13385
rect 10137 13345 10149 13379
rect 10183 13376 10195 13379
rect 12894 13376 12900 13388
rect 10183 13348 12900 13376
rect 10183 13345 10195 13348
rect 10137 13339 10195 13345
rect 12894 13336 12900 13348
rect 12952 13336 12958 13388
rect 13906 13376 13912 13388
rect 13867 13348 13912 13376
rect 13906 13336 13912 13348
rect 13964 13336 13970 13388
rect 15657 13379 15715 13385
rect 15657 13345 15669 13379
rect 15703 13376 15715 13379
rect 15930 13376 15936 13388
rect 15703 13348 15936 13376
rect 15703 13345 15715 13348
rect 15657 13339 15715 13345
rect 15930 13336 15936 13348
rect 15988 13336 15994 13388
rect 17681 13379 17739 13385
rect 17681 13345 17693 13379
rect 17727 13376 17739 13379
rect 18046 13376 18052 13388
rect 17727 13348 18052 13376
rect 17727 13345 17739 13348
rect 17681 13339 17739 13345
rect 18046 13336 18052 13348
rect 18104 13336 18110 13388
rect 19242 13376 19248 13388
rect 19203 13348 19248 13376
rect 19242 13336 19248 13348
rect 19300 13336 19306 13388
rect 3878 13268 3884 13320
rect 3936 13308 3942 13320
rect 4249 13311 4307 13317
rect 4249 13308 4261 13311
rect 3936 13280 4261 13308
rect 3936 13268 3942 13280
rect 4249 13277 4261 13280
rect 4295 13277 4307 13311
rect 4249 13271 4307 13277
rect 6086 13268 6092 13320
rect 6144 13308 6150 13320
rect 6181 13311 6239 13317
rect 6181 13308 6193 13311
rect 6144 13280 6193 13308
rect 6144 13268 6150 13280
rect 6181 13277 6193 13280
rect 6227 13308 6239 13311
rect 6362 13308 6368 13320
rect 6227 13280 6368 13308
rect 6227 13277 6239 13280
rect 6181 13271 6239 13277
rect 6362 13268 6368 13280
rect 6420 13268 6426 13320
rect 7561 13311 7619 13317
rect 7561 13277 7573 13311
rect 7607 13277 7619 13311
rect 7561 13271 7619 13277
rect 2455 13212 3464 13240
rect 5537 13243 5595 13249
rect 2455 13209 2467 13212
rect 2409 13203 2467 13209
rect 5537 13209 5549 13243
rect 5583 13240 5595 13243
rect 7576 13240 7604 13271
rect 7650 13268 7656 13320
rect 7708 13308 7714 13320
rect 7708 13280 7753 13308
rect 7708 13268 7714 13280
rect 8570 13268 8576 13320
rect 8628 13308 8634 13320
rect 9582 13308 9588 13320
rect 8628 13280 9588 13308
rect 8628 13268 8634 13280
rect 9582 13268 9588 13280
rect 9640 13308 9646 13320
rect 10229 13311 10287 13317
rect 10229 13308 10241 13311
rect 9640 13280 10241 13308
rect 9640 13268 9646 13280
rect 10229 13277 10241 13280
rect 10275 13277 10287 13311
rect 10229 13271 10287 13277
rect 12434 13268 12440 13320
rect 12492 13308 12498 13320
rect 12713 13311 12771 13317
rect 12713 13308 12725 13311
rect 12492 13280 12725 13308
rect 12492 13268 12498 13280
rect 12713 13277 12725 13280
rect 12759 13277 12771 13311
rect 12713 13271 12771 13277
rect 12805 13311 12863 13317
rect 12805 13277 12817 13311
rect 12851 13308 12863 13311
rect 14550 13308 14556 13320
rect 12851 13280 14556 13308
rect 12851 13277 12863 13280
rect 12805 13271 12863 13277
rect 5583 13212 7604 13240
rect 5583 13209 5595 13212
rect 5537 13203 5595 13209
rect 11514 13200 11520 13252
rect 11572 13240 11578 13252
rect 12820 13240 12848 13271
rect 14550 13268 14556 13280
rect 14608 13268 14614 13320
rect 15841 13311 15899 13317
rect 15841 13277 15853 13311
rect 15887 13308 15899 13311
rect 16022 13308 16028 13320
rect 15887 13280 16028 13308
rect 15887 13277 15899 13280
rect 15841 13271 15899 13277
rect 16022 13268 16028 13280
rect 16080 13268 16086 13320
rect 17494 13268 17500 13320
rect 17552 13308 17558 13320
rect 17770 13308 17776 13320
rect 17552 13280 17776 13308
rect 17552 13268 17558 13280
rect 17770 13268 17776 13280
rect 17828 13268 17834 13320
rect 17954 13308 17960 13320
rect 17915 13280 17960 13308
rect 17954 13268 17960 13280
rect 18012 13268 18018 13320
rect 19429 13311 19487 13317
rect 19429 13277 19441 13311
rect 19475 13277 19487 13311
rect 19429 13271 19487 13277
rect 11572 13212 12848 13240
rect 11572 13200 11578 13212
rect 18782 13200 18788 13252
rect 18840 13240 18846 13252
rect 19444 13240 19472 13271
rect 18840 13212 19472 13240
rect 18840 13200 18846 13212
rect 7006 13172 7012 13184
rect 1412 13144 7012 13172
rect 7006 13132 7012 13144
rect 7064 13132 7070 13184
rect 11790 13132 11796 13184
rect 11848 13172 11854 13184
rect 15102 13172 15108 13184
rect 11848 13144 15108 13172
rect 11848 13132 11854 13144
rect 15102 13132 15108 13144
rect 15160 13132 15166 13184
rect 15378 13132 15384 13184
rect 15436 13172 15442 13184
rect 17313 13175 17371 13181
rect 17313 13172 17325 13175
rect 15436 13144 17325 13172
rect 15436 13132 15442 13144
rect 17313 13141 17325 13144
rect 17359 13141 17371 13175
rect 17313 13135 17371 13141
rect 18690 13132 18696 13184
rect 18748 13172 18754 13184
rect 18877 13175 18935 13181
rect 18877 13172 18889 13175
rect 18748 13144 18889 13172
rect 18748 13132 18754 13144
rect 18877 13141 18889 13144
rect 18923 13141 18935 13175
rect 18877 13135 18935 13141
rect 1104 13082 21896 13104
rect 1104 13030 4447 13082
rect 4499 13030 4511 13082
rect 4563 13030 4575 13082
rect 4627 13030 4639 13082
rect 4691 13030 11378 13082
rect 11430 13030 11442 13082
rect 11494 13030 11506 13082
rect 11558 13030 11570 13082
rect 11622 13030 18308 13082
rect 18360 13030 18372 13082
rect 18424 13030 18436 13082
rect 18488 13030 18500 13082
rect 18552 13030 21896 13082
rect 1104 13008 21896 13030
rect 2314 12968 2320 12980
rect 2275 12940 2320 12968
rect 2314 12928 2320 12940
rect 2372 12928 2378 12980
rect 3142 12928 3148 12980
rect 3200 12968 3206 12980
rect 4065 12971 4123 12977
rect 4065 12968 4077 12971
rect 3200 12940 4077 12968
rect 3200 12928 3206 12940
rect 4065 12937 4077 12940
rect 4111 12937 4123 12971
rect 4982 12968 4988 12980
rect 4943 12940 4988 12968
rect 4065 12931 4123 12937
rect 4982 12928 4988 12940
rect 5040 12928 5046 12980
rect 6825 12971 6883 12977
rect 6825 12937 6837 12971
rect 6871 12968 6883 12971
rect 7190 12968 7196 12980
rect 6871 12940 7196 12968
rect 6871 12937 6883 12940
rect 6825 12931 6883 12937
rect 7190 12928 7196 12940
rect 7248 12928 7254 12980
rect 7742 12928 7748 12980
rect 7800 12968 7806 12980
rect 8389 12971 8447 12977
rect 8389 12968 8401 12971
rect 7800 12940 8401 12968
rect 7800 12928 7806 12940
rect 8389 12937 8401 12940
rect 8435 12937 8447 12971
rect 9214 12968 9220 12980
rect 9175 12940 9220 12968
rect 8389 12931 8447 12937
rect 9214 12928 9220 12940
rect 9272 12928 9278 12980
rect 10778 12968 10784 12980
rect 10739 12940 10784 12968
rect 10778 12928 10784 12940
rect 10836 12928 10842 12980
rect 11790 12928 11796 12980
rect 11848 12968 11854 12980
rect 11974 12968 11980 12980
rect 11848 12940 11980 12968
rect 11848 12928 11854 12940
rect 11974 12928 11980 12940
rect 12032 12928 12038 12980
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 12492 12940 12537 12968
rect 12492 12928 12498 12940
rect 12710 12928 12716 12980
rect 12768 12968 12774 12980
rect 13722 12968 13728 12980
rect 12768 12940 13728 12968
rect 12768 12928 12774 12940
rect 13722 12928 13728 12940
rect 13780 12928 13786 12980
rect 13814 12928 13820 12980
rect 13872 12968 13878 12980
rect 14001 12971 14059 12977
rect 14001 12968 14013 12971
rect 13872 12940 14013 12968
rect 13872 12928 13878 12940
rect 14001 12937 14013 12940
rect 14047 12937 14059 12971
rect 15930 12968 15936 12980
rect 15891 12940 15936 12968
rect 14001 12931 14059 12937
rect 15930 12928 15936 12940
rect 15988 12928 15994 12980
rect 17310 12928 17316 12980
rect 17368 12968 17374 12980
rect 18598 12968 18604 12980
rect 17368 12940 18604 12968
rect 17368 12928 17374 12940
rect 18598 12928 18604 12940
rect 18656 12928 18662 12980
rect 10594 12860 10600 12912
rect 10652 12900 10658 12912
rect 10652 12872 13032 12900
rect 10652 12860 10658 12872
rect 2961 12835 3019 12841
rect 2961 12801 2973 12835
rect 3007 12832 3019 12835
rect 3326 12832 3332 12844
rect 3007 12804 3332 12832
rect 3007 12801 3019 12804
rect 2961 12795 3019 12801
rect 3326 12792 3332 12804
rect 3384 12792 3390 12844
rect 5626 12832 5632 12844
rect 5587 12804 5632 12832
rect 5626 12792 5632 12804
rect 5684 12792 5690 12844
rect 7469 12835 7527 12841
rect 7469 12801 7481 12835
rect 7515 12832 7527 12835
rect 7650 12832 7656 12844
rect 7515 12804 7656 12832
rect 7515 12801 7527 12804
rect 7469 12795 7527 12801
rect 7650 12792 7656 12804
rect 7708 12792 7714 12844
rect 8496 12804 9536 12832
rect 3142 12724 3148 12776
rect 3200 12764 3206 12776
rect 3418 12764 3424 12776
rect 3200 12736 3424 12764
rect 3200 12724 3206 12736
rect 3418 12724 3424 12736
rect 3476 12724 3482 12776
rect 3881 12767 3939 12773
rect 3881 12733 3893 12767
rect 3927 12764 3939 12767
rect 8496 12764 8524 12804
rect 3927 12736 8524 12764
rect 8573 12767 8631 12773
rect 3927 12733 3939 12736
rect 3881 12727 3939 12733
rect 8573 12733 8585 12767
rect 8619 12764 8631 12767
rect 9030 12764 9036 12776
rect 8619 12736 9036 12764
rect 8619 12733 8631 12736
rect 8573 12727 8631 12733
rect 9030 12724 9036 12736
rect 9088 12724 9094 12776
rect 9508 12764 9536 12804
rect 9582 12792 9588 12844
rect 9640 12832 9646 12844
rect 11440 12841 11468 12872
rect 9769 12835 9827 12841
rect 9769 12832 9781 12835
rect 9640 12804 9781 12832
rect 9640 12792 9646 12804
rect 9769 12801 9781 12804
rect 9815 12801 9827 12835
rect 9769 12795 9827 12801
rect 11425 12835 11483 12841
rect 11425 12801 11437 12835
rect 11471 12801 11483 12835
rect 12710 12832 12716 12844
rect 11425 12795 11483 12801
rect 12544 12804 12716 12832
rect 10134 12764 10140 12776
rect 9508 12736 10140 12764
rect 10134 12724 10140 12736
rect 10192 12724 10198 12776
rect 2498 12656 2504 12708
rect 2556 12696 2562 12708
rect 2777 12699 2835 12705
rect 2777 12696 2789 12699
rect 2556 12668 2789 12696
rect 2556 12656 2562 12668
rect 2777 12665 2789 12668
rect 2823 12665 2835 12699
rect 2777 12659 2835 12665
rect 4062 12656 4068 12708
rect 4120 12696 4126 12708
rect 8478 12696 8484 12708
rect 4120 12668 8484 12696
rect 4120 12656 4126 12668
rect 8478 12656 8484 12668
rect 8536 12656 8542 12708
rect 9306 12656 9312 12708
rect 9364 12696 9370 12708
rect 9677 12699 9735 12705
rect 9677 12696 9689 12699
rect 9364 12668 9689 12696
rect 9364 12656 9370 12668
rect 9677 12665 9689 12668
rect 9723 12696 9735 12699
rect 11241 12699 11299 12705
rect 11241 12696 11253 12699
rect 9723 12668 11253 12696
rect 9723 12665 9735 12668
rect 9677 12659 9735 12665
rect 11241 12665 11253 12668
rect 11287 12665 11299 12699
rect 12544 12696 12572 12804
rect 12710 12792 12716 12804
rect 12768 12792 12774 12844
rect 12894 12832 12900 12844
rect 12855 12804 12900 12832
rect 12894 12792 12900 12804
rect 12952 12792 12958 12844
rect 13004 12841 13032 12872
rect 13078 12860 13084 12912
rect 13136 12900 13142 12912
rect 14369 12903 14427 12909
rect 14369 12900 14381 12903
rect 13136 12872 14381 12900
rect 13136 12860 13142 12872
rect 14369 12869 14381 12872
rect 14415 12869 14427 12903
rect 14369 12863 14427 12869
rect 12989 12835 13047 12841
rect 12989 12801 13001 12835
rect 13035 12832 13047 12835
rect 13446 12832 13452 12844
rect 13035 12804 13452 12832
rect 13035 12801 13047 12804
rect 12989 12795 13047 12801
rect 13446 12792 13452 12804
rect 13504 12792 13510 12844
rect 14550 12792 14556 12844
rect 14608 12832 14614 12844
rect 14921 12835 14979 12841
rect 14921 12832 14933 12835
rect 14608 12804 14933 12832
rect 14608 12792 14614 12804
rect 14921 12801 14933 12804
rect 14967 12801 14979 12835
rect 14921 12795 14979 12801
rect 16485 12835 16543 12841
rect 16485 12801 16497 12835
rect 16531 12832 16543 12835
rect 16666 12832 16672 12844
rect 16531 12804 16672 12832
rect 16531 12801 16543 12804
rect 16485 12795 16543 12801
rect 16666 12792 16672 12804
rect 16724 12792 16730 12844
rect 17126 12792 17132 12844
rect 17184 12832 17190 12844
rect 18785 12835 18843 12841
rect 18785 12832 18797 12835
rect 17184 12804 18797 12832
rect 17184 12792 17190 12804
rect 18785 12801 18797 12804
rect 18831 12801 18843 12835
rect 18785 12795 18843 12801
rect 12618 12724 12624 12776
rect 12676 12764 12682 12776
rect 14185 12767 14243 12773
rect 14185 12764 14197 12767
rect 12676 12736 14197 12764
rect 12676 12724 12682 12736
rect 14185 12733 14197 12736
rect 14231 12733 14243 12767
rect 14185 12727 14243 12733
rect 14829 12767 14887 12773
rect 14829 12733 14841 12767
rect 14875 12764 14887 12767
rect 15194 12764 15200 12776
rect 14875 12736 15200 12764
rect 14875 12733 14887 12736
rect 14829 12727 14887 12733
rect 12805 12699 12863 12705
rect 12805 12696 12817 12699
rect 12544 12668 12817 12696
rect 11241 12659 11299 12665
rect 12805 12665 12817 12668
rect 12851 12665 12863 12699
rect 12805 12659 12863 12665
rect 12986 12656 12992 12708
rect 13044 12696 13050 12708
rect 14737 12699 14795 12705
rect 14737 12696 14749 12699
rect 13044 12668 14749 12696
rect 13044 12656 13050 12668
rect 14737 12665 14749 12668
rect 14783 12665 14795 12699
rect 14737 12659 14795 12665
rect 2682 12628 2688 12640
rect 2643 12600 2688 12628
rect 2682 12588 2688 12600
rect 2740 12588 2746 12640
rect 4890 12588 4896 12640
rect 4948 12628 4954 12640
rect 5350 12628 5356 12640
rect 4948 12600 5356 12628
rect 4948 12588 4954 12600
rect 5350 12588 5356 12600
rect 5408 12588 5414 12640
rect 5445 12631 5503 12637
rect 5445 12597 5457 12631
rect 5491 12628 5503 12631
rect 6362 12628 6368 12640
rect 5491 12600 6368 12628
rect 5491 12597 5503 12600
rect 5445 12591 5503 12597
rect 6362 12588 6368 12600
rect 6420 12588 6426 12640
rect 7098 12588 7104 12640
rect 7156 12628 7162 12640
rect 7193 12631 7251 12637
rect 7193 12628 7205 12631
rect 7156 12600 7205 12628
rect 7156 12588 7162 12600
rect 7193 12597 7205 12600
rect 7239 12597 7251 12631
rect 7193 12591 7251 12597
rect 7282 12588 7288 12640
rect 7340 12628 7346 12640
rect 7340 12600 7385 12628
rect 7340 12588 7346 12600
rect 9214 12588 9220 12640
rect 9272 12628 9278 12640
rect 9585 12631 9643 12637
rect 9585 12628 9597 12631
rect 9272 12600 9597 12628
rect 9272 12588 9278 12600
rect 9585 12597 9597 12600
rect 9631 12628 9643 12631
rect 11149 12631 11207 12637
rect 11149 12628 11161 12631
rect 9631 12600 11161 12628
rect 9631 12597 9643 12600
rect 9585 12591 9643 12597
rect 11149 12597 11161 12600
rect 11195 12597 11207 12631
rect 11149 12591 11207 12597
rect 12158 12588 12164 12640
rect 12216 12628 12222 12640
rect 12894 12628 12900 12640
rect 12216 12600 12900 12628
rect 12216 12588 12222 12600
rect 12894 12588 12900 12600
rect 12952 12588 12958 12640
rect 13814 12588 13820 12640
rect 13872 12628 13878 12640
rect 14844 12628 14872 12727
rect 15194 12724 15200 12736
rect 15252 12764 15258 12776
rect 15838 12764 15844 12776
rect 15252 12736 15844 12764
rect 15252 12724 15258 12736
rect 15838 12724 15844 12736
rect 15896 12724 15902 12776
rect 16301 12767 16359 12773
rect 16301 12733 16313 12767
rect 16347 12764 16359 12767
rect 17586 12764 17592 12776
rect 16347 12736 17592 12764
rect 16347 12733 16359 12736
rect 16301 12727 16359 12733
rect 17586 12724 17592 12736
rect 17644 12724 17650 12776
rect 16393 12699 16451 12705
rect 16393 12665 16405 12699
rect 16439 12696 16451 12699
rect 16758 12696 16764 12708
rect 16439 12668 16764 12696
rect 16439 12665 16451 12668
rect 16393 12659 16451 12665
rect 16758 12656 16764 12668
rect 16816 12696 16822 12708
rect 17678 12696 17684 12708
rect 16816 12668 17684 12696
rect 16816 12656 16822 12668
rect 17678 12656 17684 12668
rect 17736 12656 17742 12708
rect 19058 12705 19064 12708
rect 19052 12659 19064 12705
rect 19116 12696 19122 12708
rect 19116 12668 19152 12696
rect 19058 12656 19064 12659
rect 19116 12656 19122 12668
rect 13872 12600 14872 12628
rect 13872 12588 13878 12600
rect 17310 12588 17316 12640
rect 17368 12628 17374 12640
rect 17494 12628 17500 12640
rect 17368 12600 17500 12628
rect 17368 12588 17374 12600
rect 17494 12588 17500 12600
rect 17552 12588 17558 12640
rect 17770 12588 17776 12640
rect 17828 12628 17834 12640
rect 18138 12628 18144 12640
rect 17828 12600 18144 12628
rect 17828 12588 17834 12600
rect 18138 12588 18144 12600
rect 18196 12588 18202 12640
rect 18782 12588 18788 12640
rect 18840 12628 18846 12640
rect 20165 12631 20223 12637
rect 20165 12628 20177 12631
rect 18840 12600 20177 12628
rect 18840 12588 18846 12600
rect 20165 12597 20177 12600
rect 20211 12597 20223 12631
rect 20165 12591 20223 12597
rect 1104 12538 21896 12560
rect 1104 12486 7912 12538
rect 7964 12486 7976 12538
rect 8028 12486 8040 12538
rect 8092 12486 8104 12538
rect 8156 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 15035 12538
rect 15087 12486 21896 12538
rect 1104 12464 21896 12486
rect 2406 12384 2412 12436
rect 2464 12424 2470 12436
rect 2685 12427 2743 12433
rect 2685 12424 2697 12427
rect 2464 12396 2697 12424
rect 2464 12384 2470 12396
rect 2685 12393 2697 12396
rect 2731 12393 2743 12427
rect 2685 12387 2743 12393
rect 5445 12427 5503 12433
rect 5445 12393 5457 12427
rect 5491 12424 5503 12427
rect 5534 12424 5540 12436
rect 5491 12396 5540 12424
rect 5491 12393 5503 12396
rect 5445 12387 5503 12393
rect 5534 12384 5540 12396
rect 5592 12424 5598 12436
rect 6914 12424 6920 12436
rect 5592 12396 6920 12424
rect 5592 12384 5598 12396
rect 6914 12384 6920 12396
rect 6972 12384 6978 12436
rect 7006 12384 7012 12436
rect 7064 12424 7070 12436
rect 7193 12427 7251 12433
rect 7193 12424 7205 12427
rect 7064 12396 7205 12424
rect 7064 12384 7070 12396
rect 7193 12393 7205 12396
rect 7239 12393 7251 12427
rect 11238 12424 11244 12436
rect 7193 12387 7251 12393
rect 7300 12396 11244 12424
rect 3878 12316 3884 12368
rect 3936 12356 3942 12368
rect 7300 12356 7328 12396
rect 11238 12384 11244 12396
rect 11296 12384 11302 12436
rect 12253 12427 12311 12433
rect 12253 12424 12265 12427
rect 11992 12396 12265 12424
rect 11992 12368 12020 12396
rect 12253 12393 12265 12396
rect 12299 12424 12311 12427
rect 12526 12424 12532 12436
rect 12299 12396 12532 12424
rect 12299 12393 12311 12396
rect 12253 12387 12311 12393
rect 12526 12384 12532 12396
rect 12584 12384 12590 12436
rect 13538 12384 13544 12436
rect 13596 12424 13602 12436
rect 13817 12427 13875 12433
rect 13817 12424 13829 12427
rect 13596 12396 13829 12424
rect 13596 12384 13602 12396
rect 13817 12393 13829 12396
rect 13863 12393 13875 12427
rect 13817 12387 13875 12393
rect 14734 12384 14740 12436
rect 14792 12424 14798 12436
rect 15657 12427 15715 12433
rect 15657 12424 15669 12427
rect 14792 12396 15669 12424
rect 14792 12384 14798 12396
rect 15657 12393 15669 12396
rect 15703 12393 15715 12427
rect 15657 12387 15715 12393
rect 16574 12384 16580 12436
rect 16632 12424 16638 12436
rect 17862 12424 17868 12436
rect 16632 12396 17868 12424
rect 16632 12384 16638 12396
rect 17862 12384 17868 12396
rect 17920 12384 17926 12436
rect 19886 12424 19892 12436
rect 19847 12396 19892 12424
rect 19886 12384 19892 12396
rect 19944 12384 19950 12436
rect 3936 12328 7328 12356
rect 3936 12316 3942 12328
rect 7650 12316 7656 12368
rect 7708 12356 7714 12368
rect 10045 12359 10103 12365
rect 10045 12356 10057 12359
rect 7708 12328 10057 12356
rect 7708 12316 7714 12328
rect 10045 12325 10057 12328
rect 10091 12325 10103 12359
rect 10045 12319 10103 12325
rect 11974 12316 11980 12368
rect 12032 12316 12038 12368
rect 13354 12316 13360 12368
rect 13412 12356 13418 12368
rect 13909 12359 13967 12365
rect 13909 12356 13921 12359
rect 13412 12328 13921 12356
rect 13412 12316 13418 12328
rect 13909 12325 13921 12328
rect 13955 12325 13967 12359
rect 13909 12319 13967 12325
rect 14366 12316 14372 12368
rect 14424 12356 14430 12368
rect 15749 12359 15807 12365
rect 15749 12356 15761 12359
rect 14424 12328 15761 12356
rect 14424 12316 14430 12328
rect 15749 12325 15761 12328
rect 15795 12325 15807 12359
rect 15749 12319 15807 12325
rect 18966 12316 18972 12368
rect 19024 12356 19030 12368
rect 19978 12356 19984 12368
rect 19024 12328 19984 12356
rect 19024 12316 19030 12328
rect 19978 12316 19984 12328
rect 20036 12316 20042 12368
rect 2593 12291 2651 12297
rect 2593 12257 2605 12291
rect 2639 12288 2651 12291
rect 4065 12291 4123 12297
rect 4065 12288 4077 12291
rect 2639 12260 4077 12288
rect 2639 12257 2651 12260
rect 2593 12251 2651 12257
rect 4065 12257 4077 12260
rect 4111 12257 4123 12291
rect 4065 12251 4123 12257
rect 6086 12248 6092 12300
rect 6144 12288 6150 12300
rect 6730 12288 6736 12300
rect 6144 12260 6736 12288
rect 6144 12248 6150 12260
rect 6730 12248 6736 12260
rect 6788 12288 6794 12300
rect 8481 12291 8539 12297
rect 8481 12288 8493 12291
rect 6788 12260 7420 12288
rect 6788 12248 6794 12260
rect 2869 12223 2927 12229
rect 2869 12189 2881 12223
rect 2915 12220 2927 12223
rect 2958 12220 2964 12232
rect 2915 12192 2964 12220
rect 2915 12189 2927 12192
rect 2869 12183 2927 12189
rect 2958 12180 2964 12192
rect 3016 12180 3022 12232
rect 5166 12180 5172 12232
rect 5224 12220 5230 12232
rect 5537 12223 5595 12229
rect 5537 12220 5549 12223
rect 5224 12192 5549 12220
rect 5224 12180 5230 12192
rect 5537 12189 5549 12192
rect 5583 12189 5595 12223
rect 5537 12183 5595 12189
rect 5629 12223 5687 12229
rect 5629 12189 5641 12223
rect 5675 12189 5687 12223
rect 5629 12183 5687 12189
rect 2225 12155 2283 12161
rect 2225 12121 2237 12155
rect 2271 12152 2283 12155
rect 2682 12152 2688 12164
rect 2271 12124 2688 12152
rect 2271 12121 2283 12124
rect 2225 12115 2283 12121
rect 2682 12112 2688 12124
rect 2740 12112 2746 12164
rect 4062 12112 4068 12164
rect 4120 12152 4126 12164
rect 4120 12124 5212 12152
rect 4120 12112 4126 12124
rect 2314 12044 2320 12096
rect 2372 12084 2378 12096
rect 5077 12087 5135 12093
rect 5077 12084 5089 12087
rect 2372 12056 5089 12084
rect 2372 12044 2378 12056
rect 5077 12053 5089 12056
rect 5123 12053 5135 12087
rect 5184 12084 5212 12124
rect 5442 12112 5448 12164
rect 5500 12152 5506 12164
rect 5644 12152 5672 12183
rect 7006 12180 7012 12232
rect 7064 12220 7070 12232
rect 7392 12229 7420 12260
rect 7668 12260 8493 12288
rect 7285 12223 7343 12229
rect 7285 12220 7297 12223
rect 7064 12192 7297 12220
rect 7064 12180 7070 12192
rect 7285 12189 7297 12192
rect 7331 12189 7343 12223
rect 7285 12183 7343 12189
rect 7377 12223 7435 12229
rect 7377 12189 7389 12223
rect 7423 12189 7435 12223
rect 7377 12183 7435 12189
rect 5500 12124 5672 12152
rect 6825 12155 6883 12161
rect 5500 12112 5506 12124
rect 6825 12121 6837 12155
rect 6871 12152 6883 12155
rect 7098 12152 7104 12164
rect 6871 12124 7104 12152
rect 6871 12121 6883 12124
rect 6825 12115 6883 12121
rect 7098 12112 7104 12124
rect 7156 12112 7162 12164
rect 7190 12112 7196 12164
rect 7248 12152 7254 12164
rect 7668 12152 7696 12260
rect 8481 12257 8493 12260
rect 8527 12288 8539 12291
rect 9950 12288 9956 12300
rect 8527 12260 9956 12288
rect 8527 12257 8539 12260
rect 8481 12251 8539 12257
rect 9950 12248 9956 12260
rect 10008 12248 10014 12300
rect 14182 12288 14188 12300
rect 10336 12260 14188 12288
rect 7742 12180 7748 12232
rect 7800 12220 7806 12232
rect 10336 12229 10364 12260
rect 10137 12223 10195 12229
rect 10137 12220 10149 12223
rect 7800 12192 10149 12220
rect 7800 12180 7806 12192
rect 10137 12189 10149 12192
rect 10183 12189 10195 12223
rect 10137 12183 10195 12189
rect 10321 12223 10379 12229
rect 10321 12189 10333 12223
rect 10367 12189 10379 12223
rect 10321 12183 10379 12189
rect 10686 12180 10692 12232
rect 10744 12220 10750 12232
rect 12452 12229 12480 12260
rect 14182 12248 14188 12260
rect 14240 12288 14246 12300
rect 14550 12288 14556 12300
rect 14240 12260 14556 12288
rect 14240 12248 14246 12260
rect 14550 12248 14556 12260
rect 14608 12248 14614 12300
rect 17126 12288 17132 12300
rect 17087 12260 17132 12288
rect 17126 12248 17132 12260
rect 17184 12248 17190 12300
rect 17218 12248 17224 12300
rect 17276 12288 17282 12300
rect 17385 12291 17443 12297
rect 17385 12288 17397 12291
rect 17276 12260 17397 12288
rect 17276 12248 17282 12260
rect 17385 12257 17397 12260
rect 17431 12257 17443 12291
rect 19702 12288 19708 12300
rect 19663 12260 19708 12288
rect 17385 12251 17443 12257
rect 19702 12248 19708 12260
rect 19760 12248 19766 12300
rect 12345 12223 12403 12229
rect 12345 12220 12357 12223
rect 10744 12192 12357 12220
rect 10744 12180 10750 12192
rect 12345 12189 12357 12192
rect 12391 12189 12403 12223
rect 12345 12183 12403 12189
rect 12437 12223 12495 12229
rect 12437 12189 12449 12223
rect 12483 12189 12495 12223
rect 13998 12220 14004 12232
rect 13959 12192 14004 12220
rect 12437 12183 12495 12189
rect 13998 12180 14004 12192
rect 14056 12180 14062 12232
rect 15933 12223 15991 12229
rect 15933 12189 15945 12223
rect 15979 12220 15991 12223
rect 16114 12220 16120 12232
rect 15979 12192 16120 12220
rect 15979 12189 15991 12192
rect 15933 12183 15991 12189
rect 16114 12180 16120 12192
rect 16172 12180 16178 12232
rect 7248 12124 7696 12152
rect 9677 12155 9735 12161
rect 7248 12112 7254 12124
rect 9677 12121 9689 12155
rect 9723 12152 9735 12155
rect 13449 12155 13507 12161
rect 9723 12124 13308 12152
rect 9723 12121 9735 12124
rect 9677 12115 9735 12121
rect 8386 12084 8392 12096
rect 5184 12056 8392 12084
rect 5077 12047 5135 12053
rect 8386 12044 8392 12056
rect 8444 12044 8450 12096
rect 8665 12087 8723 12093
rect 8665 12053 8677 12087
rect 8711 12084 8723 12087
rect 10502 12084 10508 12096
rect 8711 12056 10508 12084
rect 8711 12053 8723 12056
rect 8665 12047 8723 12053
rect 10502 12044 10508 12056
rect 10560 12044 10566 12096
rect 11885 12087 11943 12093
rect 11885 12053 11897 12087
rect 11931 12084 11943 12087
rect 12526 12084 12532 12096
rect 11931 12056 12532 12084
rect 11931 12053 11943 12056
rect 11885 12047 11943 12053
rect 12526 12044 12532 12056
rect 12584 12044 12590 12096
rect 12618 12044 12624 12096
rect 12676 12084 12682 12096
rect 12802 12084 12808 12096
rect 12676 12056 12808 12084
rect 12676 12044 12682 12056
rect 12802 12044 12808 12056
rect 12860 12044 12866 12096
rect 13280 12084 13308 12124
rect 13449 12121 13461 12155
rect 13495 12152 13507 12155
rect 13906 12152 13912 12164
rect 13495 12124 13912 12152
rect 13495 12121 13507 12124
rect 13449 12115 13507 12121
rect 13906 12112 13912 12124
rect 13964 12112 13970 12164
rect 14090 12084 14096 12096
rect 13280 12056 14096 12084
rect 14090 12044 14096 12056
rect 14148 12044 14154 12096
rect 15289 12087 15347 12093
rect 15289 12053 15301 12087
rect 15335 12084 15347 12087
rect 16298 12084 16304 12096
rect 15335 12056 16304 12084
rect 15335 12053 15347 12056
rect 15289 12047 15347 12053
rect 16298 12044 16304 12056
rect 16356 12044 16362 12096
rect 18046 12044 18052 12096
rect 18104 12084 18110 12096
rect 18509 12087 18567 12093
rect 18509 12084 18521 12087
rect 18104 12056 18521 12084
rect 18104 12044 18110 12056
rect 18509 12053 18521 12056
rect 18555 12084 18567 12087
rect 19058 12084 19064 12096
rect 18555 12056 19064 12084
rect 18555 12053 18567 12056
rect 18509 12047 18567 12053
rect 19058 12044 19064 12056
rect 19116 12044 19122 12096
rect 1104 11994 21896 12016
rect 1104 11942 4447 11994
rect 4499 11942 4511 11994
rect 4563 11942 4575 11994
rect 4627 11942 4639 11994
rect 4691 11942 11378 11994
rect 11430 11942 11442 11994
rect 11494 11942 11506 11994
rect 11558 11942 11570 11994
rect 11622 11942 18308 11994
rect 18360 11942 18372 11994
rect 18424 11942 18436 11994
rect 18488 11942 18500 11994
rect 18552 11942 21896 11994
rect 1104 11920 21896 11942
rect 2406 11840 2412 11892
rect 2464 11880 2470 11892
rect 3421 11883 3479 11889
rect 3421 11880 3433 11883
rect 2464 11852 3433 11880
rect 2464 11840 2470 11852
rect 3421 11849 3433 11852
rect 3467 11849 3479 11883
rect 3421 11843 3479 11849
rect 4985 11883 5043 11889
rect 4985 11849 4997 11883
rect 5031 11880 5043 11883
rect 5258 11880 5264 11892
rect 5031 11852 5264 11880
rect 5031 11849 5043 11852
rect 4985 11843 5043 11849
rect 5258 11840 5264 11852
rect 5316 11840 5322 11892
rect 7282 11840 7288 11892
rect 7340 11880 7346 11892
rect 7377 11883 7435 11889
rect 7377 11880 7389 11883
rect 7340 11852 7389 11880
rect 7340 11840 7346 11852
rect 7377 11849 7389 11852
rect 7423 11849 7435 11883
rect 10594 11880 10600 11892
rect 7377 11843 7435 11849
rect 7484 11852 10600 11880
rect 1857 11815 1915 11821
rect 1857 11781 1869 11815
rect 1903 11812 1915 11815
rect 4154 11812 4160 11824
rect 1903 11784 4160 11812
rect 1903 11781 1915 11784
rect 1857 11775 1915 11781
rect 4154 11772 4160 11784
rect 4212 11772 4218 11824
rect 6549 11815 6607 11821
rect 6549 11781 6561 11815
rect 6595 11812 6607 11815
rect 7484 11812 7512 11852
rect 10594 11840 10600 11852
rect 10652 11840 10658 11892
rect 12069 11883 12127 11889
rect 12069 11849 12081 11883
rect 12115 11880 12127 11883
rect 12434 11880 12440 11892
rect 12115 11852 12440 11880
rect 12115 11849 12127 11852
rect 12069 11843 12127 11849
rect 12434 11840 12440 11852
rect 12492 11840 12498 11892
rect 12820 11852 14136 11880
rect 6595 11784 7512 11812
rect 11057 11815 11115 11821
rect 6595 11781 6607 11784
rect 6549 11775 6607 11781
rect 11057 11781 11069 11815
rect 11103 11812 11115 11815
rect 12618 11812 12624 11824
rect 11103 11784 12624 11812
rect 11103 11781 11115 11784
rect 11057 11775 11115 11781
rect 12618 11772 12624 11784
rect 12676 11772 12682 11824
rect 2314 11744 2320 11756
rect 2275 11716 2320 11744
rect 2314 11704 2320 11716
rect 2372 11704 2378 11756
rect 2501 11747 2559 11753
rect 2501 11713 2513 11747
rect 2547 11744 2559 11747
rect 2958 11744 2964 11756
rect 2547 11716 2964 11744
rect 2547 11713 2559 11716
rect 2501 11707 2559 11713
rect 2958 11704 2964 11716
rect 3016 11704 3022 11756
rect 3694 11704 3700 11756
rect 3752 11744 3758 11756
rect 4065 11747 4123 11753
rect 4065 11744 4077 11747
rect 3752 11716 4077 11744
rect 3752 11704 3758 11716
rect 4065 11713 4077 11716
rect 4111 11744 4123 11747
rect 5442 11744 5448 11756
rect 4111 11716 5448 11744
rect 4111 11713 4123 11716
rect 4065 11707 4123 11713
rect 5442 11704 5448 11716
rect 5500 11744 5506 11756
rect 5537 11747 5595 11753
rect 5537 11744 5549 11747
rect 5500 11716 5549 11744
rect 5500 11704 5506 11716
rect 5537 11713 5549 11716
rect 5583 11713 5595 11747
rect 5537 11707 5595 11713
rect 6730 11704 6736 11756
rect 6788 11744 6794 11756
rect 7929 11747 7987 11753
rect 7929 11744 7941 11747
rect 6788 11716 7941 11744
rect 6788 11704 6794 11716
rect 7929 11713 7941 11716
rect 7975 11713 7987 11747
rect 7929 11707 7987 11713
rect 8662 11704 8668 11756
rect 8720 11744 8726 11756
rect 9677 11747 9735 11753
rect 9677 11744 9689 11747
rect 8720 11716 9689 11744
rect 8720 11704 8726 11716
rect 9677 11713 9689 11716
rect 9723 11713 9735 11747
rect 9677 11707 9735 11713
rect 10870 11704 10876 11756
rect 10928 11744 10934 11756
rect 12820 11744 12848 11852
rect 14108 11812 14136 11852
rect 14182 11840 14188 11892
rect 14240 11880 14246 11892
rect 14369 11883 14427 11889
rect 14369 11880 14381 11883
rect 14240 11852 14381 11880
rect 14240 11840 14246 11852
rect 14369 11849 14381 11852
rect 14415 11849 14427 11883
rect 14369 11843 14427 11849
rect 16393 11883 16451 11889
rect 16393 11849 16405 11883
rect 16439 11880 16451 11883
rect 16574 11880 16580 11892
rect 16439 11852 16580 11880
rect 16439 11849 16451 11852
rect 16393 11843 16451 11849
rect 16574 11840 16580 11852
rect 16632 11840 16638 11892
rect 19061 11883 19119 11889
rect 19061 11849 19073 11883
rect 19107 11880 19119 11883
rect 19242 11880 19248 11892
rect 19107 11852 19248 11880
rect 19107 11849 19119 11852
rect 19061 11843 19119 11849
rect 19242 11840 19248 11852
rect 19300 11840 19306 11892
rect 14108 11784 20668 11812
rect 10928 11716 12848 11744
rect 10928 11704 10934 11716
rect 12894 11704 12900 11756
rect 12952 11744 12958 11756
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 12952 11716 13001 11744
rect 12952 11704 12958 11716
rect 12989 11713 13001 11716
rect 13035 11713 13047 11747
rect 12989 11707 13047 11713
rect 17037 11747 17095 11753
rect 17037 11713 17049 11747
rect 17083 11713 17095 11747
rect 17037 11707 17095 11713
rect 1946 11636 1952 11688
rect 2004 11676 2010 11688
rect 2866 11676 2872 11688
rect 2004 11648 2872 11676
rect 2004 11636 2010 11648
rect 2866 11636 2872 11648
rect 2924 11636 2930 11688
rect 3786 11636 3792 11688
rect 3844 11676 3850 11688
rect 9766 11676 9772 11688
rect 3844 11648 9772 11676
rect 3844 11636 3850 11648
rect 9766 11636 9772 11648
rect 9824 11636 9830 11688
rect 9944 11679 10002 11685
rect 9944 11645 9956 11679
rect 9990 11676 10002 11679
rect 10318 11676 10324 11688
rect 9990 11648 10324 11676
rect 9990 11645 10002 11648
rect 9944 11639 10002 11645
rect 10318 11636 10324 11648
rect 10376 11636 10382 11688
rect 10962 11636 10968 11688
rect 11020 11676 11026 11688
rect 12253 11679 12311 11685
rect 12253 11676 12265 11679
rect 11020 11648 12265 11676
rect 11020 11636 11026 11648
rect 12253 11645 12265 11648
rect 12299 11645 12311 11679
rect 12253 11639 12311 11645
rect 15289 11679 15347 11685
rect 15289 11645 15301 11679
rect 15335 11676 15347 11679
rect 16482 11676 16488 11688
rect 15335 11648 16488 11676
rect 15335 11645 15347 11648
rect 15289 11639 15347 11645
rect 16482 11636 16488 11648
rect 16540 11636 16546 11688
rect 17052 11676 17080 11707
rect 17954 11704 17960 11756
rect 18012 11744 18018 11756
rect 18049 11747 18107 11753
rect 18049 11744 18061 11747
rect 18012 11716 18061 11744
rect 18012 11704 18018 11716
rect 18049 11713 18061 11716
rect 18095 11713 18107 11747
rect 18049 11707 18107 11713
rect 19058 11704 19064 11756
rect 19116 11744 19122 11756
rect 20640 11753 20668 11784
rect 19613 11747 19671 11753
rect 19613 11744 19625 11747
rect 19116 11716 19625 11744
rect 19116 11704 19122 11716
rect 19613 11713 19625 11716
rect 19659 11713 19671 11747
rect 19613 11707 19671 11713
rect 20625 11747 20683 11753
rect 20625 11713 20637 11747
rect 20671 11713 20683 11747
rect 20625 11707 20683 11713
rect 17052 11648 18092 11676
rect 18064 11620 18092 11648
rect 19426 11636 19432 11688
rect 19484 11676 19490 11688
rect 19521 11679 19579 11685
rect 19521 11676 19533 11679
rect 19484 11648 19533 11676
rect 19484 11636 19490 11648
rect 19521 11645 19533 11648
rect 19567 11645 19579 11679
rect 19521 11639 19579 11645
rect 2225 11611 2283 11617
rect 2225 11577 2237 11611
rect 2271 11608 2283 11611
rect 2406 11608 2412 11620
rect 2271 11580 2412 11608
rect 2271 11577 2283 11580
rect 2225 11571 2283 11577
rect 2406 11568 2412 11580
rect 2464 11568 2470 11620
rect 3881 11611 3939 11617
rect 3881 11577 3893 11611
rect 3927 11608 3939 11611
rect 4338 11608 4344 11620
rect 3927 11580 4344 11608
rect 3927 11577 3939 11580
rect 3881 11571 3939 11577
rect 4338 11568 4344 11580
rect 4396 11608 4402 11620
rect 4982 11608 4988 11620
rect 4396 11580 4988 11608
rect 4396 11568 4402 11580
rect 4982 11568 4988 11580
rect 5040 11568 5046 11620
rect 5445 11611 5503 11617
rect 5445 11577 5457 11611
rect 5491 11608 5503 11611
rect 6549 11611 6607 11617
rect 6549 11608 6561 11611
rect 5491 11580 6561 11608
rect 5491 11577 5503 11580
rect 5445 11571 5503 11577
rect 6549 11577 6561 11580
rect 6595 11577 6607 11611
rect 6549 11571 6607 11577
rect 8202 11568 8208 11620
rect 8260 11608 8266 11620
rect 13256 11611 13314 11617
rect 8260 11580 13216 11608
rect 8260 11568 8266 11580
rect 3789 11543 3847 11549
rect 3789 11509 3801 11543
rect 3835 11540 3847 11543
rect 4154 11540 4160 11552
rect 3835 11512 4160 11540
rect 3835 11509 3847 11512
rect 3789 11503 3847 11509
rect 4154 11500 4160 11512
rect 4212 11500 4218 11552
rect 4246 11500 4252 11552
rect 4304 11540 4310 11552
rect 4890 11540 4896 11552
rect 4304 11512 4896 11540
rect 4304 11500 4310 11512
rect 4890 11500 4896 11512
rect 4948 11540 4954 11552
rect 5353 11543 5411 11549
rect 5353 11540 5365 11543
rect 4948 11512 5365 11540
rect 4948 11500 4954 11512
rect 5353 11509 5365 11512
rect 5399 11509 5411 11543
rect 5353 11503 5411 11509
rect 6362 11500 6368 11552
rect 6420 11540 6426 11552
rect 7745 11543 7803 11549
rect 7745 11540 7757 11543
rect 6420 11512 7757 11540
rect 6420 11500 6426 11512
rect 7745 11509 7757 11512
rect 7791 11509 7803 11543
rect 7745 11503 7803 11509
rect 7837 11543 7895 11549
rect 7837 11509 7849 11543
rect 7883 11540 7895 11543
rect 11698 11540 11704 11552
rect 7883 11512 11704 11540
rect 7883 11509 7895 11512
rect 7837 11503 7895 11509
rect 11698 11500 11704 11512
rect 11756 11500 11762 11552
rect 13188 11540 13216 11580
rect 13256 11577 13268 11611
rect 13302 11608 13314 11611
rect 13906 11608 13912 11620
rect 13302 11580 13912 11608
rect 13302 11577 13314 11580
rect 13256 11571 13314 11577
rect 13906 11568 13912 11580
rect 13964 11568 13970 11620
rect 16853 11611 16911 11617
rect 16853 11608 16865 11611
rect 15304 11580 16865 11608
rect 15304 11540 15332 11580
rect 16853 11577 16865 11580
rect 16899 11608 16911 11611
rect 16942 11608 16948 11620
rect 16899 11580 16948 11608
rect 16899 11577 16911 11580
rect 16853 11571 16911 11577
rect 16942 11568 16948 11580
rect 17000 11568 17006 11620
rect 18046 11568 18052 11620
rect 18104 11568 18110 11620
rect 13188 11512 15332 11540
rect 15473 11543 15531 11549
rect 15473 11509 15485 11543
rect 15519 11540 15531 11543
rect 16390 11540 16396 11552
rect 15519 11512 16396 11540
rect 15519 11509 15531 11512
rect 15473 11503 15531 11509
rect 16390 11500 16396 11512
rect 16448 11500 16454 11552
rect 16666 11500 16672 11552
rect 16724 11540 16730 11552
rect 16761 11543 16819 11549
rect 16761 11540 16773 11543
rect 16724 11512 16773 11540
rect 16724 11500 16730 11512
rect 16761 11509 16773 11512
rect 16807 11509 16819 11543
rect 19426 11540 19432 11552
rect 19387 11512 19432 11540
rect 16761 11503 16819 11509
rect 19426 11500 19432 11512
rect 19484 11500 19490 11552
rect 1104 11450 21896 11472
rect 1104 11398 7912 11450
rect 7964 11398 7976 11450
rect 8028 11398 8040 11450
rect 8092 11398 8104 11450
rect 8156 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 15035 11450
rect 15087 11398 21896 11450
rect 1104 11376 21896 11398
rect 2409 11339 2467 11345
rect 2409 11305 2421 11339
rect 2455 11336 2467 11339
rect 2498 11336 2504 11348
rect 2455 11308 2504 11336
rect 2455 11305 2467 11308
rect 2409 11299 2467 11305
rect 2498 11296 2504 11308
rect 2556 11296 2562 11348
rect 2774 11296 2780 11348
rect 2832 11336 2838 11348
rect 2832 11308 2877 11336
rect 2832 11296 2838 11308
rect 3418 11296 3424 11348
rect 3476 11336 3482 11348
rect 4062 11336 4068 11348
rect 3476 11308 4068 11336
rect 3476 11296 3482 11308
rect 4062 11296 4068 11308
rect 4120 11296 4126 11348
rect 5442 11296 5448 11348
rect 5500 11336 5506 11348
rect 8757 11339 8815 11345
rect 8757 11336 8769 11339
rect 5500 11308 8769 11336
rect 5500 11296 5506 11308
rect 8757 11305 8769 11308
rect 8803 11305 8815 11339
rect 8757 11299 8815 11305
rect 12434 11296 12440 11348
rect 12492 11336 12498 11348
rect 12894 11336 12900 11348
rect 12492 11308 12900 11336
rect 12492 11296 12498 11308
rect 12894 11296 12900 11308
rect 12952 11296 12958 11348
rect 13633 11339 13691 11345
rect 13633 11305 13645 11339
rect 13679 11336 13691 11339
rect 13998 11336 14004 11348
rect 13679 11308 14004 11336
rect 13679 11305 13691 11308
rect 13633 11299 13691 11305
rect 13998 11296 14004 11308
rect 14056 11296 14062 11348
rect 14090 11296 14096 11348
rect 14148 11336 14154 11348
rect 16945 11339 17003 11345
rect 14148 11308 14193 11336
rect 14148 11296 14154 11308
rect 16945 11305 16957 11339
rect 16991 11336 17003 11339
rect 17218 11336 17224 11348
rect 16991 11308 17224 11336
rect 16991 11305 17003 11308
rect 16945 11299 17003 11305
rect 17218 11296 17224 11308
rect 17276 11296 17282 11348
rect 18138 11296 18144 11348
rect 18196 11336 18202 11348
rect 18233 11339 18291 11345
rect 18233 11336 18245 11339
rect 18196 11308 18245 11336
rect 18196 11296 18202 11308
rect 18233 11305 18245 11308
rect 18279 11305 18291 11339
rect 18233 11299 18291 11305
rect 2866 11268 2872 11280
rect 2827 11240 2872 11268
rect 2866 11228 2872 11240
rect 2924 11228 2930 11280
rect 4341 11271 4399 11277
rect 4341 11237 4353 11271
rect 4387 11268 4399 11271
rect 7006 11268 7012 11280
rect 4387 11240 7012 11268
rect 4387 11237 4399 11240
rect 4341 11231 4399 11237
rect 7006 11228 7012 11240
rect 7064 11228 7070 11280
rect 7558 11228 7564 11280
rect 7616 11277 7622 11280
rect 7616 11271 7680 11277
rect 7616 11237 7634 11271
rect 7668 11237 7680 11271
rect 10410 11268 10416 11280
rect 10371 11240 10416 11268
rect 7616 11231 7680 11237
rect 7616 11228 7622 11231
rect 10410 11228 10416 11240
rect 10468 11228 10474 11280
rect 11698 11228 11704 11280
rect 11756 11268 11762 11280
rect 12066 11268 12072 11280
rect 11756 11240 12072 11268
rect 11756 11228 11762 11240
rect 12066 11228 12072 11240
rect 12124 11228 12130 11280
rect 12520 11271 12578 11277
rect 12520 11237 12532 11271
rect 12566 11268 12578 11271
rect 12618 11268 12624 11280
rect 12566 11240 12624 11268
rect 12566 11237 12578 11240
rect 12520 11231 12578 11237
rect 12618 11228 12624 11240
rect 12676 11228 12682 11280
rect 15746 11228 15752 11280
rect 15804 11268 15810 11280
rect 15804 11240 19564 11268
rect 15804 11228 15810 11240
rect 3418 11160 3424 11212
rect 3476 11200 3482 11212
rect 4065 11203 4123 11209
rect 4065 11200 4077 11203
rect 3476 11172 4077 11200
rect 3476 11160 3482 11172
rect 4065 11169 4077 11172
rect 4111 11169 4123 11203
rect 4065 11163 4123 11169
rect 5166 11160 5172 11212
rect 5224 11200 5230 11212
rect 5721 11203 5779 11209
rect 5721 11200 5733 11203
rect 5224 11172 5733 11200
rect 5224 11160 5230 11172
rect 5721 11169 5733 11172
rect 5767 11169 5779 11203
rect 5721 11163 5779 11169
rect 6638 11160 6644 11212
rect 6696 11200 6702 11212
rect 7377 11203 7435 11209
rect 7377 11200 7389 11203
rect 6696 11172 7389 11200
rect 6696 11160 6702 11172
rect 7377 11169 7389 11172
rect 7423 11169 7435 11203
rect 7377 11163 7435 11169
rect 15470 11160 15476 11212
rect 15528 11200 15534 11212
rect 15832 11203 15890 11209
rect 15832 11200 15844 11203
rect 15528 11172 15844 11200
rect 15528 11160 15534 11172
rect 15832 11169 15844 11172
rect 15878 11200 15890 11203
rect 15878 11172 16988 11200
rect 15878 11169 15890 11172
rect 15832 11163 15890 11169
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11101 1455 11135
rect 2958 11132 2964 11144
rect 2871 11104 2964 11132
rect 1397 11095 1455 11101
rect 1412 10996 1440 11095
rect 2958 11092 2964 11104
rect 3016 11092 3022 11144
rect 5810 11132 5816 11144
rect 5771 11104 5816 11132
rect 5810 11092 5816 11104
rect 5868 11092 5874 11144
rect 5994 11132 6000 11144
rect 5955 11104 6000 11132
rect 5994 11092 6000 11104
rect 6052 11092 6058 11144
rect 12250 11132 12256 11144
rect 12211 11104 12256 11132
rect 12250 11092 12256 11104
rect 12308 11092 12314 11144
rect 13814 11092 13820 11144
rect 13872 11132 13878 11144
rect 14185 11135 14243 11141
rect 14185 11132 14197 11135
rect 13872 11104 14197 11132
rect 13872 11092 13878 11104
rect 14185 11101 14197 11104
rect 14231 11101 14243 11135
rect 14185 11095 14243 11101
rect 14274 11092 14280 11144
rect 14332 11132 14338 11144
rect 14332 11104 14377 11132
rect 14332 11092 14338 11104
rect 15286 11092 15292 11144
rect 15344 11132 15350 11144
rect 15565 11135 15623 11141
rect 15565 11132 15577 11135
rect 15344 11104 15577 11132
rect 15344 11092 15350 11104
rect 15565 11101 15577 11104
rect 15611 11101 15623 11135
rect 16960 11132 16988 11172
rect 17126 11160 17132 11212
rect 17184 11200 17190 11212
rect 19536 11209 19564 11240
rect 19702 11228 19708 11280
rect 19760 11268 19766 11280
rect 19797 11271 19855 11277
rect 19797 11268 19809 11271
rect 19760 11240 19809 11268
rect 19760 11228 19766 11240
rect 19797 11237 19809 11240
rect 19843 11237 19855 11271
rect 19797 11231 19855 11237
rect 18141 11203 18199 11209
rect 18141 11200 18153 11203
rect 17184 11172 18153 11200
rect 17184 11160 17190 11172
rect 18141 11169 18153 11172
rect 18187 11169 18199 11203
rect 18141 11163 18199 11169
rect 19521 11203 19579 11209
rect 19521 11169 19533 11203
rect 19567 11169 19579 11203
rect 19521 11163 19579 11169
rect 18325 11135 18383 11141
rect 18325 11132 18337 11135
rect 16960 11104 18337 11132
rect 15565 11095 15623 11101
rect 18325 11101 18337 11104
rect 18371 11101 18383 11135
rect 18325 11095 18383 11101
rect 2976 11064 3004 11092
rect 3878 11064 3884 11076
rect 2976 11036 3884 11064
rect 3878 11024 3884 11036
rect 3936 11024 3942 11076
rect 5353 11067 5411 11073
rect 5353 11033 5365 11067
rect 5399 11064 5411 11067
rect 5534 11064 5540 11076
rect 5399 11036 5540 11064
rect 5399 11033 5411 11036
rect 5353 11027 5411 11033
rect 5534 11024 5540 11036
rect 5592 11024 5598 11076
rect 10226 11024 10232 11076
rect 10284 11064 10290 11076
rect 10962 11064 10968 11076
rect 10284 11036 10968 11064
rect 10284 11024 10290 11036
rect 10962 11024 10968 11036
rect 11020 11064 11026 11076
rect 11701 11067 11759 11073
rect 11701 11064 11713 11067
rect 11020 11036 11713 11064
rect 11020 11024 11026 11036
rect 11701 11033 11713 11036
rect 11747 11033 11759 11067
rect 11701 11027 11759 11033
rect 13648 11036 13952 11064
rect 4246 10996 4252 11008
rect 1412 10968 4252 10996
rect 4246 10956 4252 10968
rect 4304 10956 4310 11008
rect 6914 10956 6920 11008
rect 6972 10996 6978 11008
rect 13648 10996 13676 11036
rect 6972 10968 13676 10996
rect 6972 10956 6978 10968
rect 13722 10956 13728 11008
rect 13780 10996 13786 11008
rect 13924 10996 13952 11036
rect 18138 11024 18144 11076
rect 18196 11064 18202 11076
rect 18340 11064 18368 11095
rect 18196 11036 18368 11064
rect 18196 11024 18202 11036
rect 14550 10996 14556 11008
rect 13780 10968 13825 10996
rect 13924 10968 14556 10996
rect 13780 10956 13786 10968
rect 14550 10956 14556 10968
rect 14608 10956 14614 11008
rect 17770 10996 17776 11008
rect 17731 10968 17776 10996
rect 17770 10956 17776 10968
rect 17828 10956 17834 11008
rect 1104 10906 21896 10928
rect 1104 10854 4447 10906
rect 4499 10854 4511 10906
rect 4563 10854 4575 10906
rect 4627 10854 4639 10906
rect 4691 10854 11378 10906
rect 11430 10854 11442 10906
rect 11494 10854 11506 10906
rect 11558 10854 11570 10906
rect 11622 10854 18308 10906
rect 18360 10854 18372 10906
rect 18424 10854 18436 10906
rect 18488 10854 18500 10906
rect 18552 10854 21896 10906
rect 1104 10832 21896 10854
rect 5169 10795 5227 10801
rect 5169 10792 5181 10795
rect 1596 10764 5181 10792
rect 1596 10597 1624 10764
rect 5169 10761 5181 10764
rect 5215 10761 5227 10795
rect 7558 10792 7564 10804
rect 5169 10755 5227 10761
rect 5828 10764 7564 10792
rect 3878 10684 3884 10736
rect 3936 10724 3942 10736
rect 4249 10727 4307 10733
rect 4249 10724 4261 10727
rect 3936 10696 4261 10724
rect 3936 10684 3942 10696
rect 4249 10693 4261 10696
rect 4295 10693 4307 10727
rect 4249 10687 4307 10693
rect 5828 10665 5856 10764
rect 7558 10752 7564 10764
rect 7616 10792 7622 10804
rect 8205 10795 8263 10801
rect 8205 10792 8217 10795
rect 7616 10764 8217 10792
rect 7616 10752 7622 10764
rect 8205 10761 8217 10764
rect 8251 10761 8263 10795
rect 8205 10755 8263 10761
rect 8570 10752 8576 10804
rect 8628 10792 8634 10804
rect 12618 10792 12624 10804
rect 8628 10764 12624 10792
rect 8628 10752 8634 10764
rect 12618 10752 12624 10764
rect 12676 10752 12682 10804
rect 13265 10795 13323 10801
rect 13265 10761 13277 10795
rect 13311 10792 13323 10795
rect 18509 10795 18567 10801
rect 13311 10764 17356 10792
rect 13311 10761 13323 10764
rect 13265 10755 13323 10761
rect 5902 10684 5908 10736
rect 5960 10724 5966 10736
rect 6454 10724 6460 10736
rect 5960 10696 6460 10724
rect 5960 10684 5966 10696
rect 6454 10684 6460 10696
rect 6512 10684 6518 10736
rect 7834 10684 7840 10736
rect 7892 10724 7898 10736
rect 11054 10724 11060 10736
rect 7892 10696 11060 10724
rect 7892 10684 7898 10696
rect 11054 10684 11060 10696
rect 11112 10684 11118 10736
rect 14829 10727 14887 10733
rect 14829 10693 14841 10727
rect 14875 10724 14887 10727
rect 14875 10696 16896 10724
rect 14875 10693 14887 10696
rect 14829 10687 14887 10693
rect 5813 10659 5871 10665
rect 5813 10625 5825 10659
rect 5859 10625 5871 10659
rect 5813 10619 5871 10625
rect 9950 10616 9956 10668
rect 10008 10656 10014 10668
rect 10045 10659 10103 10665
rect 10045 10656 10057 10659
rect 10008 10628 10057 10656
rect 10008 10616 10014 10628
rect 10045 10625 10057 10628
rect 10091 10625 10103 10659
rect 10045 10619 10103 10625
rect 10594 10616 10600 10668
rect 10652 10656 10658 10668
rect 11698 10656 11704 10668
rect 10652 10628 11704 10656
rect 10652 10616 10658 10628
rect 11698 10616 11704 10628
rect 11756 10616 11762 10668
rect 13722 10656 13728 10668
rect 13683 10628 13728 10656
rect 13722 10616 13728 10628
rect 13780 10616 13786 10668
rect 13906 10656 13912 10668
rect 13867 10628 13912 10656
rect 13906 10616 13912 10628
rect 13964 10616 13970 10668
rect 15194 10616 15200 10668
rect 15252 10656 15258 10668
rect 16868 10665 16896 10696
rect 15289 10659 15347 10665
rect 15289 10656 15301 10659
rect 15252 10628 15301 10656
rect 15252 10616 15258 10628
rect 15289 10625 15301 10628
rect 15335 10625 15347 10659
rect 15289 10619 15347 10625
rect 15381 10659 15439 10665
rect 15381 10625 15393 10659
rect 15427 10625 15439 10659
rect 15381 10619 15439 10625
rect 16853 10659 16911 10665
rect 16853 10625 16865 10659
rect 16899 10625 16911 10659
rect 16853 10619 16911 10625
rect 17037 10659 17095 10665
rect 17037 10625 17049 10659
rect 17083 10656 17095 10659
rect 17218 10656 17224 10668
rect 17083 10628 17224 10656
rect 17083 10625 17095 10628
rect 17037 10619 17095 10625
rect 1591 10591 1649 10597
rect 1591 10557 1603 10591
rect 1637 10557 1649 10591
rect 2866 10588 2872 10600
rect 2827 10560 2872 10588
rect 1591 10551 1649 10557
rect 2866 10548 2872 10560
rect 2924 10548 2930 10600
rect 3136 10591 3194 10597
rect 3136 10557 3148 10591
rect 3182 10588 3194 10591
rect 3694 10588 3700 10600
rect 3182 10560 3700 10588
rect 3182 10557 3194 10560
rect 3136 10551 3194 10557
rect 3694 10548 3700 10560
rect 3752 10548 3758 10600
rect 5534 10588 5540 10600
rect 5495 10560 5540 10588
rect 5534 10548 5540 10560
rect 5592 10548 5598 10600
rect 6454 10548 6460 10600
rect 6512 10588 6518 10600
rect 6825 10591 6883 10597
rect 6825 10588 6837 10591
rect 6512 10560 6837 10588
rect 6512 10548 6518 10560
rect 6825 10557 6837 10560
rect 6871 10557 6883 10591
rect 6825 10551 6883 10557
rect 9217 10591 9275 10597
rect 9217 10557 9229 10591
rect 9263 10588 9275 10591
rect 10226 10588 10232 10600
rect 9263 10560 10232 10588
rect 9263 10557 9275 10560
rect 9217 10551 9275 10557
rect 10226 10548 10232 10560
rect 10284 10548 10290 10600
rect 10321 10591 10379 10597
rect 10321 10557 10333 10591
rect 10367 10588 10379 10591
rect 11146 10588 11152 10600
rect 10367 10560 11152 10588
rect 10367 10557 10379 10560
rect 10321 10551 10379 10557
rect 11146 10548 11152 10560
rect 11204 10548 11210 10600
rect 11241 10591 11299 10597
rect 11241 10557 11253 10591
rect 11287 10588 11299 10591
rect 14734 10588 14740 10600
rect 11287 10560 14740 10588
rect 11287 10557 11299 10560
rect 11241 10551 11299 10557
rect 14734 10548 14740 10560
rect 14792 10548 14798 10600
rect 15396 10588 15424 10619
rect 17218 10616 17224 10628
rect 17276 10616 17282 10668
rect 17328 10656 17356 10764
rect 18509 10761 18521 10795
rect 18555 10792 18567 10795
rect 18874 10792 18880 10804
rect 18555 10764 18880 10792
rect 18555 10761 18567 10764
rect 18509 10755 18567 10761
rect 18874 10752 18880 10764
rect 18932 10752 18938 10804
rect 18230 10684 18236 10736
rect 18288 10724 18294 10736
rect 18782 10724 18788 10736
rect 18288 10696 18788 10724
rect 18288 10684 18294 10696
rect 18782 10684 18788 10696
rect 18840 10684 18846 10736
rect 19334 10656 19340 10668
rect 17328 10628 19340 10656
rect 19334 10616 19340 10628
rect 19392 10616 19398 10668
rect 15470 10588 15476 10600
rect 15396 10560 15476 10588
rect 15470 10548 15476 10560
rect 15528 10548 15534 10600
rect 16761 10591 16819 10597
rect 16761 10557 16773 10591
rect 16807 10588 16819 10591
rect 17770 10588 17776 10600
rect 16807 10560 17776 10588
rect 16807 10557 16819 10560
rect 16761 10551 16819 10557
rect 17770 10548 17776 10560
rect 17828 10548 17834 10600
rect 18325 10591 18383 10597
rect 18325 10557 18337 10591
rect 18371 10588 18383 10591
rect 19150 10588 19156 10600
rect 18371 10560 19156 10588
rect 18371 10557 18383 10560
rect 18325 10551 18383 10557
rect 19150 10548 19156 10560
rect 19208 10548 19214 10600
rect 19429 10591 19487 10597
rect 19429 10557 19441 10591
rect 19475 10557 19487 10591
rect 19429 10551 19487 10557
rect 1857 10523 1915 10529
rect 1857 10489 1869 10523
rect 1903 10520 1915 10523
rect 2222 10520 2228 10532
rect 1903 10492 2228 10520
rect 1903 10489 1915 10492
rect 1857 10483 1915 10489
rect 2222 10480 2228 10492
rect 2280 10480 2286 10532
rect 4062 10480 4068 10532
rect 4120 10520 4126 10532
rect 7092 10523 7150 10529
rect 4120 10492 5764 10520
rect 4120 10480 4126 10492
rect 5626 10452 5632 10464
rect 5587 10424 5632 10452
rect 5626 10412 5632 10424
rect 5684 10412 5690 10464
rect 5736 10452 5764 10492
rect 7092 10489 7104 10523
rect 7138 10520 7150 10523
rect 7374 10520 7380 10532
rect 7138 10492 7380 10520
rect 7138 10489 7150 10492
rect 7092 10483 7150 10489
rect 7374 10480 7380 10492
rect 7432 10480 7438 10532
rect 9953 10523 10011 10529
rect 9953 10520 9965 10523
rect 7484 10492 9965 10520
rect 7484 10452 7512 10492
rect 9953 10489 9965 10492
rect 9999 10489 10011 10523
rect 9953 10483 10011 10489
rect 10870 10480 10876 10532
rect 10928 10520 10934 10532
rect 15197 10523 15255 10529
rect 15197 10520 15209 10523
rect 10928 10492 15209 10520
rect 10928 10480 10934 10492
rect 15197 10489 15209 10492
rect 15243 10489 15255 10523
rect 15197 10483 15255 10489
rect 16850 10480 16856 10532
rect 16908 10520 16914 10532
rect 16908 10492 18000 10520
rect 16908 10480 16914 10492
rect 5736 10424 7512 10452
rect 8846 10412 8852 10464
rect 8904 10452 8910 10464
rect 9030 10452 9036 10464
rect 8904 10424 9036 10452
rect 8904 10412 8910 10424
rect 9030 10412 9036 10424
rect 9088 10412 9094 10464
rect 9493 10455 9551 10461
rect 9493 10421 9505 10455
rect 9539 10452 9551 10455
rect 9674 10452 9680 10464
rect 9539 10424 9680 10452
rect 9539 10421 9551 10424
rect 9493 10415 9551 10421
rect 9674 10412 9680 10424
rect 9732 10412 9738 10464
rect 9858 10452 9864 10464
rect 9819 10424 9864 10452
rect 9858 10412 9864 10424
rect 9916 10412 9922 10464
rect 10410 10412 10416 10464
rect 10468 10452 10474 10464
rect 10505 10455 10563 10461
rect 10505 10452 10517 10455
rect 10468 10424 10517 10452
rect 10468 10412 10474 10424
rect 10505 10421 10517 10424
rect 10551 10421 10563 10455
rect 11422 10452 11428 10464
rect 11383 10424 11428 10452
rect 10505 10415 10563 10421
rect 11422 10412 11428 10424
rect 11480 10412 11486 10464
rect 13630 10452 13636 10464
rect 13591 10424 13636 10452
rect 13630 10412 13636 10424
rect 13688 10412 13694 10464
rect 16393 10455 16451 10461
rect 16393 10421 16405 10455
rect 16439 10452 16451 10455
rect 17218 10452 17224 10464
rect 16439 10424 17224 10452
rect 16439 10421 16451 10424
rect 16393 10415 16451 10421
rect 17218 10412 17224 10424
rect 17276 10412 17282 10464
rect 17972 10452 18000 10492
rect 19334 10480 19340 10532
rect 19392 10520 19398 10532
rect 19444 10520 19472 10551
rect 19674 10523 19732 10529
rect 19674 10520 19686 10523
rect 19392 10492 19472 10520
rect 19536 10492 19686 10520
rect 19392 10480 19398 10492
rect 18046 10452 18052 10464
rect 17959 10424 18052 10452
rect 18046 10412 18052 10424
rect 18104 10452 18110 10464
rect 19536 10452 19564 10492
rect 19674 10489 19686 10492
rect 19720 10489 19732 10523
rect 19674 10483 19732 10489
rect 20806 10452 20812 10464
rect 18104 10424 19564 10452
rect 20767 10424 20812 10452
rect 18104 10412 18110 10424
rect 20806 10412 20812 10424
rect 20864 10412 20870 10464
rect 1104 10362 21896 10384
rect 1104 10310 7912 10362
rect 7964 10310 7976 10362
rect 8028 10310 8040 10362
rect 8092 10310 8104 10362
rect 8156 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 15035 10362
rect 15087 10310 21896 10362
rect 1104 10288 21896 10310
rect 2501 10251 2559 10257
rect 2501 10217 2513 10251
rect 2547 10248 2559 10251
rect 3050 10248 3056 10260
rect 2547 10220 3056 10248
rect 2547 10217 2559 10220
rect 2501 10211 2559 10217
rect 3050 10208 3056 10220
rect 3108 10208 3114 10260
rect 5810 10208 5816 10260
rect 5868 10248 5874 10260
rect 6733 10251 6791 10257
rect 6733 10248 6745 10251
rect 5868 10220 6745 10248
rect 5868 10208 5874 10220
rect 6733 10217 6745 10220
rect 6779 10217 6791 10251
rect 8478 10248 8484 10260
rect 8439 10220 8484 10248
rect 6733 10211 6791 10217
rect 8478 10208 8484 10220
rect 8536 10208 8542 10260
rect 12069 10251 12127 10257
rect 12069 10217 12081 10251
rect 12115 10248 12127 10251
rect 13630 10248 13636 10260
rect 12115 10220 13636 10248
rect 12115 10217 12127 10220
rect 12069 10211 12127 10217
rect 13630 10208 13636 10220
rect 13688 10208 13694 10260
rect 15838 10248 15844 10260
rect 13740 10220 15240 10248
rect 15799 10220 15844 10248
rect 7098 10180 7104 10192
rect 7059 10152 7104 10180
rect 7098 10140 7104 10152
rect 7156 10140 7162 10192
rect 7282 10140 7288 10192
rect 7340 10180 7346 10192
rect 7340 10152 13492 10180
rect 7340 10140 7346 10152
rect 1946 10072 1952 10124
rect 2004 10112 2010 10124
rect 2409 10115 2467 10121
rect 2409 10112 2421 10115
rect 2004 10084 2421 10112
rect 2004 10072 2010 10084
rect 2409 10081 2421 10084
rect 2455 10081 2467 10115
rect 2409 10075 2467 10081
rect 2866 10072 2872 10124
rect 2924 10112 2930 10124
rect 3878 10112 3884 10124
rect 2924 10084 3884 10112
rect 2924 10072 2930 10084
rect 3878 10072 3884 10084
rect 3936 10112 3942 10124
rect 4525 10115 4583 10121
rect 4525 10112 4537 10115
rect 3936 10084 4537 10112
rect 3936 10072 3942 10084
rect 4525 10081 4537 10084
rect 4571 10081 4583 10115
rect 4525 10075 4583 10081
rect 4792 10115 4850 10121
rect 4792 10081 4804 10115
rect 4838 10112 4850 10115
rect 5718 10112 5724 10124
rect 4838 10084 5724 10112
rect 4838 10081 4850 10084
rect 4792 10075 4850 10081
rect 5718 10072 5724 10084
rect 5776 10072 5782 10124
rect 7006 10072 7012 10124
rect 7064 10112 7070 10124
rect 8297 10115 8355 10121
rect 8297 10112 8309 10115
rect 7064 10084 8309 10112
rect 7064 10072 7070 10084
rect 8297 10081 8309 10084
rect 8343 10081 8355 10115
rect 8297 10075 8355 10081
rect 9677 10115 9735 10121
rect 9677 10081 9689 10115
rect 9723 10112 9735 10115
rect 9766 10112 9772 10124
rect 9723 10084 9772 10112
rect 9723 10081 9735 10084
rect 9677 10075 9735 10081
rect 9766 10072 9772 10084
rect 9824 10072 9830 10124
rect 9950 10121 9956 10124
rect 9944 10112 9956 10121
rect 9911 10084 9956 10112
rect 9944 10075 9956 10084
rect 9950 10072 9956 10075
rect 10008 10072 10014 10124
rect 12437 10115 12495 10121
rect 12437 10081 12449 10115
rect 12483 10112 12495 10115
rect 13078 10112 13084 10124
rect 12483 10084 13084 10112
rect 12483 10081 12495 10084
rect 12437 10075 12495 10081
rect 13078 10072 13084 10084
rect 13136 10072 13142 10124
rect 13464 10112 13492 10152
rect 13740 10112 13768 10220
rect 13998 10180 14004 10192
rect 13959 10152 14004 10180
rect 13998 10140 14004 10152
rect 14056 10140 14062 10192
rect 13464 10084 13768 10112
rect 14093 10115 14151 10121
rect 14093 10081 14105 10115
rect 14139 10112 14151 10115
rect 15102 10112 15108 10124
rect 14139 10084 15108 10112
rect 14139 10081 14151 10084
rect 14093 10075 14151 10081
rect 15102 10072 15108 10084
rect 15160 10072 15166 10124
rect 2685 10047 2743 10053
rect 2685 10013 2697 10047
rect 2731 10044 2743 10047
rect 4338 10044 4344 10056
rect 2731 10016 4344 10044
rect 2731 10013 2743 10016
rect 2685 10007 2743 10013
rect 4338 10004 4344 10016
rect 4396 10004 4402 10056
rect 6086 10004 6092 10056
rect 6144 10044 6150 10056
rect 6638 10044 6644 10056
rect 6144 10016 6644 10044
rect 6144 10004 6150 10016
rect 6638 10004 6644 10016
rect 6696 10044 6702 10056
rect 7193 10047 7251 10053
rect 7193 10044 7205 10047
rect 6696 10016 7205 10044
rect 6696 10004 6702 10016
rect 7193 10013 7205 10016
rect 7239 10013 7251 10047
rect 7193 10007 7251 10013
rect 7285 10047 7343 10053
rect 7285 10013 7297 10047
rect 7331 10044 7343 10047
rect 12526 10044 12532 10056
rect 7331 10016 7512 10044
rect 12487 10016 12532 10044
rect 7331 10013 7343 10016
rect 7285 10007 7343 10013
rect 5905 9979 5963 9985
rect 5905 9945 5917 9979
rect 5951 9976 5963 9979
rect 5994 9976 6000 9988
rect 5951 9948 6000 9976
rect 5951 9945 5963 9948
rect 5905 9939 5963 9945
rect 5994 9936 6000 9948
rect 6052 9976 6058 9988
rect 7374 9976 7380 9988
rect 6052 9948 7380 9976
rect 6052 9936 6058 9948
rect 7374 9936 7380 9948
rect 7432 9936 7438 9988
rect 2038 9908 2044 9920
rect 1999 9880 2044 9908
rect 2038 9868 2044 9880
rect 2096 9868 2102 9920
rect 5718 9868 5724 9920
rect 5776 9908 5782 9920
rect 6546 9908 6552 9920
rect 5776 9880 6552 9908
rect 5776 9868 5782 9880
rect 6546 9868 6552 9880
rect 6604 9908 6610 9920
rect 7484 9908 7512 10016
rect 12526 10004 12532 10016
rect 12584 10004 12590 10056
rect 12713 10047 12771 10053
rect 12713 10013 12725 10047
rect 12759 10044 12771 10047
rect 14182 10044 14188 10056
rect 12759 10016 13952 10044
rect 14143 10016 14188 10044
rect 12759 10013 12771 10016
rect 12713 10007 12771 10013
rect 13633 9979 13691 9985
rect 13633 9945 13645 9979
rect 13679 9976 13691 9979
rect 13814 9976 13820 9988
rect 13679 9948 13820 9976
rect 13679 9945 13691 9948
rect 13633 9939 13691 9945
rect 13814 9936 13820 9948
rect 13872 9936 13878 9988
rect 13924 9976 13952 10016
rect 14182 10004 14188 10016
rect 14240 10004 14246 10056
rect 15212 10044 15240 10220
rect 15838 10208 15844 10220
rect 15896 10208 15902 10260
rect 16758 10208 16764 10260
rect 16816 10248 16822 10260
rect 17586 10248 17592 10260
rect 16816 10220 17592 10248
rect 16816 10208 16822 10220
rect 17586 10208 17592 10220
rect 17644 10208 17650 10260
rect 18138 10208 18144 10260
rect 18196 10248 18202 10260
rect 18325 10251 18383 10257
rect 18325 10248 18337 10251
rect 18196 10220 18337 10248
rect 18196 10208 18202 10220
rect 18325 10217 18337 10220
rect 18371 10217 18383 10251
rect 18325 10211 18383 10217
rect 19242 10208 19248 10260
rect 19300 10248 19306 10260
rect 19705 10251 19763 10257
rect 19705 10248 19717 10251
rect 19300 10220 19717 10248
rect 19300 10208 19306 10220
rect 19705 10217 19717 10220
rect 19751 10217 19763 10251
rect 19705 10211 19763 10217
rect 15286 10140 15292 10192
rect 15344 10180 15350 10192
rect 15470 10180 15476 10192
rect 15344 10152 15476 10180
rect 15344 10140 15350 10152
rect 15470 10140 15476 10152
rect 15528 10180 15534 10192
rect 19150 10180 19156 10192
rect 15528 10152 19156 10180
rect 15528 10140 15534 10152
rect 15562 10072 15568 10124
rect 15620 10112 15626 10124
rect 15749 10115 15807 10121
rect 15749 10112 15761 10115
rect 15620 10084 15761 10112
rect 15620 10072 15626 10084
rect 15749 10081 15761 10084
rect 15795 10081 15807 10115
rect 16758 10112 16764 10124
rect 15749 10075 15807 10081
rect 15856 10084 16764 10112
rect 15856 10044 15884 10084
rect 16758 10072 16764 10084
rect 16816 10072 16822 10124
rect 16960 10121 16988 10152
rect 19150 10140 19156 10152
rect 19208 10140 19214 10192
rect 16945 10115 17003 10121
rect 16945 10081 16957 10115
rect 16991 10081 17003 10115
rect 16945 10075 17003 10081
rect 17212 10115 17270 10121
rect 17212 10081 17224 10115
rect 17258 10112 17270 10115
rect 17770 10112 17776 10124
rect 17258 10084 17776 10112
rect 17258 10081 17270 10084
rect 17212 10075 17270 10081
rect 17770 10072 17776 10084
rect 17828 10072 17834 10124
rect 19610 10112 19616 10124
rect 19571 10084 19616 10112
rect 19610 10072 19616 10084
rect 19668 10072 19674 10124
rect 16022 10044 16028 10056
rect 15212 10016 15884 10044
rect 15983 10016 16028 10044
rect 16022 10004 16028 10016
rect 16080 10004 16086 10056
rect 19889 10047 19947 10053
rect 19889 10013 19901 10047
rect 19935 10044 19947 10047
rect 20622 10044 20628 10056
rect 19935 10016 20628 10044
rect 19935 10013 19947 10016
rect 19889 10007 19947 10013
rect 20622 10004 20628 10016
rect 20680 10004 20686 10056
rect 14274 9976 14280 9988
rect 13924 9948 14280 9976
rect 14274 9936 14280 9948
rect 14332 9936 14338 9988
rect 14550 9936 14556 9988
rect 14608 9976 14614 9988
rect 14608 9948 16896 9976
rect 14608 9936 14614 9948
rect 11054 9908 11060 9920
rect 6604 9880 7512 9908
rect 11015 9880 11060 9908
rect 6604 9868 6610 9880
rect 11054 9868 11060 9880
rect 11112 9868 11118 9920
rect 15381 9911 15439 9917
rect 15381 9877 15393 9911
rect 15427 9908 15439 9911
rect 16758 9908 16764 9920
rect 15427 9880 16764 9908
rect 15427 9877 15439 9880
rect 15381 9871 15439 9877
rect 16758 9868 16764 9880
rect 16816 9868 16822 9920
rect 16868 9908 16896 9948
rect 17954 9936 17960 9988
rect 18012 9976 18018 9988
rect 20438 9976 20444 9988
rect 18012 9948 20444 9976
rect 18012 9936 18018 9948
rect 20438 9936 20444 9948
rect 20496 9936 20502 9988
rect 17862 9908 17868 9920
rect 16868 9880 17868 9908
rect 17862 9868 17868 9880
rect 17920 9868 17926 9920
rect 19245 9911 19303 9917
rect 19245 9877 19257 9911
rect 19291 9908 19303 9911
rect 20530 9908 20536 9920
rect 19291 9880 20536 9908
rect 19291 9877 19303 9880
rect 19245 9871 19303 9877
rect 20530 9868 20536 9880
rect 20588 9868 20594 9920
rect 1104 9818 21896 9840
rect 1104 9766 4447 9818
rect 4499 9766 4511 9818
rect 4563 9766 4575 9818
rect 4627 9766 4639 9818
rect 4691 9766 11378 9818
rect 11430 9766 11442 9818
rect 11494 9766 11506 9818
rect 11558 9766 11570 9818
rect 11622 9766 18308 9818
rect 18360 9766 18372 9818
rect 18424 9766 18436 9818
rect 18488 9766 18500 9818
rect 18552 9766 21896 9818
rect 1104 9744 21896 9766
rect 3234 9664 3240 9716
rect 3292 9704 3298 9716
rect 4062 9704 4068 9716
rect 3292 9676 4068 9704
rect 3292 9664 3298 9676
rect 4062 9664 4068 9676
rect 4120 9664 4126 9716
rect 5000 9676 5304 9704
rect 5000 9636 5028 9676
rect 5166 9636 5172 9648
rect 3712 9608 5028 9636
rect 5127 9608 5172 9636
rect 3712 9580 3740 9608
rect 5166 9596 5172 9608
rect 5224 9596 5230 9648
rect 5276 9636 5304 9676
rect 5626 9664 5632 9716
rect 5684 9704 5690 9716
rect 6825 9707 6883 9713
rect 6825 9704 6837 9707
rect 5684 9676 6837 9704
rect 5684 9664 5690 9676
rect 6825 9673 6837 9676
rect 6871 9673 6883 9707
rect 6825 9667 6883 9673
rect 12434 9664 12440 9716
rect 12492 9704 12498 9716
rect 12492 9676 13400 9704
rect 12492 9664 12498 9676
rect 9582 9636 9588 9648
rect 5276 9608 9588 9636
rect 9582 9596 9588 9608
rect 9640 9596 9646 9648
rect 9769 9639 9827 9645
rect 9769 9605 9781 9639
rect 9815 9636 9827 9639
rect 11238 9636 11244 9648
rect 9815 9608 11244 9636
rect 9815 9605 9827 9608
rect 9769 9599 9827 9605
rect 11238 9596 11244 9608
rect 11296 9596 11302 9648
rect 13372 9636 13400 9676
rect 13538 9664 13544 9716
rect 13596 9704 13602 9716
rect 19610 9704 19616 9716
rect 13596 9676 19616 9704
rect 13596 9664 13602 9676
rect 19610 9664 19616 9676
rect 19668 9664 19674 9716
rect 20162 9664 20168 9716
rect 20220 9704 20226 9716
rect 20438 9704 20444 9716
rect 20220 9676 20444 9704
rect 20220 9664 20226 9676
rect 20438 9664 20444 9676
rect 20496 9664 20502 9716
rect 13814 9636 13820 9648
rect 13372 9608 13492 9636
rect 13727 9608 13820 9636
rect 2501 9571 2559 9577
rect 2501 9537 2513 9571
rect 2547 9568 2559 9571
rect 2866 9568 2872 9580
rect 2547 9540 2872 9568
rect 2547 9537 2559 9540
rect 2501 9531 2559 9537
rect 2866 9528 2872 9540
rect 2924 9528 2930 9580
rect 3694 9528 3700 9580
rect 3752 9528 3758 9580
rect 4157 9571 4215 9577
rect 4157 9537 4169 9571
rect 4203 9568 4215 9571
rect 5442 9568 5448 9580
rect 4203 9540 5448 9568
rect 4203 9537 4215 9540
rect 4157 9531 4215 9537
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 5718 9568 5724 9580
rect 5679 9540 5724 9568
rect 5718 9528 5724 9540
rect 5776 9528 5782 9580
rect 7374 9568 7380 9580
rect 7335 9540 7380 9568
rect 7374 9528 7380 9540
rect 7432 9528 7438 9580
rect 10226 9568 10232 9580
rect 10187 9540 10232 9568
rect 10226 9528 10232 9540
rect 10284 9528 10290 9580
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9568 10471 9571
rect 11054 9568 11060 9580
rect 10459 9540 11060 9568
rect 10459 9537 10471 9540
rect 10413 9531 10471 9537
rect 11054 9528 11060 9540
rect 11112 9528 11118 9580
rect 13464 9568 13492 9608
rect 13814 9596 13820 9608
rect 13872 9636 13878 9648
rect 14274 9636 14280 9648
rect 13872 9608 14280 9636
rect 13872 9596 13878 9608
rect 14274 9596 14280 9608
rect 14332 9596 14338 9648
rect 16022 9636 16028 9648
rect 15488 9608 16028 9636
rect 14366 9568 14372 9580
rect 13464 9540 14372 9568
rect 14366 9528 14372 9540
rect 14424 9568 14430 9580
rect 14550 9568 14556 9580
rect 14424 9540 14556 9568
rect 14424 9528 14430 9540
rect 14550 9528 14556 9540
rect 14608 9528 14614 9580
rect 15286 9568 15292 9580
rect 15247 9540 15292 9568
rect 15286 9528 15292 9540
rect 15344 9528 15350 9580
rect 15488 9577 15516 9608
rect 16022 9596 16028 9608
rect 16080 9636 16086 9648
rect 16080 9608 17080 9636
rect 16080 9596 16086 9608
rect 15473 9571 15531 9577
rect 15473 9537 15485 9571
rect 15519 9537 15531 9571
rect 15473 9531 15531 9537
rect 16945 9571 17003 9577
rect 16945 9537 16957 9571
rect 16991 9537 17003 9571
rect 17052 9568 17080 9608
rect 17052 9540 19380 9568
rect 16945 9531 17003 9537
rect 2038 9460 2044 9512
rect 2096 9500 2102 9512
rect 2225 9503 2283 9509
rect 2225 9500 2237 9503
rect 2096 9472 2237 9500
rect 2096 9460 2102 9472
rect 2225 9469 2237 9472
rect 2271 9469 2283 9503
rect 4065 9503 4123 9509
rect 4065 9500 4077 9503
rect 2225 9463 2283 9469
rect 3712 9472 4077 9500
rect 3712 9444 3740 9472
rect 4065 9469 4077 9472
rect 4111 9469 4123 9503
rect 4065 9463 4123 9469
rect 4246 9460 4252 9512
rect 4304 9500 4310 9512
rect 5537 9503 5595 9509
rect 5537 9500 5549 9503
rect 4304 9472 5549 9500
rect 4304 9460 4310 9472
rect 5537 9469 5549 9472
rect 5583 9469 5595 9503
rect 8665 9503 8723 9509
rect 5537 9463 5595 9469
rect 5644 9472 7420 9500
rect 3694 9392 3700 9444
rect 3752 9392 3758 9444
rect 3786 9392 3792 9444
rect 3844 9432 3850 9444
rect 5644 9432 5672 9472
rect 3844 9404 5672 9432
rect 3844 9392 3850 9404
rect 6730 9392 6736 9444
rect 6788 9432 6794 9444
rect 7285 9435 7343 9441
rect 7285 9432 7297 9435
rect 6788 9404 7297 9432
rect 6788 9392 6794 9404
rect 7285 9401 7297 9404
rect 7331 9401 7343 9435
rect 7392 9432 7420 9472
rect 8665 9469 8677 9503
rect 8711 9500 8723 9503
rect 10318 9500 10324 9512
rect 8711 9472 10324 9500
rect 8711 9469 8723 9472
rect 8665 9463 8723 9469
rect 10318 9460 10324 9472
rect 10376 9460 10382 9512
rect 12342 9460 12348 9512
rect 12400 9500 12406 9512
rect 12437 9503 12495 9509
rect 12437 9500 12449 9503
rect 12400 9472 12449 9500
rect 12400 9460 12406 9472
rect 12437 9469 12449 9472
rect 12483 9469 12495 9503
rect 12437 9463 12495 9469
rect 12704 9503 12762 9509
rect 12704 9469 12716 9503
rect 12750 9500 12762 9503
rect 14182 9500 14188 9512
rect 12750 9472 14188 9500
rect 12750 9469 12762 9472
rect 12704 9463 12762 9469
rect 14182 9460 14188 9472
rect 14240 9460 14246 9512
rect 16758 9500 16764 9512
rect 16719 9472 16764 9500
rect 16758 9460 16764 9472
rect 16816 9460 16822 9512
rect 7392 9404 9536 9432
rect 7285 9395 7343 9401
rect 1854 9364 1860 9376
rect 1815 9336 1860 9364
rect 1854 9324 1860 9336
rect 1912 9324 1918 9376
rect 2314 9364 2320 9376
rect 2275 9336 2320 9364
rect 2314 9324 2320 9336
rect 2372 9324 2378 9376
rect 3602 9364 3608 9376
rect 3563 9336 3608 9364
rect 3602 9324 3608 9336
rect 3660 9324 3666 9376
rect 3973 9367 4031 9373
rect 3973 9333 3985 9367
rect 4019 9364 4031 9367
rect 4062 9364 4068 9376
rect 4019 9336 4068 9364
rect 4019 9333 4031 9336
rect 3973 9327 4031 9333
rect 4062 9324 4068 9336
rect 4120 9324 4126 9376
rect 4154 9324 4160 9376
rect 4212 9364 4218 9376
rect 5166 9364 5172 9376
rect 4212 9336 5172 9364
rect 4212 9324 4218 9336
rect 5166 9324 5172 9336
rect 5224 9364 5230 9376
rect 5629 9367 5687 9373
rect 5629 9364 5641 9367
rect 5224 9336 5641 9364
rect 5224 9324 5230 9336
rect 5629 9333 5641 9336
rect 5675 9333 5687 9367
rect 5629 9327 5687 9333
rect 6546 9324 6552 9376
rect 6604 9364 6610 9376
rect 6914 9364 6920 9376
rect 6604 9336 6920 9364
rect 6604 9324 6610 9336
rect 6914 9324 6920 9336
rect 6972 9324 6978 9376
rect 7190 9364 7196 9376
rect 7151 9336 7196 9364
rect 7190 9324 7196 9336
rect 7248 9324 7254 9376
rect 8849 9367 8907 9373
rect 8849 9333 8861 9367
rect 8895 9364 8907 9367
rect 9398 9364 9404 9376
rect 8895 9336 9404 9364
rect 8895 9333 8907 9336
rect 8849 9327 8907 9333
rect 9398 9324 9404 9336
rect 9456 9324 9462 9376
rect 9508 9364 9536 9404
rect 9674 9392 9680 9444
rect 9732 9432 9738 9444
rect 10137 9435 10195 9441
rect 10137 9432 10149 9435
rect 9732 9404 10149 9432
rect 9732 9392 9738 9404
rect 10137 9401 10149 9404
rect 10183 9401 10195 9435
rect 12158 9432 12164 9444
rect 10137 9395 10195 9401
rect 10244 9404 12164 9432
rect 10244 9364 10272 9404
rect 12158 9392 12164 9404
rect 12216 9392 12222 9444
rect 12802 9392 12808 9444
rect 12860 9432 12866 9444
rect 13998 9432 14004 9444
rect 12860 9404 14004 9432
rect 12860 9392 12866 9404
rect 13998 9392 14004 9404
rect 14056 9392 14062 9444
rect 16853 9435 16911 9441
rect 16853 9432 16865 9435
rect 14844 9404 16865 9432
rect 9508 9336 10272 9364
rect 11333 9367 11391 9373
rect 11333 9333 11345 9367
rect 11379 9364 11391 9367
rect 12986 9364 12992 9376
rect 11379 9336 12992 9364
rect 11379 9333 11391 9336
rect 11333 9327 11391 9333
rect 12986 9324 12992 9336
rect 13044 9324 13050 9376
rect 14844 9373 14872 9404
rect 16853 9401 16865 9404
rect 16899 9401 16911 9435
rect 16960 9432 16988 9531
rect 17954 9460 17960 9512
rect 18012 9500 18018 9512
rect 18049 9503 18107 9509
rect 18049 9500 18061 9503
rect 18012 9472 18061 9500
rect 18012 9460 18018 9472
rect 18049 9469 18061 9472
rect 18095 9469 18107 9503
rect 18049 9463 18107 9469
rect 19150 9460 19156 9512
rect 19208 9500 19214 9512
rect 19245 9503 19303 9509
rect 19245 9500 19257 9503
rect 19208 9472 19257 9500
rect 19208 9460 19214 9472
rect 19245 9469 19257 9472
rect 19291 9469 19303 9503
rect 19352 9500 19380 9540
rect 19512 9503 19570 9509
rect 19512 9500 19524 9503
rect 19352 9472 19524 9500
rect 19245 9463 19303 9469
rect 19512 9469 19524 9472
rect 19558 9500 19570 9503
rect 20806 9500 20812 9512
rect 19558 9472 20812 9500
rect 19558 9469 19570 9472
rect 19512 9463 19570 9469
rect 20806 9460 20812 9472
rect 20864 9460 20870 9512
rect 19702 9432 19708 9444
rect 16960 9404 19708 9432
rect 16853 9395 16911 9401
rect 19702 9392 19708 9404
rect 19760 9432 19766 9444
rect 19760 9404 20668 9432
rect 19760 9392 19766 9404
rect 14829 9367 14887 9373
rect 14829 9333 14841 9367
rect 14875 9333 14887 9367
rect 15194 9364 15200 9376
rect 15155 9336 15200 9364
rect 14829 9327 14887 9333
rect 15194 9324 15200 9336
rect 15252 9324 15258 9376
rect 16393 9367 16451 9373
rect 16393 9333 16405 9367
rect 16439 9364 16451 9367
rect 16942 9364 16948 9376
rect 16439 9336 16948 9364
rect 16439 9333 16451 9336
rect 16393 9327 16451 9333
rect 16942 9324 16948 9336
rect 17000 9324 17006 9376
rect 17494 9324 17500 9376
rect 17552 9364 17558 9376
rect 20640 9373 20668 9404
rect 18233 9367 18291 9373
rect 18233 9364 18245 9367
rect 17552 9336 18245 9364
rect 17552 9324 17558 9336
rect 18233 9333 18245 9336
rect 18279 9333 18291 9367
rect 18233 9327 18291 9333
rect 20625 9367 20683 9373
rect 20625 9333 20637 9367
rect 20671 9333 20683 9367
rect 20625 9327 20683 9333
rect 1104 9274 21896 9296
rect 1104 9222 7912 9274
rect 7964 9222 7976 9274
rect 8028 9222 8040 9274
rect 8092 9222 8104 9274
rect 8156 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 15035 9274
rect 15087 9222 21896 9274
rect 1104 9200 21896 9222
rect 3145 9163 3203 9169
rect 3145 9129 3157 9163
rect 3191 9129 3203 9163
rect 3145 9123 3203 9129
rect 2774 9052 2780 9104
rect 2832 9092 2838 9104
rect 3160 9092 3188 9123
rect 4062 9120 4068 9172
rect 4120 9160 4126 9172
rect 12434 9160 12440 9172
rect 4120 9132 12440 9160
rect 4120 9120 4126 9132
rect 12434 9120 12440 9132
rect 12492 9120 12498 9172
rect 13906 9120 13912 9172
rect 13964 9160 13970 9172
rect 14369 9163 14427 9169
rect 14369 9160 14381 9163
rect 13964 9132 14381 9160
rect 13964 9120 13970 9132
rect 14369 9129 14381 9132
rect 14415 9160 14427 9163
rect 14458 9160 14464 9172
rect 14415 9132 14464 9160
rect 14415 9129 14427 9132
rect 14369 9123 14427 9129
rect 14458 9120 14464 9132
rect 14516 9120 14522 9172
rect 15473 9163 15531 9169
rect 15473 9129 15485 9163
rect 15519 9160 15531 9163
rect 16758 9160 16764 9172
rect 15519 9132 16764 9160
rect 15519 9129 15531 9132
rect 15473 9123 15531 9129
rect 16758 9120 16764 9132
rect 16816 9120 16822 9172
rect 17770 9160 17776 9172
rect 17731 9132 17776 9160
rect 17770 9120 17776 9132
rect 17828 9120 17834 9172
rect 18138 9120 18144 9172
rect 18196 9160 18202 9172
rect 19150 9160 19156 9172
rect 18196 9132 19156 9160
rect 18196 9120 18202 9132
rect 19150 9120 19156 9132
rect 19208 9120 19214 9172
rect 4310 9095 4368 9101
rect 4310 9092 4322 9095
rect 2832 9064 4322 9092
rect 2832 9052 2838 9064
rect 4310 9061 4322 9064
rect 4356 9061 4368 9095
rect 7193 9095 7251 9101
rect 7193 9092 7205 9095
rect 4310 9055 4368 9061
rect 5644 9064 7205 9092
rect 2032 9027 2090 9033
rect 2032 8993 2044 9027
rect 2078 9024 2090 9027
rect 2866 9024 2872 9036
rect 2078 8996 2872 9024
rect 2078 8993 2090 8996
rect 2032 8987 2090 8993
rect 2866 8984 2872 8996
rect 2924 9024 2930 9036
rect 3510 9024 3516 9036
rect 2924 8996 3516 9024
rect 2924 8984 2930 8996
rect 3510 8984 3516 8996
rect 3568 8984 3574 9036
rect 3602 8984 3608 9036
rect 3660 9024 3666 9036
rect 5644 9024 5672 9064
rect 7193 9061 7205 9064
rect 7239 9061 7251 9095
rect 7193 9055 7251 9061
rect 8202 9052 8208 9104
rect 8260 9092 8266 9104
rect 10772 9095 10830 9101
rect 8260 9064 9168 9092
rect 8260 9052 8266 9064
rect 3660 8996 5672 9024
rect 6641 9027 6699 9033
rect 3660 8984 3666 8996
rect 6641 8993 6653 9027
rect 6687 9024 6699 9027
rect 6687 8996 6868 9024
rect 6687 8993 6699 8996
rect 6641 8987 6699 8993
rect 1765 8959 1823 8965
rect 1765 8925 1777 8959
rect 1811 8925 1823 8959
rect 1765 8919 1823 8925
rect 1780 8820 1808 8919
rect 3878 8916 3884 8968
rect 3936 8956 3942 8968
rect 4065 8959 4123 8965
rect 4065 8956 4077 8959
rect 3936 8928 4077 8956
rect 3936 8916 3942 8928
rect 4065 8925 4077 8928
rect 4111 8925 4123 8959
rect 4065 8919 4123 8925
rect 4080 8820 4108 8919
rect 6730 8888 6736 8900
rect 6691 8860 6736 8888
rect 6730 8848 6736 8860
rect 6788 8848 6794 8900
rect 6840 8888 6868 8996
rect 7006 8984 7012 9036
rect 7064 9024 7070 9036
rect 7101 9027 7159 9033
rect 7101 9024 7113 9027
rect 7064 8996 7113 9024
rect 7064 8984 7070 8996
rect 7101 8993 7113 8996
rect 7147 8993 7159 9027
rect 7101 8987 7159 8993
rect 8481 9027 8539 9033
rect 8481 8993 8493 9027
rect 8527 9024 8539 9027
rect 9030 9024 9036 9036
rect 8527 8996 9036 9024
rect 8527 8993 8539 8996
rect 8481 8987 8539 8993
rect 9030 8984 9036 8996
rect 9088 8984 9094 9036
rect 9140 9024 9168 9064
rect 10772 9061 10784 9095
rect 10818 9092 10830 9095
rect 11054 9092 11060 9104
rect 10818 9064 11060 9092
rect 10818 9061 10830 9064
rect 10772 9055 10830 9061
rect 11054 9052 11060 9064
rect 11112 9052 11118 9104
rect 11146 9052 11152 9104
rect 11204 9092 11210 9104
rect 17788 9092 17816 9120
rect 11204 9064 15240 9092
rect 17788 9064 19104 9092
rect 11204 9052 11210 9064
rect 12802 9024 12808 9036
rect 9140 8996 12808 9024
rect 12802 8984 12808 8996
rect 12860 8984 12866 9036
rect 12894 8984 12900 9036
rect 12952 9024 12958 9036
rect 13256 9027 13314 9033
rect 12952 8996 12997 9024
rect 12952 8984 12958 8996
rect 13256 8993 13268 9027
rect 13302 9024 13314 9027
rect 13814 9024 13820 9036
rect 13302 8996 13820 9024
rect 13302 8993 13314 8996
rect 13256 8987 13314 8993
rect 13814 8984 13820 8996
rect 13872 8984 13878 9036
rect 6914 8916 6920 8968
rect 6972 8956 6978 8968
rect 7285 8959 7343 8965
rect 7285 8956 7297 8959
rect 6972 8928 7297 8956
rect 6972 8916 6978 8928
rect 7285 8925 7297 8928
rect 7331 8925 7343 8959
rect 7285 8919 7343 8925
rect 9122 8916 9128 8968
rect 9180 8956 9186 8968
rect 9766 8956 9772 8968
rect 9180 8928 9772 8956
rect 9180 8916 9186 8928
rect 9766 8916 9772 8928
rect 9824 8956 9830 8968
rect 10505 8959 10563 8965
rect 10505 8956 10517 8959
rect 9824 8928 10517 8956
rect 9824 8916 9830 8928
rect 10505 8925 10517 8928
rect 10551 8925 10563 8959
rect 10505 8919 10563 8925
rect 12342 8916 12348 8968
rect 12400 8956 12406 8968
rect 12989 8959 13047 8965
rect 12989 8956 13001 8959
rect 12400 8928 13001 8956
rect 12400 8916 12406 8928
rect 12989 8925 13001 8928
rect 13035 8925 13047 8959
rect 15212 8956 15240 9064
rect 15289 9027 15347 9033
rect 15289 8993 15301 9027
rect 15335 9024 15347 9027
rect 15378 9024 15384 9036
rect 15335 8996 15384 9024
rect 15335 8993 15347 8996
rect 15289 8987 15347 8993
rect 15378 8984 15384 8996
rect 15436 8984 15442 9036
rect 15470 8984 15476 9036
rect 15528 9024 15534 9036
rect 16393 9027 16451 9033
rect 16393 9024 16405 9027
rect 15528 8996 16405 9024
rect 15528 8984 15534 8996
rect 16040 8968 16068 8996
rect 16393 8993 16405 8996
rect 16439 8993 16451 9027
rect 16393 8987 16451 8993
rect 16660 9027 16718 9033
rect 16660 8993 16672 9027
rect 16706 9024 16718 9027
rect 17034 9024 17040 9036
rect 16706 8996 17040 9024
rect 16706 8993 16718 8996
rect 16660 8987 16718 8993
rect 17034 8984 17040 8996
rect 17092 8984 17098 9036
rect 18046 8984 18052 9036
rect 18104 9024 18110 9036
rect 18969 9027 19027 9033
rect 18969 9024 18981 9027
rect 18104 8996 18981 9024
rect 18104 8984 18110 8996
rect 18969 8993 18981 8996
rect 19015 8993 19027 9027
rect 19076 9024 19104 9064
rect 19076 8996 19196 9024
rect 18969 8987 19027 8993
rect 15212 8928 15424 8956
rect 12989 8919 13047 8925
rect 8846 8888 8852 8900
rect 6840 8860 8852 8888
rect 8846 8848 8852 8860
rect 8904 8848 8910 8900
rect 5074 8820 5080 8832
rect 1780 8792 5080 8820
rect 5074 8780 5080 8792
rect 5132 8780 5138 8832
rect 5442 8820 5448 8832
rect 5355 8792 5448 8820
rect 5442 8780 5448 8792
rect 5500 8820 5506 8832
rect 6086 8820 6092 8832
rect 5500 8792 6092 8820
rect 5500 8780 5506 8792
rect 6086 8780 6092 8792
rect 6144 8780 6150 8832
rect 6457 8823 6515 8829
rect 6457 8789 6469 8823
rect 6503 8820 6515 8823
rect 6914 8820 6920 8832
rect 6503 8792 6920 8820
rect 6503 8789 6515 8792
rect 6457 8783 6515 8789
rect 6914 8780 6920 8792
rect 6972 8780 6978 8832
rect 8662 8820 8668 8832
rect 8623 8792 8668 8820
rect 8662 8780 8668 8792
rect 8720 8780 8726 8832
rect 11790 8780 11796 8832
rect 11848 8820 11854 8832
rect 11885 8823 11943 8829
rect 11885 8820 11897 8823
rect 11848 8792 11897 8820
rect 11848 8780 11854 8792
rect 11885 8789 11897 8792
rect 11931 8789 11943 8823
rect 11885 8783 11943 8789
rect 12250 8780 12256 8832
rect 12308 8820 12314 8832
rect 12713 8823 12771 8829
rect 12713 8820 12725 8823
rect 12308 8792 12725 8820
rect 12308 8780 12314 8792
rect 12713 8789 12725 8792
rect 12759 8820 12771 8823
rect 15286 8820 15292 8832
rect 12759 8792 15292 8820
rect 12759 8789 12771 8792
rect 12713 8783 12771 8789
rect 15286 8780 15292 8792
rect 15344 8780 15350 8832
rect 15396 8820 15424 8928
rect 16022 8916 16028 8968
rect 16080 8916 16086 8968
rect 18782 8916 18788 8968
rect 18840 8956 18846 8968
rect 19168 8965 19196 8996
rect 19061 8959 19119 8965
rect 19061 8956 19073 8959
rect 18840 8928 19073 8956
rect 18840 8916 18846 8928
rect 19061 8925 19073 8928
rect 19107 8925 19119 8959
rect 19061 8919 19119 8925
rect 19153 8959 19211 8965
rect 19153 8925 19165 8959
rect 19199 8925 19211 8959
rect 19153 8919 19211 8925
rect 18230 8848 18236 8900
rect 18288 8888 18294 8900
rect 19886 8888 19892 8900
rect 18288 8860 19892 8888
rect 18288 8848 18294 8860
rect 19886 8848 19892 8860
rect 19944 8848 19950 8900
rect 18138 8820 18144 8832
rect 15396 8792 18144 8820
rect 18138 8780 18144 8792
rect 18196 8780 18202 8832
rect 18601 8823 18659 8829
rect 18601 8789 18613 8823
rect 18647 8820 18659 8823
rect 19058 8820 19064 8832
rect 18647 8792 19064 8820
rect 18647 8789 18659 8792
rect 18601 8783 18659 8789
rect 19058 8780 19064 8792
rect 19116 8780 19122 8832
rect 1104 8730 21896 8752
rect 1104 8678 4447 8730
rect 4499 8678 4511 8730
rect 4563 8678 4575 8730
rect 4627 8678 4639 8730
rect 4691 8678 11378 8730
rect 11430 8678 11442 8730
rect 11494 8678 11506 8730
rect 11558 8678 11570 8730
rect 11622 8678 18308 8730
rect 18360 8678 18372 8730
rect 18424 8678 18436 8730
rect 18488 8678 18500 8730
rect 18552 8678 21896 8730
rect 1104 8656 21896 8678
rect 2133 8619 2191 8625
rect 2133 8585 2145 8619
rect 2179 8616 2191 8619
rect 3418 8616 3424 8628
rect 2179 8588 3424 8616
rect 2179 8585 2191 8588
rect 2133 8579 2191 8585
rect 3418 8576 3424 8588
rect 3476 8576 3482 8628
rect 5074 8576 5080 8628
rect 5132 8616 5138 8628
rect 5997 8619 6055 8625
rect 5997 8616 6009 8619
rect 5132 8588 6009 8616
rect 5132 8576 5138 8588
rect 5997 8585 6009 8588
rect 6043 8585 6055 8619
rect 5997 8579 6055 8585
rect 6086 8576 6092 8628
rect 6144 8616 6150 8628
rect 6144 8588 7880 8616
rect 6144 8576 6150 8588
rect 4338 8508 4344 8560
rect 4396 8548 4402 8560
rect 7006 8548 7012 8560
rect 4396 8520 5120 8548
rect 6967 8520 7012 8548
rect 4396 8508 4402 8520
rect 5092 8492 5120 8520
rect 7006 8508 7012 8520
rect 7064 8508 7070 8560
rect 7742 8548 7748 8560
rect 7484 8520 7748 8548
rect 1302 8440 1308 8492
rect 1360 8480 1366 8492
rect 1360 8452 2728 8480
rect 1360 8440 1366 8452
rect 1854 8372 1860 8424
rect 1912 8412 1918 8424
rect 2501 8415 2559 8421
rect 2501 8412 2513 8415
rect 1912 8384 2513 8412
rect 1912 8372 1918 8384
rect 2501 8381 2513 8384
rect 2547 8381 2559 8415
rect 2700 8412 2728 8452
rect 2774 8440 2780 8492
rect 2832 8480 2838 8492
rect 4890 8480 4896 8492
rect 2832 8452 2877 8480
rect 4851 8452 4896 8480
rect 2832 8440 2838 8452
rect 4890 8440 4896 8452
rect 4948 8440 4954 8492
rect 5074 8480 5080 8492
rect 5035 8452 5080 8480
rect 5074 8440 5080 8452
rect 5132 8440 5138 8492
rect 7098 8440 7104 8492
rect 7156 8480 7162 8492
rect 7484 8489 7512 8520
rect 7742 8508 7748 8520
rect 7800 8508 7806 8560
rect 7469 8483 7527 8489
rect 7469 8480 7481 8483
rect 7156 8452 7481 8480
rect 7156 8440 7162 8452
rect 7469 8449 7481 8452
rect 7515 8449 7527 8483
rect 7469 8443 7527 8449
rect 7653 8483 7711 8489
rect 7653 8449 7665 8483
rect 7699 8480 7711 8483
rect 7852 8480 7880 8588
rect 9950 8576 9956 8628
rect 10008 8616 10014 8628
rect 10318 8616 10324 8628
rect 10008 8588 10324 8616
rect 10008 8576 10014 8588
rect 10318 8576 10324 8588
rect 10376 8616 10382 8628
rect 10597 8619 10655 8625
rect 10597 8616 10609 8619
rect 10376 8588 10609 8616
rect 10376 8576 10382 8588
rect 10597 8585 10609 8588
rect 10643 8585 10655 8619
rect 12434 8616 12440 8628
rect 12395 8588 12440 8616
rect 10597 8579 10655 8585
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 12802 8576 12808 8628
rect 12860 8616 12866 8628
rect 16393 8619 16451 8625
rect 12860 8588 15240 8616
rect 12860 8576 12866 8588
rect 11514 8508 11520 8560
rect 11572 8548 11578 8560
rect 12069 8551 12127 8557
rect 12069 8548 12081 8551
rect 11572 8520 12081 8548
rect 11572 8508 11578 8520
rect 12069 8517 12081 8520
rect 12115 8548 12127 8551
rect 12342 8548 12348 8560
rect 12115 8520 12348 8548
rect 12115 8517 12127 8520
rect 12069 8511 12127 8517
rect 12342 8508 12348 8520
rect 12400 8548 12406 8560
rect 12400 8520 14228 8548
rect 12400 8508 12406 8520
rect 14200 8492 14228 8520
rect 7699 8452 7880 8480
rect 7699 8449 7711 8452
rect 7653 8443 7711 8449
rect 8386 8440 8392 8492
rect 8444 8480 8450 8492
rect 8444 8452 9352 8480
rect 8444 8440 8450 8452
rect 4798 8412 4804 8424
rect 2700 8384 4804 8412
rect 2501 8375 2559 8381
rect 4798 8372 4804 8384
rect 4856 8372 4862 8424
rect 6181 8415 6239 8421
rect 6181 8381 6193 8415
rect 6227 8412 6239 8415
rect 6914 8412 6920 8424
rect 6227 8384 6920 8412
rect 6227 8381 6239 8384
rect 6181 8375 6239 8381
rect 6914 8372 6920 8384
rect 6972 8412 6978 8424
rect 7742 8412 7748 8424
rect 6972 8384 7748 8412
rect 6972 8372 6978 8384
rect 7742 8372 7748 8384
rect 7800 8372 7806 8424
rect 9122 8372 9128 8424
rect 9180 8412 9186 8424
rect 9217 8415 9275 8421
rect 9217 8412 9229 8415
rect 9180 8384 9229 8412
rect 9180 8372 9186 8384
rect 9217 8381 9229 8384
rect 9263 8381 9275 8415
rect 9324 8412 9352 8452
rect 12894 8440 12900 8492
rect 12952 8480 12958 8492
rect 12989 8483 13047 8489
rect 12989 8480 13001 8483
rect 12952 8452 13001 8480
rect 12952 8440 12958 8452
rect 12989 8449 13001 8452
rect 13035 8449 13047 8483
rect 14182 8480 14188 8492
rect 14095 8452 14188 8480
rect 12989 8443 13047 8449
rect 14182 8440 14188 8452
rect 14240 8440 14246 8492
rect 15212 8480 15240 8588
rect 16393 8585 16405 8619
rect 16439 8616 16451 8619
rect 18046 8616 18052 8628
rect 16439 8588 17724 8616
rect 18007 8588 18052 8616
rect 16439 8585 16451 8588
rect 16393 8579 16451 8585
rect 15565 8551 15623 8557
rect 15565 8517 15577 8551
rect 15611 8548 15623 8551
rect 15930 8548 15936 8560
rect 15611 8520 15936 8548
rect 15611 8517 15623 8520
rect 15565 8511 15623 8517
rect 15930 8508 15936 8520
rect 15988 8508 15994 8560
rect 17696 8548 17724 8588
rect 18046 8576 18052 8588
rect 18104 8576 18110 8628
rect 18782 8576 18788 8628
rect 18840 8576 18846 8628
rect 18800 8548 18828 8576
rect 17696 8520 18828 8548
rect 17034 8480 17040 8492
rect 15212 8452 16804 8480
rect 16947 8452 17040 8480
rect 12250 8412 12256 8424
rect 9324 8384 9904 8412
rect 12211 8384 12256 8412
rect 9217 8375 9275 8381
rect 2593 8347 2651 8353
rect 2593 8313 2605 8347
rect 2639 8344 2651 8347
rect 4154 8344 4160 8356
rect 2639 8316 4160 8344
rect 2639 8313 2651 8316
rect 2593 8307 2651 8313
rect 4154 8304 4160 8316
rect 4212 8304 4218 8356
rect 4264 8316 4568 8344
rect 4062 8236 4068 8288
rect 4120 8276 4126 8288
rect 4264 8276 4292 8316
rect 4120 8248 4292 8276
rect 4120 8236 4126 8248
rect 4338 8236 4344 8288
rect 4396 8276 4402 8288
rect 4433 8279 4491 8285
rect 4433 8276 4445 8279
rect 4396 8248 4445 8276
rect 4396 8236 4402 8248
rect 4433 8245 4445 8248
rect 4479 8245 4491 8279
rect 4540 8276 4568 8316
rect 7282 8304 7288 8356
rect 7340 8344 7346 8356
rect 7377 8347 7435 8353
rect 7377 8344 7389 8347
rect 7340 8316 7389 8344
rect 7340 8304 7346 8316
rect 7377 8313 7389 8316
rect 7423 8344 7435 8347
rect 7650 8344 7656 8356
rect 7423 8316 7656 8344
rect 7423 8313 7435 8316
rect 7377 8307 7435 8313
rect 7650 8304 7656 8316
rect 7708 8304 7714 8356
rect 9484 8347 9542 8353
rect 9484 8313 9496 8347
rect 9530 8344 9542 8347
rect 9766 8344 9772 8356
rect 9530 8316 9772 8344
rect 9530 8313 9542 8316
rect 9484 8307 9542 8313
rect 9766 8304 9772 8316
rect 9824 8304 9830 8356
rect 9876 8344 9904 8384
rect 12250 8372 12256 8384
rect 12308 8372 12314 8424
rect 12805 8415 12863 8421
rect 12805 8381 12817 8415
rect 12851 8412 12863 8415
rect 14090 8412 14096 8424
rect 12851 8384 14096 8412
rect 12851 8381 12863 8384
rect 12805 8375 12863 8381
rect 14090 8372 14096 8384
rect 14148 8372 14154 8424
rect 14458 8421 14464 8424
rect 14452 8412 14464 8421
rect 14419 8384 14464 8412
rect 14452 8375 14464 8384
rect 14458 8372 14464 8375
rect 14516 8372 14522 8424
rect 16776 8421 16804 8452
rect 17034 8440 17040 8452
rect 17092 8480 17098 8492
rect 18693 8483 18751 8489
rect 18693 8480 18705 8483
rect 17092 8452 18705 8480
rect 17092 8440 17098 8452
rect 18693 8449 18705 8452
rect 18739 8480 18751 8483
rect 18782 8480 18788 8492
rect 18739 8452 18788 8480
rect 18739 8449 18751 8452
rect 18693 8443 18751 8449
rect 18782 8440 18788 8452
rect 18840 8440 18846 8492
rect 20530 8480 20536 8492
rect 20491 8452 20536 8480
rect 20530 8440 20536 8452
rect 20588 8440 20594 8492
rect 20625 8483 20683 8489
rect 20625 8449 20637 8483
rect 20671 8449 20683 8483
rect 20625 8443 20683 8449
rect 16761 8415 16819 8421
rect 16761 8381 16773 8415
rect 16807 8381 16819 8415
rect 20640 8412 20668 8443
rect 16761 8375 16819 8381
rect 20548 8384 20668 8412
rect 20548 8356 20576 8384
rect 12897 8347 12955 8353
rect 12897 8344 12909 8347
rect 9876 8316 12909 8344
rect 12897 8313 12909 8316
rect 12943 8313 12955 8347
rect 12897 8307 12955 8313
rect 13262 8304 13268 8356
rect 13320 8344 13326 8356
rect 13630 8344 13636 8356
rect 13320 8316 13636 8344
rect 13320 8304 13326 8316
rect 13630 8304 13636 8316
rect 13688 8304 13694 8356
rect 15286 8304 15292 8356
rect 15344 8344 15350 8356
rect 16574 8344 16580 8356
rect 15344 8316 16580 8344
rect 15344 8304 15350 8316
rect 16574 8304 16580 8316
rect 16632 8304 16638 8356
rect 16853 8347 16911 8353
rect 16853 8313 16865 8347
rect 16899 8344 16911 8347
rect 17862 8344 17868 8356
rect 16899 8316 17868 8344
rect 16899 8313 16911 8316
rect 16853 8307 16911 8313
rect 17862 8304 17868 8316
rect 17920 8304 17926 8356
rect 17972 8316 18552 8344
rect 11974 8276 11980 8288
rect 4540 8248 11980 8276
rect 4433 8239 4491 8245
rect 11974 8236 11980 8248
rect 12032 8276 12038 8288
rect 12158 8276 12164 8288
rect 12032 8248 12164 8276
rect 12032 8236 12038 8248
rect 12158 8236 12164 8248
rect 12216 8236 12222 8288
rect 15654 8236 15660 8288
rect 15712 8276 15718 8288
rect 16114 8276 16120 8288
rect 15712 8248 16120 8276
rect 15712 8236 15718 8248
rect 16114 8236 16120 8248
rect 16172 8236 16178 8288
rect 17586 8236 17592 8288
rect 17644 8276 17650 8288
rect 17972 8276 18000 8316
rect 17644 8248 18000 8276
rect 17644 8236 17650 8248
rect 18138 8236 18144 8288
rect 18196 8276 18202 8288
rect 18524 8285 18552 8316
rect 18966 8304 18972 8356
rect 19024 8344 19030 8356
rect 20441 8347 20499 8353
rect 20441 8344 20453 8347
rect 19024 8316 20453 8344
rect 19024 8304 19030 8316
rect 20441 8313 20453 8316
rect 20487 8313 20499 8347
rect 20441 8307 20499 8313
rect 20530 8304 20536 8356
rect 20588 8304 20594 8356
rect 18417 8279 18475 8285
rect 18417 8276 18429 8279
rect 18196 8248 18429 8276
rect 18196 8236 18202 8248
rect 18417 8245 18429 8248
rect 18463 8245 18475 8279
rect 18417 8239 18475 8245
rect 18509 8279 18567 8285
rect 18509 8245 18521 8279
rect 18555 8245 18567 8279
rect 20070 8276 20076 8288
rect 20031 8248 20076 8276
rect 18509 8239 18567 8245
rect 20070 8236 20076 8248
rect 20128 8236 20134 8288
rect 1104 8186 21896 8208
rect 1104 8134 7912 8186
rect 7964 8134 7976 8186
rect 8028 8134 8040 8186
rect 8092 8134 8104 8186
rect 8156 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 15035 8186
rect 15087 8134 21896 8186
rect 1104 8112 21896 8134
rect 1857 8075 1915 8081
rect 1857 8041 1869 8075
rect 1903 8072 1915 8075
rect 1946 8072 1952 8084
rect 1903 8044 1952 8072
rect 1903 8041 1915 8044
rect 1857 8035 1915 8041
rect 1946 8032 1952 8044
rect 2004 8032 2010 8084
rect 2133 8075 2191 8081
rect 2133 8041 2145 8075
rect 2179 8072 2191 8075
rect 2314 8072 2320 8084
rect 2179 8044 2320 8072
rect 2179 8041 2191 8044
rect 2133 8035 2191 8041
rect 2314 8032 2320 8044
rect 2372 8032 2378 8084
rect 6181 8075 6239 8081
rect 6181 8041 6193 8075
rect 6227 8072 6239 8075
rect 6546 8072 6552 8084
rect 6227 8044 6552 8072
rect 6227 8041 6239 8044
rect 6181 8035 6239 8041
rect 6546 8032 6552 8044
rect 6604 8032 6610 8084
rect 7101 8075 7159 8081
rect 7101 8041 7113 8075
rect 7147 8072 7159 8075
rect 7190 8072 7196 8084
rect 7147 8044 7196 8072
rect 7147 8041 7159 8044
rect 7101 8035 7159 8041
rect 7190 8032 7196 8044
rect 7248 8032 7254 8084
rect 7561 8075 7619 8081
rect 7561 8041 7573 8075
rect 7607 8072 7619 8075
rect 9677 8075 9735 8081
rect 7607 8044 9628 8072
rect 7607 8041 7619 8044
rect 7561 8035 7619 8041
rect 5068 8007 5126 8013
rect 5068 7973 5080 8007
rect 5114 8004 5126 8007
rect 5442 8004 5448 8016
rect 5114 7976 5448 8004
rect 5114 7973 5126 7976
rect 5068 7967 5126 7973
rect 5442 7964 5448 7976
rect 5500 7964 5506 8016
rect 9600 8004 9628 8044
rect 9677 8041 9689 8075
rect 9723 8072 9735 8075
rect 10226 8072 10232 8084
rect 9723 8044 10232 8072
rect 9723 8041 9735 8044
rect 9677 8035 9735 8041
rect 10226 8032 10232 8044
rect 10284 8032 10290 8084
rect 11146 8032 11152 8084
rect 11204 8072 11210 8084
rect 14734 8072 14740 8084
rect 11204 8044 14740 8072
rect 11204 8032 11210 8044
rect 14734 8032 14740 8044
rect 14792 8072 14798 8084
rect 15194 8072 15200 8084
rect 14792 8044 15200 8072
rect 14792 8032 14798 8044
rect 15194 8032 15200 8044
rect 15252 8032 15258 8084
rect 17497 8075 17555 8081
rect 17497 8041 17509 8075
rect 17543 8041 17555 8075
rect 17497 8035 17555 8041
rect 10502 8004 10508 8016
rect 9600 7976 10508 8004
rect 10502 7964 10508 7976
rect 10560 8004 10566 8016
rect 10686 8004 10692 8016
rect 10560 7976 10692 8004
rect 10560 7964 10566 7976
rect 10686 7964 10692 7976
rect 10744 7964 10750 8016
rect 11790 8013 11796 8016
rect 11784 8004 11796 8013
rect 11703 7976 11796 8004
rect 11784 7967 11796 7976
rect 11848 8004 11854 8016
rect 11974 8004 11980 8016
rect 11848 7976 11980 8004
rect 11790 7964 11796 7967
rect 11848 7964 11854 7976
rect 11974 7964 11980 7976
rect 12032 7964 12038 8016
rect 14274 7964 14280 8016
rect 14332 8004 14338 8016
rect 15534 8007 15592 8013
rect 15534 8004 15546 8007
rect 14332 7976 15546 8004
rect 14332 7964 14338 7976
rect 15534 7973 15546 7976
rect 15580 7973 15592 8007
rect 15534 7967 15592 7973
rect 15746 7964 15752 8016
rect 15804 8004 15810 8016
rect 16022 8004 16028 8016
rect 15804 7976 16028 8004
rect 15804 7964 15810 7976
rect 16022 7964 16028 7976
rect 16080 8004 16086 8016
rect 17512 8004 17540 8035
rect 18782 8032 18788 8084
rect 18840 8072 18846 8084
rect 19337 8075 19395 8081
rect 19337 8072 19349 8075
rect 18840 8044 19349 8072
rect 18840 8032 18846 8044
rect 19337 8041 19349 8044
rect 19383 8041 19395 8075
rect 19337 8035 19395 8041
rect 18224 8007 18282 8013
rect 16080 7976 18000 8004
rect 16080 7964 16086 7976
rect 2314 7896 2320 7948
rect 2372 7936 2378 7948
rect 2501 7939 2559 7945
rect 2501 7936 2513 7939
rect 2372 7908 2513 7936
rect 2372 7896 2378 7908
rect 2501 7905 2513 7908
rect 2547 7905 2559 7939
rect 2501 7899 2559 7905
rect 4801 7939 4859 7945
rect 4801 7905 4813 7939
rect 4847 7936 4859 7939
rect 4847 7908 6316 7936
rect 4847 7905 4859 7908
rect 4801 7899 4859 7905
rect 2406 7828 2412 7880
rect 2464 7868 2470 7880
rect 2590 7868 2596 7880
rect 2464 7840 2596 7868
rect 2464 7828 2470 7840
rect 2590 7828 2596 7840
rect 2648 7828 2654 7880
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7868 2835 7871
rect 2866 7868 2872 7880
rect 2823 7840 2872 7868
rect 2823 7837 2835 7840
rect 2777 7831 2835 7837
rect 2866 7828 2872 7840
rect 2924 7868 2930 7880
rect 4430 7868 4436 7880
rect 2924 7840 4436 7868
rect 2924 7828 2930 7840
rect 4430 7828 4436 7840
rect 4488 7828 4494 7880
rect 6288 7868 6316 7908
rect 6362 7896 6368 7948
rect 6420 7936 6426 7948
rect 7469 7939 7527 7945
rect 7469 7936 7481 7939
rect 6420 7908 7481 7936
rect 6420 7896 6426 7908
rect 7469 7905 7481 7908
rect 7515 7905 7527 7939
rect 7469 7899 7527 7905
rect 7834 7896 7840 7948
rect 7892 7936 7898 7948
rect 8849 7939 8907 7945
rect 8849 7936 8861 7939
rect 7892 7908 8861 7936
rect 7892 7896 7898 7908
rect 8849 7905 8861 7908
rect 8895 7905 8907 7939
rect 8849 7899 8907 7905
rect 9582 7896 9588 7948
rect 9640 7936 9646 7948
rect 10042 7936 10048 7948
rect 9640 7908 10048 7936
rect 9640 7896 9646 7908
rect 10042 7896 10048 7908
rect 10100 7896 10106 7948
rect 11238 7896 11244 7948
rect 11296 7936 11302 7948
rect 13909 7939 13967 7945
rect 13909 7936 13921 7939
rect 11296 7908 13921 7936
rect 11296 7896 11302 7908
rect 13909 7905 13921 7908
rect 13955 7905 13967 7939
rect 13909 7899 13967 7905
rect 14182 7896 14188 7948
rect 14240 7936 14246 7948
rect 15289 7939 15347 7945
rect 15289 7936 15301 7939
rect 14240 7908 15301 7936
rect 14240 7896 14246 7908
rect 15289 7905 15301 7908
rect 15335 7905 15347 7939
rect 15289 7899 15347 7905
rect 16574 7896 16580 7948
rect 16632 7936 16638 7948
rect 17972 7945 18000 7976
rect 18224 7973 18236 8007
rect 18270 8004 18282 8007
rect 18874 8004 18880 8016
rect 18270 7976 18880 8004
rect 18270 7973 18282 7976
rect 18224 7967 18282 7973
rect 18874 7964 18880 7976
rect 18932 7964 18938 8016
rect 17681 7939 17739 7945
rect 17681 7936 17693 7939
rect 16632 7908 17693 7936
rect 16632 7896 16638 7908
rect 17681 7905 17693 7908
rect 17727 7905 17739 7939
rect 17681 7899 17739 7905
rect 17957 7939 18015 7945
rect 17957 7905 17969 7939
rect 18003 7936 18015 7939
rect 19150 7936 19156 7948
rect 18003 7908 19156 7936
rect 18003 7905 18015 7908
rect 17957 7899 18015 7905
rect 19150 7896 19156 7908
rect 19208 7896 19214 7948
rect 6454 7868 6460 7880
rect 6288 7840 6460 7868
rect 6454 7828 6460 7840
rect 6512 7828 6518 7880
rect 6546 7828 6552 7880
rect 6604 7868 6610 7880
rect 7653 7871 7711 7877
rect 7653 7868 7665 7871
rect 6604 7840 7665 7868
rect 6604 7828 6610 7840
rect 7653 7837 7665 7840
rect 7699 7837 7711 7871
rect 10134 7868 10140 7880
rect 10095 7840 10140 7868
rect 7653 7831 7711 7837
rect 10134 7828 10140 7840
rect 10192 7828 10198 7880
rect 10318 7868 10324 7880
rect 10279 7840 10324 7868
rect 10318 7828 10324 7840
rect 10376 7828 10382 7880
rect 11514 7868 11520 7880
rect 11475 7840 11520 7868
rect 11514 7828 11520 7840
rect 11572 7828 11578 7880
rect 13078 7828 13084 7880
rect 13136 7868 13142 7880
rect 13538 7868 13544 7880
rect 13136 7840 13544 7868
rect 13136 7828 13142 7840
rect 13538 7828 13544 7840
rect 13596 7828 13602 7880
rect 13814 7828 13820 7880
rect 13872 7868 13878 7880
rect 14093 7871 14151 7877
rect 14093 7868 14105 7871
rect 13872 7840 14105 7868
rect 13872 7828 13878 7840
rect 14093 7837 14105 7840
rect 14139 7837 14151 7871
rect 14093 7831 14151 7837
rect 5902 7760 5908 7812
rect 5960 7800 5966 7812
rect 11054 7800 11060 7812
rect 5960 7772 11060 7800
rect 5960 7760 5966 7772
rect 11054 7760 11060 7772
rect 11112 7760 11118 7812
rect 14366 7800 14372 7812
rect 12728 7772 14372 7800
rect 3786 7692 3792 7744
rect 3844 7732 3850 7744
rect 8386 7732 8392 7744
rect 3844 7704 8392 7732
rect 3844 7692 3850 7704
rect 8386 7692 8392 7704
rect 8444 7692 8450 7744
rect 8665 7735 8723 7741
rect 8665 7701 8677 7735
rect 8711 7732 8723 7735
rect 9122 7732 9128 7744
rect 8711 7704 9128 7732
rect 8711 7701 8723 7704
rect 8665 7695 8723 7701
rect 9122 7692 9128 7704
rect 9180 7692 9186 7744
rect 9490 7692 9496 7744
rect 9548 7732 9554 7744
rect 10962 7732 10968 7744
rect 9548 7704 10968 7732
rect 9548 7692 9554 7704
rect 10962 7692 10968 7704
rect 11020 7692 11026 7744
rect 12158 7692 12164 7744
rect 12216 7732 12222 7744
rect 12728 7732 12756 7772
rect 14366 7760 14372 7772
rect 14424 7760 14430 7812
rect 12894 7732 12900 7744
rect 12216 7704 12756 7732
rect 12855 7704 12900 7732
rect 12216 7692 12222 7704
rect 12894 7692 12900 7704
rect 12952 7732 12958 7744
rect 13998 7732 14004 7744
rect 12952 7704 14004 7732
rect 12952 7692 12958 7704
rect 13998 7692 14004 7704
rect 14056 7692 14062 7744
rect 15470 7692 15476 7744
rect 15528 7732 15534 7744
rect 16669 7735 16727 7741
rect 16669 7732 16681 7735
rect 15528 7704 16681 7732
rect 15528 7692 15534 7704
rect 16669 7701 16681 7704
rect 16715 7701 16727 7735
rect 16669 7695 16727 7701
rect 1104 7642 21896 7664
rect 1104 7590 4447 7642
rect 4499 7590 4511 7642
rect 4563 7590 4575 7642
rect 4627 7590 4639 7642
rect 4691 7590 11378 7642
rect 11430 7590 11442 7642
rect 11494 7590 11506 7642
rect 11558 7590 11570 7642
rect 11622 7590 18308 7642
rect 18360 7590 18372 7642
rect 18424 7590 18436 7642
rect 18488 7590 18500 7642
rect 18552 7590 21896 7642
rect 1104 7568 21896 7590
rect 1394 7528 1400 7540
rect 1355 7500 1400 7528
rect 1394 7488 1400 7500
rect 1452 7488 1458 7540
rect 2130 7488 2136 7540
rect 2188 7528 2194 7540
rect 2409 7531 2467 7537
rect 2409 7528 2421 7531
rect 2188 7500 2421 7528
rect 2188 7488 2194 7500
rect 2409 7497 2421 7500
rect 2455 7497 2467 7531
rect 2409 7491 2467 7497
rect 3510 7488 3516 7540
rect 3568 7528 3574 7540
rect 3568 7500 4016 7528
rect 3568 7488 3574 7500
rect 3988 7469 4016 7500
rect 4154 7488 4160 7540
rect 4212 7528 4218 7540
rect 4801 7531 4859 7537
rect 4801 7528 4813 7531
rect 4212 7500 4813 7528
rect 4212 7488 4218 7500
rect 4801 7497 4813 7500
rect 4847 7497 4859 7531
rect 4801 7491 4859 7497
rect 7742 7488 7748 7540
rect 7800 7528 7806 7540
rect 9490 7528 9496 7540
rect 7800 7500 9496 7528
rect 7800 7488 7806 7500
rect 9490 7488 9496 7500
rect 9548 7488 9554 7540
rect 9766 7528 9772 7540
rect 9727 7500 9772 7528
rect 9766 7488 9772 7500
rect 9824 7488 9830 7540
rect 10134 7488 10140 7540
rect 10192 7528 10198 7540
rect 10597 7531 10655 7537
rect 10597 7528 10609 7531
rect 10192 7500 10609 7528
rect 10192 7488 10198 7500
rect 10597 7497 10609 7500
rect 10643 7497 10655 7531
rect 10597 7491 10655 7497
rect 12618 7488 12624 7540
rect 12676 7528 12682 7540
rect 14001 7531 14059 7537
rect 14001 7528 14013 7531
rect 12676 7500 14013 7528
rect 12676 7488 12682 7500
rect 14001 7497 14013 7500
rect 14047 7497 14059 7531
rect 14001 7491 14059 7497
rect 14182 7488 14188 7540
rect 14240 7528 14246 7540
rect 18782 7528 18788 7540
rect 14240 7500 18788 7528
rect 14240 7488 14246 7500
rect 18782 7488 18788 7500
rect 18840 7488 18846 7540
rect 19794 7528 19800 7540
rect 18883 7500 19800 7528
rect 3973 7463 4031 7469
rect 3973 7429 3985 7463
rect 4019 7429 4031 7463
rect 3973 7423 4031 7429
rect 1762 7352 1768 7404
rect 1820 7392 1826 7404
rect 1949 7395 2007 7401
rect 1949 7392 1961 7395
rect 1820 7364 1961 7392
rect 1820 7352 1826 7364
rect 1949 7361 1961 7364
rect 1995 7361 2007 7395
rect 3988 7392 4016 7423
rect 5353 7395 5411 7401
rect 5353 7392 5365 7395
rect 3988 7364 5365 7392
rect 1949 7355 2007 7361
rect 5353 7361 5365 7364
rect 5399 7361 5411 7395
rect 5353 7355 5411 7361
rect 5442 7352 5448 7404
rect 5500 7392 5506 7404
rect 7377 7395 7435 7401
rect 7377 7392 7389 7395
rect 5500 7364 7389 7392
rect 5500 7352 5506 7364
rect 7377 7361 7389 7364
rect 7423 7361 7435 7395
rect 9784 7392 9812 7488
rect 12253 7463 12311 7469
rect 12253 7429 12265 7463
rect 12299 7460 12311 7463
rect 12437 7463 12495 7469
rect 12437 7460 12449 7463
rect 12299 7432 12449 7460
rect 12299 7429 12311 7432
rect 12253 7423 12311 7429
rect 12437 7429 12449 7432
rect 12483 7429 12495 7463
rect 12437 7423 12495 7429
rect 12526 7420 12532 7472
rect 12584 7460 12590 7472
rect 12584 7432 12940 7460
rect 12584 7420 12590 7432
rect 12912 7401 12940 7432
rect 12986 7420 12992 7472
rect 13044 7460 13050 7472
rect 13044 7432 13124 7460
rect 13044 7420 13050 7432
rect 13096 7401 13124 7432
rect 17034 7420 17040 7472
rect 17092 7460 17098 7472
rect 18883 7460 18911 7500
rect 19794 7488 19800 7500
rect 19852 7488 19858 7540
rect 20622 7488 20628 7540
rect 20680 7528 20686 7540
rect 20809 7531 20867 7537
rect 20809 7528 20821 7531
rect 20680 7500 20821 7528
rect 20680 7488 20686 7500
rect 20809 7497 20821 7500
rect 20855 7497 20867 7531
rect 20809 7491 20867 7497
rect 17092 7432 18911 7460
rect 17092 7420 17098 7432
rect 11149 7395 11207 7401
rect 11149 7392 11161 7395
rect 9784 7364 11161 7392
rect 7377 7355 7435 7361
rect 11149 7361 11161 7364
rect 11195 7361 11207 7395
rect 11149 7355 11207 7361
rect 12897 7395 12955 7401
rect 12897 7361 12909 7395
rect 12943 7361 12955 7395
rect 12897 7355 12955 7361
rect 13081 7395 13139 7401
rect 13081 7361 13093 7395
rect 13127 7361 13139 7395
rect 13081 7355 13139 7361
rect 13998 7352 14004 7404
rect 14056 7392 14062 7404
rect 14553 7395 14611 7401
rect 14553 7392 14565 7395
rect 14056 7364 14565 7392
rect 14056 7352 14062 7364
rect 14553 7361 14565 7364
rect 14599 7361 14611 7395
rect 14553 7355 14611 7361
rect 15746 7352 15752 7404
rect 15804 7392 15810 7404
rect 18138 7392 18144 7404
rect 15804 7364 15849 7392
rect 18099 7364 18144 7392
rect 15804 7352 15810 7364
rect 18138 7352 18144 7364
rect 18196 7352 18202 7404
rect 19150 7352 19156 7404
rect 19208 7392 19214 7404
rect 19429 7395 19487 7401
rect 19429 7392 19441 7395
rect 19208 7364 19441 7392
rect 19208 7352 19214 7364
rect 19429 7361 19441 7364
rect 19475 7361 19487 7395
rect 19429 7355 19487 7361
rect 1578 7284 1584 7336
rect 1636 7324 1642 7336
rect 1857 7327 1915 7333
rect 1857 7324 1869 7327
rect 1636 7296 1869 7324
rect 1636 7284 1642 7296
rect 1857 7293 1869 7296
rect 1903 7293 1915 7327
rect 2222 7324 2228 7336
rect 2183 7296 2228 7324
rect 1857 7287 1915 7293
rect 2222 7284 2228 7296
rect 2280 7284 2286 7336
rect 2593 7327 2651 7333
rect 2593 7293 2605 7327
rect 2639 7324 2651 7327
rect 3878 7324 3884 7336
rect 2639 7296 3884 7324
rect 2639 7293 2651 7296
rect 2593 7287 2651 7293
rect 3878 7284 3884 7296
rect 3936 7284 3942 7336
rect 4338 7284 4344 7336
rect 4396 7324 4402 7336
rect 5169 7327 5227 7333
rect 5169 7324 5181 7327
rect 4396 7296 5181 7324
rect 4396 7284 4402 7296
rect 5169 7293 5181 7296
rect 5215 7293 5227 7327
rect 5169 7287 5227 7293
rect 6454 7284 6460 7336
rect 6512 7324 6518 7336
rect 8389 7327 8447 7333
rect 8389 7324 8401 7327
rect 6512 7296 8401 7324
rect 6512 7284 6518 7296
rect 8389 7293 8401 7296
rect 8435 7324 8447 7327
rect 9122 7324 9128 7336
rect 8435 7296 9128 7324
rect 8435 7293 8447 7296
rect 8389 7287 8447 7293
rect 9122 7284 9128 7296
rect 9180 7284 9186 7336
rect 11054 7324 11060 7336
rect 10967 7296 11060 7324
rect 11054 7284 11060 7296
rect 11112 7324 11118 7336
rect 14182 7324 14188 7336
rect 11112 7296 14188 7324
rect 11112 7284 11118 7296
rect 14182 7284 14188 7296
rect 14240 7284 14246 7336
rect 19702 7333 19708 7336
rect 19696 7324 19708 7333
rect 19663 7296 19708 7324
rect 19696 7287 19708 7296
rect 19702 7284 19708 7287
rect 19760 7284 19766 7336
rect 1765 7259 1823 7265
rect 1765 7225 1777 7259
rect 1811 7256 1823 7259
rect 2498 7256 2504 7268
rect 1811 7228 2504 7256
rect 1811 7225 1823 7228
rect 1765 7219 1823 7225
rect 2498 7216 2504 7228
rect 2556 7216 2562 7268
rect 2866 7265 2872 7268
rect 2860 7256 2872 7265
rect 2827 7228 2872 7256
rect 2860 7219 2872 7228
rect 2866 7216 2872 7219
rect 2924 7216 2930 7268
rect 5902 7216 5908 7268
rect 5960 7256 5966 7268
rect 7285 7259 7343 7265
rect 7285 7256 7297 7259
rect 5960 7228 7297 7256
rect 5960 7216 5966 7228
rect 7285 7225 7297 7228
rect 7331 7256 7343 7259
rect 7742 7256 7748 7268
rect 7331 7228 7748 7256
rect 7331 7225 7343 7228
rect 7285 7219 7343 7225
rect 7742 7216 7748 7228
rect 7800 7216 7806 7268
rect 8478 7216 8484 7268
rect 8536 7256 8542 7268
rect 8634 7259 8692 7265
rect 8634 7256 8646 7259
rect 8536 7228 8646 7256
rect 8536 7216 8542 7228
rect 8634 7225 8646 7228
rect 8680 7225 8692 7259
rect 12158 7256 12164 7268
rect 8634 7219 8692 7225
rect 8772 7228 12164 7256
rect 5261 7191 5319 7197
rect 5261 7157 5273 7191
rect 5307 7188 5319 7191
rect 6546 7188 6552 7200
rect 5307 7160 6552 7188
rect 5307 7157 5319 7160
rect 5261 7151 5319 7157
rect 6546 7148 6552 7160
rect 6604 7148 6610 7200
rect 6822 7188 6828 7200
rect 6783 7160 6828 7188
rect 6822 7148 6828 7160
rect 6880 7148 6886 7200
rect 7190 7188 7196 7200
rect 7151 7160 7196 7188
rect 7190 7148 7196 7160
rect 7248 7188 7254 7200
rect 7374 7188 7380 7200
rect 7248 7160 7380 7188
rect 7248 7148 7254 7160
rect 7374 7148 7380 7160
rect 7432 7148 7438 7200
rect 7558 7148 7564 7200
rect 7616 7188 7622 7200
rect 8772 7188 8800 7228
rect 12158 7216 12164 7228
rect 12216 7216 12222 7268
rect 12253 7259 12311 7265
rect 12253 7225 12265 7259
rect 12299 7256 12311 7259
rect 14461 7259 14519 7265
rect 14461 7256 14473 7259
rect 12299 7228 14473 7256
rect 12299 7225 12311 7228
rect 12253 7219 12311 7225
rect 14461 7225 14473 7228
rect 14507 7225 14519 7259
rect 14461 7219 14519 7225
rect 16016 7259 16074 7265
rect 16016 7225 16028 7259
rect 16062 7256 16074 7259
rect 20530 7256 20536 7268
rect 16062 7228 20536 7256
rect 16062 7225 16074 7228
rect 16016 7219 16074 7225
rect 20530 7216 20536 7228
rect 20588 7216 20594 7268
rect 7616 7160 8800 7188
rect 7616 7148 7622 7160
rect 9490 7148 9496 7200
rect 9548 7188 9554 7200
rect 10965 7191 11023 7197
rect 10965 7188 10977 7191
rect 9548 7160 10977 7188
rect 9548 7148 9554 7160
rect 10965 7157 10977 7160
rect 11011 7188 11023 7191
rect 11146 7188 11152 7200
rect 11011 7160 11152 7188
rect 11011 7157 11023 7160
rect 10965 7151 11023 7157
rect 11146 7148 11152 7160
rect 11204 7148 11210 7200
rect 12805 7191 12863 7197
rect 12805 7157 12817 7191
rect 12851 7188 12863 7191
rect 13078 7188 13084 7200
rect 12851 7160 13084 7188
rect 12851 7157 12863 7160
rect 12805 7151 12863 7157
rect 13078 7148 13084 7160
rect 13136 7148 13142 7200
rect 14366 7188 14372 7200
rect 14327 7160 14372 7188
rect 14366 7148 14372 7160
rect 14424 7148 14430 7200
rect 15286 7148 15292 7200
rect 15344 7188 15350 7200
rect 17129 7191 17187 7197
rect 17129 7188 17141 7191
rect 15344 7160 17141 7188
rect 15344 7148 15350 7160
rect 17129 7157 17141 7160
rect 17175 7157 17187 7191
rect 17129 7151 17187 7157
rect 1104 7098 21896 7120
rect 1104 7046 7912 7098
rect 7964 7046 7976 7098
rect 8028 7046 8040 7098
rect 8092 7046 8104 7098
rect 8156 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 15035 7098
rect 15087 7046 21896 7098
rect 1104 7024 21896 7046
rect 2222 6944 2228 6996
rect 2280 6984 2286 6996
rect 2317 6987 2375 6993
rect 2317 6984 2329 6987
rect 2280 6956 2329 6984
rect 2280 6944 2286 6956
rect 2317 6953 2329 6956
rect 2363 6984 2375 6987
rect 2774 6984 2780 6996
rect 2363 6956 2780 6984
rect 2363 6953 2375 6956
rect 2317 6947 2375 6953
rect 2774 6944 2780 6956
rect 2832 6944 2838 6996
rect 4890 6944 4896 6996
rect 4948 6984 4954 6996
rect 8205 6987 8263 6993
rect 8205 6984 8217 6987
rect 4948 6956 8217 6984
rect 4948 6944 4954 6956
rect 8205 6953 8217 6956
rect 8251 6953 8263 6987
rect 8205 6947 8263 6953
rect 8386 6944 8392 6996
rect 8444 6984 8450 6996
rect 12250 6984 12256 6996
rect 8444 6956 12256 6984
rect 8444 6944 8450 6956
rect 12250 6944 12256 6956
rect 12308 6944 12314 6996
rect 12437 6987 12495 6993
rect 12437 6953 12449 6987
rect 12483 6984 12495 6987
rect 12618 6984 12624 6996
rect 12483 6956 12624 6984
rect 12483 6953 12495 6956
rect 12437 6947 12495 6953
rect 12618 6944 12624 6956
rect 12676 6944 12682 6996
rect 13262 6944 13268 6996
rect 13320 6984 13326 6996
rect 14001 6987 14059 6993
rect 14001 6984 14013 6987
rect 13320 6956 14013 6984
rect 13320 6944 13326 6956
rect 14001 6953 14013 6956
rect 14047 6953 14059 6987
rect 14001 6947 14059 6953
rect 14093 6987 14151 6993
rect 14093 6953 14105 6987
rect 14139 6984 14151 6987
rect 14458 6984 14464 6996
rect 14139 6956 14464 6984
rect 14139 6953 14151 6956
rect 14093 6947 14151 6953
rect 14458 6944 14464 6956
rect 14516 6944 14522 6996
rect 15746 6944 15752 6996
rect 15804 6984 15810 6996
rect 17034 6984 17040 6996
rect 15804 6956 17040 6984
rect 15804 6944 15810 6956
rect 17034 6944 17040 6956
rect 17092 6944 17098 6996
rect 5077 6919 5135 6925
rect 5077 6885 5089 6919
rect 5123 6916 5135 6919
rect 6454 6916 6460 6928
rect 5123 6888 6460 6916
rect 5123 6885 5135 6888
rect 5077 6879 5135 6885
rect 6454 6876 6460 6888
rect 6512 6876 6518 6928
rect 6546 6876 6552 6928
rect 6604 6916 6610 6928
rect 6604 6888 6868 6916
rect 6604 6876 6610 6888
rect 2866 6848 2872 6860
rect 2827 6820 2872 6848
rect 2866 6808 2872 6820
rect 2924 6808 2930 6860
rect 4246 6808 4252 6860
rect 4304 6848 4310 6860
rect 5169 6851 5227 6857
rect 5169 6848 5181 6851
rect 4304 6820 5181 6848
rect 4304 6808 4310 6820
rect 5169 6817 5181 6820
rect 5215 6817 5227 6851
rect 5169 6811 5227 6817
rect 6641 6851 6699 6857
rect 6641 6817 6653 6851
rect 6687 6817 6699 6851
rect 6840 6848 6868 6888
rect 8128 6888 8340 6916
rect 8128 6848 8156 6888
rect 6840 6820 8156 6848
rect 8312 6848 8340 6888
rect 9766 6876 9772 6928
rect 9824 6916 9830 6928
rect 10594 6916 10600 6928
rect 9824 6888 10600 6916
rect 9824 6876 9830 6888
rect 10594 6876 10600 6888
rect 10652 6876 10658 6928
rect 10870 6876 10876 6928
rect 10928 6916 10934 6928
rect 12158 6916 12164 6928
rect 10928 6888 12164 6916
rect 10928 6876 10934 6888
rect 12158 6876 12164 6888
rect 12216 6876 12222 6928
rect 12526 6876 12532 6928
rect 12584 6916 12590 6928
rect 17954 6916 17960 6928
rect 12584 6888 17960 6916
rect 12584 6876 12590 6888
rect 17954 6876 17960 6888
rect 18012 6876 18018 6928
rect 10042 6848 10048 6860
rect 8312 6820 8524 6848
rect 10003 6820 10048 6848
rect 6641 6811 6699 6817
rect 2958 6780 2964 6792
rect 2919 6752 2964 6780
rect 2958 6740 2964 6752
rect 3016 6740 3022 6792
rect 5353 6783 5411 6789
rect 5353 6749 5365 6783
rect 5399 6780 5411 6783
rect 5442 6780 5448 6792
rect 5399 6752 5448 6780
rect 5399 6749 5411 6752
rect 5353 6743 5411 6749
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 4709 6715 4767 6721
rect 4709 6681 4721 6715
rect 4755 6712 4767 6715
rect 6656 6712 6684 6811
rect 6733 6783 6791 6789
rect 6733 6749 6745 6783
rect 6779 6780 6791 6783
rect 6822 6780 6828 6792
rect 6779 6752 6828 6780
rect 6779 6749 6791 6752
rect 6733 6743 6791 6749
rect 6822 6740 6828 6752
rect 6880 6740 6886 6792
rect 6917 6783 6975 6789
rect 6917 6749 6929 6783
rect 6963 6749 6975 6783
rect 6917 6743 6975 6749
rect 4755 6684 6684 6712
rect 6932 6712 6960 6743
rect 7006 6740 7012 6792
rect 7064 6780 7070 6792
rect 8297 6783 8355 6789
rect 8297 6780 8309 6783
rect 7064 6752 8309 6780
rect 7064 6740 7070 6752
rect 8297 6749 8309 6752
rect 8343 6749 8355 6783
rect 8297 6743 8355 6749
rect 8389 6783 8447 6789
rect 8389 6749 8401 6783
rect 8435 6749 8447 6783
rect 8389 6743 8447 6749
rect 7282 6712 7288 6724
rect 6932 6684 7288 6712
rect 4755 6681 4767 6684
rect 4709 6675 4767 6681
rect 7282 6672 7288 6684
rect 7340 6712 7346 6724
rect 8404 6712 8432 6743
rect 7340 6684 8432 6712
rect 8496 6712 8524 6820
rect 10042 6808 10048 6820
rect 10100 6808 10106 6860
rect 12345 6851 12403 6857
rect 12345 6817 12357 6851
rect 12391 6848 12403 6851
rect 12434 6848 12440 6860
rect 12391 6820 12440 6848
rect 12391 6817 12403 6820
rect 12345 6811 12403 6817
rect 12434 6808 12440 6820
rect 12492 6808 12498 6860
rect 14182 6848 14188 6860
rect 13096 6820 14188 6848
rect 10134 6780 10140 6792
rect 10095 6752 10140 6780
rect 10134 6740 10140 6752
rect 10192 6740 10198 6792
rect 10318 6780 10324 6792
rect 10279 6752 10324 6780
rect 10318 6740 10324 6752
rect 10376 6740 10382 6792
rect 12618 6780 12624 6792
rect 12579 6752 12624 6780
rect 12618 6740 12624 6752
rect 12676 6740 12682 6792
rect 9677 6715 9735 6721
rect 9677 6712 9689 6715
rect 8496 6684 9689 6712
rect 7340 6672 7346 6684
rect 9677 6681 9689 6684
rect 9723 6681 9735 6715
rect 11238 6712 11244 6724
rect 9677 6675 9735 6681
rect 9876 6684 11244 6712
rect 2406 6644 2412 6656
rect 2367 6616 2412 6644
rect 2406 6604 2412 6616
rect 2464 6604 2470 6656
rect 6270 6644 6276 6656
rect 6231 6616 6276 6644
rect 6270 6604 6276 6616
rect 6328 6604 6334 6656
rect 7742 6604 7748 6656
rect 7800 6644 7806 6656
rect 7837 6647 7895 6653
rect 7837 6644 7849 6647
rect 7800 6616 7849 6644
rect 7800 6604 7806 6616
rect 7837 6613 7849 6616
rect 7883 6613 7895 6647
rect 7837 6607 7895 6613
rect 9582 6604 9588 6656
rect 9640 6644 9646 6656
rect 9876 6644 9904 6684
rect 11238 6672 11244 6684
rect 11296 6672 11302 6724
rect 11977 6715 12035 6721
rect 11977 6681 11989 6715
rect 12023 6712 12035 6715
rect 13096 6712 13124 6820
rect 14182 6808 14188 6820
rect 14240 6808 14246 6860
rect 15562 6808 15568 6860
rect 15620 6848 15626 6860
rect 16097 6851 16155 6857
rect 16097 6848 16109 6851
rect 15620 6820 16109 6848
rect 15620 6808 15626 6820
rect 16097 6817 16109 6820
rect 16143 6817 16155 6851
rect 19521 6851 19579 6857
rect 19521 6848 19533 6851
rect 16097 6811 16155 6817
rect 17972 6820 19533 6848
rect 17972 6792 18000 6820
rect 19521 6817 19533 6820
rect 19567 6817 19579 6851
rect 19521 6811 19579 6817
rect 14277 6783 14335 6789
rect 14277 6749 14289 6783
rect 14323 6780 14335 6783
rect 14366 6780 14372 6792
rect 14323 6752 14372 6780
rect 14323 6749 14335 6752
rect 14277 6743 14335 6749
rect 14366 6740 14372 6752
rect 14424 6740 14430 6792
rect 15746 6740 15752 6792
rect 15804 6780 15810 6792
rect 15841 6783 15899 6789
rect 15841 6780 15853 6783
rect 15804 6752 15853 6780
rect 15804 6740 15810 6752
rect 15841 6749 15853 6752
rect 15887 6749 15899 6783
rect 15841 6743 15899 6749
rect 17954 6740 17960 6792
rect 18012 6740 18018 6792
rect 18138 6780 18144 6792
rect 18099 6752 18144 6780
rect 18138 6740 18144 6752
rect 18196 6740 18202 6792
rect 19613 6783 19671 6789
rect 19613 6780 19625 6783
rect 19536 6752 19625 6780
rect 19536 6724 19564 6752
rect 19613 6749 19625 6752
rect 19659 6749 19671 6783
rect 19613 6743 19671 6749
rect 19705 6783 19763 6789
rect 19705 6749 19717 6783
rect 19751 6749 19763 6783
rect 19705 6743 19763 6749
rect 14458 6712 14464 6724
rect 12023 6684 13124 6712
rect 13188 6684 14464 6712
rect 12023 6681 12035 6684
rect 11977 6675 12035 6681
rect 9640 6616 9904 6644
rect 9640 6604 9646 6616
rect 9950 6604 9956 6656
rect 10008 6644 10014 6656
rect 13188 6644 13216 6684
rect 14458 6672 14464 6684
rect 14516 6672 14522 6724
rect 18874 6672 18880 6724
rect 18932 6712 18938 6724
rect 18932 6684 19472 6712
rect 18932 6672 18938 6684
rect 10008 6616 13216 6644
rect 13633 6647 13691 6653
rect 10008 6604 10014 6616
rect 13633 6613 13645 6647
rect 13679 6644 13691 6647
rect 15746 6644 15752 6656
rect 13679 6616 15752 6644
rect 13679 6613 13691 6616
rect 13633 6607 13691 6613
rect 15746 6604 15752 6616
rect 15804 6604 15810 6656
rect 17221 6647 17279 6653
rect 17221 6613 17233 6647
rect 17267 6644 17279 6647
rect 17310 6644 17316 6656
rect 17267 6616 17316 6644
rect 17267 6613 17279 6616
rect 17221 6607 17279 6613
rect 17310 6604 17316 6616
rect 17368 6604 17374 6656
rect 19150 6644 19156 6656
rect 19111 6616 19156 6644
rect 19150 6604 19156 6616
rect 19208 6604 19214 6656
rect 19444 6644 19472 6684
rect 19518 6672 19524 6724
rect 19576 6672 19582 6724
rect 19720 6644 19748 6743
rect 19444 6616 19748 6644
rect 1104 6554 21896 6576
rect 1104 6502 4447 6554
rect 4499 6502 4511 6554
rect 4563 6502 4575 6554
rect 4627 6502 4639 6554
rect 4691 6502 11378 6554
rect 11430 6502 11442 6554
rect 11494 6502 11506 6554
rect 11558 6502 11570 6554
rect 11622 6502 18308 6554
rect 18360 6502 18372 6554
rect 18424 6502 18436 6554
rect 18488 6502 18500 6554
rect 18552 6502 21896 6554
rect 1104 6480 21896 6502
rect 5905 6443 5963 6449
rect 2424 6412 5856 6440
rect 2038 6304 2044 6316
rect 1999 6276 2044 6304
rect 2038 6264 2044 6276
rect 2096 6264 2102 6316
rect 2225 6307 2283 6313
rect 2225 6273 2237 6307
rect 2271 6273 2283 6307
rect 2225 6267 2283 6273
rect 2240 6168 2268 6267
rect 2424 6245 2452 6412
rect 2590 6372 2596 6384
rect 2551 6344 2596 6372
rect 2590 6332 2596 6344
rect 2648 6332 2654 6384
rect 5828 6372 5856 6412
rect 5905 6409 5917 6443
rect 5951 6440 5963 6443
rect 7282 6440 7288 6452
rect 5951 6412 7288 6440
rect 5951 6409 5963 6412
rect 5905 6403 5963 6409
rect 7282 6400 7288 6412
rect 7340 6400 7346 6452
rect 8389 6443 8447 6449
rect 8389 6409 8401 6443
rect 8435 6440 8447 6443
rect 8478 6440 8484 6452
rect 8435 6412 8484 6440
rect 8435 6409 8447 6412
rect 8389 6403 8447 6409
rect 8478 6400 8484 6412
rect 8536 6400 8542 6452
rect 8570 6400 8576 6452
rect 8628 6440 8634 6452
rect 10318 6440 10324 6452
rect 8628 6412 10324 6440
rect 8628 6400 8634 6412
rect 10318 6400 10324 6412
rect 10376 6440 10382 6452
rect 10781 6443 10839 6449
rect 10781 6440 10793 6443
rect 10376 6412 10793 6440
rect 10376 6400 10382 6412
rect 10781 6409 10793 6412
rect 10827 6409 10839 6443
rect 10781 6403 10839 6409
rect 12618 6400 12624 6452
rect 12676 6440 12682 6452
rect 13817 6443 13875 6449
rect 13817 6440 13829 6443
rect 12676 6412 13829 6440
rect 12676 6400 12682 6412
rect 13817 6409 13829 6412
rect 13863 6409 13875 6443
rect 13817 6403 13875 6409
rect 14550 6400 14556 6452
rect 14608 6440 14614 6452
rect 14608 6412 15700 6440
rect 14608 6400 14614 6412
rect 6917 6375 6975 6381
rect 6917 6372 6929 6375
rect 5828 6344 6929 6372
rect 6917 6341 6929 6344
rect 6963 6341 6975 6375
rect 6917 6335 6975 6341
rect 15470 6332 15476 6384
rect 15528 6332 15534 6384
rect 2774 6264 2780 6316
rect 2832 6304 2838 6316
rect 3878 6304 3884 6316
rect 2832 6276 3884 6304
rect 2832 6264 2838 6276
rect 3878 6264 3884 6276
rect 3936 6304 3942 6316
rect 4522 6304 4528 6316
rect 3936 6276 4528 6304
rect 3936 6264 3942 6276
rect 4522 6264 4528 6276
rect 4580 6264 4586 6316
rect 14366 6264 14372 6316
rect 14424 6304 14430 6316
rect 15488 6304 15516 6332
rect 15565 6307 15623 6313
rect 15565 6304 15577 6307
rect 14424 6276 15577 6304
rect 14424 6264 14430 6276
rect 15565 6273 15577 6276
rect 15611 6273 15623 6307
rect 15565 6267 15623 6273
rect 2409 6239 2467 6245
rect 2409 6205 2421 6239
rect 2455 6205 2467 6239
rect 2409 6199 2467 6205
rect 3421 6239 3479 6245
rect 3421 6205 3433 6239
rect 3467 6236 3479 6239
rect 4338 6236 4344 6248
rect 3467 6208 4344 6236
rect 3467 6205 3479 6208
rect 3421 6199 3479 6205
rect 4338 6196 4344 6208
rect 4396 6196 4402 6248
rect 4614 6196 4620 6248
rect 4672 6236 4678 6248
rect 4672 6208 6776 6236
rect 4672 6196 4678 6208
rect 2958 6168 2964 6180
rect 2240 6140 2964 6168
rect 2958 6128 2964 6140
rect 3016 6128 3022 6180
rect 4792 6171 4850 6177
rect 4792 6168 4804 6171
rect 3528 6140 4804 6168
rect 1581 6103 1639 6109
rect 1581 6069 1593 6103
rect 1627 6100 1639 6103
rect 1670 6100 1676 6112
rect 1627 6072 1676 6100
rect 1627 6069 1639 6072
rect 1581 6063 1639 6069
rect 1670 6060 1676 6072
rect 1728 6060 1734 6112
rect 1946 6100 1952 6112
rect 1907 6072 1952 6100
rect 1946 6060 1952 6072
rect 2004 6060 2010 6112
rect 2682 6060 2688 6112
rect 2740 6100 2746 6112
rect 3528 6100 3556 6140
rect 4792 6137 4804 6140
rect 4838 6137 4850 6171
rect 6748 6168 6776 6208
rect 6914 6196 6920 6248
rect 6972 6236 6978 6248
rect 7282 6245 7288 6248
rect 7009 6239 7067 6245
rect 7009 6236 7021 6239
rect 6972 6208 7021 6236
rect 6972 6196 6978 6208
rect 7009 6205 7021 6208
rect 7055 6205 7067 6239
rect 7276 6236 7288 6245
rect 7243 6208 7288 6236
rect 7009 6199 7067 6205
rect 7276 6199 7288 6208
rect 7282 6196 7288 6199
rect 7340 6196 7346 6248
rect 9122 6196 9128 6248
rect 9180 6236 9186 6248
rect 9401 6239 9459 6245
rect 9401 6236 9413 6239
rect 9180 6208 9413 6236
rect 9180 6196 9186 6208
rect 9401 6205 9413 6208
rect 9447 6205 9459 6239
rect 9950 6236 9956 6248
rect 9401 6199 9459 6205
rect 9499 6208 9956 6236
rect 9499 6168 9527 6208
rect 9950 6196 9956 6208
rect 10008 6196 10014 6248
rect 10686 6236 10692 6248
rect 10612 6208 10692 6236
rect 6748 6140 9527 6168
rect 9668 6171 9726 6177
rect 4792 6131 4850 6137
rect 9668 6137 9680 6171
rect 9714 6168 9726 6171
rect 10612 6168 10640 6208
rect 10686 6196 10692 6208
rect 10744 6196 10750 6248
rect 11974 6196 11980 6248
rect 12032 6236 12038 6248
rect 12342 6236 12348 6248
rect 12032 6208 12348 6236
rect 12032 6196 12038 6208
rect 12342 6196 12348 6208
rect 12400 6236 12406 6248
rect 12437 6239 12495 6245
rect 12437 6236 12449 6239
rect 12400 6208 12449 6236
rect 12400 6196 12406 6208
rect 12437 6205 12449 6208
rect 12483 6205 12495 6239
rect 12437 6199 12495 6205
rect 15381 6239 15439 6245
rect 15381 6205 15393 6239
rect 15427 6236 15439 6239
rect 15672 6236 15700 6412
rect 17954 6400 17960 6452
rect 18012 6440 18018 6452
rect 18049 6443 18107 6449
rect 18049 6440 18061 6443
rect 18012 6412 18061 6440
rect 18012 6400 18018 6412
rect 18049 6409 18061 6412
rect 18095 6409 18107 6443
rect 18049 6403 18107 6409
rect 17862 6332 17868 6384
rect 17920 6372 17926 6384
rect 17920 6344 18736 6372
rect 17920 6332 17926 6344
rect 16945 6307 17003 6313
rect 16945 6273 16957 6307
rect 16991 6304 17003 6307
rect 17126 6304 17132 6316
rect 16991 6276 17132 6304
rect 16991 6273 17003 6276
rect 16945 6267 17003 6273
rect 17126 6264 17132 6276
rect 17184 6264 17190 6316
rect 17310 6264 17316 6316
rect 17368 6304 17374 6316
rect 18601 6307 18659 6313
rect 18601 6304 18613 6307
rect 17368 6276 18613 6304
rect 17368 6264 17374 6276
rect 18601 6273 18613 6276
rect 18647 6273 18659 6307
rect 18601 6267 18659 6273
rect 15427 6208 15700 6236
rect 15427 6205 15439 6208
rect 15381 6199 15439 6205
rect 17402 6196 17408 6248
rect 17460 6236 17466 6248
rect 17770 6236 17776 6248
rect 17460 6208 17776 6236
rect 17460 6196 17466 6208
rect 17770 6196 17776 6208
rect 17828 6196 17834 6248
rect 18138 6196 18144 6248
rect 18196 6236 18202 6248
rect 18417 6239 18475 6245
rect 18417 6236 18429 6239
rect 18196 6208 18429 6236
rect 18196 6196 18202 6208
rect 18417 6205 18429 6208
rect 18463 6205 18475 6239
rect 18417 6199 18475 6205
rect 18509 6239 18567 6245
rect 18509 6205 18521 6239
rect 18555 6236 18567 6239
rect 18708 6236 18736 6344
rect 19426 6264 19432 6316
rect 19484 6304 19490 6316
rect 19613 6307 19671 6313
rect 19613 6304 19625 6307
rect 19484 6276 19625 6304
rect 19484 6264 19490 6276
rect 19613 6273 19625 6276
rect 19659 6273 19671 6307
rect 19613 6267 19671 6273
rect 18555 6208 18736 6236
rect 18555 6205 18567 6208
rect 18509 6199 18567 6205
rect 9714 6140 10640 6168
rect 12704 6171 12762 6177
rect 9714 6137 9726 6140
rect 9668 6131 9726 6137
rect 12704 6137 12716 6171
rect 12750 6168 12762 6171
rect 12894 6168 12900 6180
rect 12750 6140 12900 6168
rect 12750 6137 12762 6140
rect 12704 6131 12762 6137
rect 2740 6072 3556 6100
rect 2740 6060 2746 6072
rect 3602 6060 3608 6112
rect 3660 6100 3666 6112
rect 4816 6100 4844 6131
rect 12894 6128 12900 6140
rect 12952 6128 12958 6180
rect 12986 6128 12992 6180
rect 13044 6168 13050 6180
rect 15289 6171 15347 6177
rect 15289 6168 15301 6171
rect 13044 6140 15301 6168
rect 13044 6128 13050 6140
rect 15289 6137 15301 6140
rect 15335 6137 15347 6171
rect 15289 6131 15347 6137
rect 5166 6100 5172 6112
rect 3660 6072 3705 6100
rect 4816 6072 5172 6100
rect 3660 6060 3666 6072
rect 5166 6060 5172 6072
rect 5224 6100 5230 6112
rect 5442 6100 5448 6112
rect 5224 6072 5448 6100
rect 5224 6060 5230 6072
rect 5442 6060 5448 6072
rect 5500 6060 5506 6112
rect 6917 6103 6975 6109
rect 6917 6069 6929 6103
rect 6963 6100 6975 6103
rect 11698 6100 11704 6112
rect 6963 6072 11704 6100
rect 6963 6069 6975 6072
rect 6917 6063 6975 6069
rect 11698 6060 11704 6072
rect 11756 6060 11762 6112
rect 14921 6103 14979 6109
rect 14921 6069 14933 6103
rect 14967 6100 14979 6103
rect 15194 6100 15200 6112
rect 14967 6072 15200 6100
rect 14967 6069 14979 6072
rect 14921 6063 14979 6069
rect 15194 6060 15200 6072
rect 15252 6060 15258 6112
rect 15654 6060 15660 6112
rect 15712 6100 15718 6112
rect 20625 6103 20683 6109
rect 20625 6100 20637 6103
rect 15712 6072 20637 6100
rect 15712 6060 15718 6072
rect 20625 6069 20637 6072
rect 20671 6069 20683 6103
rect 20625 6063 20683 6069
rect 1104 6010 21896 6032
rect 1104 5958 7912 6010
rect 7964 5958 7976 6010
rect 8028 5958 8040 6010
rect 8092 5958 8104 6010
rect 8156 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 15035 6010
rect 15087 5958 21896 6010
rect 1104 5936 21896 5958
rect 1397 5899 1455 5905
rect 1397 5865 1409 5899
rect 1443 5865 1455 5899
rect 1397 5859 1455 5865
rect 1412 5828 1440 5859
rect 1946 5856 1952 5908
rect 2004 5896 2010 5908
rect 4065 5899 4123 5905
rect 4065 5896 4077 5899
rect 2004 5868 4077 5896
rect 2004 5856 2010 5868
rect 4065 5865 4077 5868
rect 4111 5865 4123 5899
rect 4065 5859 4123 5865
rect 4154 5856 4160 5908
rect 4212 5896 4218 5908
rect 5258 5896 5264 5908
rect 4212 5868 5264 5896
rect 4212 5856 4218 5868
rect 5258 5856 5264 5868
rect 5316 5856 5322 5908
rect 7006 5896 7012 5908
rect 5368 5868 7012 5896
rect 5368 5828 5396 5868
rect 7006 5856 7012 5868
rect 7064 5856 7070 5908
rect 7742 5856 7748 5908
rect 7800 5896 7806 5908
rect 8021 5899 8079 5905
rect 8021 5896 8033 5899
rect 7800 5868 8033 5896
rect 7800 5856 7806 5868
rect 8021 5865 8033 5868
rect 8067 5865 8079 5899
rect 10042 5896 10048 5908
rect 10003 5868 10048 5896
rect 8021 5859 8079 5865
rect 10042 5856 10048 5868
rect 10100 5856 10106 5908
rect 10413 5899 10471 5905
rect 10413 5865 10425 5899
rect 10459 5896 10471 5899
rect 10502 5896 10508 5908
rect 10459 5868 10508 5896
rect 10459 5865 10471 5868
rect 10413 5859 10471 5865
rect 10502 5856 10508 5868
rect 10560 5856 10566 5908
rect 10686 5856 10692 5908
rect 10744 5896 10750 5908
rect 10744 5868 14044 5896
rect 10744 5856 10750 5868
rect 1412 5800 5396 5828
rect 7374 5788 7380 5840
rect 7432 5828 7438 5840
rect 7929 5831 7987 5837
rect 7929 5828 7941 5831
rect 7432 5800 7941 5828
rect 7432 5788 7438 5800
rect 7929 5797 7941 5800
rect 7975 5797 7987 5831
rect 7929 5791 7987 5797
rect 8036 5800 8677 5828
rect 1762 5760 1768 5772
rect 1723 5732 1768 5760
rect 1762 5720 1768 5732
rect 1820 5720 1826 5772
rect 2777 5763 2835 5769
rect 2777 5729 2789 5763
rect 2823 5760 2835 5763
rect 4798 5760 4804 5772
rect 2823 5732 4804 5760
rect 2823 5729 2835 5732
rect 2777 5723 2835 5729
rect 4798 5720 4804 5732
rect 4856 5720 4862 5772
rect 5620 5763 5678 5769
rect 5620 5729 5632 5763
rect 5666 5760 5678 5763
rect 8036 5760 8064 5800
rect 5666 5732 8064 5760
rect 5666 5729 5678 5732
rect 5620 5723 5678 5729
rect 8386 5720 8392 5772
rect 8444 5760 8450 5772
rect 8649 5760 8677 5800
rect 8846 5788 8852 5840
rect 8904 5828 8910 5840
rect 10962 5828 10968 5840
rect 8904 5800 10968 5828
rect 8904 5788 8910 5800
rect 10962 5788 10968 5800
rect 11020 5788 11026 5840
rect 14016 5828 14044 5868
rect 14090 5856 14096 5908
rect 14148 5896 14154 5908
rect 14185 5899 14243 5905
rect 14185 5896 14197 5899
rect 14148 5868 14197 5896
rect 14148 5856 14154 5868
rect 14185 5865 14197 5868
rect 14231 5865 14243 5899
rect 14185 5859 14243 5865
rect 15194 5856 15200 5908
rect 15252 5896 15258 5908
rect 15657 5899 15715 5905
rect 15657 5896 15669 5899
rect 15252 5868 15669 5896
rect 15252 5856 15258 5868
rect 15657 5865 15669 5868
rect 15703 5865 15715 5899
rect 15657 5859 15715 5865
rect 15746 5856 15752 5908
rect 15804 5896 15810 5908
rect 15804 5868 15849 5896
rect 15804 5856 15810 5868
rect 16942 5856 16948 5908
rect 17000 5896 17006 5908
rect 18601 5899 18659 5905
rect 17000 5868 18092 5896
rect 17000 5856 17006 5868
rect 15286 5828 15292 5840
rect 11072 5800 13952 5828
rect 14016 5800 15292 5828
rect 10042 5760 10048 5772
rect 8444 5732 8616 5760
rect 8649 5732 10048 5760
rect 8444 5720 8450 5732
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5661 1915 5695
rect 1857 5655 1915 5661
rect 2041 5695 2099 5701
rect 2041 5661 2053 5695
rect 2087 5692 2099 5695
rect 2682 5692 2688 5704
rect 2087 5664 2688 5692
rect 2087 5661 2099 5664
rect 2041 5655 2099 5661
rect 1872 5624 1900 5655
rect 2682 5652 2688 5664
rect 2740 5652 2746 5704
rect 2866 5692 2872 5704
rect 2827 5664 2872 5692
rect 2866 5652 2872 5664
rect 2924 5652 2930 5704
rect 2961 5695 3019 5701
rect 2961 5661 2973 5695
rect 3007 5661 3019 5695
rect 2961 5655 3019 5661
rect 2317 5627 2375 5633
rect 2317 5624 2329 5627
rect 1872 5596 2329 5624
rect 2317 5593 2329 5596
rect 2363 5624 2375 5627
rect 2498 5624 2504 5636
rect 2363 5596 2504 5624
rect 2363 5593 2375 5596
rect 2317 5587 2375 5593
rect 2498 5584 2504 5596
rect 2556 5584 2562 5636
rect 2590 5584 2596 5636
rect 2648 5624 2654 5636
rect 2976 5624 3004 5655
rect 4522 5652 4528 5704
rect 4580 5692 4586 5704
rect 5353 5695 5411 5701
rect 5353 5692 5365 5695
rect 4580 5664 5365 5692
rect 4580 5652 4586 5664
rect 5353 5661 5365 5664
rect 5399 5661 5411 5695
rect 5353 5655 5411 5661
rect 8205 5695 8263 5701
rect 8205 5661 8217 5695
rect 8251 5692 8263 5695
rect 8478 5692 8484 5704
rect 8251 5664 8484 5692
rect 8251 5661 8263 5664
rect 8205 5655 8263 5661
rect 8478 5652 8484 5664
rect 8536 5652 8542 5704
rect 8588 5692 8616 5732
rect 10042 5720 10048 5732
rect 10100 5720 10106 5772
rect 11072 5760 11100 5800
rect 10152 5732 11100 5760
rect 12244 5763 12302 5769
rect 10152 5692 10180 5732
rect 12244 5729 12256 5763
rect 12290 5760 12302 5763
rect 12618 5760 12624 5772
rect 12290 5732 12624 5760
rect 12290 5729 12302 5732
rect 12244 5723 12302 5729
rect 12618 5720 12624 5732
rect 12676 5720 12682 5772
rect 10502 5692 10508 5704
rect 8588 5664 10180 5692
rect 10463 5664 10508 5692
rect 10502 5652 10508 5664
rect 10560 5652 10566 5704
rect 10686 5692 10692 5704
rect 10647 5664 10692 5692
rect 10686 5652 10692 5664
rect 10744 5652 10750 5704
rect 11974 5692 11980 5704
rect 11935 5664 11980 5692
rect 11974 5652 11980 5664
rect 12032 5652 12038 5704
rect 13924 5692 13952 5800
rect 15286 5788 15292 5800
rect 15344 5788 15350 5840
rect 17954 5828 17960 5840
rect 15396 5800 17960 5828
rect 15396 5692 15424 5800
rect 17954 5788 17960 5800
rect 18012 5788 18018 5840
rect 17034 5720 17040 5772
rect 17092 5760 17098 5772
rect 17221 5763 17279 5769
rect 17221 5760 17233 5763
rect 17092 5732 17233 5760
rect 17092 5720 17098 5732
rect 17221 5729 17233 5732
rect 17267 5729 17279 5763
rect 17221 5723 17279 5729
rect 17310 5720 17316 5772
rect 17368 5760 17374 5772
rect 17494 5769 17500 5772
rect 17488 5760 17500 5769
rect 17368 5732 17500 5760
rect 17368 5720 17374 5732
rect 17488 5723 17500 5732
rect 17494 5720 17500 5723
rect 17552 5720 17558 5772
rect 18064 5760 18092 5868
rect 18601 5865 18613 5899
rect 18647 5896 18659 5899
rect 18874 5896 18880 5908
rect 18647 5868 18880 5896
rect 18647 5865 18659 5868
rect 18601 5859 18659 5865
rect 18874 5856 18880 5868
rect 18932 5856 18938 5908
rect 19705 5831 19763 5837
rect 19705 5797 19717 5831
rect 19751 5828 19763 5831
rect 19886 5828 19892 5840
rect 19751 5800 19892 5828
rect 19751 5797 19763 5800
rect 19705 5791 19763 5797
rect 19886 5788 19892 5800
rect 19944 5788 19950 5840
rect 19429 5763 19487 5769
rect 19429 5760 19441 5763
rect 18064 5732 19441 5760
rect 19429 5729 19441 5732
rect 19475 5729 19487 5763
rect 19429 5723 19487 5729
rect 13924 5664 15424 5692
rect 15562 5652 15568 5704
rect 15620 5692 15626 5704
rect 15841 5695 15899 5701
rect 15841 5692 15853 5695
rect 15620 5664 15853 5692
rect 15620 5652 15626 5664
rect 15841 5661 15853 5664
rect 15887 5661 15899 5695
rect 15841 5655 15899 5661
rect 15930 5652 15936 5704
rect 15988 5692 15994 5704
rect 17126 5692 17132 5704
rect 15988 5664 17132 5692
rect 15988 5652 15994 5664
rect 17126 5652 17132 5664
rect 17184 5652 17190 5704
rect 2648 5596 3004 5624
rect 2648 5584 2654 5596
rect 3326 5584 3332 5636
rect 3384 5624 3390 5636
rect 5258 5624 5264 5636
rect 3384 5596 5264 5624
rect 3384 5584 3390 5596
rect 5258 5584 5264 5596
rect 5316 5584 5322 5636
rect 6638 5584 6644 5636
rect 6696 5624 6702 5636
rect 11606 5624 11612 5636
rect 6696 5596 11612 5624
rect 6696 5584 6702 5596
rect 11606 5584 11612 5596
rect 11664 5584 11670 5636
rect 2409 5559 2467 5565
rect 2409 5525 2421 5559
rect 2455 5556 2467 5559
rect 5994 5556 6000 5568
rect 2455 5528 6000 5556
rect 2455 5525 2467 5528
rect 2409 5519 2467 5525
rect 5994 5516 6000 5528
rect 6052 5516 6058 5568
rect 6362 5516 6368 5568
rect 6420 5556 6426 5568
rect 6733 5559 6791 5565
rect 6733 5556 6745 5559
rect 6420 5528 6745 5556
rect 6420 5516 6426 5528
rect 6733 5525 6745 5528
rect 6779 5525 6791 5559
rect 6733 5519 6791 5525
rect 7561 5559 7619 5565
rect 7561 5525 7573 5559
rect 7607 5556 7619 5559
rect 9582 5556 9588 5568
rect 7607 5528 9588 5556
rect 7607 5525 7619 5528
rect 7561 5519 7619 5525
rect 9582 5516 9588 5528
rect 9640 5516 9646 5568
rect 9950 5516 9956 5568
rect 10008 5556 10014 5568
rect 12894 5556 12900 5568
rect 10008 5528 12900 5556
rect 10008 5516 10014 5528
rect 12894 5516 12900 5528
rect 12952 5516 12958 5568
rect 13354 5556 13360 5568
rect 13315 5528 13360 5556
rect 13354 5516 13360 5528
rect 13412 5516 13418 5568
rect 15289 5559 15347 5565
rect 15289 5525 15301 5559
rect 15335 5556 15347 5559
rect 15470 5556 15476 5568
rect 15335 5528 15476 5556
rect 15335 5525 15347 5528
rect 15289 5519 15347 5525
rect 15470 5516 15476 5528
rect 15528 5516 15534 5568
rect 1104 5466 21896 5488
rect 1104 5414 4447 5466
rect 4499 5414 4511 5466
rect 4563 5414 4575 5466
rect 4627 5414 4639 5466
rect 4691 5414 11378 5466
rect 11430 5414 11442 5466
rect 11494 5414 11506 5466
rect 11558 5414 11570 5466
rect 11622 5414 18308 5466
rect 18360 5414 18372 5466
rect 18424 5414 18436 5466
rect 18488 5414 18500 5466
rect 18552 5414 21896 5466
rect 1104 5392 21896 5414
rect 9674 5352 9680 5364
rect 3344 5324 9680 5352
rect 1664 5151 1722 5157
rect 1664 5117 1676 5151
rect 1710 5148 1722 5151
rect 3344 5148 3372 5324
rect 9674 5312 9680 5324
rect 9732 5312 9738 5364
rect 9950 5352 9956 5364
rect 9784 5324 9956 5352
rect 3421 5287 3479 5293
rect 3421 5253 3433 5287
rect 3467 5284 3479 5287
rect 9784 5284 9812 5324
rect 9950 5312 9956 5324
rect 10008 5312 10014 5364
rect 14369 5355 14427 5361
rect 14369 5321 14381 5355
rect 14415 5352 14427 5355
rect 16390 5352 16396 5364
rect 14415 5324 16396 5352
rect 14415 5321 14427 5324
rect 14369 5315 14427 5321
rect 16390 5312 16396 5324
rect 16448 5312 16454 5364
rect 16850 5312 16856 5364
rect 16908 5352 16914 5364
rect 17310 5352 17316 5364
rect 16908 5324 17316 5352
rect 16908 5312 16914 5324
rect 17310 5312 17316 5324
rect 17368 5312 17374 5364
rect 20530 5312 20536 5364
rect 20588 5352 20594 5364
rect 20809 5355 20867 5361
rect 20809 5352 20821 5355
rect 20588 5324 20821 5352
rect 20588 5312 20594 5324
rect 20809 5321 20821 5324
rect 20855 5321 20867 5355
rect 20809 5315 20867 5321
rect 3467 5256 9812 5284
rect 9861 5287 9919 5293
rect 3467 5253 3479 5256
rect 3421 5247 3479 5253
rect 3786 5176 3792 5228
rect 3844 5216 3850 5228
rect 4356 5225 4384 5256
rect 9861 5253 9873 5287
rect 9907 5284 9919 5287
rect 10134 5284 10140 5296
rect 9907 5256 10140 5284
rect 9907 5253 9919 5256
rect 9861 5247 9919 5253
rect 10134 5244 10140 5256
rect 10192 5244 10198 5296
rect 12894 5244 12900 5296
rect 12952 5284 12958 5296
rect 12952 5256 16988 5284
rect 12952 5244 12958 5256
rect 16960 5228 16988 5256
rect 4157 5219 4215 5225
rect 4157 5216 4169 5219
rect 3844 5188 4169 5216
rect 3844 5176 3850 5188
rect 4157 5185 4169 5188
rect 4203 5185 4215 5219
rect 4157 5179 4215 5185
rect 4341 5219 4399 5225
rect 4341 5185 4353 5219
rect 4387 5185 4399 5219
rect 4341 5179 4399 5185
rect 5258 5176 5264 5228
rect 5316 5216 5322 5228
rect 5629 5219 5687 5225
rect 5629 5216 5641 5219
rect 5316 5188 5641 5216
rect 5316 5176 5322 5188
rect 5629 5185 5641 5188
rect 5675 5216 5687 5219
rect 6362 5216 6368 5228
rect 5675 5188 6368 5216
rect 5675 5185 5687 5188
rect 5629 5179 5687 5185
rect 6362 5176 6368 5188
rect 6420 5176 6426 5228
rect 6454 5176 6460 5228
rect 6512 5216 6518 5228
rect 6825 5219 6883 5225
rect 6825 5216 6837 5219
rect 6512 5188 6837 5216
rect 6512 5176 6518 5188
rect 6825 5185 6837 5188
rect 6871 5185 6883 5219
rect 6825 5179 6883 5185
rect 8849 5219 8907 5225
rect 8849 5185 8861 5219
rect 8895 5216 8907 5219
rect 9950 5216 9956 5228
rect 8895 5188 9956 5216
rect 8895 5185 8907 5188
rect 8849 5179 8907 5185
rect 9950 5176 9956 5188
rect 10008 5176 10014 5228
rect 10226 5176 10232 5228
rect 10284 5216 10290 5228
rect 10321 5219 10379 5225
rect 10321 5216 10333 5219
rect 10284 5188 10333 5216
rect 10284 5176 10290 5188
rect 10321 5185 10333 5188
rect 10367 5185 10379 5219
rect 10321 5179 10379 5185
rect 10505 5219 10563 5225
rect 10505 5185 10517 5219
rect 10551 5216 10563 5219
rect 10686 5216 10692 5228
rect 10551 5188 10692 5216
rect 10551 5185 10563 5188
rect 10505 5179 10563 5185
rect 1710 5120 3372 5148
rect 1710 5117 1722 5120
rect 1664 5111 1722 5117
rect 3878 5108 3884 5160
rect 3936 5148 3942 5160
rect 8021 5151 8079 5157
rect 3936 5120 5580 5148
rect 3936 5108 3942 5120
rect 3605 5083 3663 5089
rect 3605 5049 3617 5083
rect 3651 5080 3663 5083
rect 4062 5080 4068 5092
rect 3651 5052 4068 5080
rect 3651 5049 3663 5052
rect 3605 5043 3663 5049
rect 4062 5040 4068 5052
rect 4120 5040 4126 5092
rect 4798 5040 4804 5092
rect 4856 5080 4862 5092
rect 5258 5080 5264 5092
rect 4856 5052 5264 5080
rect 4856 5040 4862 5052
rect 5258 5040 5264 5052
rect 5316 5040 5322 5092
rect 5552 5089 5580 5120
rect 8021 5117 8033 5151
rect 8067 5148 8079 5151
rect 9490 5148 9496 5160
rect 8067 5120 9496 5148
rect 8067 5117 8079 5120
rect 8021 5111 8079 5117
rect 9490 5108 9496 5120
rect 9548 5108 9554 5160
rect 9582 5108 9588 5160
rect 9640 5148 9646 5160
rect 10134 5148 10140 5160
rect 9640 5120 10140 5148
rect 9640 5108 9646 5120
rect 10134 5108 10140 5120
rect 10192 5108 10198 5160
rect 5537 5083 5595 5089
rect 5537 5049 5549 5083
rect 5583 5080 5595 5083
rect 9858 5080 9864 5092
rect 5583 5052 9864 5080
rect 5583 5049 5595 5052
rect 5537 5043 5595 5049
rect 9858 5040 9864 5052
rect 9916 5040 9922 5092
rect 10336 5080 10364 5179
rect 10686 5176 10692 5188
rect 10744 5176 10750 5228
rect 11698 5176 11704 5228
rect 11756 5216 11762 5228
rect 12713 5219 12771 5225
rect 12713 5216 12725 5219
rect 11756 5188 12725 5216
rect 11756 5176 11762 5188
rect 12713 5185 12725 5188
rect 12759 5185 12771 5219
rect 15194 5216 15200 5228
rect 12713 5179 12771 5185
rect 14200 5188 15200 5216
rect 11146 5108 11152 5160
rect 11204 5148 11210 5160
rect 14200 5157 14228 5188
rect 15194 5176 15200 5188
rect 15252 5176 15258 5228
rect 16942 5216 16948 5228
rect 16855 5188 16948 5216
rect 16942 5176 16948 5188
rect 17000 5176 17006 5228
rect 18417 5219 18475 5225
rect 18417 5185 18429 5219
rect 18463 5216 18475 5219
rect 18966 5216 18972 5228
rect 18463 5188 18972 5216
rect 18463 5185 18475 5188
rect 18417 5179 18475 5185
rect 18966 5176 18972 5188
rect 19024 5176 19030 5228
rect 12529 5151 12587 5157
rect 12529 5148 12541 5151
rect 11204 5120 12541 5148
rect 11204 5108 11210 5120
rect 12529 5117 12541 5120
rect 12575 5117 12587 5151
rect 12529 5111 12587 5117
rect 14185 5151 14243 5157
rect 14185 5117 14197 5151
rect 14231 5117 14243 5151
rect 15286 5148 15292 5160
rect 15247 5120 15292 5148
rect 14185 5111 14243 5117
rect 15286 5108 15292 5120
rect 15344 5108 15350 5160
rect 15396 5120 16896 5148
rect 13630 5080 13636 5092
rect 10336 5052 13636 5080
rect 13630 5040 13636 5052
rect 13688 5040 13694 5092
rect 13906 5040 13912 5092
rect 13964 5080 13970 5092
rect 15396 5080 15424 5120
rect 13964 5052 15424 5080
rect 13964 5040 13970 5052
rect 16574 5040 16580 5092
rect 16632 5080 16638 5092
rect 16761 5083 16819 5089
rect 16761 5080 16773 5083
rect 16632 5052 16773 5080
rect 16632 5040 16638 5052
rect 16761 5049 16773 5052
rect 16807 5049 16819 5083
rect 16868 5080 16896 5120
rect 17034 5108 17040 5160
rect 17092 5148 17098 5160
rect 18138 5148 18144 5160
rect 17092 5120 18144 5148
rect 17092 5108 17098 5120
rect 18138 5108 18144 5120
rect 18196 5148 18202 5160
rect 19429 5151 19487 5157
rect 19429 5148 19441 5151
rect 18196 5120 19441 5148
rect 18196 5108 18202 5120
rect 19429 5117 19441 5120
rect 19475 5117 19487 5151
rect 19429 5111 19487 5117
rect 19696 5151 19754 5157
rect 19696 5117 19708 5151
rect 19742 5148 19754 5151
rect 20622 5148 20628 5160
rect 19742 5120 20628 5148
rect 19742 5117 19754 5120
rect 19696 5111 19754 5117
rect 20622 5108 20628 5120
rect 20680 5108 20686 5160
rect 16868 5052 19748 5080
rect 16761 5043 16819 5049
rect 19720 5024 19748 5052
rect 2777 5015 2835 5021
rect 2777 4981 2789 5015
rect 2823 5012 2835 5015
rect 3421 5015 3479 5021
rect 3421 5012 3433 5015
rect 2823 4984 3433 5012
rect 2823 4981 2835 4984
rect 2777 4975 2835 4981
rect 3421 4981 3433 4984
rect 3467 4981 3479 5015
rect 3694 5012 3700 5024
rect 3655 4984 3700 5012
rect 3421 4975 3479 4981
rect 3694 4972 3700 4984
rect 3752 4972 3758 5024
rect 4246 4972 4252 5024
rect 4304 5012 4310 5024
rect 5077 5015 5135 5021
rect 5077 5012 5089 5015
rect 4304 4984 5089 5012
rect 4304 4972 4310 4984
rect 5077 4981 5089 4984
rect 5123 4981 5135 5015
rect 5442 5012 5448 5024
rect 5403 4984 5448 5012
rect 5077 4975 5135 4981
rect 5442 4972 5448 4984
rect 5500 4972 5506 5024
rect 6914 4972 6920 5024
rect 6972 5012 6978 5024
rect 7374 5012 7380 5024
rect 6972 4984 7380 5012
rect 6972 4972 6978 4984
rect 7374 4972 7380 4984
rect 7432 5012 7438 5024
rect 9122 5012 9128 5024
rect 7432 4984 9128 5012
rect 7432 4972 7438 4984
rect 9122 4972 9128 4984
rect 9180 4972 9186 5024
rect 10229 5015 10287 5021
rect 10229 4981 10241 5015
rect 10275 5012 10287 5015
rect 10778 5012 10784 5024
rect 10275 4984 10784 5012
rect 10275 4981 10287 4984
rect 10229 4975 10287 4981
rect 10778 4972 10784 4984
rect 10836 4972 10842 5024
rect 15473 5015 15531 5021
rect 15473 4981 15485 5015
rect 15519 5012 15531 5015
rect 15930 5012 15936 5024
rect 15519 4984 15936 5012
rect 15519 4981 15531 4984
rect 15473 4975 15531 4981
rect 15930 4972 15936 4984
rect 15988 4972 15994 5024
rect 16393 5015 16451 5021
rect 16393 4981 16405 5015
rect 16439 5012 16451 5015
rect 16666 5012 16672 5024
rect 16439 4984 16672 5012
rect 16439 4981 16451 4984
rect 16393 4975 16451 4981
rect 16666 4972 16672 4984
rect 16724 4972 16730 5024
rect 16850 4972 16856 5024
rect 16908 5012 16914 5024
rect 16908 4984 16953 5012
rect 16908 4972 16914 4984
rect 19702 4972 19708 5024
rect 19760 4972 19766 5024
rect 1104 4922 21896 4944
rect 1104 4870 7912 4922
rect 7964 4870 7976 4922
rect 8028 4870 8040 4922
rect 8092 4870 8104 4922
rect 8156 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 15035 4922
rect 15087 4870 21896 4922
rect 1104 4848 21896 4870
rect 2682 4768 2688 4820
rect 2740 4808 2746 4820
rect 2777 4811 2835 4817
rect 2777 4808 2789 4811
rect 2740 4780 2789 4808
rect 2740 4768 2746 4780
rect 2777 4777 2789 4780
rect 2823 4777 2835 4811
rect 2777 4771 2835 4777
rect 2869 4811 2927 4817
rect 2869 4777 2881 4811
rect 2915 4808 2927 4811
rect 4525 4811 4583 4817
rect 4525 4808 4537 4811
rect 2915 4780 4537 4808
rect 2915 4777 2927 4780
rect 2869 4771 2927 4777
rect 4525 4777 4537 4780
rect 4571 4777 4583 4811
rect 4890 4808 4896 4820
rect 4851 4780 4896 4808
rect 4525 4771 4583 4777
rect 4890 4768 4896 4780
rect 4948 4768 4954 4820
rect 5442 4768 5448 4820
rect 5500 4808 5506 4820
rect 5721 4811 5779 4817
rect 5721 4808 5733 4811
rect 5500 4780 5733 4808
rect 5500 4768 5506 4780
rect 5721 4777 5733 4780
rect 5767 4777 5779 4811
rect 5721 4771 5779 4777
rect 7098 4768 7104 4820
rect 7156 4808 7162 4820
rect 13262 4808 13268 4820
rect 7156 4780 13268 4808
rect 7156 4768 7162 4780
rect 13262 4768 13268 4780
rect 13320 4768 13326 4820
rect 14093 4811 14151 4817
rect 14093 4777 14105 4811
rect 14139 4808 14151 4811
rect 14274 4808 14280 4820
rect 14139 4780 14280 4808
rect 14139 4777 14151 4780
rect 14093 4771 14151 4777
rect 14274 4768 14280 4780
rect 14332 4768 14338 4820
rect 16025 4811 16083 4817
rect 16025 4777 16037 4811
rect 16071 4808 16083 4811
rect 16850 4808 16856 4820
rect 16071 4780 16856 4808
rect 16071 4777 16083 4780
rect 16025 4771 16083 4777
rect 16850 4768 16856 4780
rect 16908 4768 16914 4820
rect 19610 4808 19616 4820
rect 19571 4780 19616 4808
rect 19610 4768 19616 4780
rect 19668 4808 19674 4820
rect 19797 4811 19855 4817
rect 19797 4808 19809 4811
rect 19668 4780 19809 4808
rect 19668 4768 19674 4780
rect 19797 4777 19809 4780
rect 19843 4777 19855 4811
rect 19797 4771 19855 4777
rect 198 4700 204 4752
rect 256 4740 262 4752
rect 3234 4740 3240 4752
rect 256 4712 3240 4740
rect 256 4700 262 4712
rect 3234 4700 3240 4712
rect 3292 4700 3298 4752
rect 3329 4743 3387 4749
rect 3329 4709 3341 4743
rect 3375 4709 3387 4743
rect 3329 4703 3387 4709
rect 1664 4675 1722 4681
rect 1664 4641 1676 4675
rect 1710 4672 1722 4675
rect 2590 4672 2596 4684
rect 1710 4644 2596 4672
rect 1710 4641 1722 4644
rect 1664 4635 1722 4641
rect 2590 4632 2596 4644
rect 2648 4632 2654 4684
rect 3344 4672 3372 4703
rect 3786 4700 3792 4752
rect 3844 4740 3850 4752
rect 5810 4740 5816 4752
rect 3844 4712 5816 4740
rect 3844 4700 3850 4712
rect 5810 4700 5816 4712
rect 5868 4700 5874 4752
rect 7558 4700 7564 4752
rect 7616 4740 7622 4752
rect 12980 4743 13038 4749
rect 7616 4712 11560 4740
rect 7616 4700 7622 4712
rect 4062 4672 4068 4684
rect 3344 4644 4068 4672
rect 4062 4632 4068 4644
rect 4120 4632 4126 4684
rect 4154 4632 4160 4684
rect 4212 4672 4218 4684
rect 4433 4675 4491 4681
rect 4433 4672 4445 4675
rect 4212 4644 4445 4672
rect 4212 4632 4218 4644
rect 4433 4641 4445 4644
rect 4479 4641 4491 4675
rect 5261 4675 5319 4681
rect 5261 4672 5273 4675
rect 4433 4635 4491 4641
rect 4540 4644 5273 4672
rect 2958 4564 2964 4616
rect 3016 4604 3022 4616
rect 3421 4607 3479 4613
rect 3421 4604 3433 4607
rect 3016 4576 3433 4604
rect 3016 4564 3022 4576
rect 3421 4573 3433 4576
rect 3467 4573 3479 4607
rect 3421 4567 3479 4573
rect 3786 4564 3792 4616
rect 3844 4604 3850 4616
rect 4540 4604 4568 4644
rect 5261 4641 5273 4644
rect 5307 4672 5319 4675
rect 6914 4672 6920 4684
rect 5307 4644 6920 4672
rect 5307 4641 5319 4644
rect 5261 4635 5319 4641
rect 6914 4632 6920 4644
rect 6972 4632 6978 4684
rect 7374 4672 7380 4684
rect 7335 4644 7380 4672
rect 7374 4632 7380 4644
rect 7432 4632 7438 4684
rect 7644 4675 7702 4681
rect 7644 4641 7656 4675
rect 7690 4672 7702 4675
rect 9950 4672 9956 4684
rect 7690 4644 9956 4672
rect 7690 4641 7702 4644
rect 7644 4635 7702 4641
rect 9950 4632 9956 4644
rect 10008 4632 10014 4684
rect 10045 4675 10103 4681
rect 10045 4641 10057 4675
rect 10091 4672 10103 4675
rect 10091 4644 11284 4672
rect 10091 4641 10103 4644
rect 10045 4635 10103 4641
rect 3844 4576 4568 4604
rect 4709 4607 4767 4613
rect 3844 4564 3850 4576
rect 4709 4573 4721 4607
rect 4755 4604 4767 4607
rect 4798 4604 4804 4616
rect 4755 4576 4804 4604
rect 4755 4573 4767 4576
rect 4709 4567 4767 4573
rect 4798 4564 4804 4576
rect 4856 4564 4862 4616
rect 5350 4604 5356 4616
rect 5311 4576 5356 4604
rect 5350 4564 5356 4576
rect 5408 4564 5414 4616
rect 5445 4607 5503 4613
rect 5445 4573 5457 4607
rect 5491 4573 5503 4607
rect 9674 4604 9680 4616
rect 5445 4567 5503 4573
rect 8404 4576 9680 4604
rect 2866 4496 2872 4548
rect 2924 4536 2930 4548
rect 4065 4539 4123 4545
rect 4065 4536 4077 4539
rect 2924 4508 4077 4536
rect 2924 4496 2930 4508
rect 4065 4505 4077 4508
rect 4111 4505 4123 4539
rect 4065 4499 4123 4505
rect 5166 4496 5172 4548
rect 5224 4536 5230 4548
rect 5460 4536 5488 4567
rect 5224 4508 5488 4536
rect 5224 4496 5230 4508
rect 3142 4428 3148 4480
rect 3200 4468 3206 4480
rect 3881 4471 3939 4477
rect 3881 4468 3893 4471
rect 3200 4440 3893 4468
rect 3200 4428 3206 4440
rect 3881 4437 3893 4440
rect 3927 4437 3939 4471
rect 3881 4431 3939 4437
rect 3970 4428 3976 4480
rect 4028 4468 4034 4480
rect 8404 4468 8432 4576
rect 9674 4564 9680 4576
rect 9732 4564 9738 4616
rect 10134 4604 10140 4616
rect 10095 4576 10140 4604
rect 10134 4564 10140 4576
rect 10192 4564 10198 4616
rect 10229 4607 10287 4613
rect 10229 4573 10241 4607
rect 10275 4573 10287 4607
rect 10229 4567 10287 4573
rect 8757 4539 8815 4545
rect 8757 4505 8769 4539
rect 8803 4536 8815 4539
rect 9582 4536 9588 4548
rect 8803 4508 9588 4536
rect 8803 4505 8815 4508
rect 8757 4499 8815 4505
rect 9582 4496 9588 4508
rect 9640 4536 9646 4548
rect 10244 4536 10272 4567
rect 9640 4508 10272 4536
rect 9640 4496 9646 4508
rect 4028 4440 8432 4468
rect 9677 4471 9735 4477
rect 4028 4428 4034 4440
rect 9677 4437 9689 4471
rect 9723 4468 9735 4471
rect 10594 4468 10600 4480
rect 9723 4440 10600 4468
rect 9723 4437 9735 4440
rect 9677 4431 9735 4437
rect 10594 4428 10600 4440
rect 10652 4428 10658 4480
rect 11256 4468 11284 4644
rect 11330 4632 11336 4684
rect 11388 4672 11394 4684
rect 11425 4675 11483 4681
rect 11425 4672 11437 4675
rect 11388 4644 11437 4672
rect 11388 4632 11394 4644
rect 11425 4641 11437 4644
rect 11471 4641 11483 4675
rect 11425 4635 11483 4641
rect 11532 4536 11560 4712
rect 12980 4709 12992 4743
rect 13026 4740 13038 4743
rect 13354 4740 13360 4752
rect 13026 4712 13360 4740
rect 13026 4709 13038 4712
rect 12980 4703 13038 4709
rect 13354 4700 13360 4712
rect 13412 4700 13418 4752
rect 16040 4712 16528 4740
rect 16040 4684 16068 4712
rect 11974 4632 11980 4684
rect 12032 4672 12038 4684
rect 12713 4675 12771 4681
rect 12713 4672 12725 4675
rect 12032 4644 12725 4672
rect 12032 4632 12038 4644
rect 12713 4641 12725 4644
rect 12759 4641 12771 4675
rect 12713 4635 12771 4641
rect 12802 4632 12808 4684
rect 12860 4632 12866 4684
rect 16022 4632 16028 4684
rect 16080 4632 16086 4684
rect 16500 4681 16528 4712
rect 16942 4700 16948 4752
rect 17000 4740 17006 4752
rect 17834 4743 17892 4749
rect 17834 4740 17846 4743
rect 17000 4712 17846 4740
rect 17000 4700 17006 4712
rect 17834 4709 17846 4712
rect 17880 4709 17892 4743
rect 17834 4703 17892 4709
rect 16393 4675 16451 4681
rect 16393 4641 16405 4675
rect 16439 4641 16451 4675
rect 16393 4635 16451 4641
rect 16485 4675 16543 4681
rect 16485 4641 16497 4675
rect 16531 4672 16543 4675
rect 18782 4672 18788 4684
rect 16531 4644 18788 4672
rect 16531 4641 16543 4644
rect 16485 4635 16543 4641
rect 11701 4607 11759 4613
rect 11701 4573 11713 4607
rect 11747 4604 11759 4607
rect 12526 4604 12532 4616
rect 11747 4576 12532 4604
rect 11747 4573 11759 4576
rect 11701 4567 11759 4573
rect 12526 4564 12532 4576
rect 12584 4564 12590 4616
rect 12820 4604 12848 4632
rect 12728 4576 12848 4604
rect 12728 4536 12756 4576
rect 11532 4508 12756 4536
rect 12986 4468 12992 4480
rect 11256 4440 12992 4468
rect 12986 4428 12992 4440
rect 13044 4428 13050 4480
rect 13630 4428 13636 4480
rect 13688 4468 13694 4480
rect 15746 4468 15752 4480
rect 13688 4440 15752 4468
rect 13688 4428 13694 4440
rect 15746 4428 15752 4440
rect 15804 4428 15810 4480
rect 16408 4468 16436 4635
rect 18782 4632 18788 4644
rect 18840 4632 18846 4684
rect 16669 4607 16727 4613
rect 16669 4573 16681 4607
rect 16715 4573 16727 4607
rect 16669 4567 16727 4573
rect 16684 4536 16712 4567
rect 17034 4564 17040 4616
rect 17092 4604 17098 4616
rect 17589 4607 17647 4613
rect 17589 4604 17601 4607
rect 17092 4576 17601 4604
rect 17092 4564 17098 4576
rect 17589 4573 17601 4576
rect 17635 4573 17647 4607
rect 17589 4567 17647 4573
rect 17126 4536 17132 4548
rect 16684 4508 17132 4536
rect 17126 4496 17132 4508
rect 17184 4496 17190 4548
rect 17770 4468 17776 4480
rect 16408 4440 17776 4468
rect 17770 4428 17776 4440
rect 17828 4428 17834 4480
rect 18966 4468 18972 4480
rect 18927 4440 18972 4468
rect 18966 4428 18972 4440
rect 19024 4428 19030 4480
rect 1104 4378 21896 4400
rect 1104 4326 4447 4378
rect 4499 4326 4511 4378
rect 4563 4326 4575 4378
rect 4627 4326 4639 4378
rect 4691 4326 11378 4378
rect 11430 4326 11442 4378
rect 11494 4326 11506 4378
rect 11558 4326 11570 4378
rect 11622 4326 18308 4378
rect 18360 4326 18372 4378
rect 18424 4326 18436 4378
rect 18488 4326 18500 4378
rect 18552 4326 21896 4378
rect 1104 4304 21896 4326
rect 3142 4224 3148 4276
rect 3200 4264 3206 4276
rect 4062 4264 4068 4276
rect 3200 4236 4068 4264
rect 3200 4224 3206 4236
rect 4062 4224 4068 4236
rect 4120 4224 4126 4276
rect 4798 4264 4804 4276
rect 4264 4236 4804 4264
rect 2869 4199 2927 4205
rect 2869 4165 2881 4199
rect 2915 4165 2927 4199
rect 4264 4196 4292 4236
rect 4798 4224 4804 4236
rect 4856 4224 4862 4276
rect 9490 4224 9496 4276
rect 9548 4264 9554 4276
rect 13906 4264 13912 4276
rect 9548 4236 13912 4264
rect 9548 4224 9554 4236
rect 13906 4224 13912 4236
rect 13964 4224 13970 4276
rect 17126 4264 17132 4276
rect 14016 4236 17132 4264
rect 2869 4159 2927 4165
rect 4080 4168 4292 4196
rect 4341 4199 4399 4205
rect 2884 4128 2912 4159
rect 2884 4100 3096 4128
rect 1489 4063 1547 4069
rect 1489 4029 1501 4063
rect 1535 4060 1547 4063
rect 1578 4060 1584 4072
rect 1535 4032 1584 4060
rect 1535 4029 1547 4032
rect 1489 4023 1547 4029
rect 1578 4020 1584 4032
rect 1636 4060 1642 4072
rect 2774 4060 2780 4072
rect 1636 4032 2780 4060
rect 1636 4020 1642 4032
rect 2774 4020 2780 4032
rect 2832 4060 2838 4072
rect 2961 4063 3019 4069
rect 2961 4060 2973 4063
rect 2832 4032 2973 4060
rect 2832 4020 2838 4032
rect 2961 4029 2973 4032
rect 3007 4029 3019 4063
rect 3068 4060 3096 4100
rect 4080 4060 4108 4168
rect 4341 4165 4353 4199
rect 4387 4165 4399 4199
rect 4341 4159 4399 4165
rect 4356 4128 4384 4159
rect 9582 4156 9588 4208
rect 9640 4196 9646 4208
rect 9640 4168 11008 4196
rect 9640 4156 9646 4168
rect 5721 4131 5779 4137
rect 5721 4128 5733 4131
rect 4264 4100 5733 4128
rect 4264 4060 4292 4100
rect 5721 4097 5733 4100
rect 5767 4097 5779 4131
rect 6086 4128 6092 4140
rect 5721 4091 5779 4097
rect 5828 4100 6092 4128
rect 4430 4060 4436 4072
rect 3068 4032 4108 4060
rect 4172 4032 4292 4060
rect 4391 4032 4436 4060
rect 2961 4023 3019 4029
rect 1756 3995 1814 4001
rect 1756 3961 1768 3995
rect 1802 3992 1814 3995
rect 2866 3992 2872 4004
rect 1802 3964 2872 3992
rect 1802 3961 1814 3964
rect 1756 3955 1814 3961
rect 2866 3952 2872 3964
rect 2924 3952 2930 4004
rect 3228 3995 3286 4001
rect 3228 3961 3240 3995
rect 3274 3992 3286 3995
rect 3326 3992 3332 4004
rect 3274 3964 3332 3992
rect 3274 3961 3286 3964
rect 3228 3955 3286 3961
rect 3326 3952 3332 3964
rect 3384 3952 3390 4004
rect 3602 3884 3608 3936
rect 3660 3924 3666 3936
rect 4172 3924 4200 4032
rect 4430 4020 4436 4032
rect 4488 4020 4494 4072
rect 4890 4020 4896 4072
rect 4948 4060 4954 4072
rect 5828 4060 5856 4100
rect 6086 4088 6092 4100
rect 6144 4088 6150 4140
rect 6822 4088 6828 4140
rect 6880 4128 6886 4140
rect 10502 4128 10508 4140
rect 6880 4100 10508 4128
rect 6880 4088 6886 4100
rect 10502 4088 10508 4100
rect 10560 4128 10566 4140
rect 10778 4128 10784 4140
rect 10560 4100 10784 4128
rect 10560 4088 10566 4100
rect 10778 4088 10784 4100
rect 10836 4088 10842 4140
rect 10870 4088 10876 4140
rect 10928 4088 10934 4140
rect 10980 4128 11008 4168
rect 11054 4156 11060 4208
rect 11112 4196 11118 4208
rect 12618 4196 12624 4208
rect 11112 4168 12624 4196
rect 11112 4156 11118 4168
rect 12618 4156 12624 4168
rect 12676 4196 12682 4208
rect 14016 4196 14044 4236
rect 17126 4224 17132 4236
rect 17184 4224 17190 4276
rect 14274 4196 14280 4208
rect 12676 4168 14044 4196
rect 14108 4168 14280 4196
rect 12676 4156 12682 4168
rect 11149 4131 11207 4137
rect 11149 4128 11161 4131
rect 10980 4100 11161 4128
rect 11149 4097 11161 4100
rect 11195 4097 11207 4131
rect 11149 4091 11207 4097
rect 12802 4088 12808 4140
rect 12860 4128 12866 4140
rect 14108 4137 14136 4168
rect 14274 4156 14280 4168
rect 14332 4156 14338 4208
rect 18509 4199 18567 4205
rect 18509 4196 18521 4199
rect 14936 4168 18521 4196
rect 13909 4131 13967 4137
rect 13909 4128 13921 4131
rect 12860 4100 13921 4128
rect 12860 4088 12866 4100
rect 13909 4097 13921 4100
rect 13955 4097 13967 4131
rect 13909 4091 13967 4097
rect 14093 4131 14151 4137
rect 14093 4097 14105 4131
rect 14139 4097 14151 4131
rect 14093 4091 14151 4097
rect 4948 4032 5856 4060
rect 4948 4020 4954 4032
rect 5994 4020 6000 4072
rect 6052 4060 6058 4072
rect 7469 4063 7527 4069
rect 7469 4060 7481 4063
rect 6052 4032 7481 4060
rect 6052 4020 6058 4032
rect 7469 4029 7481 4032
rect 7515 4029 7527 4063
rect 7469 4023 7527 4029
rect 9493 4063 9551 4069
rect 9493 4029 9505 4063
rect 9539 4060 9551 4063
rect 10888 4060 10916 4088
rect 9539 4032 10916 4060
rect 10965 4063 11023 4069
rect 9539 4029 9551 4032
rect 9493 4023 9551 4029
rect 10965 4029 10977 4063
rect 11011 4060 11023 4063
rect 11011 4032 12480 4060
rect 11011 4029 11023 4032
rect 10965 4023 11023 4029
rect 4338 3952 4344 4004
rect 4396 3992 4402 4004
rect 4709 3995 4767 4001
rect 4709 3992 4721 3995
rect 4396 3964 4721 3992
rect 4396 3952 4402 3964
rect 4709 3961 4721 3964
rect 4755 3961 4767 3995
rect 4709 3955 4767 3961
rect 5537 3995 5595 4001
rect 5537 3961 5549 3995
rect 5583 3992 5595 3995
rect 6638 3992 6644 4004
rect 5583 3964 6644 3992
rect 5583 3961 5595 3964
rect 5537 3955 5595 3961
rect 6638 3952 6644 3964
rect 6696 3952 6702 4004
rect 7745 3995 7803 4001
rect 7745 3961 7757 3995
rect 7791 3992 7803 3995
rect 8570 3992 8576 4004
rect 7791 3964 8576 3992
rect 7791 3961 7803 3964
rect 7745 3955 7803 3961
rect 8570 3952 8576 3964
rect 8628 3952 8634 4004
rect 8662 3952 8668 4004
rect 8720 3992 8726 4004
rect 12342 3992 12348 4004
rect 8720 3964 12348 3992
rect 8720 3952 8726 3964
rect 12342 3952 12348 3964
rect 12400 3952 12406 4004
rect 12452 3992 12480 4032
rect 12526 4020 12532 4072
rect 12584 4060 12590 4072
rect 13538 4060 13544 4072
rect 12584 4032 13544 4060
rect 12584 4020 12590 4032
rect 13538 4020 13544 4032
rect 13596 4020 13602 4072
rect 13722 4020 13728 4072
rect 13780 4060 13786 4072
rect 14936 4060 14964 4168
rect 18509 4165 18521 4168
rect 18555 4165 18567 4199
rect 18509 4159 18567 4165
rect 15194 4128 15200 4140
rect 15155 4100 15200 4128
rect 15194 4088 15200 4100
rect 15252 4088 15258 4140
rect 16298 4088 16304 4140
rect 16356 4128 16362 4140
rect 17862 4128 17868 4140
rect 16356 4100 17868 4128
rect 16356 4088 16362 4100
rect 17862 4088 17868 4100
rect 17920 4088 17926 4140
rect 18966 4088 18972 4140
rect 19024 4128 19030 4140
rect 19061 4131 19119 4137
rect 19061 4128 19073 4131
rect 19024 4100 19073 4128
rect 19024 4088 19030 4100
rect 19061 4097 19073 4100
rect 19107 4097 19119 4131
rect 19061 4091 19119 4097
rect 13780 4032 14964 4060
rect 15013 4063 15071 4069
rect 13780 4020 13786 4032
rect 15013 4029 15025 4063
rect 15059 4029 15071 4063
rect 15013 4023 15071 4029
rect 13170 3992 13176 4004
rect 12452 3964 13176 3992
rect 13170 3952 13176 3964
rect 13228 3952 13234 4004
rect 15028 3992 15056 4023
rect 17954 4020 17960 4072
rect 18012 4060 18018 4072
rect 18877 4063 18935 4069
rect 18877 4060 18889 4063
rect 18012 4032 18889 4060
rect 18012 4020 18018 4032
rect 18877 4029 18889 4032
rect 18923 4029 18935 4063
rect 20530 4060 20536 4072
rect 20491 4032 20536 4060
rect 18877 4023 18935 4029
rect 20530 4020 20536 4032
rect 20588 4020 20594 4072
rect 13464 3964 15056 3992
rect 5166 3924 5172 3936
rect 3660 3896 4200 3924
rect 5127 3896 5172 3924
rect 3660 3884 3666 3896
rect 5166 3884 5172 3896
rect 5224 3884 5230 3936
rect 5629 3927 5687 3933
rect 5629 3893 5641 3927
rect 5675 3924 5687 3927
rect 6914 3924 6920 3936
rect 5675 3896 6920 3924
rect 5675 3893 5687 3896
rect 5629 3887 5687 3893
rect 6914 3884 6920 3896
rect 6972 3884 6978 3936
rect 9677 3927 9735 3933
rect 9677 3893 9689 3927
rect 9723 3924 9735 3927
rect 10226 3924 10232 3936
rect 9723 3896 10232 3924
rect 9723 3893 9735 3896
rect 9677 3887 9735 3893
rect 10226 3884 10232 3896
rect 10284 3884 10290 3936
rect 10502 3884 10508 3936
rect 10560 3924 10566 3936
rect 10597 3927 10655 3933
rect 10597 3924 10609 3927
rect 10560 3896 10609 3924
rect 10560 3884 10566 3896
rect 10597 3893 10609 3896
rect 10643 3893 10655 3927
rect 11054 3924 11060 3936
rect 11015 3896 11060 3924
rect 10597 3887 10655 3893
rect 11054 3884 11060 3896
rect 11112 3884 11118 3936
rect 11146 3884 11152 3936
rect 11204 3924 11210 3936
rect 11790 3924 11796 3936
rect 11204 3896 11796 3924
rect 11204 3884 11210 3896
rect 11790 3884 11796 3896
rect 11848 3884 11854 3936
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 13464 3933 13492 3964
rect 15194 3952 15200 4004
rect 15252 3992 15258 4004
rect 15562 3992 15568 4004
rect 15252 3964 15568 3992
rect 15252 3952 15258 3964
rect 15562 3952 15568 3964
rect 15620 3952 15626 4004
rect 16666 3952 16672 4004
rect 16724 3992 16730 4004
rect 18969 3995 19027 4001
rect 18969 3992 18981 3995
rect 16724 3964 18981 3992
rect 16724 3952 16730 3964
rect 18969 3961 18981 3964
rect 19015 3961 19027 3995
rect 18969 3955 19027 3961
rect 13449 3927 13507 3933
rect 12492 3896 12537 3924
rect 12492 3884 12498 3896
rect 13449 3893 13461 3927
rect 13495 3893 13507 3927
rect 13449 3887 13507 3893
rect 13722 3884 13728 3936
rect 13780 3924 13786 3936
rect 13817 3927 13875 3933
rect 13817 3924 13829 3927
rect 13780 3896 13829 3924
rect 13780 3884 13786 3896
rect 13817 3893 13829 3896
rect 13863 3893 13875 3927
rect 13817 3887 13875 3893
rect 14090 3884 14096 3936
rect 14148 3924 14154 3936
rect 16022 3924 16028 3936
rect 14148 3896 16028 3924
rect 14148 3884 14154 3896
rect 16022 3884 16028 3896
rect 16080 3884 16086 3936
rect 16298 3924 16304 3936
rect 16259 3896 16304 3924
rect 16298 3884 16304 3896
rect 16356 3884 16362 3936
rect 20717 3927 20775 3933
rect 20717 3893 20729 3927
rect 20763 3924 20775 3927
rect 21726 3924 21732 3936
rect 20763 3896 21732 3924
rect 20763 3893 20775 3896
rect 20717 3887 20775 3893
rect 21726 3884 21732 3896
rect 21784 3884 21790 3936
rect 1104 3834 21896 3856
rect 1104 3782 7912 3834
rect 7964 3782 7976 3834
rect 8028 3782 8040 3834
rect 8092 3782 8104 3834
rect 8156 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 15035 3834
rect 15087 3782 21896 3834
rect 1104 3760 21896 3782
rect 2958 3720 2964 3732
rect 2919 3692 2964 3720
rect 2958 3680 2964 3692
rect 3016 3680 3022 3732
rect 3053 3723 3111 3729
rect 3053 3689 3065 3723
rect 3099 3720 3111 3723
rect 4154 3720 4160 3732
rect 3099 3692 4160 3720
rect 3099 3689 3111 3692
rect 3053 3683 3111 3689
rect 4154 3680 4160 3692
rect 4212 3680 4218 3732
rect 4338 3680 4344 3732
rect 4396 3720 4402 3732
rect 4982 3720 4988 3732
rect 4396 3692 4988 3720
rect 4396 3680 4402 3692
rect 4982 3680 4988 3692
rect 5040 3680 5046 3732
rect 5166 3680 5172 3732
rect 5224 3720 5230 3732
rect 5997 3723 6055 3729
rect 5997 3720 6009 3723
rect 5224 3692 6009 3720
rect 5224 3680 5230 3692
rect 5997 3689 6009 3692
rect 6043 3689 6055 3723
rect 6638 3720 6644 3732
rect 6599 3692 6644 3720
rect 5997 3683 6055 3689
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 7006 3720 7012 3732
rect 6919 3692 7012 3720
rect 7006 3680 7012 3692
rect 7064 3720 7070 3732
rect 8202 3720 8208 3732
rect 7064 3692 8208 3720
rect 7064 3680 7070 3692
rect 8202 3680 8208 3692
rect 8260 3680 8266 3732
rect 8573 3723 8631 3729
rect 8573 3689 8585 3723
rect 8619 3720 8631 3723
rect 9858 3720 9864 3732
rect 8619 3692 9864 3720
rect 8619 3689 8631 3692
rect 8573 3683 8631 3689
rect 9858 3680 9864 3692
rect 9916 3680 9922 3732
rect 10428 3692 10732 3720
rect 1848 3655 1906 3661
rect 1848 3621 1860 3655
rect 1894 3652 1906 3655
rect 5074 3652 5080 3664
rect 1894 3624 5080 3652
rect 1894 3621 1906 3624
rect 1848 3615 1906 3621
rect 5074 3612 5080 3624
rect 5132 3612 5138 3664
rect 5350 3612 5356 3664
rect 5408 3652 5414 3664
rect 7098 3652 7104 3664
rect 5408 3624 7104 3652
rect 5408 3612 5414 3624
rect 7098 3612 7104 3624
rect 7156 3612 7162 3664
rect 9398 3612 9404 3664
rect 9456 3652 9462 3664
rect 10428 3652 10456 3692
rect 10594 3652 10600 3664
rect 9456 3624 10456 3652
rect 10555 3624 10600 3652
rect 9456 3612 9462 3624
rect 10594 3612 10600 3624
rect 10652 3612 10658 3664
rect 10704 3652 10732 3692
rect 10778 3680 10784 3732
rect 10836 3720 10842 3732
rect 12253 3723 12311 3729
rect 12253 3720 12265 3723
rect 10836 3692 12265 3720
rect 10836 3680 10842 3692
rect 12253 3689 12265 3692
rect 12299 3689 12311 3723
rect 12253 3683 12311 3689
rect 13170 3680 13176 3732
rect 13228 3720 13234 3732
rect 13446 3720 13452 3732
rect 13228 3692 13452 3720
rect 13228 3680 13234 3692
rect 13446 3680 13452 3692
rect 13504 3680 13510 3732
rect 13541 3723 13599 3729
rect 13541 3689 13553 3723
rect 13587 3720 13599 3723
rect 13722 3720 13728 3732
rect 13587 3692 13728 3720
rect 13587 3689 13599 3692
rect 13541 3683 13599 3689
rect 13722 3680 13728 3692
rect 13780 3680 13786 3732
rect 13909 3723 13967 3729
rect 13909 3689 13921 3723
rect 13955 3720 13967 3723
rect 16298 3720 16304 3732
rect 13955 3692 16304 3720
rect 13955 3689 13967 3692
rect 13909 3683 13967 3689
rect 16298 3680 16304 3692
rect 16356 3680 16362 3732
rect 13998 3652 14004 3664
rect 10704 3624 13308 3652
rect 13959 3624 14004 3652
rect 1578 3584 1584 3596
rect 1539 3556 1584 3584
rect 1578 3544 1584 3556
rect 1636 3544 1642 3596
rect 3142 3544 3148 3596
rect 3200 3584 3206 3596
rect 3421 3587 3479 3593
rect 3421 3584 3433 3587
rect 3200 3556 3433 3584
rect 3200 3544 3206 3556
rect 3421 3553 3433 3556
rect 3467 3553 3479 3587
rect 3421 3547 3479 3553
rect 3513 3587 3571 3593
rect 3513 3553 3525 3587
rect 3559 3584 3571 3587
rect 4332 3587 4390 3593
rect 3559 3556 4108 3584
rect 3559 3553 3571 3556
rect 3513 3547 3571 3553
rect 3605 3519 3663 3525
rect 3605 3485 3617 3519
rect 3651 3485 3663 3519
rect 3605 3479 3663 3485
rect 2958 3408 2964 3460
rect 3016 3448 3022 3460
rect 3620 3448 3648 3479
rect 3016 3420 3648 3448
rect 3016 3408 3022 3420
rect 1118 3340 1124 3392
rect 1176 3380 1182 3392
rect 4080 3380 4108 3556
rect 4332 3553 4344 3587
rect 4378 3584 4390 3587
rect 5626 3584 5632 3596
rect 4378 3556 5632 3584
rect 4378 3553 4390 3556
rect 4332 3547 4390 3553
rect 5626 3544 5632 3556
rect 5684 3544 5690 3596
rect 5902 3584 5908 3596
rect 5863 3556 5908 3584
rect 5902 3544 5908 3556
rect 5960 3544 5966 3596
rect 5994 3544 6000 3596
rect 6052 3584 6058 3596
rect 9306 3584 9312 3596
rect 6052 3556 9312 3584
rect 6052 3544 6058 3556
rect 9306 3544 9312 3556
rect 9364 3544 9370 3596
rect 10502 3544 10508 3596
rect 10560 3584 10566 3596
rect 10689 3587 10747 3593
rect 10689 3584 10701 3587
rect 10560 3556 10701 3584
rect 10560 3544 10566 3556
rect 10689 3553 10701 3556
rect 10735 3553 10747 3587
rect 12161 3587 12219 3593
rect 12161 3584 12173 3587
rect 10689 3547 10747 3553
rect 10796 3556 12173 3584
rect 5074 3476 5080 3528
rect 5132 3516 5138 3528
rect 6089 3519 6147 3525
rect 6089 3516 6101 3519
rect 5132 3488 6101 3516
rect 5132 3476 5138 3488
rect 6089 3485 6101 3488
rect 6135 3485 6147 3519
rect 6089 3479 6147 3485
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 7193 3519 7251 3525
rect 7193 3516 7205 3519
rect 6512 3488 7205 3516
rect 6512 3476 6518 3488
rect 7193 3485 7205 3488
rect 7239 3485 7251 3519
rect 7193 3479 7251 3485
rect 10318 3476 10324 3528
rect 10376 3516 10382 3528
rect 10796 3516 10824 3556
rect 12161 3553 12173 3556
rect 12207 3553 12219 3587
rect 12161 3547 12219 3553
rect 10376 3488 10824 3516
rect 10376 3476 10382 3488
rect 10870 3476 10876 3528
rect 10928 3516 10934 3528
rect 12437 3519 12495 3525
rect 10928 3488 10973 3516
rect 10928 3476 10934 3488
rect 12437 3485 12449 3519
rect 12483 3516 12495 3519
rect 12618 3516 12624 3528
rect 12483 3488 12624 3516
rect 12483 3485 12495 3488
rect 12437 3479 12495 3485
rect 12618 3476 12624 3488
rect 12676 3476 12682 3528
rect 13280 3516 13308 3624
rect 13998 3612 14004 3624
rect 14056 3612 14062 3664
rect 16574 3652 16580 3664
rect 14660 3624 16580 3652
rect 13354 3544 13360 3596
rect 13412 3584 13418 3596
rect 13412 3556 14136 3584
rect 13412 3544 13418 3556
rect 13998 3516 14004 3528
rect 13280 3488 14004 3516
rect 13998 3476 14004 3488
rect 14056 3476 14062 3528
rect 14108 3525 14136 3556
rect 14093 3519 14151 3525
rect 14093 3485 14105 3519
rect 14139 3485 14151 3519
rect 14093 3479 14151 3485
rect 5000 3420 6684 3448
rect 5000 3380 5028 3420
rect 5442 3380 5448 3392
rect 1176 3352 5028 3380
rect 5403 3352 5448 3380
rect 1176 3340 1182 3352
rect 5442 3340 5448 3352
rect 5500 3340 5506 3392
rect 5537 3383 5595 3389
rect 5537 3349 5549 3383
rect 5583 3380 5595 3383
rect 6546 3380 6552 3392
rect 5583 3352 6552 3380
rect 5583 3349 5595 3352
rect 5537 3343 5595 3349
rect 6546 3340 6552 3352
rect 6604 3340 6610 3392
rect 6656 3380 6684 3420
rect 7374 3408 7380 3460
rect 7432 3448 7438 3460
rect 9858 3448 9864 3460
rect 7432 3420 9864 3448
rect 7432 3408 7438 3420
rect 9858 3408 9864 3420
rect 9916 3408 9922 3460
rect 10229 3451 10287 3457
rect 10229 3417 10241 3451
rect 10275 3448 10287 3451
rect 11238 3448 11244 3460
rect 10275 3420 11244 3448
rect 10275 3417 10287 3420
rect 10229 3411 10287 3417
rect 11238 3408 11244 3420
rect 11296 3408 11302 3460
rect 11793 3451 11851 3457
rect 11793 3417 11805 3451
rect 11839 3448 11851 3451
rect 14660 3448 14688 3624
rect 16574 3612 16580 3624
rect 16632 3612 16638 3664
rect 18868 3655 18926 3661
rect 18868 3621 18880 3655
rect 18914 3652 18926 3655
rect 18966 3652 18972 3664
rect 18914 3624 18972 3652
rect 18914 3621 18926 3624
rect 18868 3615 18926 3621
rect 18966 3612 18972 3624
rect 19024 3612 19030 3664
rect 19058 3612 19064 3664
rect 19116 3612 19122 3664
rect 14734 3544 14740 3596
rect 14792 3584 14798 3596
rect 15657 3587 15715 3593
rect 15657 3584 15669 3587
rect 14792 3556 15669 3584
rect 14792 3544 14798 3556
rect 15657 3553 15669 3556
rect 15703 3553 15715 3587
rect 15657 3547 15715 3553
rect 15746 3544 15752 3596
rect 15804 3584 15810 3596
rect 17129 3587 17187 3593
rect 15804 3556 15849 3584
rect 15804 3544 15810 3556
rect 17129 3553 17141 3587
rect 17175 3584 17187 3587
rect 19076 3584 19104 3612
rect 17175 3556 19104 3584
rect 17175 3553 17187 3556
rect 17129 3547 17187 3553
rect 15933 3519 15991 3525
rect 15933 3485 15945 3519
rect 15979 3516 15991 3519
rect 15979 3488 16436 3516
rect 15979 3485 15991 3488
rect 15933 3479 15991 3485
rect 11839 3420 14688 3448
rect 11839 3417 11851 3420
rect 11793 3411 11851 3417
rect 15010 3408 15016 3460
rect 15068 3448 15074 3460
rect 15948 3448 15976 3479
rect 15068 3420 15976 3448
rect 15068 3408 15074 3420
rect 8386 3380 8392 3392
rect 6656 3352 8392 3380
rect 8386 3340 8392 3352
rect 8444 3340 8450 3392
rect 10042 3340 10048 3392
rect 10100 3380 10106 3392
rect 10686 3380 10692 3392
rect 10100 3352 10692 3380
rect 10100 3340 10106 3352
rect 10686 3340 10692 3352
rect 10744 3380 10750 3392
rect 10870 3380 10876 3392
rect 10744 3352 10876 3380
rect 10744 3340 10750 3352
rect 10870 3340 10876 3352
rect 10928 3340 10934 3392
rect 11054 3340 11060 3392
rect 11112 3380 11118 3392
rect 15289 3383 15347 3389
rect 15289 3380 15301 3383
rect 11112 3352 15301 3380
rect 11112 3340 11118 3352
rect 15289 3349 15301 3352
rect 15335 3349 15347 3383
rect 16408 3380 16436 3488
rect 16482 3476 16488 3528
rect 16540 3516 16546 3528
rect 17313 3519 17371 3525
rect 17313 3516 17325 3519
rect 16540 3488 17325 3516
rect 16540 3476 16546 3488
rect 17313 3485 17325 3488
rect 17359 3485 17371 3519
rect 17313 3479 17371 3485
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 18601 3519 18659 3525
rect 18601 3516 18613 3519
rect 18288 3488 18613 3516
rect 18288 3476 18294 3488
rect 18601 3485 18613 3488
rect 18647 3485 18659 3519
rect 18601 3479 18659 3485
rect 19981 3383 20039 3389
rect 19981 3380 19993 3383
rect 16408 3352 19993 3380
rect 15289 3343 15347 3349
rect 19981 3349 19993 3352
rect 20027 3349 20039 3383
rect 19981 3343 20039 3349
rect 1104 3290 21896 3312
rect 1104 3238 4447 3290
rect 4499 3238 4511 3290
rect 4563 3238 4575 3290
rect 4627 3238 4639 3290
rect 4691 3238 11378 3290
rect 11430 3238 11442 3290
rect 11494 3238 11506 3290
rect 11558 3238 11570 3290
rect 11622 3238 18308 3290
rect 18360 3238 18372 3290
rect 18424 3238 18436 3290
rect 18488 3238 18500 3290
rect 18552 3238 21896 3290
rect 1104 3216 21896 3238
rect 2869 3179 2927 3185
rect 2869 3145 2881 3179
rect 2915 3176 2927 3179
rect 5902 3176 5908 3188
rect 2915 3148 5908 3176
rect 2915 3145 2927 3148
rect 2869 3139 2927 3145
rect 5902 3136 5908 3148
rect 5960 3136 5966 3188
rect 6730 3136 6736 3188
rect 6788 3176 6794 3188
rect 6825 3179 6883 3185
rect 6825 3176 6837 3179
rect 6788 3148 6837 3176
rect 6788 3136 6794 3148
rect 6825 3145 6837 3148
rect 6871 3145 6883 3179
rect 6825 3139 6883 3145
rect 8662 3136 8668 3188
rect 8720 3176 8726 3188
rect 10686 3176 10692 3188
rect 8720 3148 10548 3176
rect 10647 3148 10692 3176
rect 8720 3136 8726 3148
rect 2774 3068 2780 3120
rect 2832 3108 2838 3120
rect 2832 3080 2877 3108
rect 2832 3068 2838 3080
rect 5074 3068 5080 3120
rect 5132 3108 5138 3120
rect 5169 3111 5227 3117
rect 5169 3108 5181 3111
rect 5132 3080 5181 3108
rect 5132 3068 5138 3080
rect 5169 3077 5181 3080
rect 5215 3077 5227 3111
rect 5169 3071 5227 3077
rect 5258 3068 5264 3120
rect 5316 3108 5322 3120
rect 7742 3108 7748 3120
rect 5316 3080 5361 3108
rect 7300 3080 7748 3108
rect 5316 3068 5322 3080
rect 3513 3043 3571 3049
rect 3513 3009 3525 3043
rect 3559 3040 3571 3043
rect 3602 3040 3608 3052
rect 3559 3012 3608 3040
rect 3559 3009 3571 3012
rect 3513 3003 3571 3009
rect 3602 3000 3608 3012
rect 3660 3040 3666 3052
rect 3660 3012 3924 3040
rect 3660 3000 3666 3012
rect 1397 2975 1455 2981
rect 1397 2941 1409 2975
rect 1443 2972 1455 2975
rect 1486 2972 1492 2984
rect 1443 2944 1492 2972
rect 1443 2941 1455 2944
rect 1397 2935 1455 2941
rect 1486 2932 1492 2944
rect 1544 2972 1550 2984
rect 3789 2975 3847 2981
rect 3789 2972 3801 2975
rect 1544 2944 3801 2972
rect 1544 2932 1550 2944
rect 3789 2941 3801 2944
rect 3835 2941 3847 2975
rect 3896 2972 3924 3012
rect 4798 3000 4804 3052
rect 4856 3040 4862 3052
rect 5813 3043 5871 3049
rect 5813 3040 5825 3043
rect 4856 3012 5825 3040
rect 4856 3000 4862 3012
rect 5813 3009 5825 3012
rect 5859 3009 5871 3043
rect 6362 3040 6368 3052
rect 6323 3012 6368 3040
rect 5813 3003 5871 3009
rect 6362 3000 6368 3012
rect 6420 3000 6426 3052
rect 7300 3049 7328 3080
rect 7742 3068 7748 3080
rect 7800 3068 7806 3120
rect 10520 3108 10548 3148
rect 10686 3136 10692 3148
rect 10744 3136 10750 3188
rect 12158 3176 12164 3188
rect 10796 3148 12164 3176
rect 10796 3108 10824 3148
rect 12158 3136 12164 3148
rect 12216 3136 12222 3188
rect 12802 3176 12808 3188
rect 12763 3148 12808 3176
rect 12802 3136 12808 3148
rect 12860 3136 12866 3188
rect 13354 3136 13360 3188
rect 13412 3136 13418 3188
rect 13446 3136 13452 3188
rect 13504 3176 13510 3188
rect 14369 3179 14427 3185
rect 14369 3176 14381 3179
rect 13504 3148 14381 3176
rect 13504 3136 13510 3148
rect 14369 3145 14381 3148
rect 14415 3145 14427 3179
rect 14369 3139 14427 3145
rect 14550 3136 14556 3188
rect 14608 3176 14614 3188
rect 20714 3176 20720 3188
rect 14608 3148 20720 3176
rect 14608 3136 14614 3148
rect 20714 3136 20720 3148
rect 20772 3136 20778 3188
rect 10520 3080 10824 3108
rect 7285 3043 7343 3049
rect 7285 3009 7297 3043
rect 7331 3009 7343 3043
rect 7285 3003 7343 3009
rect 7469 3043 7527 3049
rect 7469 3009 7481 3043
rect 7515 3040 7527 3043
rect 8478 3040 8484 3052
rect 7515 3012 8484 3040
rect 7515 3009 7527 3012
rect 7469 3003 7527 3009
rect 8478 3000 8484 3012
rect 8536 3000 8542 3052
rect 13372 3049 13400 3136
rect 18046 3068 18052 3120
rect 18104 3108 18110 3120
rect 19613 3111 19671 3117
rect 18104 3080 18276 3108
rect 18104 3068 18110 3080
rect 13357 3043 13415 3049
rect 13357 3009 13369 3043
rect 13403 3009 13415 3043
rect 13357 3003 13415 3009
rect 14182 3000 14188 3052
rect 14240 3040 14246 3052
rect 15010 3040 15016 3052
rect 14240 3012 14872 3040
rect 14971 3012 15016 3040
rect 14240 3000 14246 3012
rect 4045 2975 4103 2981
rect 4045 2972 4057 2975
rect 3896 2944 4057 2972
rect 3789 2935 3847 2941
rect 4045 2941 4057 2944
rect 4091 2941 4103 2975
rect 4045 2935 4103 2941
rect 5442 2932 5448 2984
rect 5500 2972 5506 2984
rect 5500 2944 5672 2972
rect 5500 2932 5506 2944
rect 1664 2907 1722 2913
rect 1664 2873 1676 2907
rect 1710 2904 1722 2907
rect 2222 2904 2228 2916
rect 1710 2876 2228 2904
rect 1710 2873 1722 2876
rect 1664 2867 1722 2873
rect 2222 2864 2228 2876
rect 2280 2864 2286 2916
rect 3237 2907 3295 2913
rect 3237 2873 3249 2907
rect 3283 2904 3295 2907
rect 4246 2904 4252 2916
rect 3283 2876 4252 2904
rect 3283 2873 3295 2876
rect 3237 2867 3295 2873
rect 4246 2864 4252 2876
rect 4304 2864 4310 2916
rect 5534 2904 5540 2916
rect 5092 2876 5540 2904
rect 658 2796 664 2848
rect 716 2836 722 2848
rect 1762 2836 1768 2848
rect 716 2808 1768 2836
rect 716 2796 722 2808
rect 1762 2796 1768 2808
rect 1820 2796 1826 2848
rect 3329 2839 3387 2845
rect 3329 2805 3341 2839
rect 3375 2836 3387 2839
rect 5092 2836 5120 2876
rect 5534 2864 5540 2876
rect 5592 2864 5598 2916
rect 5644 2904 5672 2944
rect 5718 2932 5724 2984
rect 5776 2972 5782 2984
rect 6089 2975 6147 2981
rect 5776 2944 5821 2972
rect 5776 2932 5782 2944
rect 6089 2941 6101 2975
rect 6135 2972 6147 2975
rect 6178 2972 6184 2984
rect 6135 2944 6184 2972
rect 6135 2941 6147 2944
rect 6089 2935 6147 2941
rect 6178 2932 6184 2944
rect 6236 2932 6242 2984
rect 6546 2932 6552 2984
rect 6604 2972 6610 2984
rect 7837 2975 7895 2981
rect 7837 2972 7849 2975
rect 6604 2944 7849 2972
rect 6604 2932 6610 2944
rect 7837 2941 7849 2944
rect 7883 2941 7895 2975
rect 7837 2935 7895 2941
rect 9122 2932 9128 2984
rect 9180 2972 9186 2984
rect 9582 2981 9588 2984
rect 9309 2975 9367 2981
rect 9309 2972 9321 2975
rect 9180 2944 9321 2972
rect 9180 2932 9186 2944
rect 9309 2941 9321 2944
rect 9355 2941 9367 2975
rect 9576 2972 9588 2981
rect 9543 2944 9588 2972
rect 9309 2935 9367 2941
rect 9576 2935 9588 2944
rect 9582 2932 9588 2935
rect 9640 2932 9646 2984
rect 9858 2932 9864 2984
rect 9916 2972 9922 2984
rect 14737 2975 14795 2981
rect 14737 2972 14749 2975
rect 9916 2944 14749 2972
rect 9916 2932 9922 2944
rect 14737 2941 14749 2944
rect 14783 2941 14795 2975
rect 14844 2972 14872 3012
rect 15010 3000 15016 3012
rect 15068 3000 15074 3052
rect 15286 3000 15292 3052
rect 15344 3040 15350 3052
rect 18248 3049 18276 3080
rect 19613 3077 19625 3111
rect 19659 3108 19671 3111
rect 21266 3108 21272 3120
rect 19659 3080 21272 3108
rect 19659 3077 19671 3080
rect 19613 3071 19671 3077
rect 21266 3068 21272 3080
rect 21324 3068 21330 3120
rect 16117 3043 16175 3049
rect 16117 3040 16129 3043
rect 15344 3012 16129 3040
rect 15344 3000 15350 3012
rect 16117 3009 16129 3012
rect 16163 3009 16175 3043
rect 16117 3003 16175 3009
rect 18233 3043 18291 3049
rect 18233 3009 18245 3043
rect 18279 3009 18291 3043
rect 18233 3003 18291 3009
rect 15933 2975 15991 2981
rect 15933 2972 15945 2975
rect 14844 2944 15945 2972
rect 14737 2935 14795 2941
rect 15933 2941 15945 2944
rect 15979 2941 15991 2975
rect 15933 2935 15991 2941
rect 18049 2975 18107 2981
rect 18049 2941 18061 2975
rect 18095 2972 18107 2975
rect 19150 2972 19156 2984
rect 18095 2944 19156 2972
rect 18095 2941 18107 2944
rect 18049 2935 18107 2941
rect 19150 2932 19156 2944
rect 19208 2932 19214 2984
rect 19426 2972 19432 2984
rect 19387 2944 19432 2972
rect 19426 2932 19432 2944
rect 19484 2932 19490 2984
rect 20530 2972 20536 2984
rect 20491 2944 20536 2972
rect 20530 2932 20536 2944
rect 20588 2932 20594 2984
rect 5902 2904 5908 2916
rect 5644 2876 5908 2904
rect 5902 2864 5908 2876
rect 5960 2864 5966 2916
rect 7193 2907 7251 2913
rect 7193 2873 7205 2907
rect 7239 2904 7251 2907
rect 7742 2904 7748 2916
rect 7239 2876 7748 2904
rect 7239 2873 7251 2876
rect 7193 2867 7251 2873
rect 7742 2864 7748 2876
rect 7800 2864 7806 2916
rect 8113 2907 8171 2913
rect 8113 2873 8125 2907
rect 8159 2904 8171 2907
rect 11422 2904 11428 2916
rect 8159 2876 11428 2904
rect 8159 2873 8171 2876
rect 8113 2867 8171 2873
rect 11422 2864 11428 2876
rect 11480 2864 11486 2916
rect 13173 2907 13231 2913
rect 13173 2904 13185 2907
rect 12544 2876 13185 2904
rect 3375 2808 5120 2836
rect 3375 2805 3387 2808
rect 3329 2799 3387 2805
rect 5166 2796 5172 2848
rect 5224 2836 5230 2848
rect 5629 2839 5687 2845
rect 5629 2836 5641 2839
rect 5224 2808 5641 2836
rect 5224 2796 5230 2808
rect 5629 2805 5641 2808
rect 5675 2805 5687 2839
rect 5629 2799 5687 2805
rect 6362 2796 6368 2848
rect 6420 2836 6426 2848
rect 7466 2836 7472 2848
rect 6420 2808 7472 2836
rect 6420 2796 6426 2808
rect 7466 2796 7472 2808
rect 7524 2796 7530 2848
rect 8386 2796 8392 2848
rect 8444 2836 8450 2848
rect 12544 2836 12572 2876
rect 13173 2873 13185 2876
rect 13219 2904 13231 2907
rect 14829 2907 14887 2913
rect 14829 2904 14841 2907
rect 13219 2876 14841 2904
rect 13219 2873 13231 2876
rect 13173 2867 13231 2873
rect 14829 2873 14841 2876
rect 14875 2873 14887 2907
rect 14829 2867 14887 2873
rect 15286 2864 15292 2916
rect 15344 2904 15350 2916
rect 15838 2904 15844 2916
rect 15344 2876 15844 2904
rect 15344 2864 15350 2876
rect 15838 2864 15844 2876
rect 15896 2864 15902 2916
rect 20162 2864 20168 2916
rect 20220 2904 20226 2916
rect 22646 2904 22652 2916
rect 20220 2876 22652 2904
rect 20220 2864 20226 2876
rect 22646 2864 22652 2876
rect 22704 2864 22710 2916
rect 13262 2836 13268 2848
rect 8444 2808 12572 2836
rect 13223 2808 13268 2836
rect 8444 2796 8450 2808
rect 13262 2796 13268 2808
rect 13320 2796 13326 2848
rect 13998 2796 14004 2848
rect 14056 2836 14062 2848
rect 19334 2836 19340 2848
rect 14056 2808 19340 2836
rect 14056 2796 14062 2808
rect 19334 2796 19340 2808
rect 19392 2796 19398 2848
rect 20717 2839 20775 2845
rect 20717 2805 20729 2839
rect 20763 2836 20775 2839
rect 22186 2836 22192 2848
rect 20763 2808 22192 2836
rect 20763 2805 20775 2808
rect 20717 2799 20775 2805
rect 22186 2796 22192 2808
rect 22244 2796 22250 2848
rect 1104 2746 21896 2768
rect 1104 2694 7912 2746
rect 7964 2694 7976 2746
rect 8028 2694 8040 2746
rect 8092 2694 8104 2746
rect 8156 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 15035 2746
rect 15087 2694 21896 2746
rect 1104 2672 21896 2694
rect 2866 2632 2872 2644
rect 2827 2604 2872 2632
rect 2866 2592 2872 2604
rect 2924 2592 2930 2644
rect 3142 2592 3148 2644
rect 3200 2632 3206 2644
rect 3237 2635 3295 2641
rect 3237 2632 3249 2635
rect 3200 2604 3249 2632
rect 3200 2592 3206 2604
rect 3237 2601 3249 2604
rect 3283 2601 3295 2635
rect 3237 2595 3295 2601
rect 3329 2635 3387 2641
rect 3329 2601 3341 2635
rect 3375 2632 3387 2635
rect 3418 2632 3424 2644
rect 3375 2604 3424 2632
rect 3375 2601 3387 2604
rect 3329 2595 3387 2601
rect 3418 2592 3424 2604
rect 3476 2592 3482 2644
rect 5534 2632 5540 2644
rect 5495 2604 5540 2632
rect 5534 2592 5540 2604
rect 5592 2592 5598 2644
rect 5810 2592 5816 2644
rect 5868 2632 5874 2644
rect 5905 2635 5963 2641
rect 5905 2632 5917 2635
rect 5868 2604 5917 2632
rect 5868 2592 5874 2604
rect 5905 2601 5917 2604
rect 5951 2601 5963 2635
rect 6914 2632 6920 2644
rect 6875 2604 6920 2632
rect 5905 2595 5963 2601
rect 6914 2592 6920 2604
rect 6972 2592 6978 2644
rect 7377 2635 7435 2641
rect 7377 2601 7389 2635
rect 7423 2632 7435 2635
rect 8757 2635 8815 2641
rect 7423 2604 8708 2632
rect 7423 2601 7435 2604
rect 7377 2595 7435 2601
rect 2038 2524 2044 2576
rect 2096 2564 2102 2576
rect 3160 2564 3188 2592
rect 2096 2536 3188 2564
rect 4332 2567 4390 2573
rect 2096 2524 2102 2536
rect 4332 2533 4344 2567
rect 4378 2564 4390 2567
rect 4798 2564 4804 2576
rect 4378 2536 4804 2564
rect 4378 2533 4390 2536
rect 4332 2527 4390 2533
rect 4798 2524 4804 2536
rect 4856 2524 4862 2576
rect 7285 2567 7343 2573
rect 7285 2533 7297 2567
rect 7331 2564 7343 2567
rect 7466 2564 7472 2576
rect 7331 2536 7472 2564
rect 7331 2533 7343 2536
rect 7285 2527 7343 2533
rect 7466 2524 7472 2536
rect 7524 2524 7530 2576
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2496 1455 2499
rect 1486 2496 1492 2508
rect 1443 2468 1492 2496
rect 1443 2465 1455 2468
rect 1397 2459 1455 2465
rect 1486 2456 1492 2468
rect 1544 2456 1550 2508
rect 1664 2499 1722 2505
rect 1664 2465 1676 2499
rect 1710 2496 1722 2499
rect 3418 2496 3424 2508
rect 1710 2468 3424 2496
rect 1710 2465 1722 2468
rect 1664 2459 1722 2465
rect 3418 2456 3424 2468
rect 3476 2456 3482 2508
rect 3694 2456 3700 2508
rect 3752 2496 3758 2508
rect 5997 2499 6055 2505
rect 5997 2496 6009 2499
rect 3752 2468 6009 2496
rect 3752 2456 3758 2468
rect 5997 2465 6009 2468
rect 6043 2496 6055 2499
rect 6086 2496 6092 2508
rect 6043 2468 6092 2496
rect 6043 2465 6055 2468
rect 5997 2459 6055 2465
rect 6086 2456 6092 2468
rect 6144 2456 6150 2508
rect 6365 2499 6423 2505
rect 6365 2465 6377 2499
rect 6411 2496 6423 2499
rect 7926 2496 7932 2508
rect 6411 2468 7932 2496
rect 6411 2465 6423 2468
rect 6365 2459 6423 2465
rect 7926 2456 7932 2468
rect 7984 2456 7990 2508
rect 8110 2496 8116 2508
rect 8071 2468 8116 2496
rect 8110 2456 8116 2468
rect 8168 2456 8174 2508
rect 8570 2496 8576 2508
rect 8531 2468 8576 2496
rect 8570 2456 8576 2468
rect 8628 2456 8634 2508
rect 8680 2496 8708 2604
rect 8757 2601 8769 2635
rect 8803 2601 8815 2635
rect 8757 2595 8815 2601
rect 8772 2564 8800 2595
rect 9674 2592 9680 2644
rect 9732 2632 9738 2644
rect 10137 2635 10195 2641
rect 10137 2632 10149 2635
rect 9732 2604 10149 2632
rect 9732 2592 9738 2604
rect 10137 2601 10149 2604
rect 10183 2601 10195 2635
rect 10137 2595 10195 2601
rect 10229 2635 10287 2641
rect 10229 2601 10241 2635
rect 10275 2632 10287 2635
rect 10410 2632 10416 2644
rect 10275 2604 10416 2632
rect 10275 2601 10287 2604
rect 10229 2595 10287 2601
rect 10410 2592 10416 2604
rect 10468 2592 10474 2644
rect 12434 2592 12440 2644
rect 12492 2632 12498 2644
rect 12621 2635 12679 2641
rect 12492 2604 12572 2632
rect 12492 2592 12498 2604
rect 8772 2536 12480 2564
rect 12452 2508 12480 2536
rect 8846 2496 8852 2508
rect 8680 2468 8852 2496
rect 8846 2456 8852 2468
rect 8904 2456 8910 2508
rect 11422 2496 11428 2508
rect 11383 2468 11428 2496
rect 11422 2456 11428 2468
rect 11480 2456 11486 2508
rect 12434 2456 12440 2508
rect 12492 2456 12498 2508
rect 12544 2496 12572 2604
rect 12621 2601 12633 2635
rect 12667 2632 12679 2635
rect 12986 2632 12992 2644
rect 12667 2604 12992 2632
rect 12667 2601 12679 2604
rect 12621 2595 12679 2601
rect 12986 2592 12992 2604
rect 13044 2592 13050 2644
rect 20162 2632 20168 2644
rect 20123 2604 20168 2632
rect 20162 2592 20168 2604
rect 20220 2592 20226 2644
rect 12894 2524 12900 2576
rect 12952 2564 12958 2576
rect 13081 2567 13139 2573
rect 13081 2564 13093 2567
rect 12952 2536 13093 2564
rect 12952 2524 12958 2536
rect 13081 2533 13093 2536
rect 13127 2533 13139 2567
rect 13081 2527 13139 2533
rect 15378 2524 15384 2576
rect 15436 2564 15442 2576
rect 15749 2567 15807 2573
rect 15749 2564 15761 2567
rect 15436 2536 15761 2564
rect 15436 2524 15442 2536
rect 15749 2533 15761 2536
rect 15795 2533 15807 2567
rect 15749 2527 15807 2533
rect 17218 2524 17224 2576
rect 17276 2524 17282 2576
rect 12989 2499 13047 2505
rect 12989 2496 13001 2499
rect 12544 2468 13001 2496
rect 12989 2465 13001 2468
rect 13035 2465 13047 2499
rect 12989 2459 13047 2465
rect 13538 2456 13544 2508
rect 13596 2496 13602 2508
rect 14185 2499 14243 2505
rect 14185 2496 14197 2499
rect 13596 2468 14197 2496
rect 13596 2456 13602 2468
rect 14185 2465 14197 2468
rect 14231 2465 14243 2499
rect 14734 2496 14740 2508
rect 14185 2459 14243 2465
rect 14292 2468 14740 2496
rect 3513 2431 3571 2437
rect 3513 2397 3525 2431
rect 3559 2428 3571 2431
rect 3602 2428 3608 2440
rect 3559 2400 3608 2428
rect 3559 2397 3571 2400
rect 3513 2391 3571 2397
rect 3602 2388 3608 2400
rect 3660 2388 3666 2440
rect 6181 2431 6239 2437
rect 6181 2397 6193 2431
rect 6227 2428 6239 2431
rect 6454 2428 6460 2440
rect 6227 2400 6460 2428
rect 6227 2397 6239 2400
rect 6181 2391 6239 2397
rect 6454 2388 6460 2400
rect 6512 2428 6518 2440
rect 7469 2431 7527 2437
rect 7469 2428 7481 2431
rect 6512 2400 7481 2428
rect 6512 2388 6518 2400
rect 7469 2397 7481 2400
rect 7515 2397 7527 2431
rect 8202 2428 8208 2440
rect 8163 2400 8208 2428
rect 7469 2391 7527 2397
rect 8202 2388 8208 2400
rect 8260 2388 8266 2440
rect 8297 2431 8355 2437
rect 8297 2397 8309 2431
rect 8343 2428 8355 2431
rect 8662 2428 8668 2440
rect 8343 2400 8668 2428
rect 8343 2397 8355 2400
rect 8297 2391 8355 2397
rect 2590 2320 2596 2372
rect 2648 2360 2654 2372
rect 2648 2332 4108 2360
rect 2648 2320 2654 2332
rect 2774 2252 2780 2304
rect 2832 2292 2838 2304
rect 4080 2292 4108 2332
rect 5902 2320 5908 2372
rect 5960 2360 5966 2372
rect 5960 2332 7236 2360
rect 5960 2320 5966 2332
rect 5445 2295 5503 2301
rect 5445 2292 5457 2295
rect 2832 2264 2877 2292
rect 4080 2264 5457 2292
rect 2832 2252 2838 2264
rect 5445 2261 5457 2264
rect 5491 2261 5503 2295
rect 6546 2292 6552 2304
rect 6507 2264 6552 2292
rect 5445 2255 5503 2261
rect 6546 2252 6552 2264
rect 6604 2252 6610 2304
rect 7208 2292 7236 2332
rect 7282 2320 7288 2372
rect 7340 2360 7346 2372
rect 7745 2363 7803 2369
rect 7745 2360 7757 2363
rect 7340 2332 7757 2360
rect 7340 2320 7346 2332
rect 7745 2329 7757 2332
rect 7791 2329 7803 2363
rect 7745 2323 7803 2329
rect 8312 2292 8340 2391
rect 8662 2388 8668 2400
rect 8720 2388 8726 2440
rect 9950 2388 9956 2440
rect 10008 2428 10014 2440
rect 10413 2431 10471 2437
rect 10413 2428 10425 2431
rect 10008 2400 10425 2428
rect 10008 2388 10014 2400
rect 10413 2397 10425 2400
rect 10459 2428 10471 2431
rect 13265 2431 13323 2437
rect 13265 2428 13277 2431
rect 10459 2400 13277 2428
rect 10459 2397 10471 2400
rect 10413 2391 10471 2397
rect 13265 2397 13277 2400
rect 13311 2428 13323 2431
rect 14292 2428 14320 2468
rect 14734 2456 14740 2468
rect 14792 2456 14798 2508
rect 15470 2496 15476 2508
rect 15431 2468 15476 2496
rect 15470 2456 15476 2468
rect 15528 2456 15534 2508
rect 16853 2499 16911 2505
rect 16853 2465 16865 2499
rect 16899 2496 16911 2499
rect 17236 2496 17264 2524
rect 18690 2496 18696 2508
rect 16899 2468 17264 2496
rect 18651 2468 18696 2496
rect 16899 2465 16911 2468
rect 16853 2459 16911 2465
rect 18690 2456 18696 2468
rect 18748 2456 18754 2508
rect 19978 2496 19984 2508
rect 19939 2468 19984 2496
rect 19978 2456 19984 2468
rect 20036 2456 20042 2508
rect 13311 2400 14320 2428
rect 13311 2397 13323 2400
rect 13265 2391 13323 2397
rect 14642 2388 14648 2440
rect 14700 2428 14706 2440
rect 17037 2431 17095 2437
rect 17037 2428 17049 2431
rect 14700 2400 17049 2428
rect 14700 2388 14706 2400
rect 17037 2397 17049 2400
rect 17083 2397 17095 2431
rect 17037 2391 17095 2397
rect 17218 2388 17224 2440
rect 17276 2428 17282 2440
rect 18877 2431 18935 2437
rect 18877 2428 18889 2431
rect 17276 2400 18889 2428
rect 17276 2388 17282 2400
rect 18877 2397 18889 2400
rect 18923 2397 18935 2431
rect 18877 2391 18935 2397
rect 9769 2363 9827 2369
rect 9769 2329 9781 2363
rect 9815 2360 9827 2363
rect 10134 2360 10140 2372
rect 9815 2332 10140 2360
rect 9815 2329 9827 2332
rect 9769 2323 9827 2329
rect 10134 2320 10140 2332
rect 10192 2320 10198 2372
rect 11609 2363 11667 2369
rect 11609 2329 11621 2363
rect 11655 2360 11667 2363
rect 14090 2360 14096 2372
rect 11655 2332 14096 2360
rect 11655 2329 11667 2332
rect 11609 2323 11667 2329
rect 14090 2320 14096 2332
rect 14148 2320 14154 2372
rect 7208 2264 8340 2292
rect 12434 2252 12440 2304
rect 12492 2292 12498 2304
rect 13446 2292 13452 2304
rect 12492 2264 13452 2292
rect 12492 2252 12498 2264
rect 13446 2252 13452 2264
rect 13504 2252 13510 2304
rect 13538 2252 13544 2304
rect 13596 2292 13602 2304
rect 14369 2295 14427 2301
rect 14369 2292 14381 2295
rect 13596 2264 14381 2292
rect 13596 2252 13602 2264
rect 14369 2261 14381 2264
rect 14415 2261 14427 2295
rect 14369 2255 14427 2261
rect 1104 2202 21896 2224
rect 1104 2150 4447 2202
rect 4499 2150 4511 2202
rect 4563 2150 4575 2202
rect 4627 2150 4639 2202
rect 4691 2150 11378 2202
rect 11430 2150 11442 2202
rect 11494 2150 11506 2202
rect 11558 2150 11570 2202
rect 11622 2150 18308 2202
rect 18360 2150 18372 2202
rect 18424 2150 18436 2202
rect 18488 2150 18500 2202
rect 18552 2150 21896 2202
rect 1104 2128 21896 2150
rect 1578 2048 1584 2100
rect 1636 2088 1642 2100
rect 5350 2088 5356 2100
rect 1636 2060 5356 2088
rect 1636 2048 1642 2060
rect 5350 2048 5356 2060
rect 5408 2048 5414 2100
rect 6546 2048 6552 2100
rect 6604 2088 6610 2100
rect 15470 2088 15476 2100
rect 6604 2060 15476 2088
rect 6604 2048 6610 2060
rect 15470 2048 15476 2060
rect 15528 2048 15534 2100
rect 2590 1980 2596 2032
rect 2648 2020 2654 2032
rect 3786 2020 3792 2032
rect 2648 1992 3792 2020
rect 2648 1980 2654 1992
rect 3786 1980 3792 1992
rect 3844 1980 3850 2032
rect 8202 1980 8208 2032
rect 8260 2020 8266 2032
rect 8260 1992 13400 2020
rect 8260 1980 8266 1992
rect 2866 1912 2872 1964
rect 2924 1952 2930 1964
rect 13265 1955 13323 1961
rect 13265 1952 13277 1955
rect 2924 1924 13277 1952
rect 2924 1912 2930 1924
rect 13265 1921 13277 1924
rect 13311 1921 13323 1955
rect 13372 1952 13400 1992
rect 13446 1980 13452 2032
rect 13504 2020 13510 2032
rect 14458 2020 14464 2032
rect 13504 1992 14464 2020
rect 13504 1980 13510 1992
rect 14458 1980 14464 1992
rect 14516 1980 14522 2032
rect 16206 1952 16212 1964
rect 13372 1924 16212 1952
rect 13265 1915 13323 1921
rect 16206 1912 16212 1924
rect 16264 1912 16270 1964
rect 3326 1844 3332 1896
rect 3384 1884 3390 1896
rect 19978 1884 19984 1896
rect 3384 1856 19984 1884
rect 3384 1844 3390 1856
rect 19978 1844 19984 1856
rect 20036 1844 20042 1896
rect 8110 1776 8116 1828
rect 8168 1816 8174 1828
rect 16114 1816 16120 1828
rect 8168 1788 16120 1816
rect 8168 1776 8174 1788
rect 16114 1776 16120 1788
rect 16172 1776 16178 1828
rect 3602 1708 3608 1760
rect 3660 1748 3666 1760
rect 17494 1748 17500 1760
rect 3660 1720 17500 1748
rect 3660 1708 3666 1720
rect 17494 1708 17500 1720
rect 17552 1708 17558 1760
rect 2774 1640 2780 1692
rect 2832 1680 2838 1692
rect 15194 1680 15200 1692
rect 2832 1652 15200 1680
rect 2832 1640 2838 1652
rect 15194 1640 15200 1652
rect 15252 1640 15258 1692
rect 7926 1572 7932 1624
rect 7984 1612 7990 1624
rect 13814 1612 13820 1624
rect 7984 1584 13820 1612
rect 7984 1572 7990 1584
rect 13814 1572 13820 1584
rect 13872 1572 13878 1624
rect 9030 1504 9036 1556
rect 9088 1544 9094 1556
rect 17218 1544 17224 1556
rect 9088 1516 17224 1544
rect 9088 1504 9094 1516
rect 17218 1504 17224 1516
rect 17276 1504 17282 1556
rect 3418 1436 3424 1488
rect 3476 1476 3482 1488
rect 14366 1476 14372 1488
rect 3476 1448 14372 1476
rect 3476 1436 3482 1448
rect 14366 1436 14372 1448
rect 14424 1436 14430 1488
rect 19518 1476 19524 1488
rect 14476 1448 19524 1476
rect 13265 1411 13323 1417
rect 13265 1377 13277 1411
rect 13311 1408 13323 1411
rect 14476 1408 14504 1448
rect 19518 1436 19524 1448
rect 19576 1436 19582 1488
rect 13311 1380 14504 1408
rect 13311 1377 13323 1380
rect 13265 1371 13323 1377
rect 18322 1368 18328 1420
rect 18380 1408 18386 1420
rect 19058 1408 19064 1420
rect 18380 1380 19064 1408
rect 18380 1368 18386 1380
rect 19058 1368 19064 1380
rect 19116 1368 19122 1420
rect 12342 1300 12348 1352
rect 12400 1340 12406 1352
rect 18874 1340 18880 1352
rect 12400 1312 18880 1340
rect 12400 1300 12406 1312
rect 18874 1300 18880 1312
rect 18932 1300 18938 1352
rect 3602 280 3608 332
rect 3660 320 3666 332
rect 6270 320 6276 332
rect 3660 292 6276 320
rect 3660 280 3666 292
rect 6270 280 6276 292
rect 6328 280 6334 332
<< via1 >>
rect 3516 21292 3568 21344
rect 9312 21292 9364 21344
rect 3148 21088 3200 21140
rect 7656 21088 7708 21140
rect 4068 20816 4120 20868
rect 8208 20816 8260 20868
rect 4447 20646 4499 20698
rect 4511 20646 4563 20698
rect 4575 20646 4627 20698
rect 4639 20646 4691 20698
rect 11378 20646 11430 20698
rect 11442 20646 11494 20698
rect 11506 20646 11558 20698
rect 11570 20646 11622 20698
rect 18308 20646 18360 20698
rect 18372 20646 18424 20698
rect 18436 20646 18488 20698
rect 18500 20646 18552 20698
rect 3976 20544 4028 20596
rect 8208 20587 8260 20596
rect 8208 20553 8217 20587
rect 8217 20553 8251 20587
rect 8251 20553 8260 20587
rect 8208 20544 8260 20553
rect 18052 20544 18104 20596
rect 20168 20587 20220 20596
rect 20168 20553 20177 20587
rect 20177 20553 20211 20587
rect 20211 20553 20220 20587
rect 20168 20544 20220 20553
rect 4068 20476 4120 20528
rect 8208 20408 8260 20460
rect 12532 20408 12584 20460
rect 13636 20476 13688 20528
rect 13912 20408 13964 20460
rect 14004 20408 14056 20460
rect 18144 20476 18196 20528
rect 18236 20476 18288 20528
rect 18880 20451 18932 20460
rect 3792 20340 3844 20392
rect 5172 20383 5224 20392
rect 5172 20349 5181 20383
rect 5181 20349 5215 20383
rect 5215 20349 5224 20383
rect 5172 20340 5224 20349
rect 7196 20340 7248 20392
rect 7564 20340 7616 20392
rect 12624 20340 12676 20392
rect 5448 20272 5500 20324
rect 12164 20272 12216 20324
rect 17224 20340 17276 20392
rect 18880 20417 18889 20451
rect 18889 20417 18923 20451
rect 18923 20417 18932 20451
rect 18880 20408 18932 20417
rect 18788 20340 18840 20392
rect 1952 20247 2004 20256
rect 1952 20213 1961 20247
rect 1961 20213 1995 20247
rect 1995 20213 2004 20247
rect 1952 20204 2004 20213
rect 2872 20204 2924 20256
rect 3332 20204 3384 20256
rect 10048 20247 10100 20256
rect 10048 20213 10057 20247
rect 10057 20213 10091 20247
rect 10091 20213 10100 20247
rect 10048 20204 10100 20213
rect 11336 20247 11388 20256
rect 11336 20213 11345 20247
rect 11345 20213 11379 20247
rect 11379 20213 11388 20247
rect 11336 20204 11388 20213
rect 12440 20204 12492 20256
rect 15200 20204 15252 20256
rect 18052 20272 18104 20324
rect 15844 20247 15896 20256
rect 15844 20213 15853 20247
rect 15853 20213 15887 20247
rect 15887 20213 15896 20247
rect 15844 20204 15896 20213
rect 18604 20204 18656 20256
rect 7912 20102 7964 20154
rect 7976 20102 8028 20154
rect 8040 20102 8092 20154
rect 8104 20102 8156 20154
rect 14843 20102 14895 20154
rect 14907 20102 14959 20154
rect 14971 20102 15023 20154
rect 15035 20102 15087 20154
rect 10048 20000 10100 20052
rect 17868 20000 17920 20052
rect 19156 20000 19208 20052
rect 1768 19907 1820 19916
rect 1768 19873 1777 19907
rect 1777 19873 1811 19907
rect 1811 19873 1820 19907
rect 1768 19864 1820 19873
rect 3240 19864 3292 19916
rect 5540 19907 5592 19916
rect 5540 19873 5549 19907
rect 5549 19873 5583 19907
rect 5583 19873 5592 19907
rect 5540 19864 5592 19873
rect 5632 19839 5684 19848
rect 5632 19805 5641 19839
rect 5641 19805 5675 19839
rect 5675 19805 5684 19839
rect 5632 19796 5684 19805
rect 14372 19932 14424 19984
rect 15660 19932 15712 19984
rect 18236 19932 18288 19984
rect 7380 19864 7432 19916
rect 8576 19864 8628 19916
rect 12532 19907 12584 19916
rect 12532 19873 12566 19907
rect 12566 19873 12584 19907
rect 12532 19864 12584 19873
rect 13636 19864 13688 19916
rect 15384 19864 15436 19916
rect 19340 19864 19392 19916
rect 20076 19864 20128 19916
rect 6736 19839 6788 19848
rect 6736 19805 6745 19839
rect 6745 19805 6779 19839
rect 6779 19805 6788 19839
rect 6736 19796 6788 19805
rect 9680 19839 9732 19848
rect 9680 19805 9689 19839
rect 9689 19805 9723 19839
rect 9723 19805 9732 19839
rect 9680 19796 9732 19805
rect 11888 19796 11940 19848
rect 18144 19839 18196 19848
rect 5724 19728 5776 19780
rect 11336 19728 11388 19780
rect 11980 19728 12032 19780
rect 2780 19660 2832 19712
rect 3056 19703 3108 19712
rect 3056 19669 3065 19703
rect 3065 19669 3099 19703
rect 3099 19669 3108 19703
rect 3056 19660 3108 19669
rect 4160 19660 4212 19712
rect 4804 19660 4856 19712
rect 12164 19660 12216 19712
rect 13912 19660 13964 19712
rect 18144 19805 18153 19839
rect 18153 19805 18187 19839
rect 18187 19805 18196 19839
rect 18144 19796 18196 19805
rect 18880 19796 18932 19848
rect 20168 19796 20220 19848
rect 16396 19660 16448 19712
rect 16672 19703 16724 19712
rect 16672 19669 16681 19703
rect 16681 19669 16715 19703
rect 16715 19669 16724 19703
rect 16672 19660 16724 19669
rect 16764 19660 16816 19712
rect 4447 19558 4499 19610
rect 4511 19558 4563 19610
rect 4575 19558 4627 19610
rect 4639 19558 4691 19610
rect 11378 19558 11430 19610
rect 11442 19558 11494 19610
rect 11506 19558 11558 19610
rect 11570 19558 11622 19610
rect 18308 19558 18360 19610
rect 18372 19558 18424 19610
rect 18436 19558 18488 19610
rect 18500 19558 18552 19610
rect 5540 19456 5592 19508
rect 19340 19456 19392 19508
rect 5172 19320 5224 19372
rect 2688 19252 2740 19304
rect 4804 19295 4856 19304
rect 3516 19184 3568 19236
rect 4804 19261 4813 19295
rect 4813 19261 4847 19295
rect 4847 19261 4856 19295
rect 4804 19252 4856 19261
rect 5816 19320 5868 19372
rect 7380 19363 7432 19372
rect 7380 19329 7389 19363
rect 7389 19329 7423 19363
rect 7423 19329 7432 19363
rect 7380 19320 7432 19329
rect 10784 19363 10836 19372
rect 10784 19329 10793 19363
rect 10793 19329 10827 19363
rect 10827 19329 10836 19363
rect 10784 19320 10836 19329
rect 15384 19320 15436 19372
rect 18144 19320 18196 19372
rect 20168 19363 20220 19372
rect 20168 19329 20177 19363
rect 20177 19329 20211 19363
rect 20211 19329 20220 19363
rect 20168 19320 20220 19329
rect 2964 19116 3016 19168
rect 3148 19116 3200 19168
rect 7104 19184 7156 19236
rect 8852 19252 8904 19304
rect 12808 19252 12860 19304
rect 8576 19184 8628 19236
rect 5540 19116 5592 19168
rect 10416 19184 10468 19236
rect 10600 19227 10652 19236
rect 10600 19193 10609 19227
rect 10609 19193 10643 19227
rect 10643 19193 10652 19227
rect 10600 19184 10652 19193
rect 11888 19184 11940 19236
rect 15200 19252 15252 19304
rect 13912 19227 13964 19236
rect 13912 19193 13946 19227
rect 13946 19193 13964 19227
rect 13912 19184 13964 19193
rect 15292 19184 15344 19236
rect 17132 19184 17184 19236
rect 18604 19184 18656 19236
rect 18972 19184 19024 19236
rect 8760 19116 8812 19168
rect 10232 19159 10284 19168
rect 10232 19125 10241 19159
rect 10241 19125 10275 19159
rect 10275 19125 10284 19159
rect 10232 19116 10284 19125
rect 10692 19159 10744 19168
rect 10692 19125 10701 19159
rect 10701 19125 10735 19159
rect 10735 19125 10744 19159
rect 10692 19116 10744 19125
rect 12716 19159 12768 19168
rect 12716 19125 12725 19159
rect 12725 19125 12759 19159
rect 12759 19125 12768 19159
rect 12716 19116 12768 19125
rect 15384 19116 15436 19168
rect 15752 19116 15804 19168
rect 18052 19159 18104 19168
rect 18052 19125 18061 19159
rect 18061 19125 18095 19159
rect 18095 19125 18104 19159
rect 18052 19116 18104 19125
rect 19064 19116 19116 19168
rect 7912 19014 7964 19066
rect 7976 19014 8028 19066
rect 8040 19014 8092 19066
rect 8104 19014 8156 19066
rect 14843 19014 14895 19066
rect 14907 19014 14959 19066
rect 14971 19014 15023 19066
rect 15035 19014 15087 19066
rect 2688 18912 2740 18964
rect 5172 18912 5224 18964
rect 6736 18912 6788 18964
rect 7380 18912 7432 18964
rect 8208 18912 8260 18964
rect 8576 18912 8628 18964
rect 10140 18912 10192 18964
rect 4068 18819 4120 18828
rect 4068 18785 4077 18819
rect 4077 18785 4111 18819
rect 4111 18785 4120 18819
rect 4068 18776 4120 18785
rect 7748 18844 7800 18896
rect 13636 18912 13688 18964
rect 15292 18955 15344 18964
rect 15292 18921 15301 18955
rect 15301 18921 15335 18955
rect 15335 18921 15344 18955
rect 15292 18912 15344 18921
rect 18052 18912 18104 18964
rect 19248 18912 19300 18964
rect 6736 18776 6788 18828
rect 7472 18776 7524 18828
rect 3700 18708 3752 18760
rect 4804 18708 4856 18760
rect 11152 18844 11204 18896
rect 9956 18819 10008 18828
rect 9956 18785 9990 18819
rect 9990 18785 10008 18819
rect 9956 18776 10008 18785
rect 9680 18751 9732 18760
rect 9680 18717 9689 18751
rect 9689 18717 9723 18751
rect 9723 18717 9732 18751
rect 11888 18751 11940 18760
rect 9680 18708 9732 18717
rect 11888 18717 11897 18751
rect 11897 18717 11931 18751
rect 11931 18717 11940 18751
rect 12072 18844 12124 18896
rect 12348 18844 12400 18896
rect 17132 18844 17184 18896
rect 17316 18844 17368 18896
rect 18972 18844 19024 18896
rect 12164 18819 12216 18828
rect 12164 18785 12198 18819
rect 12198 18785 12216 18819
rect 12164 18776 12216 18785
rect 14004 18776 14056 18828
rect 16764 18776 16816 18828
rect 16856 18776 16908 18828
rect 17040 18776 17092 18828
rect 19432 18776 19484 18828
rect 11888 18708 11940 18717
rect 13912 18708 13964 18760
rect 19340 18708 19392 18760
rect 1032 18640 1084 18692
rect 17776 18640 17828 18692
rect 18144 18640 18196 18692
rect 19984 18640 20036 18692
rect 3332 18572 3384 18624
rect 4160 18572 4212 18624
rect 7288 18572 7340 18624
rect 8208 18572 8260 18624
rect 12900 18572 12952 18624
rect 17868 18572 17920 18624
rect 18052 18615 18104 18624
rect 18052 18581 18061 18615
rect 18061 18581 18095 18615
rect 18095 18581 18104 18615
rect 18052 18572 18104 18581
rect 4447 18470 4499 18522
rect 4511 18470 4563 18522
rect 4575 18470 4627 18522
rect 4639 18470 4691 18522
rect 11378 18470 11430 18522
rect 11442 18470 11494 18522
rect 11506 18470 11558 18522
rect 11570 18470 11622 18522
rect 18308 18470 18360 18522
rect 18372 18470 18424 18522
rect 18436 18470 18488 18522
rect 18500 18470 18552 18522
rect 5632 18368 5684 18420
rect 7472 18368 7524 18420
rect 4068 18300 4120 18352
rect 6920 18300 6972 18352
rect 12716 18368 12768 18420
rect 18604 18368 18656 18420
rect 5724 18275 5776 18284
rect 5724 18241 5733 18275
rect 5733 18241 5767 18275
rect 5767 18241 5776 18275
rect 5724 18232 5776 18241
rect 7380 18275 7432 18284
rect 7380 18241 7389 18275
rect 7389 18241 7423 18275
rect 7423 18241 7432 18275
rect 7380 18232 7432 18241
rect 11152 18275 11204 18284
rect 11152 18241 11161 18275
rect 11161 18241 11195 18275
rect 11195 18241 11204 18275
rect 11152 18232 11204 18241
rect 4804 18164 4856 18216
rect 6828 18164 6880 18216
rect 7288 18207 7340 18216
rect 7288 18173 7297 18207
rect 7297 18173 7331 18207
rect 7331 18173 7340 18207
rect 7288 18164 7340 18173
rect 8392 18207 8444 18216
rect 8392 18173 8401 18207
rect 8401 18173 8435 18207
rect 8435 18173 8444 18207
rect 8392 18164 8444 18173
rect 9680 18164 9732 18216
rect 10232 18164 10284 18216
rect 2780 18028 2832 18080
rect 3608 18096 3660 18148
rect 8668 18139 8720 18148
rect 8668 18105 8702 18139
rect 8702 18105 8720 18139
rect 12440 18164 12492 18216
rect 12716 18164 12768 18216
rect 13820 18300 13872 18352
rect 18052 18343 18104 18352
rect 14556 18232 14608 18284
rect 16212 18232 16264 18284
rect 18052 18309 18061 18343
rect 18061 18309 18095 18343
rect 18095 18309 18104 18343
rect 18052 18300 18104 18309
rect 19340 18232 19392 18284
rect 18788 18164 18840 18216
rect 8668 18096 8720 18105
rect 3884 18028 3936 18080
rect 4068 18071 4120 18080
rect 4068 18037 4077 18071
rect 4077 18037 4111 18071
rect 4111 18037 4120 18071
rect 4068 18028 4120 18037
rect 9772 18071 9824 18080
rect 9772 18037 9781 18071
rect 9781 18037 9815 18071
rect 9815 18037 9824 18071
rect 9772 18028 9824 18037
rect 11152 18096 11204 18148
rect 12992 18096 13044 18148
rect 13912 18096 13964 18148
rect 12348 18028 12400 18080
rect 13268 18028 13320 18080
rect 14372 18071 14424 18080
rect 14372 18037 14381 18071
rect 14381 18037 14415 18071
rect 14415 18037 14424 18071
rect 14372 18028 14424 18037
rect 15936 18028 15988 18080
rect 16120 18028 16172 18080
rect 16580 18096 16632 18148
rect 18236 18096 18288 18148
rect 19984 18139 20036 18148
rect 19984 18105 19993 18139
rect 19993 18105 20027 18139
rect 20027 18105 20036 18139
rect 19984 18096 20036 18105
rect 20168 18096 20220 18148
rect 20444 18096 20496 18148
rect 16764 18028 16816 18080
rect 17040 18028 17092 18080
rect 17592 18028 17644 18080
rect 18512 18071 18564 18080
rect 18512 18037 18521 18071
rect 18521 18037 18555 18071
rect 18555 18037 18564 18071
rect 18512 18028 18564 18037
rect 19064 18028 19116 18080
rect 19248 18028 19300 18080
rect 7912 17926 7964 17978
rect 7976 17926 8028 17978
rect 8040 17926 8092 17978
rect 8104 17926 8156 17978
rect 14843 17926 14895 17978
rect 14907 17926 14959 17978
rect 14971 17926 15023 17978
rect 15035 17926 15087 17978
rect 3148 17824 3200 17876
rect 7104 17867 7156 17876
rect 1768 17756 1820 17808
rect 4896 17756 4948 17808
rect 7104 17833 7113 17867
rect 7113 17833 7147 17867
rect 7147 17833 7156 17867
rect 7104 17824 7156 17833
rect 11152 17824 11204 17876
rect 13820 17824 13872 17876
rect 18696 17824 18748 17876
rect 10416 17756 10468 17808
rect 6644 17688 6696 17740
rect 10876 17731 10928 17740
rect 10876 17697 10885 17731
rect 10885 17697 10919 17731
rect 10919 17697 10928 17731
rect 10876 17688 10928 17697
rect 10968 17731 11020 17740
rect 10968 17697 10977 17731
rect 10977 17697 11011 17731
rect 11011 17697 11020 17731
rect 10968 17688 11020 17697
rect 4804 17620 4856 17672
rect 6092 17620 6144 17672
rect 7748 17663 7800 17672
rect 7748 17629 7757 17663
rect 7757 17629 7791 17663
rect 7791 17629 7800 17663
rect 7748 17620 7800 17629
rect 10784 17620 10836 17672
rect 11704 17620 11756 17672
rect 15844 17756 15896 17808
rect 16856 17756 16908 17808
rect 13176 17688 13228 17740
rect 15384 17731 15436 17740
rect 15384 17697 15393 17731
rect 15393 17697 15427 17731
rect 15427 17697 15436 17731
rect 15384 17688 15436 17697
rect 17040 17688 17092 17740
rect 19800 17688 19852 17740
rect 12716 17663 12768 17672
rect 12716 17629 12725 17663
rect 12725 17629 12759 17663
rect 12759 17629 12768 17663
rect 12716 17620 12768 17629
rect 14096 17663 14148 17672
rect 14096 17629 14105 17663
rect 14105 17629 14139 17663
rect 14139 17629 14148 17663
rect 14096 17620 14148 17629
rect 14556 17620 14608 17672
rect 16488 17663 16540 17672
rect 16488 17629 16497 17663
rect 16497 17629 16531 17663
rect 16531 17629 16540 17663
rect 16488 17620 16540 17629
rect 19340 17620 19392 17672
rect 1768 17484 1820 17536
rect 6368 17484 6420 17536
rect 9128 17484 9180 17536
rect 11888 17484 11940 17536
rect 12992 17484 13044 17536
rect 14740 17484 14792 17536
rect 17500 17552 17552 17604
rect 17408 17484 17460 17536
rect 17868 17527 17920 17536
rect 17868 17493 17877 17527
rect 17877 17493 17911 17527
rect 17911 17493 17920 17527
rect 17868 17484 17920 17493
rect 4447 17382 4499 17434
rect 4511 17382 4563 17434
rect 4575 17382 4627 17434
rect 4639 17382 4691 17434
rect 11378 17382 11430 17434
rect 11442 17382 11494 17434
rect 11506 17382 11558 17434
rect 11570 17382 11622 17434
rect 18308 17382 18360 17434
rect 18372 17382 18424 17434
rect 18436 17382 18488 17434
rect 18500 17382 18552 17434
rect 6828 17280 6880 17332
rect 7196 17212 7248 17264
rect 11796 17280 11848 17332
rect 11888 17280 11940 17332
rect 14096 17280 14148 17332
rect 16580 17280 16632 17332
rect 6000 17144 6052 17196
rect 7656 17144 7708 17196
rect 9864 17212 9916 17264
rect 9772 17144 9824 17196
rect 11244 17144 11296 17196
rect 12624 17187 12676 17196
rect 12624 17153 12633 17187
rect 12633 17153 12667 17187
rect 12667 17153 12676 17187
rect 12624 17144 12676 17153
rect 3056 17076 3108 17128
rect 1492 17008 1544 17060
rect 4068 17076 4120 17128
rect 11704 17076 11756 17128
rect 12532 17076 12584 17128
rect 4804 17008 4856 17060
rect 5356 17008 5408 17060
rect 6460 17008 6512 17060
rect 6736 17008 6788 17060
rect 7196 17051 7248 17060
rect 4896 16983 4948 16992
rect 4896 16949 4905 16983
rect 4905 16949 4939 16983
rect 4939 16949 4948 16983
rect 4896 16940 4948 16949
rect 6828 16983 6880 16992
rect 6828 16949 6837 16983
rect 6837 16949 6871 16983
rect 6871 16949 6880 16983
rect 6828 16940 6880 16949
rect 7196 17017 7205 17051
rect 7205 17017 7239 17051
rect 7239 17017 7248 17051
rect 7196 17008 7248 17017
rect 8208 17008 8260 17060
rect 9036 17008 9088 17060
rect 13176 17144 13228 17196
rect 16488 17212 16540 17264
rect 17132 17212 17184 17264
rect 14280 17187 14332 17196
rect 14280 17153 14289 17187
rect 14289 17153 14323 17187
rect 14323 17153 14332 17187
rect 14280 17144 14332 17153
rect 17040 17187 17092 17196
rect 17040 17153 17049 17187
rect 17049 17153 17083 17187
rect 17083 17153 17092 17187
rect 17040 17144 17092 17153
rect 17868 17076 17920 17128
rect 14464 17008 14516 17060
rect 8300 16940 8352 16992
rect 8944 16940 8996 16992
rect 11704 16940 11756 16992
rect 13728 16983 13780 16992
rect 13728 16949 13737 16983
rect 13737 16949 13771 16983
rect 13771 16949 13780 16983
rect 13728 16940 13780 16949
rect 14188 16983 14240 16992
rect 14188 16949 14197 16983
rect 14197 16949 14231 16983
rect 14231 16949 14240 16983
rect 14188 16940 14240 16949
rect 16028 16940 16080 16992
rect 16580 16940 16632 16992
rect 16948 16940 17000 16992
rect 17408 16940 17460 16992
rect 19708 17008 19760 17060
rect 18604 16940 18656 16992
rect 7912 16838 7964 16890
rect 7976 16838 8028 16890
rect 8040 16838 8092 16890
rect 8104 16838 8156 16890
rect 14843 16838 14895 16890
rect 14907 16838 14959 16890
rect 14971 16838 15023 16890
rect 15035 16838 15087 16890
rect 3424 16736 3476 16788
rect 4160 16779 4212 16788
rect 4160 16745 4169 16779
rect 4169 16745 4203 16779
rect 4203 16745 4212 16779
rect 4160 16736 4212 16745
rect 5540 16736 5592 16788
rect 8208 16736 8260 16788
rect 9680 16736 9732 16788
rect 9864 16779 9916 16788
rect 9864 16745 9873 16779
rect 9873 16745 9907 16779
rect 9907 16745 9916 16779
rect 9864 16736 9916 16745
rect 6736 16668 6788 16720
rect 4344 16600 4396 16652
rect 5540 16600 5592 16652
rect 2412 16532 2464 16584
rect 2596 16464 2648 16516
rect 2780 16464 2832 16516
rect 4068 16464 4120 16516
rect 5356 16532 5408 16584
rect 6000 16643 6052 16652
rect 6000 16609 6034 16643
rect 6034 16609 6052 16643
rect 6000 16600 6052 16609
rect 6552 16600 6604 16652
rect 9036 16668 9088 16720
rect 9220 16600 9272 16652
rect 10048 16600 10100 16652
rect 12072 16736 12124 16788
rect 12624 16736 12676 16788
rect 12532 16668 12584 16720
rect 13360 16736 13412 16788
rect 11244 16643 11296 16652
rect 11244 16609 11278 16643
rect 11278 16609 11296 16643
rect 11244 16600 11296 16609
rect 13544 16668 13596 16720
rect 13728 16736 13780 16788
rect 14188 16736 14240 16788
rect 16028 16779 16080 16788
rect 16028 16745 16037 16779
rect 16037 16745 16071 16779
rect 16071 16745 16080 16779
rect 16028 16736 16080 16745
rect 18604 16736 18656 16788
rect 19984 16736 20036 16788
rect 14464 16668 14516 16720
rect 15936 16711 15988 16720
rect 15936 16677 15945 16711
rect 15945 16677 15979 16711
rect 15979 16677 15988 16711
rect 15936 16668 15988 16677
rect 16580 16668 16632 16720
rect 17316 16668 17368 16720
rect 17408 16668 17460 16720
rect 17868 16668 17920 16720
rect 19616 16668 19668 16720
rect 13452 16600 13504 16652
rect 16948 16600 17000 16652
rect 19156 16600 19208 16652
rect 19708 16643 19760 16652
rect 19708 16609 19717 16643
rect 19717 16609 19751 16643
rect 19751 16609 19760 16643
rect 19708 16600 19760 16609
rect 8668 16575 8720 16584
rect 8668 16541 8677 16575
rect 8677 16541 8711 16575
rect 8711 16541 8720 16575
rect 8668 16532 8720 16541
rect 14280 16575 14332 16584
rect 14280 16541 14289 16575
rect 14289 16541 14323 16575
rect 14323 16541 14332 16575
rect 14280 16532 14332 16541
rect 9772 16464 9824 16516
rect 10968 16464 11020 16516
rect 1952 16396 2004 16448
rect 6092 16396 6144 16448
rect 7012 16396 7064 16448
rect 10324 16396 10376 16448
rect 10784 16396 10836 16448
rect 12164 16396 12216 16448
rect 13176 16396 13228 16448
rect 16212 16396 16264 16448
rect 17132 16532 17184 16584
rect 18788 16464 18840 16516
rect 19248 16464 19300 16516
rect 16580 16396 16632 16448
rect 17684 16396 17736 16448
rect 4447 16294 4499 16346
rect 4511 16294 4563 16346
rect 4575 16294 4627 16346
rect 4639 16294 4691 16346
rect 11378 16294 11430 16346
rect 11442 16294 11494 16346
rect 11506 16294 11558 16346
rect 11570 16294 11622 16346
rect 18308 16294 18360 16346
rect 18372 16294 18424 16346
rect 18436 16294 18488 16346
rect 18500 16294 18552 16346
rect 3056 16235 3108 16244
rect 3056 16201 3065 16235
rect 3065 16201 3099 16235
rect 3099 16201 3108 16235
rect 3056 16192 3108 16201
rect 4344 16192 4396 16244
rect 6736 16192 6788 16244
rect 1952 16099 2004 16108
rect 1952 16065 1961 16099
rect 1961 16065 1995 16099
rect 1995 16065 2004 16099
rect 1952 16056 2004 16065
rect 2136 16099 2188 16108
rect 2136 16065 2145 16099
rect 2145 16065 2179 16099
rect 2179 16065 2188 16099
rect 2136 16056 2188 16065
rect 2964 16056 3016 16108
rect 3608 16056 3660 16108
rect 4896 16056 4948 16108
rect 7012 16056 7064 16108
rect 8576 16192 8628 16244
rect 8668 16192 8720 16244
rect 10048 16192 10100 16244
rect 14280 16167 14332 16176
rect 14280 16133 14289 16167
rect 14289 16133 14323 16167
rect 14323 16133 14332 16167
rect 16212 16192 16264 16244
rect 20720 16235 20772 16244
rect 20720 16201 20729 16235
rect 20729 16201 20763 16235
rect 20763 16201 20772 16235
rect 20720 16192 20772 16201
rect 14280 16124 14332 16133
rect 11428 16099 11480 16108
rect 2596 15988 2648 16040
rect 3424 16031 3476 16040
rect 3424 15997 3433 16031
rect 3433 15997 3467 16031
rect 3467 15997 3476 16031
rect 3424 15988 3476 15997
rect 4160 15988 4212 16040
rect 8392 16031 8444 16040
rect 8392 15997 8401 16031
rect 8401 15997 8435 16031
rect 8435 15997 8444 16031
rect 8392 15988 8444 15997
rect 11428 16065 11437 16099
rect 11437 16065 11471 16099
rect 11471 16065 11480 16099
rect 11428 16056 11480 16065
rect 1952 15852 2004 15904
rect 2044 15852 2096 15904
rect 11888 15988 11940 16040
rect 12624 15988 12676 16040
rect 13176 16031 13228 16040
rect 13176 15997 13210 16031
rect 13210 15997 13228 16031
rect 13176 15988 13228 15997
rect 14188 15988 14240 16040
rect 11060 15920 11112 15972
rect 11520 15920 11572 15972
rect 11980 15920 12032 15972
rect 17776 16124 17828 16176
rect 15200 15988 15252 16040
rect 3424 15852 3476 15904
rect 8392 15852 8444 15904
rect 8944 15852 8996 15904
rect 10784 15895 10836 15904
rect 10784 15861 10793 15895
rect 10793 15861 10827 15895
rect 10827 15861 10836 15895
rect 10784 15852 10836 15861
rect 11152 15895 11204 15904
rect 11152 15861 11161 15895
rect 11161 15861 11195 15895
rect 11195 15861 11204 15895
rect 11152 15852 11204 15861
rect 15568 15920 15620 15972
rect 19432 15920 19484 15972
rect 18604 15852 18656 15904
rect 18880 15852 18932 15904
rect 7912 15750 7964 15802
rect 7976 15750 8028 15802
rect 8040 15750 8092 15802
rect 8104 15750 8156 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 15035 15750 15087 15802
rect 2044 15648 2096 15700
rect 2412 15691 2464 15700
rect 2412 15657 2421 15691
rect 2421 15657 2455 15691
rect 2455 15657 2464 15691
rect 2412 15648 2464 15657
rect 1400 15512 1452 15564
rect 2596 15512 2648 15564
rect 4160 15512 4212 15564
rect 5356 15648 5408 15700
rect 5540 15648 5592 15700
rect 6828 15648 6880 15700
rect 8300 15648 8352 15700
rect 9496 15648 9548 15700
rect 9680 15691 9732 15700
rect 9680 15657 9689 15691
rect 9689 15657 9723 15691
rect 9723 15657 9732 15691
rect 9680 15648 9732 15657
rect 10048 15691 10100 15700
rect 10048 15657 10057 15691
rect 10057 15657 10091 15691
rect 10091 15657 10100 15691
rect 10048 15648 10100 15657
rect 10784 15648 10836 15700
rect 15200 15648 15252 15700
rect 15660 15648 15712 15700
rect 17500 15648 17552 15700
rect 19892 15691 19944 15700
rect 19892 15657 19901 15691
rect 19901 15657 19935 15691
rect 19935 15657 19944 15691
rect 19892 15648 19944 15657
rect 2964 15487 3016 15496
rect 2964 15453 2973 15487
rect 2973 15453 3007 15487
rect 3007 15453 3016 15487
rect 4896 15512 4948 15564
rect 6184 15512 6236 15564
rect 6552 15512 6604 15564
rect 6920 15512 6972 15564
rect 7012 15487 7064 15496
rect 2964 15444 3016 15453
rect 1584 15308 1636 15360
rect 7012 15453 7021 15487
rect 7021 15453 7055 15487
rect 7055 15453 7064 15487
rect 7012 15444 7064 15453
rect 8300 15512 8352 15564
rect 8668 15487 8720 15496
rect 8668 15453 8677 15487
rect 8677 15453 8711 15487
rect 8711 15453 8720 15487
rect 8668 15444 8720 15453
rect 11428 15512 11480 15564
rect 6000 15376 6052 15428
rect 8576 15376 8628 15428
rect 12072 15444 12124 15496
rect 12164 15487 12216 15496
rect 12164 15453 12173 15487
rect 12173 15453 12207 15487
rect 12207 15453 12216 15487
rect 12532 15512 12584 15564
rect 13544 15555 13596 15564
rect 13544 15521 13553 15555
rect 13553 15521 13587 15555
rect 13587 15521 13596 15555
rect 18052 15555 18104 15564
rect 13544 15512 13596 15521
rect 18052 15521 18061 15555
rect 18061 15521 18095 15555
rect 18095 15521 18104 15555
rect 18052 15512 18104 15521
rect 19800 15512 19852 15564
rect 12164 15444 12216 15453
rect 16396 15444 16448 15496
rect 16580 15444 16632 15496
rect 18144 15487 18196 15496
rect 18144 15453 18153 15487
rect 18153 15453 18187 15487
rect 18187 15453 18196 15487
rect 18144 15444 18196 15453
rect 10416 15376 10468 15428
rect 13452 15376 13504 15428
rect 15568 15308 15620 15360
rect 15660 15308 15712 15360
rect 17408 15376 17460 15428
rect 18328 15376 18380 15428
rect 19340 15376 19392 15428
rect 18052 15308 18104 15360
rect 4447 15206 4499 15258
rect 4511 15206 4563 15258
rect 4575 15206 4627 15258
rect 4639 15206 4691 15258
rect 11378 15206 11430 15258
rect 11442 15206 11494 15258
rect 11506 15206 11558 15258
rect 11570 15206 11622 15258
rect 18308 15206 18360 15258
rect 18372 15206 18424 15258
rect 18436 15206 18488 15258
rect 18500 15206 18552 15258
rect 10416 15147 10468 15156
rect 10416 15113 10425 15147
rect 10425 15113 10459 15147
rect 10459 15113 10468 15147
rect 10416 15104 10468 15113
rect 12256 15104 12308 15156
rect 2872 15036 2924 15088
rect 10508 15036 10560 15088
rect 18696 15104 18748 15156
rect 20720 15147 20772 15156
rect 20720 15113 20729 15147
rect 20729 15113 20763 15147
rect 20763 15113 20772 15147
rect 20720 15104 20772 15113
rect 12440 15036 12492 15088
rect 13084 15036 13136 15088
rect 2136 14968 2188 15020
rect 8484 14968 8536 15020
rect 10140 14968 10192 15020
rect 10416 14968 10468 15020
rect 3332 14900 3384 14952
rect 5356 14900 5408 14952
rect 10048 14900 10100 14952
rect 10600 14900 10652 14952
rect 15292 14943 15344 14952
rect 15292 14909 15301 14943
rect 15301 14909 15335 14943
rect 15335 14909 15344 14943
rect 15292 14900 15344 14909
rect 2228 14832 2280 14884
rect 3056 14764 3108 14816
rect 3976 14832 4028 14884
rect 6920 14832 6972 14884
rect 7196 14832 7248 14884
rect 12440 14832 12492 14884
rect 4896 14807 4948 14816
rect 4896 14773 4905 14807
rect 4905 14773 4939 14807
rect 4939 14773 4948 14807
rect 4896 14764 4948 14773
rect 7748 14764 7800 14816
rect 8208 14807 8260 14816
rect 8208 14773 8217 14807
rect 8217 14773 8251 14807
rect 8251 14773 8260 14807
rect 8208 14764 8260 14773
rect 9956 14764 10008 14816
rect 12532 14764 12584 14816
rect 14556 14832 14608 14884
rect 19248 14900 19300 14952
rect 17500 14832 17552 14884
rect 16120 14764 16172 14816
rect 16488 14764 16540 14816
rect 18696 14764 18748 14816
rect 19248 14807 19300 14816
rect 19248 14773 19257 14807
rect 19257 14773 19291 14807
rect 19291 14773 19300 14807
rect 19248 14764 19300 14773
rect 7912 14662 7964 14714
rect 7976 14662 8028 14714
rect 8040 14662 8092 14714
rect 8104 14662 8156 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 15035 14662 15087 14714
rect 3424 14560 3476 14612
rect 7196 14603 7248 14612
rect 7196 14569 7205 14603
rect 7205 14569 7239 14603
rect 7239 14569 7248 14603
rect 7196 14560 7248 14569
rect 7656 14560 7708 14612
rect 8300 14560 8352 14612
rect 9864 14603 9916 14612
rect 9864 14569 9873 14603
rect 9873 14569 9907 14603
rect 9907 14569 9916 14603
rect 9864 14560 9916 14569
rect 12440 14603 12492 14612
rect 12440 14569 12449 14603
rect 12449 14569 12483 14603
rect 12483 14569 12492 14603
rect 12440 14560 12492 14569
rect 14648 14560 14700 14612
rect 15384 14560 15436 14612
rect 16212 14560 16264 14612
rect 19248 14560 19300 14612
rect 19616 14560 19668 14612
rect 3148 14424 3200 14476
rect 3516 14424 3568 14476
rect 4804 14424 4856 14476
rect 6368 14424 6420 14476
rect 7748 14424 7800 14476
rect 16672 14492 16724 14544
rect 9312 14424 9364 14476
rect 11336 14467 11388 14476
rect 11336 14433 11370 14467
rect 11370 14433 11388 14467
rect 11336 14424 11388 14433
rect 13820 14424 13872 14476
rect 15292 14467 15344 14476
rect 15292 14433 15301 14467
rect 15301 14433 15335 14467
rect 15335 14433 15344 14467
rect 15292 14424 15344 14433
rect 17132 14424 17184 14476
rect 19432 14492 19484 14544
rect 19340 14424 19392 14476
rect 2136 14356 2188 14408
rect 3700 14356 3752 14408
rect 4160 14356 4212 14408
rect 3976 14288 4028 14340
rect 5356 14356 5408 14408
rect 2412 14263 2464 14272
rect 2412 14229 2421 14263
rect 2421 14229 2455 14263
rect 2455 14229 2464 14263
rect 2412 14220 2464 14229
rect 4068 14263 4120 14272
rect 4068 14229 4077 14263
rect 4077 14229 4111 14263
rect 4111 14229 4120 14263
rect 4068 14220 4120 14229
rect 6920 14356 6972 14408
rect 8576 14399 8628 14408
rect 8576 14365 8585 14399
rect 8585 14365 8619 14399
rect 8619 14365 8628 14399
rect 8576 14356 8628 14365
rect 6552 14220 6604 14272
rect 12164 14356 12216 14408
rect 12624 14356 12676 14408
rect 12900 14356 12952 14408
rect 13268 14356 13320 14408
rect 12164 14220 12216 14272
rect 12624 14220 12676 14272
rect 13452 14220 13504 14272
rect 19432 14356 19484 14408
rect 19340 14288 19392 14340
rect 16028 14220 16080 14272
rect 18604 14263 18656 14272
rect 18604 14229 18613 14263
rect 18613 14229 18647 14263
rect 18647 14229 18656 14263
rect 18604 14220 18656 14229
rect 4447 14118 4499 14170
rect 4511 14118 4563 14170
rect 4575 14118 4627 14170
rect 4639 14118 4691 14170
rect 11378 14118 11430 14170
rect 11442 14118 11494 14170
rect 11506 14118 11558 14170
rect 11570 14118 11622 14170
rect 18308 14118 18360 14170
rect 18372 14118 18424 14170
rect 18436 14118 18488 14170
rect 18500 14118 18552 14170
rect 1676 14059 1728 14068
rect 1676 14025 1685 14059
rect 1685 14025 1719 14059
rect 1719 14025 1728 14059
rect 1676 14016 1728 14025
rect 3332 14016 3384 14068
rect 4804 14059 4856 14068
rect 4804 14025 4813 14059
rect 4813 14025 4847 14059
rect 4847 14025 4856 14059
rect 4804 14016 4856 14025
rect 6368 14016 6420 14068
rect 6276 13948 6328 14000
rect 1492 13855 1544 13864
rect 1492 13821 1501 13855
rect 1501 13821 1535 13855
rect 1535 13821 1544 13855
rect 1492 13812 1544 13821
rect 8208 13880 8260 13932
rect 5264 13855 5316 13864
rect 5264 13821 5273 13855
rect 5273 13821 5307 13855
rect 5307 13821 5316 13855
rect 5264 13812 5316 13821
rect 7748 13812 7800 13864
rect 8944 14016 8996 14068
rect 9404 13880 9456 13932
rect 13728 14016 13780 14068
rect 17500 14016 17552 14068
rect 18144 14016 18196 14068
rect 11520 13991 11572 14000
rect 11520 13957 11529 13991
rect 11529 13957 11563 13991
rect 11563 13957 11572 13991
rect 11520 13948 11572 13957
rect 12900 13948 12952 14000
rect 16120 13948 16172 14000
rect 12440 13880 12492 13932
rect 14556 13923 14608 13932
rect 14556 13889 14565 13923
rect 14565 13889 14599 13923
rect 14599 13889 14608 13923
rect 14556 13880 14608 13889
rect 16212 13880 16264 13932
rect 16672 13880 16724 13932
rect 18696 13923 18748 13932
rect 18696 13889 18705 13923
rect 18705 13889 18739 13923
rect 18739 13889 18748 13923
rect 18696 13880 18748 13889
rect 2964 13744 3016 13796
rect 6920 13744 6972 13796
rect 7564 13744 7616 13796
rect 8208 13744 8260 13796
rect 8760 13787 8812 13796
rect 8760 13753 8769 13787
rect 8769 13753 8803 13787
rect 8803 13753 8812 13787
rect 8760 13744 8812 13753
rect 9128 13744 9180 13796
rect 3332 13676 3384 13728
rect 3976 13719 4028 13728
rect 3976 13685 3985 13719
rect 3985 13685 4019 13719
rect 4019 13685 4028 13719
rect 3976 13676 4028 13685
rect 4988 13676 5040 13728
rect 6552 13676 6604 13728
rect 6644 13676 6696 13728
rect 7196 13719 7248 13728
rect 7196 13685 7205 13719
rect 7205 13685 7239 13719
rect 7239 13685 7248 13719
rect 7196 13676 7248 13685
rect 7288 13719 7340 13728
rect 7288 13685 7297 13719
rect 7297 13685 7331 13719
rect 7331 13685 7340 13719
rect 8392 13719 8444 13728
rect 7288 13676 7340 13685
rect 8392 13685 8401 13719
rect 8401 13685 8435 13719
rect 8435 13685 8444 13719
rect 8392 13676 8444 13685
rect 8944 13676 8996 13728
rect 13912 13812 13964 13864
rect 15292 13812 15344 13864
rect 17960 13812 18012 13864
rect 19248 13812 19300 13864
rect 19984 13812 20036 13864
rect 20352 13812 20404 13864
rect 10600 13744 10652 13796
rect 10784 13744 10836 13796
rect 16212 13744 16264 13796
rect 18788 13744 18840 13796
rect 12808 13719 12860 13728
rect 12808 13685 12817 13719
rect 12817 13685 12851 13719
rect 12851 13685 12860 13719
rect 12808 13676 12860 13685
rect 12900 13719 12952 13728
rect 12900 13685 12909 13719
rect 12909 13685 12943 13719
rect 12943 13685 12952 13719
rect 15936 13719 15988 13728
rect 12900 13676 12952 13685
rect 15936 13685 15945 13719
rect 15945 13685 15979 13719
rect 15979 13685 15988 13719
rect 15936 13676 15988 13685
rect 20720 13719 20772 13728
rect 20720 13685 20729 13719
rect 20729 13685 20763 13719
rect 20763 13685 20772 13719
rect 20720 13676 20772 13685
rect 7912 13574 7964 13626
rect 7976 13574 8028 13626
rect 8040 13574 8092 13626
rect 8104 13574 8156 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 15035 13574 15087 13626
rect 4068 13472 4120 13524
rect 6920 13472 6972 13524
rect 7288 13472 7340 13524
rect 8392 13472 8444 13524
rect 8484 13472 8536 13524
rect 8668 13515 8720 13524
rect 8668 13481 8677 13515
rect 8677 13481 8711 13515
rect 8711 13481 8720 13515
rect 8668 13472 8720 13481
rect 9404 13472 9456 13524
rect 9496 13472 9548 13524
rect 11152 13472 11204 13524
rect 12808 13472 12860 13524
rect 12992 13472 13044 13524
rect 13360 13472 13412 13524
rect 15292 13515 15344 13524
rect 15292 13481 15301 13515
rect 15301 13481 15335 13515
rect 15335 13481 15344 13515
rect 15292 13472 15344 13481
rect 15936 13472 15988 13524
rect 2320 13336 2372 13388
rect 4896 13404 4948 13456
rect 5356 13404 5408 13456
rect 12624 13447 12676 13456
rect 12624 13413 12633 13447
rect 12633 13413 12667 13447
rect 12667 13413 12676 13447
rect 12624 13404 12676 13413
rect 19156 13472 19208 13524
rect 17868 13404 17920 13456
rect 5816 13336 5868 13388
rect 6552 13336 6604 13388
rect 7748 13336 7800 13388
rect 12900 13336 12952 13388
rect 13912 13379 13964 13388
rect 13912 13345 13921 13379
rect 13921 13345 13955 13379
rect 13955 13345 13964 13379
rect 13912 13336 13964 13345
rect 15936 13336 15988 13388
rect 18052 13336 18104 13388
rect 19248 13379 19300 13388
rect 19248 13345 19257 13379
rect 19257 13345 19291 13379
rect 19291 13345 19300 13379
rect 19248 13336 19300 13345
rect 3884 13268 3936 13320
rect 6092 13268 6144 13320
rect 6368 13268 6420 13320
rect 7656 13311 7708 13320
rect 7656 13277 7665 13311
rect 7665 13277 7699 13311
rect 7699 13277 7708 13311
rect 7656 13268 7708 13277
rect 8576 13268 8628 13320
rect 9588 13268 9640 13320
rect 12440 13268 12492 13320
rect 11520 13200 11572 13252
rect 14556 13268 14608 13320
rect 16028 13268 16080 13320
rect 17500 13268 17552 13320
rect 17776 13311 17828 13320
rect 17776 13277 17785 13311
rect 17785 13277 17819 13311
rect 17819 13277 17828 13311
rect 17776 13268 17828 13277
rect 17960 13311 18012 13320
rect 17960 13277 17969 13311
rect 17969 13277 18003 13311
rect 18003 13277 18012 13311
rect 17960 13268 18012 13277
rect 18788 13200 18840 13252
rect 7012 13132 7064 13184
rect 11796 13132 11848 13184
rect 15108 13132 15160 13184
rect 15384 13132 15436 13184
rect 18696 13132 18748 13184
rect 4447 13030 4499 13082
rect 4511 13030 4563 13082
rect 4575 13030 4627 13082
rect 4639 13030 4691 13082
rect 11378 13030 11430 13082
rect 11442 13030 11494 13082
rect 11506 13030 11558 13082
rect 11570 13030 11622 13082
rect 18308 13030 18360 13082
rect 18372 13030 18424 13082
rect 18436 13030 18488 13082
rect 18500 13030 18552 13082
rect 2320 12971 2372 12980
rect 2320 12937 2329 12971
rect 2329 12937 2363 12971
rect 2363 12937 2372 12971
rect 2320 12928 2372 12937
rect 3148 12928 3200 12980
rect 4988 12971 5040 12980
rect 4988 12937 4997 12971
rect 4997 12937 5031 12971
rect 5031 12937 5040 12971
rect 4988 12928 5040 12937
rect 7196 12928 7248 12980
rect 7748 12928 7800 12980
rect 9220 12971 9272 12980
rect 9220 12937 9229 12971
rect 9229 12937 9263 12971
rect 9263 12937 9272 12971
rect 9220 12928 9272 12937
rect 10784 12971 10836 12980
rect 10784 12937 10793 12971
rect 10793 12937 10827 12971
rect 10827 12937 10836 12971
rect 10784 12928 10836 12937
rect 11796 12928 11848 12980
rect 11980 12928 12032 12980
rect 12440 12971 12492 12980
rect 12440 12937 12449 12971
rect 12449 12937 12483 12971
rect 12483 12937 12492 12971
rect 12440 12928 12492 12937
rect 12716 12928 12768 12980
rect 13728 12928 13780 12980
rect 13820 12928 13872 12980
rect 15936 12971 15988 12980
rect 15936 12937 15945 12971
rect 15945 12937 15979 12971
rect 15979 12937 15988 12971
rect 15936 12928 15988 12937
rect 17316 12928 17368 12980
rect 18604 12928 18656 12980
rect 10600 12860 10652 12912
rect 3332 12792 3384 12844
rect 5632 12835 5684 12844
rect 5632 12801 5641 12835
rect 5641 12801 5675 12835
rect 5675 12801 5684 12835
rect 5632 12792 5684 12801
rect 7656 12792 7708 12844
rect 3148 12724 3200 12776
rect 3424 12724 3476 12776
rect 9036 12724 9088 12776
rect 9588 12792 9640 12844
rect 10140 12724 10192 12776
rect 2504 12656 2556 12708
rect 4068 12656 4120 12708
rect 8484 12656 8536 12708
rect 9312 12656 9364 12708
rect 12716 12792 12768 12844
rect 12900 12835 12952 12844
rect 12900 12801 12909 12835
rect 12909 12801 12943 12835
rect 12943 12801 12952 12835
rect 12900 12792 12952 12801
rect 13084 12860 13136 12912
rect 13452 12792 13504 12844
rect 14556 12792 14608 12844
rect 16672 12792 16724 12844
rect 17132 12792 17184 12844
rect 12624 12724 12676 12776
rect 12992 12656 13044 12708
rect 2688 12631 2740 12640
rect 2688 12597 2697 12631
rect 2697 12597 2731 12631
rect 2731 12597 2740 12631
rect 2688 12588 2740 12597
rect 4896 12588 4948 12640
rect 5356 12631 5408 12640
rect 5356 12597 5365 12631
rect 5365 12597 5399 12631
rect 5399 12597 5408 12631
rect 5356 12588 5408 12597
rect 6368 12588 6420 12640
rect 7104 12588 7156 12640
rect 7288 12631 7340 12640
rect 7288 12597 7297 12631
rect 7297 12597 7331 12631
rect 7331 12597 7340 12631
rect 7288 12588 7340 12597
rect 9220 12588 9272 12640
rect 12164 12588 12216 12640
rect 12900 12588 12952 12640
rect 13820 12588 13872 12640
rect 15200 12724 15252 12776
rect 15844 12724 15896 12776
rect 17592 12724 17644 12776
rect 16764 12656 16816 12708
rect 17684 12656 17736 12708
rect 19064 12699 19116 12708
rect 19064 12665 19098 12699
rect 19098 12665 19116 12699
rect 19064 12656 19116 12665
rect 17316 12588 17368 12640
rect 17500 12588 17552 12640
rect 17776 12588 17828 12640
rect 18144 12588 18196 12640
rect 18788 12588 18840 12640
rect 7912 12486 7964 12538
rect 7976 12486 8028 12538
rect 8040 12486 8092 12538
rect 8104 12486 8156 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 15035 12486 15087 12538
rect 2412 12384 2464 12436
rect 5540 12384 5592 12436
rect 6920 12384 6972 12436
rect 7012 12384 7064 12436
rect 3884 12316 3936 12368
rect 11244 12384 11296 12436
rect 12532 12384 12584 12436
rect 13544 12384 13596 12436
rect 14740 12384 14792 12436
rect 16580 12384 16632 12436
rect 17868 12384 17920 12436
rect 19892 12427 19944 12436
rect 19892 12393 19901 12427
rect 19901 12393 19935 12427
rect 19935 12393 19944 12427
rect 19892 12384 19944 12393
rect 7656 12316 7708 12368
rect 11980 12316 12032 12368
rect 13360 12316 13412 12368
rect 14372 12316 14424 12368
rect 18972 12316 19024 12368
rect 19984 12316 20036 12368
rect 6092 12248 6144 12300
rect 6736 12248 6788 12300
rect 2964 12180 3016 12232
rect 5172 12180 5224 12232
rect 2688 12112 2740 12164
rect 4068 12112 4120 12164
rect 2320 12044 2372 12096
rect 5448 12112 5500 12164
rect 7012 12180 7064 12232
rect 7104 12112 7156 12164
rect 7196 12112 7248 12164
rect 9956 12248 10008 12300
rect 7748 12180 7800 12232
rect 10692 12180 10744 12232
rect 14188 12248 14240 12300
rect 14556 12248 14608 12300
rect 17132 12291 17184 12300
rect 17132 12257 17141 12291
rect 17141 12257 17175 12291
rect 17175 12257 17184 12291
rect 17132 12248 17184 12257
rect 17224 12248 17276 12300
rect 19708 12291 19760 12300
rect 19708 12257 19717 12291
rect 19717 12257 19751 12291
rect 19751 12257 19760 12291
rect 19708 12248 19760 12257
rect 14004 12223 14056 12232
rect 14004 12189 14013 12223
rect 14013 12189 14047 12223
rect 14047 12189 14056 12223
rect 14004 12180 14056 12189
rect 16120 12180 16172 12232
rect 8392 12044 8444 12096
rect 10508 12044 10560 12096
rect 12532 12044 12584 12096
rect 12624 12044 12676 12096
rect 12808 12044 12860 12096
rect 13912 12112 13964 12164
rect 14096 12044 14148 12096
rect 16304 12044 16356 12096
rect 18052 12044 18104 12096
rect 19064 12044 19116 12096
rect 4447 11942 4499 11994
rect 4511 11942 4563 11994
rect 4575 11942 4627 11994
rect 4639 11942 4691 11994
rect 11378 11942 11430 11994
rect 11442 11942 11494 11994
rect 11506 11942 11558 11994
rect 11570 11942 11622 11994
rect 18308 11942 18360 11994
rect 18372 11942 18424 11994
rect 18436 11942 18488 11994
rect 18500 11942 18552 11994
rect 2412 11840 2464 11892
rect 5264 11840 5316 11892
rect 7288 11840 7340 11892
rect 4160 11772 4212 11824
rect 10600 11840 10652 11892
rect 12440 11840 12492 11892
rect 12624 11772 12676 11824
rect 2320 11747 2372 11756
rect 2320 11713 2329 11747
rect 2329 11713 2363 11747
rect 2363 11713 2372 11747
rect 2320 11704 2372 11713
rect 2964 11704 3016 11756
rect 3700 11704 3752 11756
rect 5448 11704 5500 11756
rect 6736 11704 6788 11756
rect 8668 11704 8720 11756
rect 10876 11704 10928 11756
rect 14188 11840 14240 11892
rect 16580 11840 16632 11892
rect 19248 11840 19300 11892
rect 12900 11704 12952 11756
rect 1952 11636 2004 11688
rect 2872 11636 2924 11688
rect 3792 11636 3844 11688
rect 9772 11636 9824 11688
rect 10324 11636 10376 11688
rect 10968 11636 11020 11688
rect 16488 11636 16540 11688
rect 17960 11704 18012 11756
rect 19064 11704 19116 11756
rect 19432 11636 19484 11688
rect 2412 11568 2464 11620
rect 4344 11568 4396 11620
rect 4988 11568 5040 11620
rect 8208 11568 8260 11620
rect 4160 11500 4212 11552
rect 4252 11500 4304 11552
rect 4896 11500 4948 11552
rect 6368 11500 6420 11552
rect 11704 11500 11756 11552
rect 13912 11568 13964 11620
rect 16948 11568 17000 11620
rect 18052 11568 18104 11620
rect 16396 11500 16448 11552
rect 16672 11500 16724 11552
rect 19432 11543 19484 11552
rect 19432 11509 19441 11543
rect 19441 11509 19475 11543
rect 19475 11509 19484 11543
rect 19432 11500 19484 11509
rect 7912 11398 7964 11450
rect 7976 11398 8028 11450
rect 8040 11398 8092 11450
rect 8104 11398 8156 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 15035 11398 15087 11450
rect 2504 11296 2556 11348
rect 2780 11339 2832 11348
rect 2780 11305 2789 11339
rect 2789 11305 2823 11339
rect 2823 11305 2832 11339
rect 2780 11296 2832 11305
rect 3424 11296 3476 11348
rect 4068 11296 4120 11348
rect 5448 11296 5500 11348
rect 12440 11296 12492 11348
rect 12900 11296 12952 11348
rect 14004 11296 14056 11348
rect 14096 11339 14148 11348
rect 14096 11305 14105 11339
rect 14105 11305 14139 11339
rect 14139 11305 14148 11339
rect 14096 11296 14148 11305
rect 17224 11296 17276 11348
rect 18144 11296 18196 11348
rect 2872 11271 2924 11280
rect 2872 11237 2881 11271
rect 2881 11237 2915 11271
rect 2915 11237 2924 11271
rect 2872 11228 2924 11237
rect 7012 11228 7064 11280
rect 7564 11228 7616 11280
rect 10416 11271 10468 11280
rect 10416 11237 10425 11271
rect 10425 11237 10459 11271
rect 10459 11237 10468 11271
rect 10416 11228 10468 11237
rect 11704 11228 11756 11280
rect 12072 11228 12124 11280
rect 12624 11228 12676 11280
rect 15752 11228 15804 11280
rect 3424 11160 3476 11212
rect 5172 11160 5224 11212
rect 6644 11160 6696 11212
rect 15476 11160 15528 11212
rect 2964 11135 3016 11144
rect 2964 11101 2973 11135
rect 2973 11101 3007 11135
rect 3007 11101 3016 11135
rect 2964 11092 3016 11101
rect 5816 11135 5868 11144
rect 5816 11101 5825 11135
rect 5825 11101 5859 11135
rect 5859 11101 5868 11135
rect 5816 11092 5868 11101
rect 6000 11135 6052 11144
rect 6000 11101 6009 11135
rect 6009 11101 6043 11135
rect 6043 11101 6052 11135
rect 6000 11092 6052 11101
rect 12256 11135 12308 11144
rect 12256 11101 12265 11135
rect 12265 11101 12299 11135
rect 12299 11101 12308 11135
rect 12256 11092 12308 11101
rect 13820 11092 13872 11144
rect 14280 11135 14332 11144
rect 14280 11101 14289 11135
rect 14289 11101 14323 11135
rect 14323 11101 14332 11135
rect 14280 11092 14332 11101
rect 15292 11092 15344 11144
rect 17132 11160 17184 11212
rect 19708 11228 19760 11280
rect 3884 11024 3936 11076
rect 5540 11024 5592 11076
rect 10232 11024 10284 11076
rect 10968 11024 11020 11076
rect 4252 10956 4304 11008
rect 6920 10956 6972 11008
rect 13728 10999 13780 11008
rect 13728 10965 13737 10999
rect 13737 10965 13771 10999
rect 13771 10965 13780 10999
rect 18144 11024 18196 11076
rect 13728 10956 13780 10965
rect 14556 10956 14608 11008
rect 17776 10999 17828 11008
rect 17776 10965 17785 10999
rect 17785 10965 17819 10999
rect 17819 10965 17828 10999
rect 17776 10956 17828 10965
rect 4447 10854 4499 10906
rect 4511 10854 4563 10906
rect 4575 10854 4627 10906
rect 4639 10854 4691 10906
rect 11378 10854 11430 10906
rect 11442 10854 11494 10906
rect 11506 10854 11558 10906
rect 11570 10854 11622 10906
rect 18308 10854 18360 10906
rect 18372 10854 18424 10906
rect 18436 10854 18488 10906
rect 18500 10854 18552 10906
rect 3884 10684 3936 10736
rect 7564 10752 7616 10804
rect 8576 10752 8628 10804
rect 12624 10752 12676 10804
rect 5908 10684 5960 10736
rect 6460 10684 6512 10736
rect 7840 10684 7892 10736
rect 11060 10684 11112 10736
rect 9956 10616 10008 10668
rect 10600 10616 10652 10668
rect 11704 10616 11756 10668
rect 13728 10659 13780 10668
rect 13728 10625 13737 10659
rect 13737 10625 13771 10659
rect 13771 10625 13780 10659
rect 13728 10616 13780 10625
rect 13912 10659 13964 10668
rect 13912 10625 13921 10659
rect 13921 10625 13955 10659
rect 13955 10625 13964 10659
rect 13912 10616 13964 10625
rect 15200 10616 15252 10668
rect 2872 10591 2924 10600
rect 2872 10557 2881 10591
rect 2881 10557 2915 10591
rect 2915 10557 2924 10591
rect 2872 10548 2924 10557
rect 3700 10548 3752 10600
rect 5540 10591 5592 10600
rect 5540 10557 5549 10591
rect 5549 10557 5583 10591
rect 5583 10557 5592 10591
rect 5540 10548 5592 10557
rect 6460 10548 6512 10600
rect 10232 10548 10284 10600
rect 11152 10548 11204 10600
rect 14740 10548 14792 10600
rect 17224 10616 17276 10668
rect 18880 10752 18932 10804
rect 18236 10684 18288 10736
rect 18788 10684 18840 10736
rect 19340 10616 19392 10668
rect 15476 10548 15528 10600
rect 17776 10548 17828 10600
rect 19156 10548 19208 10600
rect 2228 10480 2280 10532
rect 4068 10480 4120 10532
rect 5632 10455 5684 10464
rect 5632 10421 5641 10455
rect 5641 10421 5675 10455
rect 5675 10421 5684 10455
rect 5632 10412 5684 10421
rect 7380 10480 7432 10532
rect 10876 10480 10928 10532
rect 16856 10480 16908 10532
rect 8852 10412 8904 10464
rect 9036 10455 9088 10464
rect 9036 10421 9045 10455
rect 9045 10421 9079 10455
rect 9079 10421 9088 10455
rect 9036 10412 9088 10421
rect 9680 10412 9732 10464
rect 9864 10455 9916 10464
rect 9864 10421 9873 10455
rect 9873 10421 9907 10455
rect 9907 10421 9916 10455
rect 9864 10412 9916 10421
rect 10416 10412 10468 10464
rect 11428 10455 11480 10464
rect 11428 10421 11437 10455
rect 11437 10421 11471 10455
rect 11471 10421 11480 10455
rect 11428 10412 11480 10421
rect 13636 10455 13688 10464
rect 13636 10421 13645 10455
rect 13645 10421 13679 10455
rect 13679 10421 13688 10455
rect 13636 10412 13688 10421
rect 17224 10412 17276 10464
rect 19340 10480 19392 10532
rect 18052 10412 18104 10464
rect 20812 10455 20864 10464
rect 20812 10421 20821 10455
rect 20821 10421 20855 10455
rect 20855 10421 20864 10455
rect 20812 10412 20864 10421
rect 7912 10310 7964 10362
rect 7976 10310 8028 10362
rect 8040 10310 8092 10362
rect 8104 10310 8156 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 15035 10310 15087 10362
rect 3056 10208 3108 10260
rect 5816 10208 5868 10260
rect 8484 10251 8536 10260
rect 8484 10217 8493 10251
rect 8493 10217 8527 10251
rect 8527 10217 8536 10251
rect 8484 10208 8536 10217
rect 13636 10208 13688 10260
rect 15844 10251 15896 10260
rect 7104 10183 7156 10192
rect 7104 10149 7113 10183
rect 7113 10149 7147 10183
rect 7147 10149 7156 10183
rect 7104 10140 7156 10149
rect 7288 10140 7340 10192
rect 1952 10072 2004 10124
rect 2872 10072 2924 10124
rect 3884 10072 3936 10124
rect 5724 10072 5776 10124
rect 7012 10072 7064 10124
rect 9772 10072 9824 10124
rect 9956 10115 10008 10124
rect 9956 10081 9990 10115
rect 9990 10081 10008 10115
rect 9956 10072 10008 10081
rect 13084 10072 13136 10124
rect 14004 10183 14056 10192
rect 14004 10149 14013 10183
rect 14013 10149 14047 10183
rect 14047 10149 14056 10183
rect 14004 10140 14056 10149
rect 15108 10072 15160 10124
rect 4344 10004 4396 10056
rect 6092 10004 6144 10056
rect 6644 10004 6696 10056
rect 12532 10047 12584 10056
rect 6000 9936 6052 9988
rect 7380 9936 7432 9988
rect 2044 9911 2096 9920
rect 2044 9877 2053 9911
rect 2053 9877 2087 9911
rect 2087 9877 2096 9911
rect 2044 9868 2096 9877
rect 5724 9868 5776 9920
rect 6552 9868 6604 9920
rect 12532 10013 12541 10047
rect 12541 10013 12575 10047
rect 12575 10013 12584 10047
rect 12532 10004 12584 10013
rect 14188 10047 14240 10056
rect 13820 9936 13872 9988
rect 14188 10013 14197 10047
rect 14197 10013 14231 10047
rect 14231 10013 14240 10047
rect 14188 10004 14240 10013
rect 15844 10217 15853 10251
rect 15853 10217 15887 10251
rect 15887 10217 15896 10251
rect 15844 10208 15896 10217
rect 16764 10208 16816 10260
rect 17592 10208 17644 10260
rect 18144 10208 18196 10260
rect 19248 10208 19300 10260
rect 15292 10140 15344 10192
rect 15476 10140 15528 10192
rect 15568 10072 15620 10124
rect 16764 10072 16816 10124
rect 19156 10140 19208 10192
rect 17776 10072 17828 10124
rect 19616 10115 19668 10124
rect 19616 10081 19625 10115
rect 19625 10081 19659 10115
rect 19659 10081 19668 10115
rect 19616 10072 19668 10081
rect 16028 10047 16080 10056
rect 16028 10013 16037 10047
rect 16037 10013 16071 10047
rect 16071 10013 16080 10047
rect 16028 10004 16080 10013
rect 20628 10004 20680 10056
rect 14280 9936 14332 9988
rect 14556 9936 14608 9988
rect 11060 9911 11112 9920
rect 11060 9877 11069 9911
rect 11069 9877 11103 9911
rect 11103 9877 11112 9911
rect 11060 9868 11112 9877
rect 16764 9868 16816 9920
rect 17960 9936 18012 9988
rect 20444 9936 20496 9988
rect 17868 9868 17920 9920
rect 20536 9868 20588 9920
rect 4447 9766 4499 9818
rect 4511 9766 4563 9818
rect 4575 9766 4627 9818
rect 4639 9766 4691 9818
rect 11378 9766 11430 9818
rect 11442 9766 11494 9818
rect 11506 9766 11558 9818
rect 11570 9766 11622 9818
rect 18308 9766 18360 9818
rect 18372 9766 18424 9818
rect 18436 9766 18488 9818
rect 18500 9766 18552 9818
rect 3240 9664 3292 9716
rect 4068 9664 4120 9716
rect 5172 9639 5224 9648
rect 5172 9605 5181 9639
rect 5181 9605 5215 9639
rect 5215 9605 5224 9639
rect 5172 9596 5224 9605
rect 5632 9664 5684 9716
rect 12440 9664 12492 9716
rect 9588 9596 9640 9648
rect 11244 9596 11296 9648
rect 13544 9664 13596 9716
rect 19616 9664 19668 9716
rect 20168 9664 20220 9716
rect 20444 9664 20496 9716
rect 13820 9639 13872 9648
rect 2872 9528 2924 9580
rect 3700 9528 3752 9580
rect 5448 9528 5500 9580
rect 5724 9571 5776 9580
rect 5724 9537 5733 9571
rect 5733 9537 5767 9571
rect 5767 9537 5776 9571
rect 5724 9528 5776 9537
rect 7380 9571 7432 9580
rect 7380 9537 7389 9571
rect 7389 9537 7423 9571
rect 7423 9537 7432 9571
rect 7380 9528 7432 9537
rect 10232 9571 10284 9580
rect 10232 9537 10241 9571
rect 10241 9537 10275 9571
rect 10275 9537 10284 9571
rect 10232 9528 10284 9537
rect 11060 9528 11112 9580
rect 13820 9605 13829 9639
rect 13829 9605 13863 9639
rect 13863 9605 13872 9639
rect 13820 9596 13872 9605
rect 14280 9596 14332 9648
rect 14372 9528 14424 9580
rect 14556 9528 14608 9580
rect 15292 9571 15344 9580
rect 15292 9537 15301 9571
rect 15301 9537 15335 9571
rect 15335 9537 15344 9571
rect 15292 9528 15344 9537
rect 16028 9596 16080 9648
rect 2044 9460 2096 9512
rect 4252 9460 4304 9512
rect 3700 9392 3752 9444
rect 3792 9392 3844 9444
rect 6736 9392 6788 9444
rect 10324 9460 10376 9512
rect 12348 9460 12400 9512
rect 14188 9460 14240 9512
rect 16764 9503 16816 9512
rect 16764 9469 16773 9503
rect 16773 9469 16807 9503
rect 16807 9469 16816 9503
rect 16764 9460 16816 9469
rect 1860 9367 1912 9376
rect 1860 9333 1869 9367
rect 1869 9333 1903 9367
rect 1903 9333 1912 9367
rect 1860 9324 1912 9333
rect 2320 9367 2372 9376
rect 2320 9333 2329 9367
rect 2329 9333 2363 9367
rect 2363 9333 2372 9367
rect 2320 9324 2372 9333
rect 3608 9367 3660 9376
rect 3608 9333 3617 9367
rect 3617 9333 3651 9367
rect 3651 9333 3660 9367
rect 3608 9324 3660 9333
rect 4068 9324 4120 9376
rect 4160 9324 4212 9376
rect 5172 9324 5224 9376
rect 6552 9324 6604 9376
rect 6920 9324 6972 9376
rect 7196 9367 7248 9376
rect 7196 9333 7205 9367
rect 7205 9333 7239 9367
rect 7239 9333 7248 9367
rect 7196 9324 7248 9333
rect 9404 9324 9456 9376
rect 9680 9392 9732 9444
rect 12164 9392 12216 9444
rect 12808 9392 12860 9444
rect 14004 9392 14056 9444
rect 12992 9324 13044 9376
rect 17960 9460 18012 9512
rect 19156 9460 19208 9512
rect 20812 9460 20864 9512
rect 19708 9392 19760 9444
rect 15200 9367 15252 9376
rect 15200 9333 15209 9367
rect 15209 9333 15243 9367
rect 15243 9333 15252 9367
rect 15200 9324 15252 9333
rect 16948 9324 17000 9376
rect 17500 9324 17552 9376
rect 7912 9222 7964 9274
rect 7976 9222 8028 9274
rect 8040 9222 8092 9274
rect 8104 9222 8156 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 15035 9222 15087 9274
rect 2780 9052 2832 9104
rect 4068 9120 4120 9172
rect 12440 9120 12492 9172
rect 13912 9120 13964 9172
rect 14464 9120 14516 9172
rect 16764 9120 16816 9172
rect 17776 9163 17828 9172
rect 17776 9129 17785 9163
rect 17785 9129 17819 9163
rect 17819 9129 17828 9163
rect 17776 9120 17828 9129
rect 18144 9120 18196 9172
rect 19156 9120 19208 9172
rect 2872 8984 2924 9036
rect 3516 8984 3568 9036
rect 3608 8984 3660 9036
rect 8208 9052 8260 9104
rect 3884 8916 3936 8968
rect 6736 8891 6788 8900
rect 6736 8857 6745 8891
rect 6745 8857 6779 8891
rect 6779 8857 6788 8891
rect 6736 8848 6788 8857
rect 7012 8984 7064 9036
rect 9036 8984 9088 9036
rect 11060 9052 11112 9104
rect 11152 9052 11204 9104
rect 12808 8984 12860 9036
rect 12900 9027 12952 9036
rect 12900 8993 12909 9027
rect 12909 8993 12943 9027
rect 12943 8993 12952 9027
rect 12900 8984 12952 8993
rect 13820 8984 13872 9036
rect 6920 8916 6972 8968
rect 9128 8916 9180 8968
rect 9772 8916 9824 8968
rect 12348 8916 12400 8968
rect 15384 8984 15436 9036
rect 15476 8984 15528 9036
rect 17040 8984 17092 9036
rect 18052 8984 18104 9036
rect 8852 8848 8904 8900
rect 5080 8780 5132 8832
rect 5448 8823 5500 8832
rect 5448 8789 5457 8823
rect 5457 8789 5491 8823
rect 5491 8789 5500 8823
rect 5448 8780 5500 8789
rect 6092 8780 6144 8832
rect 6920 8780 6972 8832
rect 8668 8823 8720 8832
rect 8668 8789 8677 8823
rect 8677 8789 8711 8823
rect 8711 8789 8720 8823
rect 8668 8780 8720 8789
rect 11796 8780 11848 8832
rect 12256 8780 12308 8832
rect 15292 8780 15344 8832
rect 16028 8916 16080 8968
rect 18788 8916 18840 8968
rect 18236 8848 18288 8900
rect 19892 8848 19944 8900
rect 18144 8780 18196 8832
rect 19064 8780 19116 8832
rect 4447 8678 4499 8730
rect 4511 8678 4563 8730
rect 4575 8678 4627 8730
rect 4639 8678 4691 8730
rect 11378 8678 11430 8730
rect 11442 8678 11494 8730
rect 11506 8678 11558 8730
rect 11570 8678 11622 8730
rect 18308 8678 18360 8730
rect 18372 8678 18424 8730
rect 18436 8678 18488 8730
rect 18500 8678 18552 8730
rect 3424 8576 3476 8628
rect 5080 8576 5132 8628
rect 6092 8576 6144 8628
rect 4344 8508 4396 8560
rect 7012 8551 7064 8560
rect 7012 8517 7021 8551
rect 7021 8517 7055 8551
rect 7055 8517 7064 8551
rect 7012 8508 7064 8517
rect 1308 8440 1360 8492
rect 1860 8372 1912 8424
rect 2780 8483 2832 8492
rect 2780 8449 2789 8483
rect 2789 8449 2823 8483
rect 2823 8449 2832 8483
rect 4896 8483 4948 8492
rect 2780 8440 2832 8449
rect 4896 8449 4905 8483
rect 4905 8449 4939 8483
rect 4939 8449 4948 8483
rect 4896 8440 4948 8449
rect 5080 8483 5132 8492
rect 5080 8449 5089 8483
rect 5089 8449 5123 8483
rect 5123 8449 5132 8483
rect 5080 8440 5132 8449
rect 7104 8440 7156 8492
rect 7748 8508 7800 8560
rect 9956 8576 10008 8628
rect 10324 8576 10376 8628
rect 12440 8619 12492 8628
rect 12440 8585 12449 8619
rect 12449 8585 12483 8619
rect 12483 8585 12492 8619
rect 12440 8576 12492 8585
rect 12808 8576 12860 8628
rect 11520 8508 11572 8560
rect 12348 8508 12400 8560
rect 8392 8440 8444 8492
rect 4804 8415 4856 8424
rect 4804 8381 4813 8415
rect 4813 8381 4847 8415
rect 4847 8381 4856 8415
rect 4804 8372 4856 8381
rect 6920 8372 6972 8424
rect 7748 8372 7800 8424
rect 9128 8372 9180 8424
rect 12900 8440 12952 8492
rect 14188 8483 14240 8492
rect 14188 8449 14197 8483
rect 14197 8449 14231 8483
rect 14231 8449 14240 8483
rect 14188 8440 14240 8449
rect 18052 8619 18104 8628
rect 15936 8508 15988 8560
rect 18052 8585 18061 8619
rect 18061 8585 18095 8619
rect 18095 8585 18104 8619
rect 18052 8576 18104 8585
rect 18788 8576 18840 8628
rect 17040 8483 17092 8492
rect 12256 8415 12308 8424
rect 4160 8304 4212 8356
rect 4068 8236 4120 8288
rect 4344 8236 4396 8288
rect 7288 8304 7340 8356
rect 7656 8304 7708 8356
rect 9772 8304 9824 8356
rect 12256 8381 12265 8415
rect 12265 8381 12299 8415
rect 12299 8381 12308 8415
rect 12256 8372 12308 8381
rect 14096 8372 14148 8424
rect 14464 8415 14516 8424
rect 14464 8381 14498 8415
rect 14498 8381 14516 8415
rect 14464 8372 14516 8381
rect 17040 8449 17049 8483
rect 17049 8449 17083 8483
rect 17083 8449 17092 8483
rect 17040 8440 17092 8449
rect 18788 8440 18840 8492
rect 20536 8483 20588 8492
rect 20536 8449 20545 8483
rect 20545 8449 20579 8483
rect 20579 8449 20588 8483
rect 20536 8440 20588 8449
rect 13268 8304 13320 8356
rect 13636 8304 13688 8356
rect 15292 8304 15344 8356
rect 16580 8304 16632 8356
rect 17868 8304 17920 8356
rect 11980 8236 12032 8288
rect 12164 8236 12216 8288
rect 15660 8236 15712 8288
rect 16120 8236 16172 8288
rect 17592 8236 17644 8288
rect 18144 8236 18196 8288
rect 18972 8304 19024 8356
rect 20536 8304 20588 8356
rect 20076 8279 20128 8288
rect 20076 8245 20085 8279
rect 20085 8245 20119 8279
rect 20119 8245 20128 8279
rect 20076 8236 20128 8245
rect 7912 8134 7964 8186
rect 7976 8134 8028 8186
rect 8040 8134 8092 8186
rect 8104 8134 8156 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 15035 8134 15087 8186
rect 1952 8032 2004 8084
rect 2320 8032 2372 8084
rect 6552 8032 6604 8084
rect 7196 8032 7248 8084
rect 5448 7964 5500 8016
rect 10232 8032 10284 8084
rect 11152 8032 11204 8084
rect 14740 8032 14792 8084
rect 15200 8032 15252 8084
rect 10508 7964 10560 8016
rect 10692 7964 10744 8016
rect 11796 8007 11848 8016
rect 11796 7973 11830 8007
rect 11830 7973 11848 8007
rect 11796 7964 11848 7973
rect 11980 7964 12032 8016
rect 14280 7964 14332 8016
rect 15752 7964 15804 8016
rect 16028 7964 16080 8016
rect 18788 8032 18840 8084
rect 2320 7896 2372 7948
rect 2412 7828 2464 7880
rect 2596 7871 2648 7880
rect 2596 7837 2605 7871
rect 2605 7837 2639 7871
rect 2639 7837 2648 7871
rect 2596 7828 2648 7837
rect 2872 7828 2924 7880
rect 4436 7828 4488 7880
rect 6368 7896 6420 7948
rect 7840 7896 7892 7948
rect 9588 7896 9640 7948
rect 10048 7939 10100 7948
rect 10048 7905 10057 7939
rect 10057 7905 10091 7939
rect 10091 7905 10100 7939
rect 10048 7896 10100 7905
rect 11244 7896 11296 7948
rect 14188 7896 14240 7948
rect 16580 7896 16632 7948
rect 18880 7964 18932 8016
rect 19156 7896 19208 7948
rect 6460 7828 6512 7880
rect 6552 7828 6604 7880
rect 10140 7871 10192 7880
rect 10140 7837 10149 7871
rect 10149 7837 10183 7871
rect 10183 7837 10192 7871
rect 10140 7828 10192 7837
rect 10324 7871 10376 7880
rect 10324 7837 10333 7871
rect 10333 7837 10367 7871
rect 10367 7837 10376 7871
rect 10324 7828 10376 7837
rect 11520 7871 11572 7880
rect 11520 7837 11529 7871
rect 11529 7837 11563 7871
rect 11563 7837 11572 7871
rect 11520 7828 11572 7837
rect 13084 7828 13136 7880
rect 13544 7828 13596 7880
rect 13820 7828 13872 7880
rect 5908 7760 5960 7812
rect 11060 7760 11112 7812
rect 3792 7692 3844 7744
rect 8392 7692 8444 7744
rect 9128 7692 9180 7744
rect 9496 7692 9548 7744
rect 10968 7692 11020 7744
rect 12164 7692 12216 7744
rect 14372 7760 14424 7812
rect 12900 7735 12952 7744
rect 12900 7701 12909 7735
rect 12909 7701 12943 7735
rect 12943 7701 12952 7735
rect 12900 7692 12952 7701
rect 14004 7692 14056 7744
rect 15476 7692 15528 7744
rect 4447 7590 4499 7642
rect 4511 7590 4563 7642
rect 4575 7590 4627 7642
rect 4639 7590 4691 7642
rect 11378 7590 11430 7642
rect 11442 7590 11494 7642
rect 11506 7590 11558 7642
rect 11570 7590 11622 7642
rect 18308 7590 18360 7642
rect 18372 7590 18424 7642
rect 18436 7590 18488 7642
rect 18500 7590 18552 7642
rect 1400 7531 1452 7540
rect 1400 7497 1409 7531
rect 1409 7497 1443 7531
rect 1443 7497 1452 7531
rect 1400 7488 1452 7497
rect 2136 7488 2188 7540
rect 3516 7488 3568 7540
rect 4160 7488 4212 7540
rect 7748 7488 7800 7540
rect 9496 7488 9548 7540
rect 9772 7531 9824 7540
rect 9772 7497 9781 7531
rect 9781 7497 9815 7531
rect 9815 7497 9824 7531
rect 9772 7488 9824 7497
rect 10140 7488 10192 7540
rect 12624 7488 12676 7540
rect 14188 7488 14240 7540
rect 18788 7488 18840 7540
rect 1768 7352 1820 7404
rect 5448 7352 5500 7404
rect 12532 7420 12584 7472
rect 12992 7420 13044 7472
rect 17040 7420 17092 7472
rect 19800 7488 19852 7540
rect 20628 7488 20680 7540
rect 14004 7352 14056 7404
rect 15752 7395 15804 7404
rect 15752 7361 15761 7395
rect 15761 7361 15795 7395
rect 15795 7361 15804 7395
rect 18144 7395 18196 7404
rect 15752 7352 15804 7361
rect 18144 7361 18153 7395
rect 18153 7361 18187 7395
rect 18187 7361 18196 7395
rect 18144 7352 18196 7361
rect 19156 7352 19208 7404
rect 1584 7284 1636 7336
rect 2228 7327 2280 7336
rect 2228 7293 2237 7327
rect 2237 7293 2271 7327
rect 2271 7293 2280 7327
rect 2228 7284 2280 7293
rect 3884 7284 3936 7336
rect 4344 7284 4396 7336
rect 6460 7284 6512 7336
rect 9128 7284 9180 7336
rect 11060 7327 11112 7336
rect 11060 7293 11069 7327
rect 11069 7293 11103 7327
rect 11103 7293 11112 7327
rect 11060 7284 11112 7293
rect 14188 7284 14240 7336
rect 19708 7327 19760 7336
rect 19708 7293 19742 7327
rect 19742 7293 19760 7327
rect 19708 7284 19760 7293
rect 2504 7216 2556 7268
rect 2872 7259 2924 7268
rect 2872 7225 2906 7259
rect 2906 7225 2924 7259
rect 2872 7216 2924 7225
rect 5908 7216 5960 7268
rect 7748 7216 7800 7268
rect 8484 7216 8536 7268
rect 6552 7148 6604 7200
rect 6828 7191 6880 7200
rect 6828 7157 6837 7191
rect 6837 7157 6871 7191
rect 6871 7157 6880 7191
rect 6828 7148 6880 7157
rect 7196 7191 7248 7200
rect 7196 7157 7205 7191
rect 7205 7157 7239 7191
rect 7239 7157 7248 7191
rect 7196 7148 7248 7157
rect 7380 7148 7432 7200
rect 7564 7148 7616 7200
rect 12164 7216 12216 7268
rect 20536 7216 20588 7268
rect 9496 7148 9548 7200
rect 11152 7148 11204 7200
rect 13084 7148 13136 7200
rect 14372 7191 14424 7200
rect 14372 7157 14381 7191
rect 14381 7157 14415 7191
rect 14415 7157 14424 7191
rect 14372 7148 14424 7157
rect 15292 7148 15344 7200
rect 7912 7046 7964 7098
rect 7976 7046 8028 7098
rect 8040 7046 8092 7098
rect 8104 7046 8156 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 15035 7046 15087 7098
rect 2228 6944 2280 6996
rect 2780 6987 2832 6996
rect 2780 6953 2789 6987
rect 2789 6953 2823 6987
rect 2823 6953 2832 6987
rect 2780 6944 2832 6953
rect 4896 6944 4948 6996
rect 8392 6944 8444 6996
rect 12256 6944 12308 6996
rect 12624 6944 12676 6996
rect 13268 6944 13320 6996
rect 14464 6944 14516 6996
rect 15752 6944 15804 6996
rect 17040 6944 17092 6996
rect 6460 6876 6512 6928
rect 6552 6876 6604 6928
rect 2872 6851 2924 6860
rect 2872 6817 2881 6851
rect 2881 6817 2915 6851
rect 2915 6817 2924 6851
rect 2872 6808 2924 6817
rect 4252 6808 4304 6860
rect 9772 6876 9824 6928
rect 10600 6876 10652 6928
rect 10876 6876 10928 6928
rect 12164 6876 12216 6928
rect 12532 6876 12584 6928
rect 17960 6876 18012 6928
rect 10048 6851 10100 6860
rect 2964 6783 3016 6792
rect 2964 6749 2973 6783
rect 2973 6749 3007 6783
rect 3007 6749 3016 6783
rect 2964 6740 3016 6749
rect 5448 6740 5500 6792
rect 6828 6740 6880 6792
rect 7012 6740 7064 6792
rect 7288 6672 7340 6724
rect 10048 6817 10057 6851
rect 10057 6817 10091 6851
rect 10091 6817 10100 6851
rect 10048 6808 10100 6817
rect 12440 6808 12492 6860
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 10324 6783 10376 6792
rect 10324 6749 10333 6783
rect 10333 6749 10367 6783
rect 10367 6749 10376 6783
rect 10324 6740 10376 6749
rect 12624 6783 12676 6792
rect 12624 6749 12633 6783
rect 12633 6749 12667 6783
rect 12667 6749 12676 6783
rect 12624 6740 12676 6749
rect 2412 6647 2464 6656
rect 2412 6613 2421 6647
rect 2421 6613 2455 6647
rect 2455 6613 2464 6647
rect 2412 6604 2464 6613
rect 6276 6647 6328 6656
rect 6276 6613 6285 6647
rect 6285 6613 6319 6647
rect 6319 6613 6328 6647
rect 6276 6604 6328 6613
rect 7748 6604 7800 6656
rect 9588 6604 9640 6656
rect 11244 6672 11296 6724
rect 14188 6808 14240 6860
rect 15568 6808 15620 6860
rect 14372 6740 14424 6792
rect 15752 6740 15804 6792
rect 17960 6740 18012 6792
rect 18144 6783 18196 6792
rect 18144 6749 18153 6783
rect 18153 6749 18187 6783
rect 18187 6749 18196 6783
rect 18144 6740 18196 6749
rect 9956 6604 10008 6656
rect 14464 6672 14516 6724
rect 18880 6672 18932 6724
rect 15752 6604 15804 6656
rect 17316 6604 17368 6656
rect 19156 6647 19208 6656
rect 19156 6613 19165 6647
rect 19165 6613 19199 6647
rect 19199 6613 19208 6647
rect 19156 6604 19208 6613
rect 19524 6672 19576 6724
rect 4447 6502 4499 6554
rect 4511 6502 4563 6554
rect 4575 6502 4627 6554
rect 4639 6502 4691 6554
rect 11378 6502 11430 6554
rect 11442 6502 11494 6554
rect 11506 6502 11558 6554
rect 11570 6502 11622 6554
rect 18308 6502 18360 6554
rect 18372 6502 18424 6554
rect 18436 6502 18488 6554
rect 18500 6502 18552 6554
rect 2044 6307 2096 6316
rect 2044 6273 2053 6307
rect 2053 6273 2087 6307
rect 2087 6273 2096 6307
rect 2044 6264 2096 6273
rect 2596 6375 2648 6384
rect 2596 6341 2605 6375
rect 2605 6341 2639 6375
rect 2639 6341 2648 6375
rect 2596 6332 2648 6341
rect 7288 6400 7340 6452
rect 8484 6400 8536 6452
rect 8576 6400 8628 6452
rect 10324 6400 10376 6452
rect 12624 6400 12676 6452
rect 14556 6400 14608 6452
rect 15476 6332 15528 6384
rect 2780 6264 2832 6316
rect 3884 6264 3936 6316
rect 4528 6307 4580 6316
rect 4528 6273 4537 6307
rect 4537 6273 4571 6307
rect 4571 6273 4580 6307
rect 4528 6264 4580 6273
rect 14372 6264 14424 6316
rect 4344 6196 4396 6248
rect 4620 6196 4672 6248
rect 2964 6128 3016 6180
rect 1676 6060 1728 6112
rect 1952 6103 2004 6112
rect 1952 6069 1961 6103
rect 1961 6069 1995 6103
rect 1995 6069 2004 6103
rect 1952 6060 2004 6069
rect 2688 6060 2740 6112
rect 6920 6196 6972 6248
rect 7288 6239 7340 6248
rect 7288 6205 7322 6239
rect 7322 6205 7340 6239
rect 7288 6196 7340 6205
rect 9128 6196 9180 6248
rect 9956 6196 10008 6248
rect 10692 6196 10744 6248
rect 11980 6196 12032 6248
rect 12348 6196 12400 6248
rect 17960 6400 18012 6452
rect 17868 6332 17920 6384
rect 17132 6264 17184 6316
rect 17316 6264 17368 6316
rect 17408 6196 17460 6248
rect 17776 6196 17828 6248
rect 18144 6196 18196 6248
rect 19432 6264 19484 6316
rect 3608 6103 3660 6112
rect 3608 6069 3617 6103
rect 3617 6069 3651 6103
rect 3651 6069 3660 6103
rect 12900 6128 12952 6180
rect 12992 6128 13044 6180
rect 3608 6060 3660 6069
rect 5172 6060 5224 6112
rect 5448 6060 5500 6112
rect 11704 6060 11756 6112
rect 15200 6060 15252 6112
rect 15660 6060 15712 6112
rect 7912 5958 7964 6010
rect 7976 5958 8028 6010
rect 8040 5958 8092 6010
rect 8104 5958 8156 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 15035 5958 15087 6010
rect 1952 5856 2004 5908
rect 4160 5856 4212 5908
rect 5264 5856 5316 5908
rect 7012 5856 7064 5908
rect 7748 5856 7800 5908
rect 10048 5899 10100 5908
rect 10048 5865 10057 5899
rect 10057 5865 10091 5899
rect 10091 5865 10100 5899
rect 10048 5856 10100 5865
rect 10508 5856 10560 5908
rect 10692 5856 10744 5908
rect 7380 5788 7432 5840
rect 1768 5763 1820 5772
rect 1768 5729 1777 5763
rect 1777 5729 1811 5763
rect 1811 5729 1820 5763
rect 1768 5720 1820 5729
rect 4804 5720 4856 5772
rect 8392 5720 8444 5772
rect 8852 5788 8904 5840
rect 10968 5788 11020 5840
rect 14096 5856 14148 5908
rect 15200 5856 15252 5908
rect 15752 5899 15804 5908
rect 15752 5865 15761 5899
rect 15761 5865 15795 5899
rect 15795 5865 15804 5899
rect 15752 5856 15804 5865
rect 16948 5856 17000 5908
rect 2688 5652 2740 5704
rect 2872 5695 2924 5704
rect 2872 5661 2881 5695
rect 2881 5661 2915 5695
rect 2915 5661 2924 5695
rect 2872 5652 2924 5661
rect 2504 5584 2556 5636
rect 2596 5584 2648 5636
rect 4528 5652 4580 5704
rect 8484 5652 8536 5704
rect 10048 5720 10100 5772
rect 12624 5720 12676 5772
rect 10508 5695 10560 5704
rect 10508 5661 10517 5695
rect 10517 5661 10551 5695
rect 10551 5661 10560 5695
rect 10508 5652 10560 5661
rect 10692 5695 10744 5704
rect 10692 5661 10701 5695
rect 10701 5661 10735 5695
rect 10735 5661 10744 5695
rect 10692 5652 10744 5661
rect 11980 5695 12032 5704
rect 11980 5661 11989 5695
rect 11989 5661 12023 5695
rect 12023 5661 12032 5695
rect 11980 5652 12032 5661
rect 15292 5788 15344 5840
rect 17960 5788 18012 5840
rect 17040 5720 17092 5772
rect 17316 5720 17368 5772
rect 17500 5763 17552 5772
rect 17500 5729 17534 5763
rect 17534 5729 17552 5763
rect 17500 5720 17552 5729
rect 18880 5856 18932 5908
rect 19892 5788 19944 5840
rect 15568 5652 15620 5704
rect 15936 5652 15988 5704
rect 17132 5652 17184 5704
rect 3332 5584 3384 5636
rect 5264 5584 5316 5636
rect 6644 5584 6696 5636
rect 11612 5584 11664 5636
rect 6000 5516 6052 5568
rect 6368 5516 6420 5568
rect 9588 5516 9640 5568
rect 9956 5516 10008 5568
rect 12900 5516 12952 5568
rect 13360 5559 13412 5568
rect 13360 5525 13369 5559
rect 13369 5525 13403 5559
rect 13403 5525 13412 5559
rect 13360 5516 13412 5525
rect 15476 5516 15528 5568
rect 4447 5414 4499 5466
rect 4511 5414 4563 5466
rect 4575 5414 4627 5466
rect 4639 5414 4691 5466
rect 11378 5414 11430 5466
rect 11442 5414 11494 5466
rect 11506 5414 11558 5466
rect 11570 5414 11622 5466
rect 18308 5414 18360 5466
rect 18372 5414 18424 5466
rect 18436 5414 18488 5466
rect 18500 5414 18552 5466
rect 9680 5312 9732 5364
rect 9956 5312 10008 5364
rect 16396 5312 16448 5364
rect 16856 5312 16908 5364
rect 17316 5312 17368 5364
rect 20536 5312 20588 5364
rect 3792 5176 3844 5228
rect 10140 5244 10192 5296
rect 12900 5244 12952 5296
rect 5264 5176 5316 5228
rect 6368 5176 6420 5228
rect 6460 5176 6512 5228
rect 9956 5176 10008 5228
rect 10232 5176 10284 5228
rect 3884 5108 3936 5160
rect 4068 5083 4120 5092
rect 4068 5049 4077 5083
rect 4077 5049 4111 5083
rect 4111 5049 4120 5083
rect 4068 5040 4120 5049
rect 4804 5040 4856 5092
rect 5264 5040 5316 5092
rect 9496 5108 9548 5160
rect 9588 5108 9640 5160
rect 10140 5108 10192 5160
rect 9864 5040 9916 5092
rect 10692 5176 10744 5228
rect 11704 5176 11756 5228
rect 11152 5108 11204 5160
rect 15200 5176 15252 5228
rect 16948 5219 17000 5228
rect 16948 5185 16957 5219
rect 16957 5185 16991 5219
rect 16991 5185 17000 5219
rect 16948 5176 17000 5185
rect 18972 5176 19024 5228
rect 15292 5151 15344 5160
rect 15292 5117 15301 5151
rect 15301 5117 15335 5151
rect 15335 5117 15344 5151
rect 15292 5108 15344 5117
rect 13636 5040 13688 5092
rect 13912 5040 13964 5092
rect 16580 5040 16632 5092
rect 17040 5108 17092 5160
rect 18144 5108 18196 5160
rect 20628 5108 20680 5160
rect 3700 5015 3752 5024
rect 3700 4981 3709 5015
rect 3709 4981 3743 5015
rect 3743 4981 3752 5015
rect 3700 4972 3752 4981
rect 4252 4972 4304 5024
rect 5448 5015 5500 5024
rect 5448 4981 5457 5015
rect 5457 4981 5491 5015
rect 5491 4981 5500 5015
rect 5448 4972 5500 4981
rect 6920 4972 6972 5024
rect 7380 4972 7432 5024
rect 9128 4972 9180 5024
rect 10784 4972 10836 5024
rect 15936 4972 15988 5024
rect 16672 4972 16724 5024
rect 16856 5015 16908 5024
rect 16856 4981 16865 5015
rect 16865 4981 16899 5015
rect 16899 4981 16908 5015
rect 16856 4972 16908 4981
rect 19708 4972 19760 5024
rect 7912 4870 7964 4922
rect 7976 4870 8028 4922
rect 8040 4870 8092 4922
rect 8104 4870 8156 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 15035 4870 15087 4922
rect 2688 4768 2740 4820
rect 4896 4811 4948 4820
rect 4896 4777 4905 4811
rect 4905 4777 4939 4811
rect 4939 4777 4948 4811
rect 4896 4768 4948 4777
rect 5448 4768 5500 4820
rect 7104 4768 7156 4820
rect 13268 4768 13320 4820
rect 14280 4768 14332 4820
rect 16856 4768 16908 4820
rect 19616 4811 19668 4820
rect 19616 4777 19625 4811
rect 19625 4777 19659 4811
rect 19659 4777 19668 4811
rect 19616 4768 19668 4777
rect 204 4700 256 4752
rect 3240 4743 3292 4752
rect 3240 4709 3249 4743
rect 3249 4709 3283 4743
rect 3283 4709 3292 4743
rect 3240 4700 3292 4709
rect 2596 4632 2648 4684
rect 3792 4700 3844 4752
rect 5816 4700 5868 4752
rect 7564 4700 7616 4752
rect 4068 4632 4120 4684
rect 4160 4632 4212 4684
rect 2964 4564 3016 4616
rect 3792 4564 3844 4616
rect 6920 4632 6972 4684
rect 7380 4675 7432 4684
rect 7380 4641 7389 4675
rect 7389 4641 7423 4675
rect 7423 4641 7432 4675
rect 7380 4632 7432 4641
rect 9956 4632 10008 4684
rect 4804 4564 4856 4616
rect 5356 4607 5408 4616
rect 5356 4573 5365 4607
rect 5365 4573 5399 4607
rect 5399 4573 5408 4607
rect 5356 4564 5408 4573
rect 2872 4496 2924 4548
rect 5172 4496 5224 4548
rect 3148 4428 3200 4480
rect 3976 4428 4028 4480
rect 9680 4564 9732 4616
rect 10140 4607 10192 4616
rect 10140 4573 10149 4607
rect 10149 4573 10183 4607
rect 10183 4573 10192 4607
rect 10140 4564 10192 4573
rect 9588 4496 9640 4548
rect 10600 4428 10652 4480
rect 11336 4632 11388 4684
rect 13360 4700 13412 4752
rect 11980 4632 12032 4684
rect 12808 4632 12860 4684
rect 16028 4632 16080 4684
rect 16948 4700 17000 4752
rect 12532 4564 12584 4616
rect 12992 4428 13044 4480
rect 13636 4428 13688 4480
rect 15752 4428 15804 4480
rect 18788 4632 18840 4684
rect 17040 4564 17092 4616
rect 17132 4496 17184 4548
rect 17776 4428 17828 4480
rect 18972 4471 19024 4480
rect 18972 4437 18981 4471
rect 18981 4437 19015 4471
rect 19015 4437 19024 4471
rect 18972 4428 19024 4437
rect 4447 4326 4499 4378
rect 4511 4326 4563 4378
rect 4575 4326 4627 4378
rect 4639 4326 4691 4378
rect 11378 4326 11430 4378
rect 11442 4326 11494 4378
rect 11506 4326 11558 4378
rect 11570 4326 11622 4378
rect 18308 4326 18360 4378
rect 18372 4326 18424 4378
rect 18436 4326 18488 4378
rect 18500 4326 18552 4378
rect 3148 4224 3200 4276
rect 4068 4224 4120 4276
rect 4804 4224 4856 4276
rect 9496 4224 9548 4276
rect 13912 4224 13964 4276
rect 1584 4020 1636 4072
rect 2780 4020 2832 4072
rect 9588 4156 9640 4208
rect 4436 4063 4488 4072
rect 2872 3952 2924 4004
rect 3332 3952 3384 4004
rect 3608 3884 3660 3936
rect 4436 4029 4445 4063
rect 4445 4029 4479 4063
rect 4479 4029 4488 4063
rect 4436 4020 4488 4029
rect 4896 4020 4948 4072
rect 6092 4088 6144 4140
rect 6828 4088 6880 4140
rect 10508 4088 10560 4140
rect 10784 4088 10836 4140
rect 10876 4088 10928 4140
rect 11060 4156 11112 4208
rect 12624 4156 12676 4208
rect 17132 4224 17184 4276
rect 12808 4088 12860 4140
rect 14280 4156 14332 4208
rect 6000 4020 6052 4072
rect 4344 3952 4396 4004
rect 6644 3952 6696 4004
rect 8576 3952 8628 4004
rect 8668 3952 8720 4004
rect 12348 3952 12400 4004
rect 12532 4020 12584 4072
rect 13544 4020 13596 4072
rect 13728 4020 13780 4072
rect 15200 4131 15252 4140
rect 15200 4097 15209 4131
rect 15209 4097 15243 4131
rect 15243 4097 15252 4131
rect 15200 4088 15252 4097
rect 16304 4088 16356 4140
rect 17868 4088 17920 4140
rect 18972 4088 19024 4140
rect 13176 3952 13228 4004
rect 17960 4020 18012 4072
rect 20536 4063 20588 4072
rect 20536 4029 20545 4063
rect 20545 4029 20579 4063
rect 20579 4029 20588 4063
rect 20536 4020 20588 4029
rect 5172 3927 5224 3936
rect 5172 3893 5181 3927
rect 5181 3893 5215 3927
rect 5215 3893 5224 3927
rect 5172 3884 5224 3893
rect 6920 3884 6972 3936
rect 10232 3884 10284 3936
rect 10508 3884 10560 3936
rect 11060 3927 11112 3936
rect 11060 3893 11069 3927
rect 11069 3893 11103 3927
rect 11103 3893 11112 3927
rect 11060 3884 11112 3893
rect 11152 3884 11204 3936
rect 11796 3884 11848 3936
rect 12440 3927 12492 3936
rect 12440 3893 12449 3927
rect 12449 3893 12483 3927
rect 12483 3893 12492 3927
rect 15200 3952 15252 4004
rect 15568 3952 15620 4004
rect 16672 3952 16724 4004
rect 12440 3884 12492 3893
rect 13728 3884 13780 3936
rect 14096 3884 14148 3936
rect 16028 3884 16080 3936
rect 16304 3927 16356 3936
rect 16304 3893 16313 3927
rect 16313 3893 16347 3927
rect 16347 3893 16356 3927
rect 16304 3884 16356 3893
rect 21732 3884 21784 3936
rect 7912 3782 7964 3834
rect 7976 3782 8028 3834
rect 8040 3782 8092 3834
rect 8104 3782 8156 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 15035 3782 15087 3834
rect 2964 3723 3016 3732
rect 2964 3689 2973 3723
rect 2973 3689 3007 3723
rect 3007 3689 3016 3723
rect 2964 3680 3016 3689
rect 4160 3680 4212 3732
rect 4344 3680 4396 3732
rect 4988 3680 5040 3732
rect 5172 3680 5224 3732
rect 6644 3723 6696 3732
rect 6644 3689 6653 3723
rect 6653 3689 6687 3723
rect 6687 3689 6696 3723
rect 6644 3680 6696 3689
rect 7012 3723 7064 3732
rect 7012 3689 7021 3723
rect 7021 3689 7055 3723
rect 7055 3689 7064 3723
rect 7012 3680 7064 3689
rect 8208 3680 8260 3732
rect 9864 3680 9916 3732
rect 5080 3612 5132 3664
rect 5356 3612 5408 3664
rect 7104 3655 7156 3664
rect 7104 3621 7113 3655
rect 7113 3621 7147 3655
rect 7147 3621 7156 3655
rect 7104 3612 7156 3621
rect 9404 3612 9456 3664
rect 10600 3655 10652 3664
rect 10600 3621 10609 3655
rect 10609 3621 10643 3655
rect 10643 3621 10652 3655
rect 10600 3612 10652 3621
rect 10784 3680 10836 3732
rect 13176 3680 13228 3732
rect 13452 3680 13504 3732
rect 13728 3680 13780 3732
rect 16304 3680 16356 3732
rect 14004 3655 14056 3664
rect 1584 3587 1636 3596
rect 1584 3553 1593 3587
rect 1593 3553 1627 3587
rect 1627 3553 1636 3587
rect 1584 3544 1636 3553
rect 3148 3544 3200 3596
rect 2964 3408 3016 3460
rect 1124 3340 1176 3392
rect 5632 3544 5684 3596
rect 5908 3587 5960 3596
rect 5908 3553 5917 3587
rect 5917 3553 5951 3587
rect 5951 3553 5960 3587
rect 5908 3544 5960 3553
rect 6000 3544 6052 3596
rect 9312 3544 9364 3596
rect 10508 3544 10560 3596
rect 5080 3476 5132 3528
rect 6460 3476 6512 3528
rect 10324 3476 10376 3528
rect 10876 3519 10928 3528
rect 10876 3485 10885 3519
rect 10885 3485 10919 3519
rect 10919 3485 10928 3519
rect 10876 3476 10928 3485
rect 12624 3476 12676 3528
rect 14004 3621 14013 3655
rect 14013 3621 14047 3655
rect 14047 3621 14056 3655
rect 14004 3612 14056 3621
rect 13360 3544 13412 3596
rect 14004 3476 14056 3528
rect 5448 3383 5500 3392
rect 5448 3349 5457 3383
rect 5457 3349 5491 3383
rect 5491 3349 5500 3383
rect 5448 3340 5500 3349
rect 6552 3340 6604 3392
rect 7380 3408 7432 3460
rect 9864 3408 9916 3460
rect 11244 3408 11296 3460
rect 16580 3612 16632 3664
rect 18972 3612 19024 3664
rect 19064 3612 19116 3664
rect 14740 3544 14792 3596
rect 15752 3587 15804 3596
rect 15752 3553 15761 3587
rect 15761 3553 15795 3587
rect 15795 3553 15804 3587
rect 15752 3544 15804 3553
rect 15016 3408 15068 3460
rect 8392 3340 8444 3392
rect 10048 3340 10100 3392
rect 10692 3340 10744 3392
rect 10876 3340 10928 3392
rect 11060 3340 11112 3392
rect 16488 3476 16540 3528
rect 18236 3476 18288 3528
rect 4447 3238 4499 3290
rect 4511 3238 4563 3290
rect 4575 3238 4627 3290
rect 4639 3238 4691 3290
rect 11378 3238 11430 3290
rect 11442 3238 11494 3290
rect 11506 3238 11558 3290
rect 11570 3238 11622 3290
rect 18308 3238 18360 3290
rect 18372 3238 18424 3290
rect 18436 3238 18488 3290
rect 18500 3238 18552 3290
rect 5908 3136 5960 3188
rect 6736 3136 6788 3188
rect 8668 3136 8720 3188
rect 10692 3179 10744 3188
rect 2780 3111 2832 3120
rect 2780 3077 2789 3111
rect 2789 3077 2823 3111
rect 2823 3077 2832 3111
rect 2780 3068 2832 3077
rect 5080 3068 5132 3120
rect 5264 3111 5316 3120
rect 5264 3077 5273 3111
rect 5273 3077 5307 3111
rect 5307 3077 5316 3111
rect 5264 3068 5316 3077
rect 3608 3000 3660 3052
rect 1492 2932 1544 2984
rect 4804 3000 4856 3052
rect 6368 3043 6420 3052
rect 6368 3009 6377 3043
rect 6377 3009 6411 3043
rect 6411 3009 6420 3043
rect 6368 3000 6420 3009
rect 7748 3068 7800 3120
rect 10692 3145 10701 3179
rect 10701 3145 10735 3179
rect 10735 3145 10744 3179
rect 10692 3136 10744 3145
rect 12164 3136 12216 3188
rect 12808 3179 12860 3188
rect 12808 3145 12817 3179
rect 12817 3145 12851 3179
rect 12851 3145 12860 3179
rect 12808 3136 12860 3145
rect 13360 3136 13412 3188
rect 13452 3136 13504 3188
rect 14556 3136 14608 3188
rect 20720 3136 20772 3188
rect 8484 3000 8536 3052
rect 18052 3068 18104 3120
rect 14188 3000 14240 3052
rect 15016 3043 15068 3052
rect 5448 2932 5500 2984
rect 2228 2864 2280 2916
rect 4252 2864 4304 2916
rect 664 2796 716 2848
rect 1768 2796 1820 2848
rect 5540 2864 5592 2916
rect 5724 2975 5776 2984
rect 5724 2941 5733 2975
rect 5733 2941 5767 2975
rect 5767 2941 5776 2975
rect 5724 2932 5776 2941
rect 6184 2932 6236 2984
rect 6552 2932 6604 2984
rect 9128 2932 9180 2984
rect 9588 2975 9640 2984
rect 9588 2941 9622 2975
rect 9622 2941 9640 2975
rect 9588 2932 9640 2941
rect 9864 2932 9916 2984
rect 15016 3009 15025 3043
rect 15025 3009 15059 3043
rect 15059 3009 15068 3043
rect 15016 3000 15068 3009
rect 15292 3000 15344 3052
rect 21272 3068 21324 3120
rect 19156 2932 19208 2984
rect 19432 2975 19484 2984
rect 19432 2941 19441 2975
rect 19441 2941 19475 2975
rect 19475 2941 19484 2975
rect 19432 2932 19484 2941
rect 20536 2975 20588 2984
rect 20536 2941 20545 2975
rect 20545 2941 20579 2975
rect 20579 2941 20588 2975
rect 20536 2932 20588 2941
rect 5908 2864 5960 2916
rect 7748 2907 7800 2916
rect 7748 2873 7757 2907
rect 7757 2873 7791 2907
rect 7791 2873 7800 2907
rect 7748 2864 7800 2873
rect 11428 2864 11480 2916
rect 5172 2796 5224 2848
rect 6368 2796 6420 2848
rect 7472 2796 7524 2848
rect 8392 2796 8444 2848
rect 15292 2864 15344 2916
rect 15844 2864 15896 2916
rect 20168 2864 20220 2916
rect 22652 2864 22704 2916
rect 13268 2839 13320 2848
rect 13268 2805 13277 2839
rect 13277 2805 13311 2839
rect 13311 2805 13320 2839
rect 13268 2796 13320 2805
rect 14004 2796 14056 2848
rect 19340 2796 19392 2848
rect 22192 2796 22244 2848
rect 7912 2694 7964 2746
rect 7976 2694 8028 2746
rect 8040 2694 8092 2746
rect 8104 2694 8156 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 15035 2694 15087 2746
rect 2872 2635 2924 2644
rect 2872 2601 2881 2635
rect 2881 2601 2915 2635
rect 2915 2601 2924 2635
rect 2872 2592 2924 2601
rect 3148 2592 3200 2644
rect 3424 2592 3476 2644
rect 5540 2635 5592 2644
rect 5540 2601 5549 2635
rect 5549 2601 5583 2635
rect 5583 2601 5592 2635
rect 5540 2592 5592 2601
rect 5816 2592 5868 2644
rect 6920 2635 6972 2644
rect 6920 2601 6929 2635
rect 6929 2601 6963 2635
rect 6963 2601 6972 2635
rect 6920 2592 6972 2601
rect 2044 2524 2096 2576
rect 4804 2524 4856 2576
rect 7472 2524 7524 2576
rect 1492 2456 1544 2508
rect 3424 2456 3476 2508
rect 3700 2456 3752 2508
rect 6092 2456 6144 2508
rect 7932 2456 7984 2508
rect 8116 2499 8168 2508
rect 8116 2465 8125 2499
rect 8125 2465 8159 2499
rect 8159 2465 8168 2499
rect 8116 2456 8168 2465
rect 8576 2499 8628 2508
rect 8576 2465 8585 2499
rect 8585 2465 8619 2499
rect 8619 2465 8628 2499
rect 8576 2456 8628 2465
rect 9680 2592 9732 2644
rect 10416 2592 10468 2644
rect 12440 2592 12492 2644
rect 8852 2456 8904 2508
rect 11428 2499 11480 2508
rect 11428 2465 11437 2499
rect 11437 2465 11471 2499
rect 11471 2465 11480 2499
rect 11428 2456 11480 2465
rect 12440 2456 12492 2508
rect 12992 2592 13044 2644
rect 20168 2635 20220 2644
rect 20168 2601 20177 2635
rect 20177 2601 20211 2635
rect 20211 2601 20220 2635
rect 20168 2592 20220 2601
rect 12900 2524 12952 2576
rect 15384 2524 15436 2576
rect 17224 2524 17276 2576
rect 13544 2456 13596 2508
rect 3608 2388 3660 2440
rect 6460 2388 6512 2440
rect 8208 2431 8260 2440
rect 8208 2397 8217 2431
rect 8217 2397 8251 2431
rect 8251 2397 8260 2431
rect 8208 2388 8260 2397
rect 2596 2320 2648 2372
rect 2780 2295 2832 2304
rect 2780 2261 2789 2295
rect 2789 2261 2823 2295
rect 2823 2261 2832 2295
rect 5908 2320 5960 2372
rect 2780 2252 2832 2261
rect 6552 2295 6604 2304
rect 6552 2261 6561 2295
rect 6561 2261 6595 2295
rect 6595 2261 6604 2295
rect 6552 2252 6604 2261
rect 7288 2320 7340 2372
rect 8668 2388 8720 2440
rect 9956 2388 10008 2440
rect 14740 2456 14792 2508
rect 15476 2499 15528 2508
rect 15476 2465 15485 2499
rect 15485 2465 15519 2499
rect 15519 2465 15528 2499
rect 15476 2456 15528 2465
rect 18696 2499 18748 2508
rect 18696 2465 18705 2499
rect 18705 2465 18739 2499
rect 18739 2465 18748 2499
rect 18696 2456 18748 2465
rect 19984 2499 20036 2508
rect 19984 2465 19993 2499
rect 19993 2465 20027 2499
rect 20027 2465 20036 2499
rect 19984 2456 20036 2465
rect 14648 2388 14700 2440
rect 17224 2388 17276 2440
rect 10140 2320 10192 2372
rect 14096 2320 14148 2372
rect 12440 2252 12492 2304
rect 13452 2252 13504 2304
rect 13544 2252 13596 2304
rect 4447 2150 4499 2202
rect 4511 2150 4563 2202
rect 4575 2150 4627 2202
rect 4639 2150 4691 2202
rect 11378 2150 11430 2202
rect 11442 2150 11494 2202
rect 11506 2150 11558 2202
rect 11570 2150 11622 2202
rect 18308 2150 18360 2202
rect 18372 2150 18424 2202
rect 18436 2150 18488 2202
rect 18500 2150 18552 2202
rect 1584 2048 1636 2100
rect 5356 2048 5408 2100
rect 6552 2048 6604 2100
rect 15476 2048 15528 2100
rect 2596 1980 2648 2032
rect 3792 1980 3844 2032
rect 8208 1980 8260 2032
rect 2872 1912 2924 1964
rect 13452 1980 13504 2032
rect 14464 1980 14516 2032
rect 16212 1912 16264 1964
rect 3332 1844 3384 1896
rect 19984 1844 20036 1896
rect 8116 1776 8168 1828
rect 16120 1776 16172 1828
rect 3608 1708 3660 1760
rect 17500 1708 17552 1760
rect 2780 1640 2832 1692
rect 15200 1640 15252 1692
rect 7932 1572 7984 1624
rect 13820 1572 13872 1624
rect 9036 1504 9088 1556
rect 17224 1504 17276 1556
rect 3424 1436 3476 1488
rect 14372 1436 14424 1488
rect 19524 1436 19576 1488
rect 18328 1368 18380 1420
rect 19064 1368 19116 1420
rect 12348 1300 12400 1352
rect 18880 1300 18932 1352
rect 3608 280 3660 332
rect 6276 280 6328 332
<< metal2 >>
rect 2870 22520 2926 23000
rect 3882 22672 3938 22681
rect 3882 22607 3938 22616
rect 2884 20346 2912 22520
rect 3514 22264 3570 22273
rect 3514 22199 3570 22208
rect 3528 21350 3556 22199
rect 3516 21344 3568 21350
rect 3146 21312 3202 21321
rect 3516 21286 3568 21292
rect 3146 21247 3202 21256
rect 3160 21146 3188 21247
rect 3148 21140 3200 21146
rect 3148 21082 3200 21088
rect 3792 20392 3844 20398
rect 2884 20318 3188 20346
rect 3896 20380 3924 22607
rect 8574 22520 8630 23000
rect 14370 22520 14426 23000
rect 18970 22672 19026 22681
rect 18970 22607 19026 22616
rect 4250 21856 4306 21865
rect 4250 21791 4306 21800
rect 4066 20904 4122 20913
rect 4066 20839 4068 20848
rect 4120 20839 4122 20848
rect 4068 20810 4120 20816
rect 3976 20596 4028 20602
rect 3976 20538 4028 20544
rect 3988 20505 4016 20538
rect 4068 20528 4120 20534
rect 3974 20496 4030 20505
rect 4068 20470 4120 20476
rect 3974 20431 4030 20440
rect 3896 20352 4016 20380
rect 3792 20334 3844 20340
rect 1952 20256 2004 20262
rect 1952 20198 2004 20204
rect 2872 20256 2924 20262
rect 2872 20198 2924 20204
rect 1768 19916 1820 19922
rect 1768 19858 1820 19864
rect 1032 18692 1084 18698
rect 1032 18634 1084 18640
rect 1044 15065 1072 18634
rect 1780 17814 1808 19858
rect 1768 17808 1820 17814
rect 1964 17785 1992 20198
rect 2780 19712 2832 19718
rect 2780 19654 2832 19660
rect 2688 19304 2740 19310
rect 2688 19246 2740 19252
rect 2700 18970 2728 19246
rect 2688 18964 2740 18970
rect 2688 18906 2740 18912
rect 2792 18170 2820 19654
rect 2884 18601 2912 20198
rect 3056 19712 3108 19718
rect 3056 19654 3108 19660
rect 2964 19168 3016 19174
rect 2964 19110 3016 19116
rect 2870 18592 2926 18601
rect 2870 18527 2926 18536
rect 2792 18142 2912 18170
rect 2780 18080 2832 18086
rect 2780 18022 2832 18028
rect 1768 17750 1820 17756
rect 1950 17776 2006 17785
rect 1950 17711 2006 17720
rect 1768 17536 1820 17542
rect 1768 17478 1820 17484
rect 1492 17060 1544 17066
rect 1492 17002 1544 17008
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1030 15056 1086 15065
rect 1030 14991 1086 15000
rect 1308 8492 1360 8498
rect 1308 8434 1360 8440
rect 204 4752 256 4758
rect 204 4694 256 4700
rect 216 480 244 4694
rect 1124 3392 1176 3398
rect 1124 3334 1176 3340
rect 664 2848 716 2854
rect 664 2790 716 2796
rect 676 480 704 2790
rect 1136 480 1164 3334
rect 1320 649 1348 8434
rect 1412 7546 1440 15506
rect 1504 13870 1532 17002
rect 1584 15360 1636 15366
rect 1584 15302 1636 15308
rect 1492 13864 1544 13870
rect 1492 13806 1544 13812
rect 1400 7540 1452 7546
rect 1400 7482 1452 7488
rect 1596 7342 1624 15302
rect 1674 14648 1730 14657
rect 1674 14583 1730 14592
rect 1688 14074 1716 14583
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 1780 7410 1808 17478
rect 2792 16946 2820 18022
rect 2608 16918 2820 16946
rect 2412 16584 2464 16590
rect 2412 16526 2464 16532
rect 1952 16448 2004 16454
rect 1952 16390 2004 16396
rect 1964 16114 1992 16390
rect 1952 16108 2004 16114
rect 1952 16050 2004 16056
rect 2136 16108 2188 16114
rect 2136 16050 2188 16056
rect 1952 15904 2004 15910
rect 1952 15846 2004 15852
rect 2044 15904 2096 15910
rect 2044 15846 2096 15852
rect 1964 11694 1992 15846
rect 2056 15706 2084 15846
rect 2044 15700 2096 15706
rect 2044 15642 2096 15648
rect 2148 15026 2176 16050
rect 2424 15706 2452 16526
rect 2608 16522 2636 16918
rect 2884 16810 2912 18142
rect 2976 16833 3004 19110
rect 3068 18193 3096 19654
rect 3160 19174 3188 20318
rect 3332 20256 3384 20262
rect 3332 20198 3384 20204
rect 3240 19916 3292 19922
rect 3240 19858 3292 19864
rect 3148 19168 3200 19174
rect 3148 19110 3200 19116
rect 3054 18184 3110 18193
rect 3054 18119 3110 18128
rect 3148 17876 3200 17882
rect 3148 17818 3200 17824
rect 3056 17128 3108 17134
rect 3056 17070 3108 17076
rect 2700 16782 2912 16810
rect 2962 16824 3018 16833
rect 2596 16516 2648 16522
rect 2596 16458 2648 16464
rect 2700 16425 2728 16782
rect 2962 16759 3018 16768
rect 2780 16516 2832 16522
rect 2780 16458 2832 16464
rect 2686 16416 2742 16425
rect 2686 16351 2742 16360
rect 2596 16040 2648 16046
rect 2596 15982 2648 15988
rect 2412 15700 2464 15706
rect 2412 15642 2464 15648
rect 2608 15570 2636 15982
rect 2596 15564 2648 15570
rect 2596 15506 2648 15512
rect 2136 15020 2188 15026
rect 2136 14962 2188 14968
rect 2148 14414 2176 14962
rect 2228 14884 2280 14890
rect 2228 14826 2280 14832
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 2134 13288 2190 13297
rect 2134 13223 2190 13232
rect 1952 11688 2004 11694
rect 1952 11630 2004 11636
rect 1952 10124 2004 10130
rect 1952 10066 2004 10072
rect 1860 9376 1912 9382
rect 1860 9318 1912 9324
rect 1872 8430 1900 9318
rect 1860 8424 1912 8430
rect 1860 8366 1912 8372
rect 1964 8090 1992 10066
rect 2044 9920 2096 9926
rect 2044 9862 2096 9868
rect 2056 9518 2084 9862
rect 2044 9512 2096 9518
rect 2044 9454 2096 9460
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 2148 7546 2176 13223
rect 2240 10690 2268 14826
rect 2412 14272 2464 14278
rect 2412 14214 2464 14220
rect 2320 13388 2372 13394
rect 2320 13330 2372 13336
rect 2332 12986 2360 13330
rect 2320 12980 2372 12986
rect 2320 12922 2372 12928
rect 2424 12442 2452 14214
rect 2504 12708 2556 12714
rect 2504 12650 2556 12656
rect 2412 12436 2464 12442
rect 2412 12378 2464 12384
rect 2320 12096 2372 12102
rect 2320 12038 2372 12044
rect 2332 11762 2360 12038
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 2320 11756 2372 11762
rect 2320 11698 2372 11704
rect 2424 11626 2452 11834
rect 2412 11620 2464 11626
rect 2412 11562 2464 11568
rect 2516 11354 2544 12650
rect 2504 11348 2556 11354
rect 2504 11290 2556 11296
rect 2240 10662 2452 10690
rect 2228 10532 2280 10538
rect 2228 10474 2280 10480
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 1768 7404 1820 7410
rect 1768 7346 1820 7352
rect 2240 7342 2268 10474
rect 2320 9376 2372 9382
rect 2320 9318 2372 9324
rect 2332 8090 2360 9318
rect 2320 8084 2372 8090
rect 2320 8026 2372 8032
rect 2424 7970 2452 10662
rect 2332 7954 2452 7970
rect 2320 7948 2452 7954
rect 2372 7942 2452 7948
rect 2320 7890 2372 7896
rect 1584 7336 1636 7342
rect 1584 7278 1636 7284
rect 2228 7336 2280 7342
rect 2228 7278 2280 7284
rect 2332 7188 2360 7890
rect 2608 7886 2636 15506
rect 2792 13705 2820 16458
rect 3068 16250 3096 17070
rect 3056 16244 3108 16250
rect 3056 16186 3108 16192
rect 2964 16108 3016 16114
rect 2964 16050 3016 16056
rect 2976 15502 3004 16050
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 2872 15088 2924 15094
rect 2872 15030 2924 15036
rect 2778 13696 2834 13705
rect 2778 13631 2834 13640
rect 2884 13546 2912 15030
rect 3056 14816 3108 14822
rect 3056 14758 3108 14764
rect 2964 13796 3016 13802
rect 2964 13738 3016 13744
rect 2792 13518 2912 13546
rect 2688 12640 2740 12646
rect 2688 12582 2740 12588
rect 2700 12170 2728 12582
rect 2688 12164 2740 12170
rect 2688 12106 2740 12112
rect 2792 11354 2820 13518
rect 2976 12238 3004 13738
rect 2964 12232 3016 12238
rect 2964 12174 3016 12180
rect 2976 11762 3004 12174
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 2872 11688 2924 11694
rect 2872 11630 2924 11636
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2884 11286 2912 11630
rect 2872 11280 2924 11286
rect 2872 11222 2924 11228
rect 2976 11150 3004 11698
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2872 10600 2924 10606
rect 2872 10542 2924 10548
rect 2884 10130 2912 10542
rect 3068 10418 3096 14758
rect 3160 14482 3188 17818
rect 3148 14476 3200 14482
rect 3148 14418 3200 14424
rect 3146 14104 3202 14113
rect 3146 14039 3202 14048
rect 3160 12986 3188 14039
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 3148 12776 3200 12782
rect 3148 12718 3200 12724
rect 2976 10390 3096 10418
rect 2976 10305 3004 10390
rect 2962 10296 3018 10305
rect 3160 10282 3188 12718
rect 3252 10713 3280 19858
rect 3344 19553 3372 20198
rect 3330 19544 3386 19553
rect 3330 19479 3386 19488
rect 3516 19236 3568 19242
rect 3516 19178 3568 19184
rect 3332 18624 3384 18630
rect 3332 18566 3384 18572
rect 3344 15881 3372 18566
rect 3424 16788 3476 16794
rect 3424 16730 3476 16736
rect 3436 16046 3464 16730
rect 3424 16040 3476 16046
rect 3424 15982 3476 15988
rect 3424 15904 3476 15910
rect 3330 15872 3386 15881
rect 3424 15846 3476 15852
rect 3330 15807 3386 15816
rect 3332 14952 3384 14958
rect 3332 14894 3384 14900
rect 3344 14074 3372 14894
rect 3436 14618 3464 15846
rect 3528 15473 3556 19178
rect 3700 18760 3752 18766
rect 3700 18702 3752 18708
rect 3608 18148 3660 18154
rect 3608 18090 3660 18096
rect 3620 16114 3648 18090
rect 3608 16108 3660 16114
rect 3608 16050 3660 16056
rect 3712 15994 3740 18702
rect 3620 15966 3740 15994
rect 3514 15464 3570 15473
rect 3514 15399 3570 15408
rect 3424 14612 3476 14618
rect 3424 14554 3476 14560
rect 3332 14068 3384 14074
rect 3332 14010 3384 14016
rect 3332 13728 3384 13734
rect 3332 13670 3384 13676
rect 3344 12850 3372 13670
rect 3332 12844 3384 12850
rect 3332 12786 3384 12792
rect 3436 12782 3464 14554
rect 3516 14476 3568 14482
rect 3516 14418 3568 14424
rect 3424 12776 3476 12782
rect 3424 12718 3476 12724
rect 3528 12458 3556 14418
rect 3436 12430 3556 12458
rect 3436 11354 3464 12430
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3424 11212 3476 11218
rect 3424 11154 3476 11160
rect 3238 10704 3294 10713
rect 3238 10639 3294 10648
rect 3068 10266 3188 10282
rect 2962 10231 3018 10240
rect 3056 10260 3188 10266
rect 2872 10124 2924 10130
rect 2872 10066 2924 10072
rect 2976 9761 3004 10231
rect 3108 10254 3188 10260
rect 3056 10202 3108 10208
rect 2962 9752 3018 9761
rect 2962 9687 3018 9696
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 2780 9104 2832 9110
rect 2780 9046 2832 9052
rect 2792 8498 2820 9046
rect 2884 9042 2912 9522
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2596 7880 2648 7886
rect 2596 7822 2648 7828
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 2148 7160 2360 7188
rect 2042 6896 2098 6905
rect 2042 6831 2098 6840
rect 2056 6322 2084 6831
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 1676 6112 1728 6118
rect 1676 6054 1728 6060
rect 1952 6112 2004 6118
rect 1952 6054 2004 6060
rect 1584 4072 1636 4078
rect 1584 4014 1636 4020
rect 1596 3602 1624 4014
rect 1584 3596 1636 3602
rect 1584 3538 1636 3544
rect 1492 2984 1544 2990
rect 1596 2972 1624 3538
rect 1688 3505 1716 6054
rect 1964 5914 1992 6054
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 1768 5772 1820 5778
rect 1768 5714 1820 5720
rect 1674 3496 1730 3505
rect 1674 3431 1730 3440
rect 1544 2944 1624 2972
rect 1492 2926 1544 2932
rect 1504 2514 1532 2926
rect 1780 2854 1808 5714
rect 1768 2848 1820 2854
rect 1768 2790 1820 2796
rect 1780 2689 1808 2790
rect 1766 2680 1822 2689
rect 1766 2615 1822 2624
rect 2044 2576 2096 2582
rect 2044 2518 2096 2524
rect 1492 2508 1544 2514
rect 1492 2450 1544 2456
rect 1584 2100 1636 2106
rect 1584 2042 1636 2048
rect 1306 640 1362 649
rect 1306 575 1362 584
rect 1596 480 1624 2042
rect 2056 480 2084 2518
rect 2148 2417 2176 7160
rect 2228 6996 2280 7002
rect 2228 6938 2280 6944
rect 2240 6089 2268 6938
rect 2424 6916 2452 7822
rect 2884 7274 2912 7822
rect 2504 7268 2556 7274
rect 2504 7210 2556 7216
rect 2872 7268 2924 7274
rect 2872 7210 2924 7216
rect 2332 6888 2452 6916
rect 2226 6080 2282 6089
rect 2226 6015 2282 6024
rect 2226 2952 2282 2961
rect 2226 2887 2228 2896
rect 2280 2887 2282 2896
rect 2228 2858 2280 2864
rect 2332 2802 2360 6888
rect 2412 6656 2464 6662
rect 2412 6598 2464 6604
rect 2424 5001 2452 6598
rect 2516 6089 2544 7210
rect 2778 7168 2834 7177
rect 2778 7103 2834 7112
rect 2792 7002 2820 7103
rect 2780 6996 2832 7002
rect 2780 6938 2832 6944
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 2884 6769 2912 6802
rect 2964 6792 3016 6798
rect 2870 6760 2926 6769
rect 2964 6734 3016 6740
rect 2870 6695 2926 6704
rect 2596 6384 2648 6390
rect 2594 6352 2596 6361
rect 2648 6352 2650 6361
rect 2594 6287 2650 6296
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 2688 6112 2740 6118
rect 2502 6080 2558 6089
rect 2688 6054 2740 6060
rect 2502 6015 2558 6024
rect 2700 5710 2728 6054
rect 2688 5704 2740 5710
rect 2502 5672 2558 5681
rect 2688 5646 2740 5652
rect 2502 5607 2504 5616
rect 2556 5607 2558 5616
rect 2596 5636 2648 5642
rect 2504 5578 2556 5584
rect 2596 5578 2648 5584
rect 2410 4992 2466 5001
rect 2410 4927 2466 4936
rect 2608 4690 2636 5578
rect 2700 4826 2728 5646
rect 2688 4820 2740 4826
rect 2688 4762 2740 4768
rect 2596 4684 2648 4690
rect 2596 4626 2648 4632
rect 2240 2774 2360 2802
rect 2134 2408 2190 2417
rect 2134 2343 2190 2352
rect 2240 1465 2268 2774
rect 2608 2378 2636 4626
rect 2792 4078 2820 6258
rect 2976 6186 3004 6734
rect 2964 6180 3016 6186
rect 2964 6122 3016 6128
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 2884 4554 2912 5646
rect 2976 4622 3004 6122
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 2872 4548 2924 4554
rect 2872 4490 2924 4496
rect 2780 4072 2832 4078
rect 2976 4026 3004 4558
rect 2780 4014 2832 4020
rect 2884 4010 3004 4026
rect 2872 4004 3004 4010
rect 2924 3998 3004 4004
rect 2872 3946 2924 3952
rect 2976 3738 3004 3998
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 2976 3466 3004 3674
rect 2964 3460 3016 3466
rect 2964 3402 3016 3408
rect 3068 3369 3096 10202
rect 3252 9722 3280 10639
rect 3330 9752 3386 9761
rect 3240 9716 3292 9722
rect 3330 9687 3386 9696
rect 3240 9658 3292 9664
rect 3252 6066 3280 9658
rect 3344 6202 3372 9687
rect 3436 8634 3464 11154
rect 3620 9466 3648 15966
rect 3700 14408 3752 14414
rect 3700 14350 3752 14356
rect 3712 11762 3740 14350
rect 3804 11778 3832 20334
rect 3884 18080 3936 18086
rect 3884 18022 3936 18028
rect 3896 13326 3924 18022
rect 3988 15008 4016 20352
rect 4080 19961 4108 20470
rect 4066 19952 4122 19961
rect 4066 19887 4122 19896
rect 4160 19712 4212 19718
rect 4160 19654 4212 19660
rect 4066 19136 4122 19145
rect 4172 19122 4200 19654
rect 4122 19094 4200 19122
rect 4066 19071 4122 19080
rect 4068 18828 4120 18834
rect 4068 18770 4120 18776
rect 4080 18358 4108 18770
rect 4160 18624 4212 18630
rect 4160 18566 4212 18572
rect 4068 18352 4120 18358
rect 4068 18294 4120 18300
rect 4068 18080 4120 18086
rect 4068 18022 4120 18028
rect 4080 17134 4108 18022
rect 4172 17241 4200 18566
rect 4158 17232 4214 17241
rect 4158 17167 4214 17176
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 4080 16522 4108 17070
rect 4160 16788 4212 16794
rect 4160 16730 4212 16736
rect 4068 16516 4120 16522
rect 4068 16458 4120 16464
rect 4172 16046 4200 16730
rect 4160 16040 4212 16046
rect 4160 15982 4212 15988
rect 4160 15564 4212 15570
rect 4264 15552 4292 21791
rect 7656 21140 7708 21146
rect 7656 21082 7708 21088
rect 4421 20700 4717 20720
rect 4477 20698 4501 20700
rect 4557 20698 4581 20700
rect 4637 20698 4661 20700
rect 4499 20646 4501 20698
rect 4563 20646 4575 20698
rect 4637 20646 4639 20698
rect 4477 20644 4501 20646
rect 4557 20644 4581 20646
rect 4637 20644 4661 20646
rect 4421 20624 4717 20644
rect 5172 20392 5224 20398
rect 5172 20334 5224 20340
rect 7196 20392 7248 20398
rect 7196 20334 7248 20340
rect 7564 20392 7616 20398
rect 7564 20334 7616 20340
rect 4804 19712 4856 19718
rect 4804 19654 4856 19660
rect 4421 19612 4717 19632
rect 4477 19610 4501 19612
rect 4557 19610 4581 19612
rect 4637 19610 4661 19612
rect 4499 19558 4501 19610
rect 4563 19558 4575 19610
rect 4637 19558 4639 19610
rect 4477 19556 4501 19558
rect 4557 19556 4581 19558
rect 4637 19556 4661 19558
rect 4421 19536 4717 19556
rect 4816 19310 4844 19654
rect 5184 19378 5212 20334
rect 5448 20324 5500 20330
rect 5448 20266 5500 20272
rect 5172 19372 5224 19378
rect 5172 19314 5224 19320
rect 4804 19304 4856 19310
rect 4804 19246 4856 19252
rect 5172 18964 5224 18970
rect 5172 18906 5224 18912
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 4421 18524 4717 18544
rect 4477 18522 4501 18524
rect 4557 18522 4581 18524
rect 4637 18522 4661 18524
rect 4499 18470 4501 18522
rect 4563 18470 4575 18522
rect 4637 18470 4639 18522
rect 4477 18468 4501 18470
rect 4557 18468 4581 18470
rect 4637 18468 4661 18470
rect 4421 18448 4717 18468
rect 4816 18222 4844 18702
rect 4804 18216 4856 18222
rect 4804 18158 4856 18164
rect 4816 17678 4844 18158
rect 4896 17808 4948 17814
rect 4896 17750 4948 17756
rect 4804 17672 4856 17678
rect 4804 17614 4856 17620
rect 4421 17436 4717 17456
rect 4477 17434 4501 17436
rect 4557 17434 4581 17436
rect 4637 17434 4661 17436
rect 4499 17382 4501 17434
rect 4563 17382 4575 17434
rect 4637 17382 4639 17434
rect 4477 17380 4501 17382
rect 4557 17380 4581 17382
rect 4637 17380 4661 17382
rect 4421 17360 4717 17380
rect 4816 17066 4844 17614
rect 4804 17060 4856 17066
rect 4804 17002 4856 17008
rect 4908 16998 4936 17750
rect 4896 16992 4948 16998
rect 4896 16934 4948 16940
rect 4344 16652 4396 16658
rect 4344 16594 4396 16600
rect 4356 16250 4384 16594
rect 4421 16348 4717 16368
rect 4477 16346 4501 16348
rect 4557 16346 4581 16348
rect 4637 16346 4661 16348
rect 4499 16294 4501 16346
rect 4563 16294 4575 16346
rect 4637 16294 4639 16346
rect 4477 16292 4501 16294
rect 4557 16292 4581 16294
rect 4637 16292 4661 16294
rect 4421 16272 4717 16292
rect 4344 16244 4396 16250
rect 4344 16186 4396 16192
rect 4908 16114 4936 16934
rect 4896 16108 4948 16114
rect 4896 16050 4948 16056
rect 4896 15564 4948 15570
rect 4212 15524 4384 15552
rect 4160 15506 4212 15512
rect 3988 14980 4292 15008
rect 3976 14884 4028 14890
rect 3976 14826 4028 14832
rect 3988 14346 4016 14826
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 3976 14340 4028 14346
rect 3976 14282 4028 14288
rect 3988 13734 4016 14282
rect 4068 14272 4120 14278
rect 4068 14214 4120 14220
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3974 13560 4030 13569
rect 4080 13530 4108 14214
rect 3974 13495 4030 13504
rect 4068 13524 4120 13530
rect 3884 13320 3936 13326
rect 3884 13262 3936 13268
rect 3884 12368 3936 12374
rect 3884 12310 3936 12316
rect 3896 11937 3924 12310
rect 3882 11928 3938 11937
rect 3882 11863 3938 11872
rect 3700 11756 3752 11762
rect 3804 11750 3924 11778
rect 3700 11698 3752 11704
rect 3712 10606 3740 11698
rect 3792 11688 3844 11694
rect 3792 11630 3844 11636
rect 3804 11393 3832 11630
rect 3790 11384 3846 11393
rect 3790 11319 3846 11328
rect 3896 11234 3924 11750
rect 3804 11206 3924 11234
rect 3700 10600 3752 10606
rect 3700 10542 3752 10548
rect 3804 9704 3832 11206
rect 3884 11076 3936 11082
rect 3884 11018 3936 11024
rect 3896 10742 3924 11018
rect 3884 10736 3936 10742
rect 3884 10678 3936 10684
rect 3884 10124 3936 10130
rect 3884 10066 3936 10072
rect 3712 9676 3832 9704
rect 3712 9586 3740 9676
rect 3790 9616 3846 9625
rect 3700 9580 3752 9586
rect 3790 9551 3846 9560
rect 3700 9522 3752 9528
rect 3620 9450 3740 9466
rect 3804 9450 3832 9551
rect 3620 9444 3752 9450
rect 3620 9438 3700 9444
rect 3700 9386 3752 9392
rect 3792 9444 3844 9450
rect 3792 9386 3844 9392
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3620 9042 3648 9318
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 3608 9036 3660 9042
rect 3608 8978 3660 8984
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 3528 7546 3556 8978
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 3712 7313 3740 9386
rect 3896 8974 3924 10066
rect 3884 8968 3936 8974
rect 3884 8910 3936 8916
rect 3790 8256 3846 8265
rect 3790 8191 3846 8200
rect 3804 7750 3832 8191
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 3698 7304 3754 7313
rect 3698 7239 3754 7248
rect 3344 6174 3556 6202
rect 3252 6038 3464 6066
rect 3332 5636 3384 5642
rect 3332 5578 3384 5584
rect 3238 5264 3294 5273
rect 3238 5199 3294 5208
rect 3252 4758 3280 5199
rect 3240 4752 3292 4758
rect 3240 4694 3292 4700
rect 3148 4480 3200 4486
rect 3148 4422 3200 4428
rect 3160 4282 3188 4422
rect 3148 4276 3200 4282
rect 3148 4218 3200 4224
rect 3146 4040 3202 4049
rect 3344 4010 3372 5578
rect 3146 3975 3202 3984
rect 3332 4004 3384 4010
rect 3160 3602 3188 3975
rect 3332 3946 3384 3952
rect 3330 3632 3386 3641
rect 3148 3596 3200 3602
rect 3330 3567 3386 3576
rect 3148 3538 3200 3544
rect 3054 3360 3110 3369
rect 3054 3295 3110 3304
rect 3054 3224 3110 3233
rect 3054 3159 3110 3168
rect 2780 3120 2832 3126
rect 2778 3088 2780 3097
rect 2832 3088 2834 3097
rect 2778 3023 2834 3032
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 2596 2372 2648 2378
rect 2596 2314 2648 2320
rect 2780 2304 2832 2310
rect 2780 2246 2832 2252
rect 2596 2032 2648 2038
rect 2596 1974 2648 1980
rect 2226 1456 2282 1465
rect 2226 1391 2282 1400
rect 2608 480 2636 1974
rect 2792 1698 2820 2246
rect 2884 1970 2912 2586
rect 2872 1964 2924 1970
rect 2872 1906 2924 1912
rect 2780 1692 2832 1698
rect 2780 1634 2832 1640
rect 3068 480 3096 3159
rect 3160 2650 3188 3538
rect 3148 2644 3200 2650
rect 3148 2586 3200 2592
rect 3344 1902 3372 3567
rect 3436 2650 3464 6038
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 3424 2508 3476 2514
rect 3424 2450 3476 2456
rect 3332 1896 3384 1902
rect 3332 1838 3384 1844
rect 3436 1494 3464 2450
rect 3528 2009 3556 6174
rect 3608 6112 3660 6118
rect 3608 6054 3660 6060
rect 3620 4729 3648 6054
rect 3804 5234 3832 7686
rect 3896 7342 3924 8910
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 3896 6322 3924 7278
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 3882 5536 3938 5545
rect 3882 5471 3938 5480
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 3896 5166 3924 5471
rect 3884 5160 3936 5166
rect 3790 5128 3846 5137
rect 3884 5102 3936 5108
rect 3790 5063 3846 5072
rect 3700 5024 3752 5030
rect 3700 4966 3752 4972
rect 3606 4720 3662 4729
rect 3606 4655 3662 4664
rect 3608 3936 3660 3942
rect 3608 3878 3660 3884
rect 3620 3058 3648 3878
rect 3712 3641 3740 4966
rect 3804 4758 3832 5063
rect 3792 4752 3844 4758
rect 3792 4694 3844 4700
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3882 4584 3938 4593
rect 3698 3632 3754 3641
rect 3698 3567 3754 3576
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 3700 2508 3752 2514
rect 3700 2450 3752 2456
rect 3608 2440 3660 2446
rect 3608 2382 3660 2388
rect 3514 2000 3570 2009
rect 3514 1935 3570 1944
rect 3620 1766 3648 2382
rect 3608 1760 3660 1766
rect 3608 1702 3660 1708
rect 3712 1612 3740 2450
rect 3804 2038 3832 4558
rect 3988 4570 4016 13495
rect 4068 13466 4120 13472
rect 4066 12744 4122 12753
rect 4066 12679 4068 12688
rect 4120 12679 4122 12688
rect 4068 12650 4120 12656
rect 4066 12336 4122 12345
rect 4066 12271 4122 12280
rect 4080 12170 4108 12271
rect 4068 12164 4120 12170
rect 4068 12106 4120 12112
rect 4172 11830 4200 14350
rect 4264 13569 4292 14980
rect 4250 13560 4306 13569
rect 4250 13495 4306 13504
rect 4356 13308 4384 15524
rect 4896 15506 4948 15512
rect 4421 15260 4717 15280
rect 4477 15258 4501 15260
rect 4557 15258 4581 15260
rect 4637 15258 4661 15260
rect 4499 15206 4501 15258
rect 4563 15206 4575 15258
rect 4637 15206 4639 15258
rect 4477 15204 4501 15206
rect 4557 15204 4581 15206
rect 4637 15204 4661 15206
rect 4421 15184 4717 15204
rect 4908 14822 4936 15506
rect 4896 14816 4948 14822
rect 4896 14758 4948 14764
rect 4804 14476 4856 14482
rect 4804 14418 4856 14424
rect 4421 14172 4717 14192
rect 4477 14170 4501 14172
rect 4557 14170 4581 14172
rect 4637 14170 4661 14172
rect 4499 14118 4501 14170
rect 4563 14118 4575 14170
rect 4637 14118 4639 14170
rect 4477 14116 4501 14118
rect 4557 14116 4581 14118
rect 4637 14116 4661 14118
rect 4421 14096 4717 14116
rect 4816 14074 4844 14418
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4434 13968 4490 13977
rect 4434 13903 4490 13912
rect 4264 13280 4384 13308
rect 4160 11824 4212 11830
rect 4160 11766 4212 11772
rect 4264 11558 4292 13280
rect 4448 13172 4476 13903
rect 4908 13462 4936 14758
rect 4988 13728 5040 13734
rect 4988 13670 5040 13676
rect 4896 13456 4948 13462
rect 4896 13398 4948 13404
rect 4356 13144 4476 13172
rect 4356 11626 4384 13144
rect 4421 13084 4717 13104
rect 4477 13082 4501 13084
rect 4557 13082 4581 13084
rect 4637 13082 4661 13084
rect 4499 13030 4501 13082
rect 4563 13030 4575 13082
rect 4637 13030 4639 13082
rect 4477 13028 4501 13030
rect 4557 13028 4581 13030
rect 4637 13028 4661 13030
rect 4421 13008 4717 13028
rect 5000 12986 5028 13670
rect 4988 12980 5040 12986
rect 4988 12922 5040 12928
rect 4896 12640 4948 12646
rect 4896 12582 4948 12588
rect 4421 11996 4717 12016
rect 4477 11994 4501 11996
rect 4557 11994 4581 11996
rect 4637 11994 4661 11996
rect 4499 11942 4501 11994
rect 4563 11942 4575 11994
rect 4637 11942 4639 11994
rect 4477 11940 4501 11942
rect 4557 11940 4581 11942
rect 4637 11940 4661 11942
rect 4421 11920 4717 11940
rect 4908 11914 4936 12582
rect 5184 12238 5212 18906
rect 5356 17060 5408 17066
rect 5356 17002 5408 17008
rect 5368 16590 5396 17002
rect 5356 16584 5408 16590
rect 5356 16526 5408 16532
rect 5368 15706 5396 16526
rect 5356 15700 5408 15706
rect 5356 15642 5408 15648
rect 5368 14958 5396 15642
rect 5356 14952 5408 14958
rect 5356 14894 5408 14900
rect 5368 14414 5396 14894
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 5264 13864 5316 13870
rect 5264 13806 5316 13812
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 4816 11886 4936 11914
rect 4344 11620 4396 11626
rect 4344 11562 4396 11568
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4172 11370 4200 11494
rect 4068 11348 4120 11354
rect 4172 11342 4384 11370
rect 4068 11290 4120 11296
rect 4080 11234 4108 11290
rect 4080 11206 4200 11234
rect 4066 10568 4122 10577
rect 4066 10503 4068 10512
rect 4120 10503 4122 10512
rect 4068 10474 4120 10480
rect 4068 9716 4120 9722
rect 4068 9658 4120 9664
rect 4080 9382 4108 9658
rect 4172 9382 4200 11206
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 4264 9518 4292 10950
rect 4356 10577 4384 11342
rect 4421 10908 4717 10928
rect 4477 10906 4501 10908
rect 4557 10906 4581 10908
rect 4637 10906 4661 10908
rect 4499 10854 4501 10906
rect 4563 10854 4575 10906
rect 4637 10854 4639 10906
rect 4477 10852 4501 10854
rect 4557 10852 4581 10854
rect 4637 10852 4661 10854
rect 4421 10832 4717 10852
rect 4342 10568 4398 10577
rect 4342 10503 4398 10512
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 4066 9208 4122 9217
rect 4066 9143 4068 9152
rect 4120 9143 4122 9152
rect 4068 9114 4120 9120
rect 4066 8664 4122 8673
rect 4122 8622 4292 8650
rect 4066 8599 4122 8608
rect 4160 8356 4212 8362
rect 4160 8298 4212 8304
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 4080 7857 4108 8230
rect 4066 7848 4122 7857
rect 4066 7783 4122 7792
rect 4172 7546 4200 8298
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 4264 6866 4292 8622
rect 4356 8566 4384 9998
rect 4421 9820 4717 9840
rect 4477 9818 4501 9820
rect 4557 9818 4581 9820
rect 4637 9818 4661 9820
rect 4499 9766 4501 9818
rect 4563 9766 4575 9818
rect 4637 9766 4639 9818
rect 4477 9764 4501 9766
rect 4557 9764 4581 9766
rect 4637 9764 4661 9766
rect 4421 9744 4717 9764
rect 4421 8732 4717 8752
rect 4477 8730 4501 8732
rect 4557 8730 4581 8732
rect 4637 8730 4661 8732
rect 4499 8678 4501 8730
rect 4563 8678 4575 8730
rect 4637 8678 4639 8730
rect 4477 8676 4501 8678
rect 4557 8676 4581 8678
rect 4637 8676 4661 8678
rect 4421 8656 4717 8676
rect 4344 8560 4396 8566
rect 4396 8520 4476 8548
rect 4344 8502 4396 8508
rect 4344 8288 4396 8294
rect 4344 8230 4396 8236
rect 4356 7342 4384 8230
rect 4448 7886 4476 8520
rect 4816 8430 4844 11886
rect 5184 11778 5212 12174
rect 5276 11898 5304 13806
rect 5356 13456 5408 13462
rect 5356 13398 5408 13404
rect 5368 12646 5396 13398
rect 5356 12640 5408 12646
rect 5356 12582 5408 12588
rect 5460 12458 5488 20266
rect 5540 19916 5592 19922
rect 5540 19858 5592 19864
rect 5552 19514 5580 19858
rect 5632 19848 5684 19854
rect 5632 19790 5684 19796
rect 6736 19848 6788 19854
rect 6736 19790 6788 19796
rect 5540 19508 5592 19514
rect 5540 19450 5592 19456
rect 5540 19168 5592 19174
rect 5540 19110 5592 19116
rect 5552 16794 5580 19110
rect 5644 18426 5672 19790
rect 5724 19780 5776 19786
rect 5724 19722 5776 19728
rect 5632 18420 5684 18426
rect 5632 18362 5684 18368
rect 5736 18290 5764 19722
rect 5816 19372 5868 19378
rect 5816 19314 5868 19320
rect 5724 18284 5776 18290
rect 5724 18226 5776 18232
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 5540 16652 5592 16658
rect 5540 16594 5592 16600
rect 5552 15706 5580 16594
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 5828 13394 5856 19314
rect 6748 18970 6776 19790
rect 7104 19236 7156 19242
rect 7104 19178 7156 19184
rect 6736 18964 6788 18970
rect 6736 18906 6788 18912
rect 6736 18828 6788 18834
rect 6736 18770 6788 18776
rect 6644 17740 6696 17746
rect 6644 17682 6696 17688
rect 6092 17672 6144 17678
rect 6092 17614 6144 17620
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 6012 16658 6040 17138
rect 6000 16652 6052 16658
rect 6000 16594 6052 16600
rect 6012 15434 6040 16594
rect 6104 16454 6132 17614
rect 6368 17536 6420 17542
rect 6368 17478 6420 17484
rect 6092 16448 6144 16454
rect 6092 16390 6144 16396
rect 6000 15428 6052 15434
rect 6000 15370 6052 15376
rect 6104 15314 6132 16390
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 6012 15286 6132 15314
rect 5816 13388 5868 13394
rect 5816 13330 5868 13336
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5460 12442 5580 12458
rect 5460 12436 5592 12442
rect 5460 12430 5540 12436
rect 5540 12378 5592 12384
rect 5644 12322 5672 12786
rect 5460 12294 5672 12322
rect 5460 12170 5488 12294
rect 5448 12164 5500 12170
rect 5448 12106 5500 12112
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 5184 11750 5304 11778
rect 5460 11762 5488 12106
rect 4988 11620 5040 11626
rect 4988 11562 5040 11568
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4908 8498 4936 11494
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 4804 8424 4856 8430
rect 4804 8366 4856 8372
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 4421 7644 4717 7664
rect 4477 7642 4501 7644
rect 4557 7642 4581 7644
rect 4637 7642 4661 7644
rect 4499 7590 4501 7642
rect 4563 7590 4575 7642
rect 4637 7590 4639 7642
rect 4477 7588 4501 7590
rect 4557 7588 4581 7590
rect 4637 7588 4661 7590
rect 4421 7568 4717 7588
rect 4344 7336 4396 7342
rect 4344 7278 4396 7284
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 4421 6556 4717 6576
rect 4477 6554 4501 6556
rect 4557 6554 4581 6556
rect 4637 6554 4661 6556
rect 4499 6502 4501 6554
rect 4563 6502 4575 6554
rect 4637 6502 4639 6554
rect 4477 6500 4501 6502
rect 4557 6500 4581 6502
rect 4637 6500 4661 6502
rect 4421 6480 4717 6500
rect 4618 6352 4674 6361
rect 4528 6316 4580 6322
rect 4618 6287 4674 6296
rect 4528 6258 4580 6264
rect 4344 6248 4396 6254
rect 4344 6190 4396 6196
rect 4160 5908 4212 5914
rect 4160 5850 4212 5856
rect 4066 5128 4122 5137
rect 4066 5063 4068 5072
rect 4120 5063 4122 5072
rect 4068 5034 4120 5040
rect 4172 4808 4200 5850
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 4080 4780 4200 4808
rect 4080 4690 4108 4780
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 3988 4542 4108 4570
rect 3882 4519 3938 4528
rect 3896 3754 3924 4519
rect 3976 4480 4028 4486
rect 3976 4422 4028 4428
rect 3988 4321 4016 4422
rect 3974 4312 4030 4321
rect 4080 4282 4108 4542
rect 3974 4247 4030 4256
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 4066 3904 4122 3913
rect 4066 3839 4122 3848
rect 3896 3726 4016 3754
rect 3792 2032 3844 2038
rect 3792 1974 3844 1980
rect 3528 1584 3740 1612
rect 3424 1488 3476 1494
rect 3424 1430 3476 1436
rect 3528 480 3556 1584
rect 3988 480 4016 3726
rect 4080 2825 4108 3839
rect 4172 3738 4200 4626
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 4264 2922 4292 4966
rect 4356 4010 4384 6190
rect 4540 5710 4568 6258
rect 4632 6254 4660 6287
rect 4620 6248 4672 6254
rect 4620 6190 4672 6196
rect 4804 5772 4856 5778
rect 4804 5714 4856 5720
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4421 5468 4717 5488
rect 4477 5466 4501 5468
rect 4557 5466 4581 5468
rect 4637 5466 4661 5468
rect 4499 5414 4501 5466
rect 4563 5414 4575 5466
rect 4637 5414 4639 5466
rect 4477 5412 4501 5414
rect 4557 5412 4581 5414
rect 4637 5412 4661 5414
rect 4421 5392 4717 5412
rect 4816 5098 4844 5714
rect 4804 5092 4856 5098
rect 4804 5034 4856 5040
rect 4908 4826 4936 6938
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4421 4380 4717 4400
rect 4477 4378 4501 4380
rect 4557 4378 4581 4380
rect 4637 4378 4661 4380
rect 4499 4326 4501 4378
rect 4563 4326 4575 4378
rect 4637 4326 4639 4378
rect 4477 4324 4501 4326
rect 4557 4324 4581 4326
rect 4637 4324 4661 4326
rect 4421 4304 4717 4324
rect 4816 4282 4844 4558
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 4436 4072 4488 4078
rect 4434 4040 4436 4049
rect 4488 4040 4490 4049
rect 4344 4004 4396 4010
rect 4434 3975 4490 3984
rect 4344 3946 4396 3952
rect 4344 3732 4396 3738
rect 4344 3674 4396 3680
rect 4252 2916 4304 2922
rect 4252 2858 4304 2864
rect 4066 2816 4122 2825
rect 4066 2751 4122 2760
rect 4356 2088 4384 3674
rect 4421 3292 4717 3312
rect 4477 3290 4501 3292
rect 4557 3290 4581 3292
rect 4637 3290 4661 3292
rect 4499 3238 4501 3290
rect 4563 3238 4575 3290
rect 4637 3238 4639 3290
rect 4477 3236 4501 3238
rect 4557 3236 4581 3238
rect 4637 3236 4661 3238
rect 4421 3216 4717 3236
rect 4816 3058 4844 4218
rect 4896 4072 4948 4078
rect 4896 4014 4948 4020
rect 4908 3618 4936 4014
rect 5000 3738 5028 11562
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 5184 9654 5212 11154
rect 5172 9648 5224 9654
rect 5172 9590 5224 9596
rect 5172 9376 5224 9382
rect 5172 9318 5224 9324
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 5092 8634 5120 8774
rect 5080 8628 5132 8634
rect 5080 8570 5132 8576
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 5092 8401 5120 8434
rect 5078 8392 5134 8401
rect 5078 8327 5134 8336
rect 5184 6202 5212 9318
rect 5092 6174 5212 6202
rect 5092 3913 5120 6174
rect 5172 6112 5224 6118
rect 5172 6054 5224 6060
rect 5184 4554 5212 6054
rect 5276 5914 5304 11750
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5460 11354 5488 11698
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 6012 11234 6040 15286
rect 6092 13320 6144 13326
rect 6092 13262 6144 13268
rect 6104 12306 6132 13262
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 6012 11206 6132 11234
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 6000 11144 6052 11150
rect 6000 11086 6052 11092
rect 5540 11076 5592 11082
rect 5540 11018 5592 11024
rect 5552 10606 5580 11018
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5644 9722 5672 10406
rect 5828 10266 5856 11086
rect 5908 10736 5960 10742
rect 5908 10678 5960 10684
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 5920 10146 5948 10678
rect 5724 10124 5776 10130
rect 5724 10066 5776 10072
rect 5828 10118 5948 10146
rect 5736 9926 5764 10066
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 5632 9716 5684 9722
rect 5632 9658 5684 9664
rect 5736 9586 5764 9862
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5460 8838 5488 9522
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 5460 8022 5488 8774
rect 5448 8016 5500 8022
rect 5448 7958 5500 7964
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5460 6798 5488 7346
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5460 6118 5488 6734
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5276 5817 5304 5850
rect 5262 5808 5318 5817
rect 5262 5743 5318 5752
rect 5828 5681 5856 10118
rect 5906 10024 5962 10033
rect 6012 9994 6040 11086
rect 6104 10062 6132 11206
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 5906 9959 5962 9968
rect 6000 9988 6052 9994
rect 5920 7818 5948 9959
rect 6000 9930 6052 9936
rect 6092 8832 6144 8838
rect 6092 8774 6144 8780
rect 6104 8634 6132 8774
rect 6092 8628 6144 8634
rect 6092 8570 6144 8576
rect 6196 7834 6224 15506
rect 6380 14482 6408 17478
rect 6460 17060 6512 17066
rect 6460 17002 6512 17008
rect 6368 14476 6420 14482
rect 6368 14418 6420 14424
rect 6380 14074 6408 14418
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6276 14000 6328 14006
rect 6276 13942 6328 13948
rect 5908 7812 5960 7818
rect 5908 7754 5960 7760
rect 6104 7806 6224 7834
rect 5908 7268 5960 7274
rect 5908 7210 5960 7216
rect 5814 5672 5870 5681
rect 5264 5636 5316 5642
rect 5814 5607 5870 5616
rect 5264 5578 5316 5584
rect 5276 5234 5304 5578
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5264 5092 5316 5098
rect 5264 5034 5316 5040
rect 5172 4548 5224 4554
rect 5172 4490 5224 4496
rect 5172 3936 5224 3942
rect 5078 3904 5134 3913
rect 5172 3878 5224 3884
rect 5078 3839 5134 3848
rect 5184 3738 5212 3878
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5080 3664 5132 3670
rect 4908 3590 5028 3618
rect 5080 3606 5132 3612
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 4816 2582 4844 2994
rect 4804 2576 4856 2582
rect 4804 2518 4856 2524
rect 4421 2204 4717 2224
rect 4477 2202 4501 2204
rect 4557 2202 4581 2204
rect 4637 2202 4661 2204
rect 4499 2150 4501 2202
rect 4563 2150 4575 2202
rect 4637 2150 4639 2202
rect 4477 2148 4501 2150
rect 4557 2148 4581 2150
rect 4637 2148 4661 2150
rect 4421 2128 4717 2148
rect 4356 2060 4476 2088
rect 4448 480 4476 2060
rect 5000 480 5028 3590
rect 5092 3534 5120 3606
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 5170 3496 5226 3505
rect 5092 3126 5120 3470
rect 5170 3431 5226 3440
rect 5080 3120 5132 3126
rect 5080 3062 5132 3068
rect 5184 2854 5212 3431
rect 5276 3126 5304 5034
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5722 4992 5778 5001
rect 5460 4826 5488 4966
rect 5722 4927 5778 4936
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5368 3670 5396 4558
rect 5356 3664 5408 3670
rect 5356 3606 5408 3612
rect 5264 3120 5316 3126
rect 5264 3062 5316 3068
rect 5172 2848 5224 2854
rect 5172 2790 5224 2796
rect 5368 2106 5396 3606
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5460 2990 5488 3334
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 5446 2816 5502 2825
rect 5446 2751 5502 2760
rect 5356 2100 5408 2106
rect 5356 2042 5408 2048
rect 5460 480 5488 2751
rect 5552 2650 5580 2858
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 5644 2417 5672 3538
rect 5736 2990 5764 4927
rect 5816 4752 5868 4758
rect 5816 4694 5868 4700
rect 5724 2984 5776 2990
rect 5724 2926 5776 2932
rect 5828 2650 5856 4694
rect 5920 3924 5948 7210
rect 6000 5568 6052 5574
rect 6000 5510 6052 5516
rect 6012 4078 6040 5510
rect 6104 4146 6132 7806
rect 6288 7698 6316 13942
rect 6380 13326 6408 14010
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6380 11558 6408 12582
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6380 7954 6408 11494
rect 6472 10742 6500 17002
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 6564 15570 6592 16594
rect 6552 15564 6604 15570
rect 6552 15506 6604 15512
rect 6552 14272 6604 14278
rect 6552 14214 6604 14220
rect 6564 13734 6592 14214
rect 6656 13734 6684 17682
rect 6748 17066 6776 18770
rect 6920 18352 6972 18358
rect 6920 18294 6972 18300
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 6840 17338 6868 18158
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 6736 17060 6788 17066
rect 6736 17002 6788 17008
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6736 16720 6788 16726
rect 6736 16662 6788 16668
rect 6748 16250 6776 16662
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 6840 15706 6868 16934
rect 6828 15700 6880 15706
rect 6828 15642 6880 15648
rect 6826 15600 6882 15609
rect 6932 15570 6960 18294
rect 7116 17882 7144 19178
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 7208 17270 7236 20334
rect 7380 19916 7432 19922
rect 7380 19858 7432 19864
rect 7392 19378 7420 19858
rect 7380 19372 7432 19378
rect 7380 19314 7432 19320
rect 7392 18970 7420 19314
rect 7380 18964 7432 18970
rect 7380 18906 7432 18912
rect 7288 18624 7340 18630
rect 7288 18566 7340 18572
rect 7300 18222 7328 18566
rect 7392 18290 7420 18906
rect 7472 18828 7524 18834
rect 7472 18770 7524 18776
rect 7484 18426 7512 18770
rect 7472 18420 7524 18426
rect 7472 18362 7524 18368
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 7288 18216 7340 18222
rect 7288 18158 7340 18164
rect 7196 17264 7248 17270
rect 7196 17206 7248 17212
rect 7208 17066 7236 17206
rect 7196 17060 7248 17066
rect 7196 17002 7248 17008
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 7024 16114 7052 16390
rect 7012 16108 7064 16114
rect 7012 16050 7064 16056
rect 6826 15535 6882 15544
rect 6920 15564 6972 15570
rect 6552 13728 6604 13734
rect 6552 13670 6604 13676
rect 6644 13728 6696 13734
rect 6644 13670 6696 13676
rect 6564 13546 6592 13670
rect 6564 13518 6684 13546
rect 6552 13388 6604 13394
rect 6552 13330 6604 13336
rect 6460 10736 6512 10742
rect 6460 10678 6512 10684
rect 6460 10600 6512 10606
rect 6460 10542 6512 10548
rect 6368 7948 6420 7954
rect 6368 7890 6420 7896
rect 6196 7670 6316 7698
rect 6092 4140 6144 4146
rect 6092 4082 6144 4088
rect 6000 4072 6052 4078
rect 6000 4014 6052 4020
rect 5920 3896 6132 3924
rect 5908 3596 5960 3602
rect 5908 3538 5960 3544
rect 6000 3596 6052 3602
rect 6000 3538 6052 3544
rect 5920 3194 5948 3538
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 5908 2916 5960 2922
rect 5908 2858 5960 2864
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 5630 2408 5686 2417
rect 5920 2378 5948 2858
rect 5630 2343 5686 2352
rect 5908 2372 5960 2378
rect 5908 2314 5960 2320
rect 6012 2258 6040 3538
rect 6104 2514 6132 3896
rect 6196 2990 6224 7670
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6288 5953 6316 6598
rect 6274 5944 6330 5953
rect 6274 5879 6330 5888
rect 6380 5658 6408 7890
rect 6472 7886 6500 10542
rect 6564 10033 6592 13330
rect 6656 11218 6684 13518
rect 6736 12300 6788 12306
rect 6736 12242 6788 12248
rect 6748 11762 6776 12242
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6644 10056 6696 10062
rect 6550 10024 6606 10033
rect 6644 9998 6696 10004
rect 6550 9959 6606 9968
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 6564 9382 6592 9862
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6564 8090 6592 9318
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 6564 7886 6592 8026
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6472 7342 6500 7822
rect 6460 7336 6512 7342
rect 6460 7278 6512 7284
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6564 6934 6592 7142
rect 6460 6928 6512 6934
rect 6460 6870 6512 6876
rect 6552 6928 6604 6934
rect 6552 6870 6604 6876
rect 6288 5630 6408 5658
rect 6184 2984 6236 2990
rect 6184 2926 6236 2932
rect 6092 2508 6144 2514
rect 6092 2450 6144 2456
rect 5920 2230 6040 2258
rect 5920 480 5948 2230
rect 202 0 258 480
rect 662 0 718 480
rect 1122 0 1178 480
rect 1582 0 1638 480
rect 2042 0 2098 480
rect 2594 0 2650 480
rect 3054 0 3110 480
rect 3514 0 3570 480
rect 3608 332 3660 338
rect 3608 274 3660 280
rect 3620 241 3648 274
rect 3606 232 3662 241
rect 3606 167 3662 176
rect 3974 0 4030 480
rect 4434 0 4490 480
rect 4986 0 5042 480
rect 5446 0 5502 480
rect 5906 0 5962 480
rect 6288 338 6316 5630
rect 6368 5568 6420 5574
rect 6368 5510 6420 5516
rect 6380 5234 6408 5510
rect 6472 5234 6500 6870
rect 6656 5760 6684 9998
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6748 8906 6776 9386
rect 6736 8900 6788 8906
rect 6736 8842 6788 8848
rect 6840 7290 6868 15535
rect 6920 15506 6972 15512
rect 7024 15502 7052 16050
rect 7012 15496 7064 15502
rect 7012 15438 7064 15444
rect 6920 14884 6972 14890
rect 6920 14826 6972 14832
rect 7196 14884 7248 14890
rect 7196 14826 7248 14832
rect 6932 14414 6960 14826
rect 7208 14618 7236 14826
rect 7196 14612 7248 14618
rect 7196 14554 7248 14560
rect 6920 14408 6972 14414
rect 6920 14350 6972 14356
rect 6920 13796 6972 13802
rect 6920 13738 6972 13744
rect 6932 13530 6960 13738
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 7288 13728 7340 13734
rect 7288 13670 7340 13676
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 7012 13184 7064 13190
rect 7012 13126 7064 13132
rect 7024 12442 7052 13126
rect 7208 12986 7236 13670
rect 7300 13530 7328 13670
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 6932 11014 6960 12378
rect 7012 12232 7064 12238
rect 7012 12174 7064 12180
rect 7024 12050 7052 12174
rect 7116 12170 7144 12582
rect 7104 12164 7156 12170
rect 7104 12106 7156 12112
rect 7196 12164 7248 12170
rect 7196 12106 7248 12112
rect 7024 12022 7144 12050
rect 7012 11280 7064 11286
rect 7012 11222 7064 11228
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 7024 10130 7052 11222
rect 7116 10305 7144 12022
rect 7102 10296 7158 10305
rect 7102 10231 7158 10240
rect 7116 10198 7144 10231
rect 7104 10192 7156 10198
rect 7104 10134 7156 10140
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 7208 9466 7236 12106
rect 7300 11898 7328 12582
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7380 10532 7432 10538
rect 7380 10474 7432 10480
rect 7288 10192 7340 10198
rect 7286 10160 7288 10169
rect 7340 10160 7342 10169
rect 7286 10095 7342 10104
rect 7392 9994 7420 10474
rect 7380 9988 7432 9994
rect 7380 9930 7432 9936
rect 7392 9586 7420 9930
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7208 9438 7420 9466
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 6932 8974 6960 9318
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6932 8430 6960 8774
rect 7024 8566 7052 8978
rect 7012 8560 7064 8566
rect 7012 8502 7064 8508
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 6564 5732 6684 5760
rect 6748 7262 6868 7290
rect 6368 5228 6420 5234
rect 6368 5170 6420 5176
rect 6460 5228 6512 5234
rect 6460 5170 6512 5176
rect 6380 3618 6408 5170
rect 6380 3590 6500 3618
rect 6472 3534 6500 3590
rect 6460 3528 6512 3534
rect 6366 3496 6422 3505
rect 6460 3470 6512 3476
rect 6564 3482 6592 5732
rect 6642 5672 6698 5681
rect 6642 5607 6644 5616
rect 6696 5607 6698 5616
rect 6644 5578 6696 5584
rect 6644 4004 6696 4010
rect 6644 3946 6696 3952
rect 6656 3738 6684 3946
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6366 3431 6422 3440
rect 6380 3058 6408 3431
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 6368 2848 6420 2854
rect 6368 2790 6420 2796
rect 6380 480 6408 2790
rect 6472 2446 6500 3470
rect 6564 3454 6684 3482
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 6564 2990 6592 3334
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 6552 2304 6604 2310
rect 6552 2246 6604 2252
rect 6564 2106 6592 2246
rect 6552 2100 6604 2106
rect 6552 2042 6604 2048
rect 6656 1057 6684 3454
rect 6748 3194 6776 7262
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 6840 6798 6868 7142
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 6932 5030 6960 6190
rect 7024 5914 7052 6734
rect 7012 5908 7064 5914
rect 7012 5850 7064 5856
rect 7116 5794 7144 8434
rect 7208 8090 7236 9318
rect 7288 8356 7340 8362
rect 7288 8298 7340 8304
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 7208 7041 7236 7142
rect 7194 7032 7250 7041
rect 7194 6967 7250 6976
rect 7300 6916 7328 8298
rect 7392 7206 7420 9438
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 7024 5766 7144 5794
rect 7208 6888 7328 6916
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 6932 4434 6960 4626
rect 7024 4593 7052 5766
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 7010 4584 7066 4593
rect 7010 4519 7066 4528
rect 6932 4406 7052 4434
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 6642 1048 6698 1057
rect 6642 983 6698 992
rect 6840 480 6868 4082
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 6932 2650 6960 3878
rect 7024 3738 7052 4406
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 7116 3670 7144 4762
rect 7104 3664 7156 3670
rect 7104 3606 7156 3612
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 7208 2258 7236 6888
rect 7288 6724 7340 6730
rect 7288 6666 7340 6672
rect 7300 6458 7328 6666
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 7300 6254 7328 6394
rect 7288 6248 7340 6254
rect 7288 6190 7340 6196
rect 7286 6080 7342 6089
rect 7286 6015 7342 6024
rect 7300 2378 7328 6015
rect 7378 5944 7434 5953
rect 7378 5879 7434 5888
rect 7392 5846 7420 5879
rect 7380 5840 7432 5846
rect 7380 5782 7432 5788
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7392 4690 7420 4966
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7378 4176 7434 4185
rect 7378 4111 7434 4120
rect 7392 3466 7420 4111
rect 7380 3460 7432 3466
rect 7380 3402 7432 3408
rect 7378 3360 7434 3369
rect 7378 3295 7434 3304
rect 7392 2961 7420 3295
rect 7378 2952 7434 2961
rect 7378 2887 7434 2896
rect 7484 2854 7512 18362
rect 7576 13802 7604 20334
rect 7668 17202 7696 21082
rect 8208 20868 8260 20874
rect 8208 20810 8260 20816
rect 8220 20602 8248 20810
rect 8208 20596 8260 20602
rect 8208 20538 8260 20544
rect 8208 20460 8260 20466
rect 8208 20402 8260 20408
rect 7886 20156 8182 20176
rect 7942 20154 7966 20156
rect 8022 20154 8046 20156
rect 8102 20154 8126 20156
rect 7964 20102 7966 20154
rect 8028 20102 8040 20154
rect 8102 20102 8104 20154
rect 7942 20100 7966 20102
rect 8022 20100 8046 20102
rect 8102 20100 8126 20102
rect 7886 20080 8182 20100
rect 7886 19068 8182 19088
rect 7942 19066 7966 19068
rect 8022 19066 8046 19068
rect 8102 19066 8126 19068
rect 7964 19014 7966 19066
rect 8028 19014 8040 19066
rect 8102 19014 8104 19066
rect 7942 19012 7966 19014
rect 8022 19012 8046 19014
rect 8102 19012 8126 19014
rect 7886 18992 8182 19012
rect 8220 18970 8248 20402
rect 8588 19922 8616 22520
rect 9312 21344 9364 21350
rect 9312 21286 9364 21292
rect 8576 19916 8628 19922
rect 8576 19858 8628 19864
rect 8852 19304 8904 19310
rect 8852 19246 8904 19252
rect 8576 19236 8628 19242
rect 8576 19178 8628 19184
rect 8588 18970 8616 19178
rect 8760 19168 8812 19174
rect 8760 19110 8812 19116
rect 8208 18964 8260 18970
rect 8208 18906 8260 18912
rect 8576 18964 8628 18970
rect 8576 18906 8628 18912
rect 7748 18896 7800 18902
rect 7748 18838 7800 18844
rect 7760 17678 7788 18838
rect 8220 18630 8248 18906
rect 8208 18624 8260 18630
rect 8208 18566 8260 18572
rect 8392 18216 8444 18222
rect 8392 18158 8444 18164
rect 7886 17980 8182 18000
rect 7942 17978 7966 17980
rect 8022 17978 8046 17980
rect 8102 17978 8126 17980
rect 7964 17926 7966 17978
rect 8028 17926 8040 17978
rect 8102 17926 8104 17978
rect 7942 17924 7966 17926
rect 8022 17924 8046 17926
rect 8102 17924 8126 17926
rect 7886 17904 8182 17924
rect 7748 17672 7800 17678
rect 7748 17614 7800 17620
rect 7656 17196 7708 17202
rect 7656 17138 7708 17144
rect 8208 17060 8260 17066
rect 8208 17002 8260 17008
rect 7886 16892 8182 16912
rect 7942 16890 7966 16892
rect 8022 16890 8046 16892
rect 8102 16890 8126 16892
rect 7964 16838 7966 16890
rect 8028 16838 8040 16890
rect 8102 16838 8104 16890
rect 7942 16836 7966 16838
rect 8022 16836 8046 16838
rect 8102 16836 8126 16838
rect 7886 16816 8182 16836
rect 8220 16794 8248 17002
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 8208 16788 8260 16794
rect 8208 16730 8260 16736
rect 7886 15804 8182 15824
rect 7942 15802 7966 15804
rect 8022 15802 8046 15804
rect 8102 15802 8126 15804
rect 7964 15750 7966 15802
rect 8028 15750 8040 15802
rect 8102 15750 8104 15802
rect 7942 15748 7966 15750
rect 8022 15748 8046 15750
rect 8102 15748 8126 15750
rect 7886 15728 8182 15748
rect 8312 15706 8340 16934
rect 8404 16046 8432 18158
rect 8668 18148 8720 18154
rect 8668 18090 8720 18096
rect 8680 16590 8708 18090
rect 8668 16584 8720 16590
rect 8668 16526 8720 16532
rect 8680 16250 8708 16526
rect 8576 16244 8628 16250
rect 8576 16186 8628 16192
rect 8668 16244 8720 16250
rect 8668 16186 8720 16192
rect 8392 16040 8444 16046
rect 8444 16000 8524 16028
rect 8392 15982 8444 15988
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8300 15700 8352 15706
rect 8300 15642 8352 15648
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 7748 14816 7800 14822
rect 7748 14758 7800 14764
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 7564 13796 7616 13802
rect 7564 13738 7616 13744
rect 7668 13326 7696 14554
rect 7760 14482 7788 14758
rect 7886 14716 8182 14736
rect 7942 14714 7966 14716
rect 8022 14714 8046 14716
rect 8102 14714 8126 14716
rect 7964 14662 7966 14714
rect 8028 14662 8040 14714
rect 8102 14662 8104 14714
rect 7942 14660 7966 14662
rect 8022 14660 8046 14662
rect 8102 14660 8126 14662
rect 7886 14640 8182 14660
rect 7748 14476 7800 14482
rect 7748 14418 7800 14424
rect 8220 13938 8248 14758
rect 8312 14618 8340 15506
rect 8300 14612 8352 14618
rect 8300 14554 8352 14560
rect 8404 14498 8432 15846
rect 8496 15026 8524 16000
rect 8588 15434 8616 16186
rect 8680 15502 8708 16186
rect 8668 15496 8720 15502
rect 8668 15438 8720 15444
rect 8576 15428 8628 15434
rect 8576 15370 8628 15376
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 8312 14470 8432 14498
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 7748 13864 7800 13870
rect 7748 13806 7800 13812
rect 7760 13394 7788 13806
rect 8208 13796 8260 13802
rect 8208 13738 8260 13744
rect 7886 13628 8182 13648
rect 7942 13626 7966 13628
rect 8022 13626 8046 13628
rect 8102 13626 8126 13628
rect 7964 13574 7966 13626
rect 8028 13574 8040 13626
rect 8102 13574 8104 13626
rect 7942 13572 7966 13574
rect 8022 13572 8046 13574
rect 8102 13572 8126 13574
rect 7886 13552 8182 13572
rect 7748 13388 7800 13394
rect 7748 13330 7800 13336
rect 7656 13320 7708 13326
rect 7656 13262 7708 13268
rect 7668 12850 7696 13262
rect 7760 12986 7788 13330
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 7886 12540 8182 12560
rect 7942 12538 7966 12540
rect 8022 12538 8046 12540
rect 8102 12538 8126 12540
rect 7964 12486 7966 12538
rect 8028 12486 8040 12538
rect 8102 12486 8104 12538
rect 7942 12484 7966 12486
rect 8022 12484 8046 12486
rect 8102 12484 8126 12486
rect 7886 12464 8182 12484
rect 7656 12368 7708 12374
rect 7656 12310 7708 12316
rect 7564 11280 7616 11286
rect 7564 11222 7616 11228
rect 7576 10810 7604 11222
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 7562 10568 7618 10577
rect 7562 10503 7618 10512
rect 7576 8242 7604 10503
rect 7668 8362 7696 12310
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 7760 8566 7788 12174
rect 8220 11626 8248 13738
rect 8208 11620 8260 11626
rect 8208 11562 8260 11568
rect 7886 11452 8182 11472
rect 7942 11450 7966 11452
rect 8022 11450 8046 11452
rect 8102 11450 8126 11452
rect 7964 11398 7966 11450
rect 8028 11398 8040 11450
rect 8102 11398 8104 11450
rect 7942 11396 7966 11398
rect 8022 11396 8046 11398
rect 8102 11396 8126 11398
rect 7886 11376 8182 11396
rect 7838 11112 7894 11121
rect 7838 11047 7894 11056
rect 7852 10742 7880 11047
rect 7840 10736 7892 10742
rect 7840 10678 7892 10684
rect 7886 10364 8182 10384
rect 7942 10362 7966 10364
rect 8022 10362 8046 10364
rect 8102 10362 8126 10364
rect 7964 10310 7966 10362
rect 8028 10310 8040 10362
rect 8102 10310 8104 10362
rect 7942 10308 7966 10310
rect 8022 10308 8046 10310
rect 8102 10308 8126 10310
rect 7886 10288 8182 10308
rect 7886 9276 8182 9296
rect 7942 9274 7966 9276
rect 8022 9274 8046 9276
rect 8102 9274 8126 9276
rect 7964 9222 7966 9274
rect 8028 9222 8040 9274
rect 8102 9222 8104 9274
rect 7942 9220 7966 9222
rect 8022 9220 8046 9222
rect 8102 9220 8126 9222
rect 7886 9200 8182 9220
rect 8208 9104 8260 9110
rect 8208 9046 8260 9052
rect 7748 8560 7800 8566
rect 7748 8502 7800 8508
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 7656 8356 7708 8362
rect 7656 8298 7708 8304
rect 7576 8214 7696 8242
rect 7564 7200 7616 7206
rect 7562 7168 7564 7177
rect 7616 7168 7618 7177
rect 7562 7103 7618 7112
rect 7564 4752 7616 4758
rect 7564 4694 7616 4700
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 7470 2680 7526 2689
rect 7576 2666 7604 4694
rect 7526 2638 7604 2666
rect 7470 2615 7526 2624
rect 7484 2582 7512 2615
rect 7472 2576 7524 2582
rect 7472 2518 7524 2524
rect 7288 2372 7340 2378
rect 7288 2314 7340 2320
rect 7208 2230 7420 2258
rect 7392 480 7420 2230
rect 7668 1442 7696 8214
rect 7760 7936 7788 8366
rect 7886 8188 8182 8208
rect 7942 8186 7966 8188
rect 8022 8186 8046 8188
rect 8102 8186 8126 8188
rect 7964 8134 7966 8186
rect 8028 8134 8040 8186
rect 8102 8134 8104 8186
rect 7942 8132 7966 8134
rect 8022 8132 8046 8134
rect 8102 8132 8126 8134
rect 7886 8112 8182 8132
rect 7840 7948 7892 7954
rect 7760 7908 7840 7936
rect 7840 7890 7892 7896
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7760 7274 7788 7482
rect 7748 7268 7800 7274
rect 7748 7210 7800 7216
rect 7886 7100 8182 7120
rect 7942 7098 7966 7100
rect 8022 7098 8046 7100
rect 8102 7098 8126 7100
rect 7964 7046 7966 7098
rect 8028 7046 8040 7098
rect 8102 7046 8104 7098
rect 7942 7044 7966 7046
rect 8022 7044 8046 7046
rect 8102 7044 8126 7046
rect 7886 7024 8182 7044
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7760 5914 7788 6598
rect 7886 6012 8182 6032
rect 7942 6010 7966 6012
rect 8022 6010 8046 6012
rect 8102 6010 8126 6012
rect 7964 5958 7966 6010
rect 8028 5958 8040 6010
rect 8102 5958 8104 6010
rect 7942 5956 7966 5958
rect 8022 5956 8046 5958
rect 8102 5956 8126 5958
rect 7886 5936 8182 5956
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 7886 4924 8182 4944
rect 7942 4922 7966 4924
rect 8022 4922 8046 4924
rect 8102 4922 8126 4924
rect 7964 4870 7966 4922
rect 8028 4870 8040 4922
rect 8102 4870 8104 4922
rect 7942 4868 7966 4870
rect 8022 4868 8046 4870
rect 8102 4868 8126 4870
rect 7886 4848 8182 4868
rect 7930 4720 7986 4729
rect 8114 4720 8170 4729
rect 7986 4678 8114 4706
rect 7930 4655 7986 4664
rect 8114 4655 8170 4664
rect 7886 3836 8182 3856
rect 7942 3834 7966 3836
rect 8022 3834 8046 3836
rect 8102 3834 8126 3836
rect 7964 3782 7966 3834
rect 8028 3782 8040 3834
rect 8102 3782 8104 3834
rect 7942 3780 7966 3782
rect 8022 3780 8046 3782
rect 8102 3780 8126 3782
rect 7886 3760 8182 3780
rect 8220 3738 8248 9046
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 7748 3120 7800 3126
rect 7746 3088 7748 3097
rect 7800 3088 7802 3097
rect 7746 3023 7802 3032
rect 7746 2952 7802 2961
rect 7746 2887 7748 2896
rect 7800 2887 7802 2896
rect 7748 2858 7800 2864
rect 7886 2748 8182 2768
rect 7942 2746 7966 2748
rect 8022 2746 8046 2748
rect 8102 2746 8126 2748
rect 7964 2694 7966 2746
rect 8028 2694 8040 2746
rect 8102 2694 8104 2746
rect 7942 2692 7966 2694
rect 8022 2692 8046 2694
rect 8102 2692 8126 2694
rect 7886 2672 8182 2692
rect 7932 2508 7984 2514
rect 7932 2450 7984 2456
rect 8116 2508 8168 2514
rect 8116 2450 8168 2456
rect 7944 1630 7972 2450
rect 8128 1834 8156 2450
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 8220 2038 8248 2382
rect 8208 2032 8260 2038
rect 8208 1974 8260 1980
rect 8116 1828 8168 1834
rect 8116 1770 8168 1776
rect 7932 1624 7984 1630
rect 7932 1566 7984 1572
rect 7668 1414 7880 1442
rect 7852 480 7880 1414
rect 8312 480 8340 14470
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 8404 13530 8432 13670
rect 8496 13530 8524 14962
rect 8588 14414 8616 15370
rect 8576 14408 8628 14414
rect 8576 14350 8628 14356
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 8588 13326 8616 14350
rect 8772 13977 8800 19110
rect 8758 13968 8814 13977
rect 8758 13903 8814 13912
rect 8760 13796 8812 13802
rect 8760 13738 8812 13744
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 8484 12708 8536 12714
rect 8484 12650 8536 12656
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8404 8498 8432 12038
rect 8496 10266 8524 12650
rect 8680 11762 8708 13466
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 8588 10713 8616 10746
rect 8574 10704 8630 10713
rect 8574 10639 8630 10648
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8574 8392 8630 8401
rect 8574 8327 8630 8336
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8404 7002 8432 7686
rect 8484 7268 8536 7274
rect 8484 7210 8536 7216
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8496 6458 8524 7210
rect 8588 6458 8616 8327
rect 8484 6452 8536 6458
rect 8484 6394 8536 6400
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 8390 5808 8446 5817
rect 8390 5743 8392 5752
rect 8444 5743 8446 5752
rect 8392 5714 8444 5720
rect 8496 5710 8524 6394
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 8680 4010 8708 8774
rect 8576 4004 8628 4010
rect 8576 3946 8628 3952
rect 8668 4004 8720 4010
rect 8668 3946 8720 3952
rect 8392 3392 8444 3398
rect 8392 3334 8444 3340
rect 8404 2854 8432 3334
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 8496 2417 8524 2994
rect 8588 2514 8616 3946
rect 8668 3188 8720 3194
rect 8668 3130 8720 3136
rect 8576 2508 8628 2514
rect 8576 2450 8628 2456
rect 8680 2446 8708 3130
rect 8668 2440 8720 2446
rect 8482 2408 8538 2417
rect 8668 2382 8720 2388
rect 8482 2343 8538 2352
rect 8772 480 8800 13738
rect 8864 10577 8892 19246
rect 9128 17536 9180 17542
rect 9128 17478 9180 17484
rect 9036 17060 9088 17066
rect 9036 17002 9088 17008
rect 8944 16992 8996 16998
rect 8944 16934 8996 16940
rect 8956 15910 8984 16934
rect 9048 16726 9076 17002
rect 9036 16720 9088 16726
rect 9036 16662 9088 16668
rect 8944 15904 8996 15910
rect 8944 15846 8996 15852
rect 8944 14068 8996 14074
rect 8944 14010 8996 14016
rect 8956 13734 8984 14010
rect 9140 13802 9168 17478
rect 9220 16652 9272 16658
rect 9220 16594 9272 16600
rect 9128 13796 9180 13802
rect 9128 13738 9180 13744
rect 8944 13728 8996 13734
rect 8944 13670 8996 13676
rect 8850 10568 8906 10577
rect 8850 10503 8906 10512
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8864 8906 8892 10406
rect 8852 8900 8904 8906
rect 8852 8842 8904 8848
rect 8850 6760 8906 6769
rect 8850 6695 8906 6704
rect 8864 5846 8892 6695
rect 8852 5840 8904 5846
rect 8852 5782 8904 5788
rect 8850 5672 8906 5681
rect 8850 5607 8906 5616
rect 8864 2514 8892 5607
rect 8956 2825 8984 13670
rect 9232 12986 9260 16594
rect 9324 14482 9352 21286
rect 11352 20700 11648 20720
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11430 20646 11432 20698
rect 11494 20646 11506 20698
rect 11568 20646 11570 20698
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11352 20624 11648 20644
rect 13636 20528 13688 20534
rect 13636 20470 13688 20476
rect 12532 20460 12584 20466
rect 12532 20402 12584 20408
rect 12164 20324 12216 20330
rect 12164 20266 12216 20272
rect 10048 20256 10100 20262
rect 10048 20198 10100 20204
rect 11336 20256 11388 20262
rect 11336 20198 11388 20204
rect 10060 20058 10088 20198
rect 10048 20052 10100 20058
rect 10048 19994 10100 20000
rect 9680 19848 9732 19854
rect 9680 19790 9732 19796
rect 9692 18766 9720 19790
rect 11348 19786 11376 20198
rect 11888 19848 11940 19854
rect 11888 19790 11940 19796
rect 11336 19780 11388 19786
rect 11336 19722 11388 19728
rect 11352 19612 11648 19632
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11430 19558 11432 19610
rect 11494 19558 11506 19610
rect 11568 19558 11570 19610
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11352 19536 11648 19556
rect 10784 19372 10836 19378
rect 10784 19314 10836 19320
rect 10416 19236 10468 19242
rect 10416 19178 10468 19184
rect 10600 19236 10652 19242
rect 10600 19178 10652 19184
rect 10232 19168 10284 19174
rect 10230 19136 10232 19145
rect 10284 19136 10286 19145
rect 10230 19071 10286 19080
rect 10140 18964 10192 18970
rect 10140 18906 10192 18912
rect 9956 18828 10008 18834
rect 9956 18770 10008 18776
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9692 18222 9720 18702
rect 9680 18216 9732 18222
rect 9680 18158 9732 18164
rect 9772 18080 9824 18086
rect 9968 18068 9996 18770
rect 9824 18040 9996 18068
rect 9772 18022 9824 18028
rect 9784 17202 9812 18022
rect 9864 17264 9916 17270
rect 9864 17206 9916 17212
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 9876 16794 9904 17206
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 9692 15706 9720 16730
rect 10048 16652 10100 16658
rect 10048 16594 10100 16600
rect 9772 16516 9824 16522
rect 9772 16458 9824 16464
rect 9496 15700 9548 15706
rect 9496 15642 9548 15648
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9312 14476 9364 14482
rect 9312 14418 9364 14424
rect 9404 13932 9456 13938
rect 9404 13874 9456 13880
rect 9416 13530 9444 13874
rect 9508 13530 9536 15642
rect 9404 13524 9456 13530
rect 9404 13466 9456 13472
rect 9496 13524 9548 13530
rect 9496 13466 9548 13472
rect 9588 13320 9640 13326
rect 9588 13262 9640 13268
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9600 12850 9628 13262
rect 9588 12844 9640 12850
rect 9588 12786 9640 12792
rect 9036 12776 9088 12782
rect 9036 12718 9088 12724
rect 9048 10470 9076 12718
rect 9312 12708 9364 12714
rect 9312 12650 9364 12656
rect 9220 12640 9272 12646
rect 9220 12582 9272 12588
rect 9036 10464 9088 10470
rect 9036 10406 9088 10412
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 8942 2816 8998 2825
rect 8942 2751 8998 2760
rect 8852 2508 8904 2514
rect 8852 2450 8904 2456
rect 9048 1562 9076 8978
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 9140 8430 9168 8910
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 9140 7750 9168 8366
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 9140 7342 9168 7686
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9140 6254 9168 7278
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 9140 5030 9168 6190
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9140 2990 9168 4966
rect 9128 2984 9180 2990
rect 9128 2926 9180 2932
rect 9036 1556 9088 1562
rect 9036 1498 9088 1504
rect 9232 480 9260 12582
rect 9324 3602 9352 12650
rect 9784 11694 9812 16458
rect 10060 16250 10088 16594
rect 10048 16244 10100 16250
rect 10048 16186 10100 16192
rect 9862 16144 9918 16153
rect 9862 16079 9918 16088
rect 9876 14618 9904 16079
rect 10060 15706 10088 16186
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 10152 15026 10180 18906
rect 10232 18216 10284 18222
rect 10232 18158 10284 18164
rect 10140 15020 10192 15026
rect 10140 14962 10192 14968
rect 10048 14952 10100 14958
rect 10048 14894 10100 14900
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9968 12306 9996 14758
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9588 9648 9640 9654
rect 9588 9590 9640 9596
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9600 9330 9628 9590
rect 9692 9450 9720 10406
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9680 9444 9732 9450
rect 9680 9386 9732 9392
rect 9416 3670 9444 9318
rect 9600 9302 9720 9330
rect 9692 9081 9720 9302
rect 9678 9072 9734 9081
rect 9678 9007 9734 9016
rect 9784 8974 9812 10066
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9772 8356 9824 8362
rect 9772 8298 9824 8304
rect 9588 7948 9640 7954
rect 9588 7890 9640 7896
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9508 7546 9536 7686
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9600 7449 9628 7890
rect 9784 7546 9812 8298
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9586 7440 9642 7449
rect 9586 7375 9642 7384
rect 9586 7304 9642 7313
rect 9586 7239 9642 7248
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9508 5273 9536 7142
rect 9600 6662 9628 7239
rect 9772 6928 9824 6934
rect 9772 6870 9824 6876
rect 9588 6656 9640 6662
rect 9588 6598 9640 6604
rect 9600 5681 9628 6598
rect 9586 5672 9642 5681
rect 9586 5607 9642 5616
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 9494 5264 9550 5273
rect 9494 5199 9550 5208
rect 9600 5166 9628 5510
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9692 5273 9720 5306
rect 9678 5264 9734 5273
rect 9678 5199 9734 5208
rect 9496 5160 9548 5166
rect 9496 5102 9548 5108
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9508 4282 9536 5102
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9588 4548 9640 4554
rect 9588 4490 9640 4496
rect 9496 4276 9548 4282
rect 9496 4218 9548 4224
rect 9600 4214 9628 4490
rect 9588 4208 9640 4214
rect 9588 4150 9640 4156
rect 9404 3664 9456 3670
rect 9404 3606 9456 3612
rect 9312 3596 9364 3602
rect 9312 3538 9364 3544
rect 9310 3224 9366 3233
rect 9310 3159 9366 3168
rect 9324 2961 9352 3159
rect 9600 2990 9628 4150
rect 9588 2984 9640 2990
rect 9310 2952 9366 2961
rect 9588 2926 9640 2932
rect 9310 2887 9366 2896
rect 9692 2650 9720 4558
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9784 480 9812 6870
rect 9876 5545 9904 10406
rect 9968 10130 9996 10610
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9968 8634 9996 10066
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 10060 7954 10088 14894
rect 10140 12776 10192 12782
rect 10140 12718 10192 12724
rect 10152 7970 10180 12718
rect 10244 11540 10272 18158
rect 10428 17814 10456 19178
rect 10416 17808 10468 17814
rect 10416 17750 10468 17756
rect 10324 16448 10376 16454
rect 10324 16390 10376 16396
rect 10336 11694 10364 16390
rect 10416 15428 10468 15434
rect 10416 15370 10468 15376
rect 10428 15162 10456 15370
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 10508 15088 10560 15094
rect 10508 15030 10560 15036
rect 10416 15020 10468 15026
rect 10416 14962 10468 14968
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10244 11512 10364 11540
rect 10232 11076 10284 11082
rect 10232 11018 10284 11024
rect 10244 10606 10272 11018
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 10336 10554 10364 11512
rect 10428 11286 10456 14962
rect 10520 12102 10548 15030
rect 10612 14958 10640 19178
rect 10692 19168 10744 19174
rect 10692 19110 10744 19116
rect 10600 14952 10652 14958
rect 10600 14894 10652 14900
rect 10600 13796 10652 13802
rect 10600 13738 10652 13744
rect 10612 12918 10640 13738
rect 10600 12912 10652 12918
rect 10600 12854 10652 12860
rect 10704 12322 10732 19110
rect 10796 17678 10824 19314
rect 11900 19242 11928 19790
rect 11980 19780 12032 19786
rect 11980 19722 12032 19728
rect 11888 19236 11940 19242
rect 11888 19178 11940 19184
rect 11152 18896 11204 18902
rect 11152 18838 11204 18844
rect 11164 18290 11192 18838
rect 11900 18766 11928 19178
rect 11888 18760 11940 18766
rect 11888 18702 11940 18708
rect 11352 18524 11648 18544
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11430 18470 11432 18522
rect 11494 18470 11506 18522
rect 11568 18470 11570 18522
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11352 18448 11648 18468
rect 11152 18284 11204 18290
rect 11152 18226 11204 18232
rect 11152 18148 11204 18154
rect 11152 18090 11204 18096
rect 11164 17882 11192 18090
rect 11152 17876 11204 17882
rect 11152 17818 11204 17824
rect 10876 17740 10928 17746
rect 10876 17682 10928 17688
rect 10968 17740 11020 17746
rect 10968 17682 11020 17688
rect 10784 17672 10836 17678
rect 10784 17614 10836 17620
rect 10796 16454 10824 17614
rect 10784 16448 10836 16454
rect 10784 16390 10836 16396
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 10796 15706 10824 15846
rect 10784 15700 10836 15706
rect 10784 15642 10836 15648
rect 10784 13796 10836 13802
rect 10784 13738 10836 13744
rect 10796 12986 10824 13738
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 10612 12294 10732 12322
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 10612 11898 10640 12294
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 10416 11280 10468 11286
rect 10416 11222 10468 11228
rect 10612 10674 10640 11834
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10336 10526 10640 10554
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 10244 8090 10272 9522
rect 10324 9512 10376 9518
rect 10322 9480 10324 9489
rect 10376 9480 10378 9489
rect 10322 9415 10378 9424
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 10048 7948 10100 7954
rect 10152 7942 10272 7970
rect 10048 7890 10100 7896
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10152 7546 10180 7822
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 9968 6254 9996 6598
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 10060 5914 10088 6802
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 9956 5568 10008 5574
rect 9862 5536 9918 5545
rect 9956 5510 10008 5516
rect 9862 5471 9918 5480
rect 9968 5370 9996 5510
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 9956 5228 10008 5234
rect 9956 5170 10008 5176
rect 9864 5092 9916 5098
rect 9864 5034 9916 5040
rect 9876 4729 9904 5034
rect 9968 5001 9996 5170
rect 9954 4992 10010 5001
rect 9954 4927 10010 4936
rect 9862 4720 9918 4729
rect 9862 4655 9918 4664
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 9862 3904 9918 3913
rect 9862 3839 9918 3848
rect 9876 3738 9904 3839
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9864 3460 9916 3466
rect 9864 3402 9916 3408
rect 9876 2990 9904 3402
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 9968 2446 9996 4626
rect 10060 3398 10088 5714
rect 10152 5302 10180 6734
rect 10140 5296 10192 5302
rect 10140 5238 10192 5244
rect 10244 5234 10272 7942
rect 10336 7886 10364 8570
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10336 6458 10364 6734
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10428 6338 10456 10406
rect 10508 8016 10560 8022
rect 10508 7958 10560 7964
rect 10520 6780 10548 7958
rect 10612 6934 10640 10526
rect 10704 8022 10732 12174
rect 10888 11762 10916 17682
rect 10980 16522 11008 17682
rect 11704 17672 11756 17678
rect 11704 17614 11756 17620
rect 11352 17436 11648 17456
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11430 17382 11432 17434
rect 11494 17382 11506 17434
rect 11568 17382 11570 17434
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11352 17360 11648 17380
rect 11244 17196 11296 17202
rect 11244 17138 11296 17144
rect 11256 16658 11284 17138
rect 11716 17134 11744 17614
rect 11888 17536 11940 17542
rect 11888 17478 11940 17484
rect 11900 17338 11928 17478
rect 11796 17332 11848 17338
rect 11796 17274 11848 17280
rect 11888 17332 11940 17338
rect 11888 17274 11940 17280
rect 11704 17128 11756 17134
rect 11704 17070 11756 17076
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 10968 16516 11020 16522
rect 10968 16458 11020 16464
rect 10980 15473 11008 16458
rect 11256 16130 11284 16594
rect 11352 16348 11648 16368
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11430 16294 11432 16346
rect 11494 16294 11506 16346
rect 11568 16294 11570 16346
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11352 16272 11648 16292
rect 11256 16114 11468 16130
rect 11256 16108 11480 16114
rect 11256 16102 11428 16108
rect 11428 16050 11480 16056
rect 11060 15972 11112 15978
rect 11060 15914 11112 15920
rect 10966 15464 11022 15473
rect 10966 15399 11022 15408
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 10980 11082 11008 11630
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 11072 10742 11100 15914
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 11164 13530 11192 15846
rect 11440 15570 11468 16050
rect 11518 16008 11574 16017
rect 11518 15943 11520 15952
rect 11572 15943 11574 15952
rect 11520 15914 11572 15920
rect 11428 15564 11480 15570
rect 11428 15506 11480 15512
rect 11352 15260 11648 15280
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11430 15206 11432 15258
rect 11494 15206 11506 15258
rect 11568 15206 11570 15258
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11352 15184 11648 15204
rect 11336 14476 11388 14482
rect 11256 14436 11336 14464
rect 11256 13988 11284 14436
rect 11336 14418 11388 14424
rect 11352 14172 11648 14192
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11430 14118 11432 14170
rect 11494 14118 11506 14170
rect 11568 14118 11570 14170
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11352 14096 11648 14116
rect 11520 14000 11572 14006
rect 11256 13960 11520 13988
rect 11520 13942 11572 13948
rect 11152 13524 11204 13530
rect 11152 13466 11204 13472
rect 11532 13258 11560 13942
rect 11520 13252 11572 13258
rect 11520 13194 11572 13200
rect 11352 13084 11648 13104
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11430 13030 11432 13082
rect 11494 13030 11506 13082
rect 11568 13030 11570 13082
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11352 13008 11648 13028
rect 11242 12608 11298 12617
rect 11242 12543 11298 12552
rect 11256 12442 11284 12543
rect 11244 12436 11296 12442
rect 11244 12378 11296 12384
rect 11352 11996 11648 12016
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11430 11942 11432 11994
rect 11494 11942 11506 11994
rect 11568 11942 11570 11994
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11352 11920 11648 11940
rect 11716 11558 11744 16934
rect 11808 13190 11836 17274
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11900 15337 11928 15982
rect 11992 15978 12020 19722
rect 12176 19718 12204 20266
rect 12440 20256 12492 20262
rect 12440 20198 12492 20204
rect 12164 19712 12216 19718
rect 12164 19654 12216 19660
rect 12072 18896 12124 18902
rect 12072 18838 12124 18844
rect 12084 16794 12112 18838
rect 12176 18834 12204 19654
rect 12348 18896 12400 18902
rect 12348 18838 12400 18844
rect 12164 18828 12216 18834
rect 12164 18770 12216 18776
rect 12360 18086 12388 18838
rect 12452 18222 12480 20198
rect 12544 19922 12572 20402
rect 12624 20392 12676 20398
rect 12624 20334 12676 20340
rect 12532 19916 12584 19922
rect 12532 19858 12584 19864
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 12348 18080 12400 18086
rect 12348 18022 12400 18028
rect 12254 17232 12310 17241
rect 12254 17167 12310 17176
rect 12072 16788 12124 16794
rect 12072 16730 12124 16736
rect 12164 16448 12216 16454
rect 12164 16390 12216 16396
rect 11980 15972 12032 15978
rect 11980 15914 12032 15920
rect 11886 15328 11942 15337
rect 11886 15263 11942 15272
rect 11796 13184 11848 13190
rect 11796 13126 11848 13132
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11716 11286 11744 11494
rect 11704 11280 11756 11286
rect 11704 11222 11756 11228
rect 11352 10908 11648 10928
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11430 10854 11432 10906
rect 11494 10854 11506 10906
rect 11568 10854 11570 10906
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11352 10832 11648 10852
rect 11060 10736 11112 10742
rect 11060 10678 11112 10684
rect 11704 10668 11756 10674
rect 11704 10610 11756 10616
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 11426 10568 11482 10577
rect 10876 10532 10928 10538
rect 10876 10474 10928 10480
rect 10782 9072 10838 9081
rect 10782 9007 10838 9016
rect 10692 8016 10744 8022
rect 10692 7958 10744 7964
rect 10600 6928 10652 6934
rect 10600 6870 10652 6876
rect 10520 6752 10640 6780
rect 10336 6310 10456 6338
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 10140 5160 10192 5166
rect 10192 5108 10272 5114
rect 10140 5102 10272 5108
rect 10152 5086 10272 5102
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 10152 2378 10180 4558
rect 10244 4457 10272 5086
rect 10230 4448 10286 4457
rect 10230 4383 10286 4392
rect 10230 4176 10286 4185
rect 10230 4111 10286 4120
rect 10244 3942 10272 4111
rect 10232 3936 10284 3942
rect 10336 3913 10364 6310
rect 10508 5908 10560 5914
rect 10428 5868 10508 5896
rect 10232 3878 10284 3884
rect 10322 3904 10378 3913
rect 10322 3839 10378 3848
rect 10324 3528 10376 3534
rect 10244 3488 10324 3516
rect 10140 2372 10192 2378
rect 10140 2314 10192 2320
rect 10244 480 10272 3488
rect 10428 3516 10456 5868
rect 10508 5850 10560 5856
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 10520 4146 10548 5646
rect 10612 5114 10640 6752
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 10704 5914 10732 6190
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10704 5710 10732 5850
rect 10692 5704 10744 5710
rect 10692 5646 10744 5652
rect 10704 5234 10732 5646
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10612 5086 10732 5114
rect 10600 4480 10652 4486
rect 10600 4422 10652 4428
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10520 3602 10548 3878
rect 10612 3670 10640 4422
rect 10600 3664 10652 3670
rect 10600 3606 10652 3612
rect 10704 3618 10732 5086
rect 10796 5030 10824 9007
rect 10888 7018 10916 10474
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 11072 9586 11100 9862
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 11072 9110 11100 9522
rect 11164 9110 11192 10542
rect 11426 10503 11482 10512
rect 11440 10470 11468 10503
rect 11428 10464 11480 10470
rect 11428 10406 11480 10412
rect 11352 9820 11648 9840
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11430 9766 11432 9818
rect 11494 9766 11506 9818
rect 11568 9766 11570 9818
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11352 9744 11648 9764
rect 11244 9648 11296 9654
rect 11244 9590 11296 9596
rect 11060 9104 11112 9110
rect 11060 9046 11112 9052
rect 11152 9104 11204 9110
rect 11152 9046 11204 9052
rect 10966 8936 11022 8945
rect 10966 8871 11022 8880
rect 10980 7750 11008 8871
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 11060 7812 11112 7818
rect 11060 7754 11112 7760
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 11072 7342 11100 7754
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 11164 7206 11192 8026
rect 11256 7954 11284 9590
rect 11352 8732 11648 8752
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11430 8678 11432 8730
rect 11494 8678 11506 8730
rect 11568 8678 11570 8730
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11352 8656 11648 8676
rect 11520 8560 11572 8566
rect 11520 8502 11572 8508
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 11532 7886 11560 8502
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 11352 7644 11648 7664
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11430 7590 11432 7642
rect 11494 7590 11506 7642
rect 11568 7590 11570 7642
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11352 7568 11648 7588
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 10888 6990 11008 7018
rect 10876 6928 10928 6934
rect 10876 6870 10928 6876
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 10888 4146 10916 6870
rect 10980 5846 11008 6990
rect 11244 6724 11296 6730
rect 11244 6666 11296 6672
rect 10968 5840 11020 5846
rect 10968 5782 11020 5788
rect 10784 4140 10836 4146
rect 10784 4082 10836 4088
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 10796 3738 10824 4082
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 10508 3596 10560 3602
rect 10704 3590 10824 3618
rect 10508 3538 10560 3544
rect 10376 3488 10456 3516
rect 10324 3470 10376 3476
rect 10692 3392 10744 3398
rect 10692 3334 10744 3340
rect 10414 3224 10470 3233
rect 10704 3194 10732 3334
rect 10414 3159 10470 3168
rect 10692 3188 10744 3194
rect 10428 2650 10456 3159
rect 10692 3130 10744 3136
rect 10796 3074 10824 3590
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10888 3398 10916 3470
rect 10876 3392 10928 3398
rect 10876 3334 10928 3340
rect 10980 3233 11008 5782
rect 11256 5681 11284 6666
rect 11352 6556 11648 6576
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11430 6502 11432 6554
rect 11494 6502 11506 6554
rect 11568 6502 11570 6554
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11352 6480 11648 6500
rect 11610 6352 11666 6361
rect 11610 6287 11666 6296
rect 11242 5672 11298 5681
rect 11624 5642 11652 6287
rect 11716 6202 11744 10610
rect 11808 9217 11836 12922
rect 11794 9208 11850 9217
rect 11794 9143 11850 9152
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11808 8022 11836 8774
rect 11796 8016 11848 8022
rect 11796 7958 11848 7964
rect 11716 6174 11836 6202
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11242 5607 11298 5616
rect 11612 5636 11664 5642
rect 11612 5578 11664 5584
rect 11352 5468 11648 5488
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11430 5414 11432 5466
rect 11494 5414 11506 5466
rect 11568 5414 11570 5466
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11352 5392 11648 5412
rect 11058 5264 11114 5273
rect 11716 5234 11744 6054
rect 11058 5199 11114 5208
rect 11704 5228 11756 5234
rect 11072 4214 11100 5199
rect 11704 5170 11756 5176
rect 11152 5160 11204 5166
rect 11152 5102 11204 5108
rect 11164 4457 11192 5102
rect 11336 4684 11388 4690
rect 11256 4644 11336 4672
rect 11150 4448 11206 4457
rect 11150 4383 11206 4392
rect 11060 4208 11112 4214
rect 11060 4150 11112 4156
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 11072 3398 11100 3878
rect 11060 3392 11112 3398
rect 11060 3334 11112 3340
rect 10966 3224 11022 3233
rect 10966 3159 11022 3168
rect 10704 3046 10824 3074
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 10704 480 10732 3046
rect 11164 480 11192 3878
rect 11256 3466 11284 4644
rect 11336 4626 11388 4632
rect 11352 4380 11648 4400
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11430 4326 11432 4378
rect 11494 4326 11506 4378
rect 11568 4326 11570 4378
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11352 4304 11648 4324
rect 11808 3942 11836 6174
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11900 3754 11928 15263
rect 11992 12986 12020 15914
rect 12176 15502 12204 16390
rect 12072 15496 12124 15502
rect 12072 15438 12124 15444
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 12084 14498 12112 15438
rect 12268 15162 12296 17167
rect 12256 15156 12308 15162
rect 12256 15098 12308 15104
rect 12452 15094 12480 18158
rect 12636 17202 12664 20334
rect 13648 19922 13676 20470
rect 13912 20460 13964 20466
rect 13912 20402 13964 20408
rect 14004 20460 14056 20466
rect 14004 20402 14056 20408
rect 13636 19916 13688 19922
rect 13636 19858 13688 19864
rect 12808 19304 12860 19310
rect 12808 19246 12860 19252
rect 12716 19168 12768 19174
rect 12716 19110 12768 19116
rect 12728 18426 12756 19110
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 12716 18216 12768 18222
rect 12716 18158 12768 18164
rect 12728 17678 12756 18158
rect 12716 17672 12768 17678
rect 12716 17614 12768 17620
rect 12624 17196 12676 17202
rect 12624 17138 12676 17144
rect 12532 17128 12584 17134
rect 12532 17070 12584 17076
rect 12544 16726 12572 17070
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12532 16720 12584 16726
rect 12532 16662 12584 16668
rect 12636 16046 12664 16730
rect 12624 16040 12676 16046
rect 12624 15982 12676 15988
rect 12532 15564 12584 15570
rect 12532 15506 12584 15512
rect 12440 15088 12492 15094
rect 12440 15030 12492 15036
rect 12440 14884 12492 14890
rect 12440 14826 12492 14832
rect 12452 14618 12480 14826
rect 12544 14822 12572 15506
rect 12532 14816 12584 14822
rect 12532 14758 12584 14764
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12084 14470 12296 14498
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 12176 14278 12204 14350
rect 12164 14272 12216 14278
rect 12164 14214 12216 14220
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 12176 12646 12204 14214
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 11980 12368 12032 12374
rect 11980 12310 12032 12316
rect 11992 8294 12020 12310
rect 12268 12084 12296 14470
rect 12452 13938 12480 14554
rect 12530 14512 12586 14521
rect 12530 14447 12586 14456
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 12438 13832 12494 13841
rect 12438 13767 12494 13776
rect 12452 13410 12480 13767
rect 12360 13382 12480 13410
rect 12360 12209 12388 13382
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 12452 12986 12480 13262
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12544 12442 12572 14447
rect 12636 14414 12664 15982
rect 12624 14408 12676 14414
rect 12624 14350 12676 14356
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12636 13462 12664 14214
rect 12624 13456 12676 13462
rect 12624 13398 12676 13404
rect 12728 13410 12756 17614
rect 12820 13841 12848 19246
rect 12990 19136 13046 19145
rect 12990 19071 13046 19080
rect 12900 18624 12952 18630
rect 12900 18566 12952 18572
rect 12912 14414 12940 18566
rect 13004 18154 13032 19071
rect 13648 18970 13676 19858
rect 13924 19718 13952 20402
rect 13912 19712 13964 19718
rect 13912 19654 13964 19660
rect 13924 19242 13952 19654
rect 13912 19236 13964 19242
rect 13912 19178 13964 19184
rect 13636 18964 13688 18970
rect 13636 18906 13688 18912
rect 13924 18766 13952 19178
rect 14016 18834 14044 20402
rect 14384 19990 14412 22520
rect 18050 20904 18106 20913
rect 18050 20839 18106 20848
rect 18064 20602 18092 20839
rect 18282 20700 18578 20720
rect 18338 20698 18362 20700
rect 18418 20698 18442 20700
rect 18498 20698 18522 20700
rect 18360 20646 18362 20698
rect 18424 20646 18436 20698
rect 18498 20646 18500 20698
rect 18338 20644 18362 20646
rect 18418 20644 18442 20646
rect 18498 20644 18522 20646
rect 18282 20624 18578 20644
rect 18052 20596 18104 20602
rect 18052 20538 18104 20544
rect 18144 20528 18196 20534
rect 18144 20470 18196 20476
rect 18236 20528 18288 20534
rect 18236 20470 18288 20476
rect 17224 20392 17276 20398
rect 17224 20334 17276 20340
rect 17958 20360 18014 20369
rect 15200 20256 15252 20262
rect 15200 20198 15252 20204
rect 15844 20256 15896 20262
rect 15844 20198 15896 20204
rect 14817 20156 15113 20176
rect 14873 20154 14897 20156
rect 14953 20154 14977 20156
rect 15033 20154 15057 20156
rect 14895 20102 14897 20154
rect 14959 20102 14971 20154
rect 15033 20102 15035 20154
rect 14873 20100 14897 20102
rect 14953 20100 14977 20102
rect 15033 20100 15057 20102
rect 14817 20080 15113 20100
rect 14372 19984 14424 19990
rect 14372 19926 14424 19932
rect 15212 19310 15240 20198
rect 15660 19984 15712 19990
rect 15660 19926 15712 19932
rect 15384 19916 15436 19922
rect 15384 19858 15436 19864
rect 15396 19378 15424 19858
rect 15384 19372 15436 19378
rect 15384 19314 15436 19320
rect 15200 19304 15252 19310
rect 15200 19246 15252 19252
rect 15292 19236 15344 19242
rect 15292 19178 15344 19184
rect 14817 19068 15113 19088
rect 14873 19066 14897 19068
rect 14953 19066 14977 19068
rect 15033 19066 15057 19068
rect 14895 19014 14897 19066
rect 14959 19014 14971 19066
rect 15033 19014 15035 19066
rect 14873 19012 14897 19014
rect 14953 19012 14977 19014
rect 15033 19012 15057 19014
rect 14817 18992 15113 19012
rect 15304 18970 15332 19178
rect 15396 19174 15424 19314
rect 15384 19168 15436 19174
rect 15384 19110 15436 19116
rect 15292 18964 15344 18970
rect 15292 18906 15344 18912
rect 14004 18828 14056 18834
rect 14004 18770 14056 18776
rect 13912 18760 13964 18766
rect 13912 18702 13964 18708
rect 13820 18352 13872 18358
rect 13820 18294 13872 18300
rect 12992 18148 13044 18154
rect 12992 18090 13044 18096
rect 13268 18080 13320 18086
rect 13268 18022 13320 18028
rect 13176 17740 13228 17746
rect 13176 17682 13228 17688
rect 12992 17536 13044 17542
rect 12992 17478 13044 17484
rect 12900 14408 12952 14414
rect 12900 14350 12952 14356
rect 12900 14000 12952 14006
rect 12900 13942 12952 13948
rect 12806 13832 12862 13841
rect 12806 13767 12862 13776
rect 12912 13734 12940 13942
rect 12808 13728 12860 13734
rect 12808 13670 12860 13676
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12820 13530 12848 13670
rect 13004 13530 13032 17478
rect 13188 17202 13216 17682
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 13176 16448 13228 16454
rect 13176 16390 13228 16396
rect 13188 16046 13216 16390
rect 13176 16040 13228 16046
rect 13176 15982 13228 15988
rect 13084 15088 13136 15094
rect 13136 15048 13216 15076
rect 13084 15030 13136 15036
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12992 13524 13044 13530
rect 12992 13466 13044 13472
rect 12728 13382 12848 13410
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 12728 12850 12756 12922
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12624 12776 12676 12782
rect 12624 12718 12676 12724
rect 12714 12744 12770 12753
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12346 12200 12402 12209
rect 12636 12186 12664 12718
rect 12714 12679 12770 12688
rect 12346 12135 12402 12144
rect 12452 12158 12664 12186
rect 12268 12056 12388 12084
rect 12072 11280 12124 11286
rect 12072 11222 12124 11228
rect 11980 8288 12032 8294
rect 11980 8230 12032 8236
rect 11980 8016 12032 8022
rect 11980 7958 12032 7964
rect 11992 7857 12020 7958
rect 11978 7848 12034 7857
rect 11978 7783 12034 7792
rect 11980 6248 12032 6254
rect 11980 6190 12032 6196
rect 11992 5710 12020 6190
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 11992 4690 12020 5646
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 11716 3726 11928 3754
rect 11244 3460 11296 3466
rect 11244 3402 11296 3408
rect 11352 3292 11648 3312
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11430 3238 11432 3290
rect 11494 3238 11506 3290
rect 11568 3238 11570 3290
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11352 3216 11648 3236
rect 11428 2916 11480 2922
rect 11428 2858 11480 2864
rect 11440 2514 11468 2858
rect 11428 2508 11480 2514
rect 11428 2450 11480 2456
rect 11352 2204 11648 2224
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11430 2150 11432 2202
rect 11494 2150 11506 2202
rect 11568 2150 11570 2202
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11352 2128 11648 2148
rect 11716 480 11744 3726
rect 11794 3632 11850 3641
rect 11794 3567 11850 3576
rect 11808 3369 11836 3567
rect 11794 3360 11850 3369
rect 11794 3295 11850 3304
rect 12084 1952 12112 11222
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 12268 9908 12296 11086
rect 12360 10010 12388 12056
rect 12452 11898 12480 12158
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12452 11354 12480 11834
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12544 10062 12572 12038
rect 12636 11830 12664 12038
rect 12624 11824 12676 11830
rect 12624 11766 12676 11772
rect 12636 11286 12664 11766
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12532 10056 12584 10062
rect 12360 9982 12480 10010
rect 12532 9998 12584 10004
rect 12268 9880 12388 9908
rect 12162 9752 12218 9761
rect 12162 9687 12218 9696
rect 12176 9450 12204 9687
rect 12360 9518 12388 9880
rect 12452 9874 12480 9982
rect 12636 9897 12664 10746
rect 12622 9888 12678 9897
rect 12452 9846 12572 9874
rect 12440 9716 12492 9722
rect 12440 9658 12492 9664
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12164 9444 12216 9450
rect 12164 9386 12216 9392
rect 12360 8974 12388 9454
rect 12452 9178 12480 9658
rect 12440 9172 12492 9178
rect 12440 9114 12492 9120
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12256 8832 12308 8838
rect 12256 8774 12308 8780
rect 12268 8430 12296 8774
rect 12360 8566 12388 8910
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12348 8560 12400 8566
rect 12348 8502 12400 8508
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 12176 7750 12204 8230
rect 12164 7744 12216 7750
rect 12164 7686 12216 7692
rect 12162 7304 12218 7313
rect 12162 7239 12164 7248
rect 12216 7239 12218 7248
rect 12164 7210 12216 7216
rect 12254 7168 12310 7177
rect 12254 7103 12310 7112
rect 12268 7002 12296 7103
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 12164 6928 12216 6934
rect 12162 6896 12164 6905
rect 12216 6896 12218 6905
rect 12162 6831 12218 6840
rect 12162 6760 12218 6769
rect 12162 6695 12218 6704
rect 12176 3194 12204 6695
rect 12360 6254 12388 8502
rect 12452 6866 12480 8570
rect 12544 7993 12572 9846
rect 12622 9823 12678 9832
rect 12530 7984 12586 7993
rect 12530 7919 12586 7928
rect 12544 7478 12572 7919
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12532 7472 12584 7478
rect 12532 7414 12584 7420
rect 12636 7002 12664 7482
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 12532 6928 12584 6934
rect 12530 6896 12532 6905
rect 12584 6896 12586 6905
rect 12440 6860 12492 6866
rect 12530 6831 12586 6840
rect 12440 6802 12492 6808
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12636 6458 12664 6734
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 12636 5778 12664 6394
rect 12624 5772 12676 5778
rect 12624 5714 12676 5720
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 12544 4078 12572 4558
rect 12624 4208 12676 4214
rect 12624 4150 12676 4156
rect 12532 4072 12584 4078
rect 12532 4014 12584 4020
rect 12348 4004 12400 4010
rect 12348 3946 12400 3952
rect 12164 3188 12216 3194
rect 12164 3130 12216 3136
rect 12084 1924 12204 1952
rect 12176 480 12204 1924
rect 12360 1358 12388 3946
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12452 2650 12480 3878
rect 12636 3534 12664 4150
rect 12624 3528 12676 3534
rect 12624 3470 12676 3476
rect 12440 2644 12492 2650
rect 12728 2632 12756 12679
rect 12820 12102 12848 13382
rect 12900 13388 12952 13394
rect 12900 13330 12952 13336
rect 12912 12850 12940 13330
rect 13084 12912 13136 12918
rect 13084 12854 13136 12860
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12912 12753 12940 12786
rect 12898 12744 12954 12753
rect 12898 12679 12954 12688
rect 12992 12708 13044 12714
rect 12992 12650 13044 12656
rect 12900 12640 12952 12646
rect 12900 12582 12952 12588
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12806 11928 12862 11937
rect 12806 11863 12862 11872
rect 12820 9450 12848 11863
rect 12912 11762 12940 12582
rect 12900 11756 12952 11762
rect 12900 11698 12952 11704
rect 12900 11348 12952 11354
rect 12900 11290 12952 11296
rect 12808 9444 12860 9450
rect 12808 9386 12860 9392
rect 12912 9042 12940 11290
rect 13004 9382 13032 12650
rect 13096 10130 13124 12854
rect 13084 10124 13136 10130
rect 13084 10066 13136 10072
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 12808 9036 12860 9042
rect 12808 8978 12860 8984
rect 12900 9036 12952 9042
rect 12900 8978 12952 8984
rect 12820 8634 12848 8978
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 12912 7750 12940 8434
rect 13084 7880 13136 7886
rect 12990 7848 13046 7857
rect 13084 7822 13136 7828
rect 12990 7783 13046 7792
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 12912 6186 12940 7686
rect 13004 7478 13032 7783
rect 12992 7472 13044 7478
rect 12992 7414 13044 7420
rect 13096 7206 13124 7822
rect 13084 7200 13136 7206
rect 13084 7142 13136 7148
rect 12900 6180 12952 6186
rect 12900 6122 12952 6128
rect 12992 6180 13044 6186
rect 12992 6122 13044 6128
rect 12900 5568 12952 5574
rect 12900 5510 12952 5516
rect 12912 5302 12940 5510
rect 12900 5296 12952 5302
rect 12900 5238 12952 5244
rect 13004 5001 13032 6122
rect 12990 4992 13046 5001
rect 12990 4927 13046 4936
rect 13096 4706 13124 7142
rect 12820 4690 13124 4706
rect 12808 4684 13124 4690
rect 12860 4678 13124 4684
rect 12808 4626 12860 4632
rect 13188 4604 13216 15048
rect 13280 14634 13308 18022
rect 13832 17882 13860 18294
rect 13912 18148 13964 18154
rect 13912 18090 13964 18096
rect 13820 17876 13872 17882
rect 13820 17818 13872 17824
rect 13728 16992 13780 16998
rect 13728 16934 13780 16940
rect 13740 16794 13768 16934
rect 13360 16788 13412 16794
rect 13360 16730 13412 16736
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 13372 14770 13400 16730
rect 13544 16720 13596 16726
rect 13544 16662 13596 16668
rect 13452 16652 13504 16658
rect 13452 16594 13504 16600
rect 13464 15434 13492 16594
rect 13556 16266 13584 16662
rect 13556 16238 13860 16266
rect 13544 15564 13596 15570
rect 13544 15506 13596 15512
rect 13452 15428 13504 15434
rect 13452 15370 13504 15376
rect 13556 15337 13584 15506
rect 13542 15328 13598 15337
rect 13542 15263 13598 15272
rect 13372 14742 13676 14770
rect 13280 14606 13584 14634
rect 13268 14408 13320 14414
rect 13268 14350 13320 14356
rect 13280 8362 13308 14350
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13360 13524 13412 13530
rect 13360 13466 13412 13472
rect 13372 12374 13400 13466
rect 13464 12850 13492 14214
rect 13452 12844 13504 12850
rect 13452 12786 13504 12792
rect 13450 12472 13506 12481
rect 13556 12442 13584 14606
rect 13450 12407 13506 12416
rect 13544 12436 13596 12442
rect 13360 12368 13412 12374
rect 13360 12310 13412 12316
rect 13268 8356 13320 8362
rect 13268 8298 13320 8304
rect 13268 6996 13320 7002
rect 13268 6938 13320 6944
rect 13280 4826 13308 6938
rect 13360 5568 13412 5574
rect 13360 5510 13412 5516
rect 13268 4820 13320 4826
rect 13268 4762 13320 4768
rect 13372 4758 13400 5510
rect 13464 4865 13492 12407
rect 13544 12378 13596 12384
rect 13648 10554 13676 14742
rect 13832 14482 13860 16238
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13740 12986 13768 14010
rect 13832 12986 13860 14418
rect 13924 13870 13952 18090
rect 14016 15892 14044 18770
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 14372 18080 14424 18086
rect 14372 18022 14424 18028
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14108 17338 14136 17614
rect 14096 17332 14148 17338
rect 14096 17274 14148 17280
rect 14280 17196 14332 17202
rect 14280 17138 14332 17144
rect 14188 16992 14240 16998
rect 14188 16934 14240 16940
rect 14200 16794 14228 16934
rect 14188 16788 14240 16794
rect 14188 16730 14240 16736
rect 14292 16674 14320 17138
rect 14200 16646 14320 16674
rect 14200 16046 14228 16646
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14292 16182 14320 16526
rect 14280 16176 14332 16182
rect 14280 16118 14332 16124
rect 14188 16040 14240 16046
rect 14188 15982 14240 15988
rect 14016 15864 14320 15892
rect 13912 13864 13964 13870
rect 13912 13806 13964 13812
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 13728 12980 13780 12986
rect 13728 12922 13780 12928
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13740 12481 13768 12922
rect 13820 12640 13872 12646
rect 13818 12608 13820 12617
rect 13872 12608 13874 12617
rect 13818 12543 13874 12552
rect 13726 12472 13782 12481
rect 13726 12407 13782 12416
rect 13924 12170 13952 13330
rect 14188 12300 14240 12306
rect 14188 12242 14240 12248
rect 14004 12232 14056 12238
rect 14004 12174 14056 12180
rect 13912 12164 13964 12170
rect 13912 12106 13964 12112
rect 14016 11642 14044 12174
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 13924 11626 14044 11642
rect 13912 11620 14044 11626
rect 13964 11614 14044 11620
rect 13912 11562 13964 11568
rect 14016 11354 14044 11614
rect 14108 11354 14136 12038
rect 14200 11898 14228 12242
rect 14292 12220 14320 15864
rect 14384 12374 14412 18022
rect 14568 17678 14596 18226
rect 14817 17980 15113 18000
rect 14873 17978 14897 17980
rect 14953 17978 14977 17980
rect 15033 17978 15057 17980
rect 14895 17926 14897 17978
rect 14959 17926 14971 17978
rect 15033 17926 15035 17978
rect 14873 17924 14897 17926
rect 14953 17924 14977 17926
rect 15033 17924 15057 17926
rect 14817 17904 15113 17924
rect 15384 17740 15436 17746
rect 15384 17682 15436 17688
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 14464 17060 14516 17066
rect 14464 17002 14516 17008
rect 14476 16726 14504 17002
rect 14464 16720 14516 16726
rect 14464 16662 14516 16668
rect 14568 14890 14596 17614
rect 14740 17536 14792 17542
rect 14740 17478 14792 17484
rect 14556 14884 14608 14890
rect 14556 14826 14608 14832
rect 14648 14612 14700 14618
rect 14648 14554 14700 14560
rect 14556 13932 14608 13938
rect 14556 13874 14608 13880
rect 14568 13326 14596 13874
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14372 12368 14424 12374
rect 14372 12310 14424 12316
rect 14568 12306 14596 12786
rect 14556 12300 14608 12306
rect 14556 12242 14608 12248
rect 14292 12192 14412 12220
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 14096 11348 14148 11354
rect 14096 11290 14148 11296
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 13728 11008 13780 11014
rect 13728 10950 13780 10956
rect 13740 10674 13768 10950
rect 13728 10668 13780 10674
rect 13728 10610 13780 10616
rect 13648 10526 13768 10554
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 13648 10266 13676 10406
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13544 9716 13596 9722
rect 13544 9658 13596 9664
rect 13556 7886 13584 9658
rect 13634 8392 13690 8401
rect 13634 8327 13636 8336
rect 13688 8327 13690 8336
rect 13636 8298 13688 8304
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13648 7698 13676 8298
rect 13556 7670 13676 7698
rect 13450 4856 13506 4865
rect 13450 4791 13506 4800
rect 13360 4752 13412 4758
rect 13266 4720 13322 4729
rect 13556 4729 13584 7670
rect 13636 5092 13688 5098
rect 13636 5034 13688 5040
rect 13360 4694 13412 4700
rect 13542 4720 13598 4729
rect 13266 4655 13322 4664
rect 13096 4576 13216 4604
rect 12992 4480 13044 4486
rect 12898 4448 12954 4457
rect 12992 4422 13044 4428
rect 12898 4383 12954 4392
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 12820 3194 12848 4082
rect 12808 3188 12860 3194
rect 12808 3130 12860 3136
rect 12440 2586 12492 2592
rect 12636 2604 12756 2632
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 12452 2310 12480 2450
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 12348 1352 12400 1358
rect 12348 1294 12400 1300
rect 12636 480 12664 2604
rect 12912 2582 12940 4383
rect 13004 2650 13032 4422
rect 12992 2644 13044 2650
rect 12992 2586 13044 2592
rect 12900 2576 12952 2582
rect 12900 2518 12952 2524
rect 13096 480 13124 4576
rect 13176 4004 13228 4010
rect 13176 3946 13228 3952
rect 13188 3738 13216 3946
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 13280 2854 13308 4655
rect 13372 3602 13400 4694
rect 13542 4655 13598 4664
rect 13648 4486 13676 5034
rect 13636 4480 13688 4486
rect 13636 4422 13688 4428
rect 13740 4078 13768 10526
rect 13832 9994 13860 11086
rect 13912 10668 13964 10674
rect 13912 10610 13964 10616
rect 13820 9988 13872 9994
rect 13820 9930 13872 9936
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13832 9042 13860 9590
rect 13924 9178 13952 10610
rect 14004 10192 14056 10198
rect 14002 10160 14004 10169
rect 14056 10160 14058 10169
rect 14002 10095 14058 10104
rect 14200 10062 14228 11834
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14200 9518 14228 9998
rect 14292 9994 14320 11086
rect 14280 9988 14332 9994
rect 14280 9930 14332 9936
rect 14292 9654 14320 9930
rect 14280 9648 14332 9654
rect 14280 9590 14332 9596
rect 14384 9586 14412 12192
rect 14556 11008 14608 11014
rect 14556 10950 14608 10956
rect 14568 9994 14596 10950
rect 14556 9988 14608 9994
rect 14556 9930 14608 9936
rect 14660 9761 14688 14554
rect 14752 12442 14780 17478
rect 14817 16892 15113 16912
rect 14873 16890 14897 16892
rect 14953 16890 14977 16892
rect 15033 16890 15057 16892
rect 14895 16838 14897 16890
rect 14959 16838 14971 16890
rect 15033 16838 15035 16890
rect 14873 16836 14897 16838
rect 14953 16836 14977 16838
rect 15033 16836 15057 16838
rect 14817 16816 15113 16836
rect 15200 16040 15252 16046
rect 15252 16000 15332 16028
rect 15200 15982 15252 15988
rect 14817 15804 15113 15824
rect 14873 15802 14897 15804
rect 14953 15802 14977 15804
rect 15033 15802 15057 15804
rect 14895 15750 14897 15802
rect 14959 15750 14971 15802
rect 15033 15750 15035 15802
rect 14873 15748 14897 15750
rect 14953 15748 14977 15750
rect 15033 15748 15057 15750
rect 14817 15728 15113 15748
rect 15200 15700 15252 15706
rect 15200 15642 15252 15648
rect 14817 14716 15113 14736
rect 14873 14714 14897 14716
rect 14953 14714 14977 14716
rect 15033 14714 15057 14716
rect 14895 14662 14897 14714
rect 14959 14662 14971 14714
rect 15033 14662 15035 14714
rect 14873 14660 14897 14662
rect 14953 14660 14977 14662
rect 15033 14660 15057 14662
rect 14817 14640 15113 14660
rect 14817 13628 15113 13648
rect 14873 13626 14897 13628
rect 14953 13626 14977 13628
rect 15033 13626 15057 13628
rect 14895 13574 14897 13626
rect 14959 13574 14971 13626
rect 15033 13574 15035 13626
rect 14873 13572 14897 13574
rect 14953 13572 14977 13574
rect 15033 13572 15057 13574
rect 14817 13552 15113 13572
rect 15108 13184 15160 13190
rect 15108 13126 15160 13132
rect 15120 12628 15148 13126
rect 15212 12782 15240 15642
rect 15304 14958 15332 16000
rect 15292 14952 15344 14958
rect 15292 14894 15344 14900
rect 15304 14482 15332 14894
rect 15396 14618 15424 17682
rect 15568 15972 15620 15978
rect 15568 15914 15620 15920
rect 15580 15366 15608 15914
rect 15672 15706 15700 19926
rect 15752 19168 15804 19174
rect 15752 19110 15804 19116
rect 15660 15700 15712 15706
rect 15660 15642 15712 15648
rect 15568 15360 15620 15366
rect 15568 15302 15620 15308
rect 15660 15360 15712 15366
rect 15660 15302 15712 15308
rect 15384 14612 15436 14618
rect 15384 14554 15436 14560
rect 15292 14476 15344 14482
rect 15292 14418 15344 14424
rect 15292 13864 15344 13870
rect 15292 13806 15344 13812
rect 15304 13530 15332 13806
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 15120 12600 15240 12628
rect 14817 12540 15113 12560
rect 14873 12538 14897 12540
rect 14953 12538 14977 12540
rect 15033 12538 15057 12540
rect 14895 12486 14897 12538
rect 14959 12486 14971 12538
rect 15033 12486 15035 12538
rect 14873 12484 14897 12486
rect 14953 12484 14977 12486
rect 15033 12484 15057 12486
rect 14817 12464 15113 12484
rect 14740 12436 14792 12442
rect 14740 12378 14792 12384
rect 14817 11452 15113 11472
rect 14873 11450 14897 11452
rect 14953 11450 14977 11452
rect 15033 11450 15057 11452
rect 14895 11398 14897 11450
rect 14959 11398 14971 11450
rect 15033 11398 15035 11450
rect 14873 11396 14897 11398
rect 14953 11396 14977 11398
rect 15033 11396 15057 11398
rect 14817 11376 15113 11396
rect 15212 11257 15240 12600
rect 15198 11248 15254 11257
rect 15198 11183 15254 11192
rect 15212 10674 15240 11183
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 15200 10668 15252 10674
rect 15200 10610 15252 10616
rect 14740 10600 14792 10606
rect 14740 10542 14792 10548
rect 14646 9752 14702 9761
rect 14646 9687 14702 9696
rect 14372 9580 14424 9586
rect 14372 9522 14424 9528
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 14188 9512 14240 9518
rect 14188 9454 14240 9460
rect 14004 9444 14056 9450
rect 14004 9386 14056 9392
rect 13912 9172 13964 9178
rect 13912 9114 13964 9120
rect 14016 9058 14044 9386
rect 14464 9172 14516 9178
rect 14464 9114 14516 9120
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13924 9030 14044 9058
rect 14370 9072 14426 9081
rect 13820 7880 13872 7886
rect 13820 7822 13872 7828
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 13728 4072 13780 4078
rect 13728 4014 13780 4020
rect 13452 3732 13504 3738
rect 13452 3674 13504 3680
rect 13360 3596 13412 3602
rect 13360 3538 13412 3544
rect 13372 3194 13400 3538
rect 13464 3194 13492 3674
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 13556 2514 13584 4014
rect 13728 3936 13780 3942
rect 13728 3878 13780 3884
rect 13740 3738 13768 3878
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13544 2508 13596 2514
rect 13544 2450 13596 2456
rect 13452 2304 13504 2310
rect 13452 2246 13504 2252
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 13464 2038 13492 2246
rect 13452 2032 13504 2038
rect 13452 1974 13504 1980
rect 13556 480 13584 2246
rect 13832 1630 13860 7822
rect 13924 7177 13952 9030
rect 14370 9007 14426 9016
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 14016 7410 14044 7686
rect 14004 7404 14056 7410
rect 14004 7346 14056 7352
rect 13910 7168 13966 7177
rect 13910 7103 13966 7112
rect 13924 6644 13952 7103
rect 13924 6616 14044 6644
rect 13912 5092 13964 5098
rect 13912 5034 13964 5040
rect 13924 4282 13952 5034
rect 13912 4276 13964 4282
rect 13912 4218 13964 4224
rect 14016 3670 14044 6616
rect 14108 5914 14136 8366
rect 14200 7954 14228 8434
rect 14280 8016 14332 8022
rect 14280 7958 14332 7964
rect 14188 7948 14240 7954
rect 14188 7890 14240 7896
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 14200 7342 14228 7482
rect 14188 7336 14240 7342
rect 14188 7278 14240 7284
rect 14188 6860 14240 6866
rect 14188 6802 14240 6808
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 14096 3936 14148 3942
rect 14096 3878 14148 3884
rect 14004 3664 14056 3670
rect 14004 3606 14056 3612
rect 14004 3528 14056 3534
rect 14108 3505 14136 3878
rect 14004 3470 14056 3476
rect 14094 3496 14150 3505
rect 14016 2854 14044 3470
rect 14094 3431 14150 3440
rect 14200 3058 14228 6802
rect 14292 4826 14320 7958
rect 14384 7936 14412 9007
rect 14476 8430 14504 9114
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 14384 7908 14504 7936
rect 14372 7812 14424 7818
rect 14372 7754 14424 7760
rect 14384 7206 14412 7754
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 14476 7002 14504 7908
rect 14464 6996 14516 7002
rect 14464 6938 14516 6944
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 14384 6322 14412 6734
rect 14464 6724 14516 6730
rect 14464 6666 14516 6672
rect 14372 6316 14424 6322
rect 14372 6258 14424 6264
rect 14280 4820 14332 4826
rect 14280 4762 14332 4768
rect 14292 4214 14320 4762
rect 14280 4208 14332 4214
rect 14280 4150 14332 4156
rect 14278 4040 14334 4049
rect 14278 3975 14334 3984
rect 14292 3505 14320 3975
rect 14278 3496 14334 3505
rect 14278 3431 14334 3440
rect 14188 3052 14240 3058
rect 14188 2994 14240 3000
rect 14004 2848 14056 2854
rect 14004 2790 14056 2796
rect 14096 2372 14148 2378
rect 14096 2314 14148 2320
rect 13820 1624 13872 1630
rect 13820 1566 13872 1572
rect 14108 480 14136 2314
rect 14384 1494 14412 6258
rect 14476 2122 14504 6666
rect 14568 6458 14596 9522
rect 14660 8537 14688 9687
rect 14752 9058 14780 10542
rect 14817 10364 15113 10384
rect 14873 10362 14897 10364
rect 14953 10362 14977 10364
rect 15033 10362 15057 10364
rect 14895 10310 14897 10362
rect 14959 10310 14971 10362
rect 15033 10310 15035 10362
rect 14873 10308 14897 10310
rect 14953 10308 14977 10310
rect 15033 10308 15057 10310
rect 14817 10288 15113 10308
rect 15304 10198 15332 11086
rect 15292 10192 15344 10198
rect 15292 10134 15344 10140
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 15120 10033 15148 10066
rect 15106 10024 15162 10033
rect 15106 9959 15162 9968
rect 15292 9580 15344 9586
rect 15396 9568 15424 13126
rect 15476 11212 15528 11218
rect 15476 11154 15528 11160
rect 15488 10606 15516 11154
rect 15476 10600 15528 10606
rect 15476 10542 15528 10548
rect 15476 10192 15528 10198
rect 15476 10134 15528 10140
rect 15344 9540 15424 9568
rect 15292 9522 15344 9528
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 14817 9276 15113 9296
rect 14873 9274 14897 9276
rect 14953 9274 14977 9276
rect 15033 9274 15057 9276
rect 14895 9222 14897 9274
rect 14959 9222 14971 9274
rect 15033 9222 15035 9274
rect 14873 9220 14897 9222
rect 14953 9220 14977 9222
rect 15033 9220 15057 9222
rect 14817 9200 15113 9220
rect 14752 9030 14872 9058
rect 14646 8528 14702 8537
rect 14646 8463 14702 8472
rect 14844 8276 14872 9030
rect 14660 8248 14872 8276
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14554 4176 14610 4185
rect 14554 4111 14610 4120
rect 14568 3194 14596 4111
rect 14556 3188 14608 3194
rect 14556 3130 14608 3136
rect 14660 2446 14688 8248
rect 14817 8188 15113 8208
rect 14873 8186 14897 8188
rect 14953 8186 14977 8188
rect 15033 8186 15057 8188
rect 14895 8134 14897 8186
rect 14959 8134 14971 8186
rect 15033 8134 15035 8186
rect 14873 8132 14897 8134
rect 14953 8132 14977 8134
rect 15033 8132 15057 8134
rect 14817 8112 15113 8132
rect 15212 8090 15240 9318
rect 15488 9042 15516 10134
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 15384 9036 15436 9042
rect 15384 8978 15436 8984
rect 15476 9036 15528 9042
rect 15476 8978 15528 8984
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 15304 8362 15332 8774
rect 15292 8356 15344 8362
rect 15292 8298 15344 8304
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 15200 8084 15252 8090
rect 15200 8026 15252 8032
rect 14752 3602 14780 8026
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 14817 7100 15113 7120
rect 14873 7098 14897 7100
rect 14953 7098 14977 7100
rect 15033 7098 15057 7100
rect 14895 7046 14897 7098
rect 14959 7046 14971 7098
rect 15033 7046 15035 7098
rect 14873 7044 14897 7046
rect 14953 7044 14977 7046
rect 15033 7044 15057 7046
rect 14817 7024 15113 7044
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 14817 6012 15113 6032
rect 14873 6010 14897 6012
rect 14953 6010 14977 6012
rect 15033 6010 15057 6012
rect 14895 5958 14897 6010
rect 14959 5958 14971 6010
rect 15033 5958 15035 6010
rect 14873 5956 14897 5958
rect 14953 5956 14977 5958
rect 15033 5956 15057 5958
rect 14817 5936 15113 5956
rect 15212 5914 15240 6054
rect 15200 5908 15252 5914
rect 15200 5850 15252 5856
rect 15304 5846 15332 7142
rect 15292 5840 15344 5846
rect 15292 5782 15344 5788
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 14817 4924 15113 4944
rect 14873 4922 14897 4924
rect 14953 4922 14977 4924
rect 15033 4922 15057 4924
rect 14895 4870 14897 4922
rect 14959 4870 14971 4922
rect 15033 4870 15035 4922
rect 14873 4868 14897 4870
rect 14953 4868 14977 4870
rect 15033 4868 15057 4870
rect 14817 4848 15113 4868
rect 15212 4146 15240 5170
rect 15292 5160 15344 5166
rect 15292 5102 15344 5108
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15200 4004 15252 4010
rect 15200 3946 15252 3952
rect 14817 3836 15113 3856
rect 14873 3834 14897 3836
rect 14953 3834 14977 3836
rect 15033 3834 15057 3836
rect 14895 3782 14897 3834
rect 14959 3782 14971 3834
rect 15033 3782 15035 3834
rect 14873 3780 14897 3782
rect 14953 3780 14977 3782
rect 15033 3780 15057 3782
rect 14817 3760 15113 3780
rect 14740 3596 14792 3602
rect 14740 3538 14792 3544
rect 15016 3460 15068 3466
rect 15016 3402 15068 3408
rect 15028 3058 15056 3402
rect 15016 3052 15068 3058
rect 15016 2994 15068 3000
rect 15028 2836 15056 2994
rect 14752 2808 15056 2836
rect 14752 2514 14780 2808
rect 14817 2748 15113 2768
rect 14873 2746 14897 2748
rect 14953 2746 14977 2748
rect 15033 2746 15057 2748
rect 14895 2694 14897 2746
rect 14959 2694 14971 2746
rect 15033 2694 15035 2746
rect 14873 2692 14897 2694
rect 14953 2692 14977 2694
rect 15033 2692 15057 2694
rect 14817 2672 15113 2692
rect 14740 2508 14792 2514
rect 14740 2450 14792 2456
rect 14648 2440 14700 2446
rect 14648 2382 14700 2388
rect 14476 2094 15056 2122
rect 14464 2032 14516 2038
rect 14464 1974 14516 1980
rect 14372 1488 14424 1494
rect 14372 1430 14424 1436
rect 14476 1306 14504 1974
rect 14476 1278 14596 1306
rect 14568 480 14596 1278
rect 15028 480 15056 2094
rect 15212 1698 15240 3946
rect 15304 3058 15332 5102
rect 15292 3052 15344 3058
rect 15292 2994 15344 3000
rect 15292 2916 15344 2922
rect 15292 2858 15344 2864
rect 15304 2417 15332 2858
rect 15396 2582 15424 8978
rect 15476 7744 15528 7750
rect 15476 7686 15528 7692
rect 15488 6390 15516 7686
rect 15580 6984 15608 10066
rect 15672 8294 15700 15302
rect 15764 11286 15792 19110
rect 15856 17814 15884 20198
rect 16396 19712 16448 19718
rect 16396 19654 16448 19660
rect 16672 19712 16724 19718
rect 16672 19654 16724 19660
rect 16764 19712 16816 19718
rect 16764 19654 16816 19660
rect 16212 18284 16264 18290
rect 16212 18226 16264 18232
rect 15936 18080 15988 18086
rect 15936 18022 15988 18028
rect 16120 18080 16172 18086
rect 16120 18022 16172 18028
rect 15844 17808 15896 17814
rect 15844 17750 15896 17756
rect 15948 16726 15976 18022
rect 16028 16992 16080 16998
rect 16028 16934 16080 16940
rect 16040 16794 16068 16934
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 15936 16720 15988 16726
rect 15934 16688 15936 16697
rect 15988 16688 15990 16697
rect 15934 16623 15990 16632
rect 16132 14906 16160 18022
rect 16224 16454 16252 18226
rect 16408 17660 16436 19654
rect 16580 18148 16632 18154
rect 16580 18090 16632 18096
rect 16488 17672 16540 17678
rect 16408 17632 16488 17660
rect 16488 17614 16540 17620
rect 16500 17270 16528 17614
rect 16592 17338 16620 18090
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 16488 17264 16540 17270
rect 16488 17206 16540 17212
rect 16580 16992 16632 16998
rect 16580 16934 16632 16940
rect 16592 16726 16620 16934
rect 16580 16720 16632 16726
rect 16580 16662 16632 16668
rect 16212 16448 16264 16454
rect 16212 16390 16264 16396
rect 16580 16448 16632 16454
rect 16580 16390 16632 16396
rect 16224 16250 16252 16390
rect 16212 16244 16264 16250
rect 16212 16186 16264 16192
rect 16592 15586 16620 16390
rect 16408 15558 16620 15586
rect 16408 15502 16436 15558
rect 16396 15496 16448 15502
rect 16580 15496 16632 15502
rect 16396 15438 16448 15444
rect 16500 15456 16580 15484
rect 16132 14878 16252 14906
rect 16120 14816 16172 14822
rect 16120 14758 16172 14764
rect 16028 14272 16080 14278
rect 16028 14214 16080 14220
rect 15936 13728 15988 13734
rect 15936 13670 15988 13676
rect 15948 13530 15976 13670
rect 15936 13524 15988 13530
rect 15936 13466 15988 13472
rect 15936 13388 15988 13394
rect 15936 13330 15988 13336
rect 15948 12986 15976 13330
rect 16040 13326 16068 14214
rect 16132 14006 16160 14758
rect 16224 14618 16252 14878
rect 16500 14822 16528 15456
rect 16580 15438 16632 15444
rect 16488 14816 16540 14822
rect 16488 14758 16540 14764
rect 16212 14612 16264 14618
rect 16212 14554 16264 14560
rect 16120 14000 16172 14006
rect 16120 13942 16172 13948
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 15936 12980 15988 12986
rect 15936 12922 15988 12928
rect 15844 12776 15896 12782
rect 15844 12718 15896 12724
rect 15752 11280 15804 11286
rect 15752 11222 15804 11228
rect 15856 10266 15884 12718
rect 16132 12238 16160 13942
rect 16224 13938 16252 14554
rect 16684 14550 16712 19654
rect 16776 18834 16804 19654
rect 17132 19236 17184 19242
rect 17132 19178 17184 19184
rect 17144 18902 17172 19178
rect 17132 18896 17184 18902
rect 17132 18838 17184 18844
rect 16764 18828 16816 18834
rect 16764 18770 16816 18776
rect 16856 18828 16908 18834
rect 16856 18770 16908 18776
rect 17040 18828 17092 18834
rect 17040 18770 17092 18776
rect 16764 18080 16816 18086
rect 16764 18022 16816 18028
rect 16672 14544 16724 14550
rect 16672 14486 16724 14492
rect 16684 13938 16712 14486
rect 16212 13932 16264 13938
rect 16212 13874 16264 13880
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 16212 13796 16264 13802
rect 16212 13738 16264 13744
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 15844 10260 15896 10266
rect 15844 10202 15896 10208
rect 16132 10146 16160 12174
rect 15856 10118 16160 10146
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 15752 8016 15804 8022
rect 15752 7958 15804 7964
rect 15764 7410 15792 7958
rect 15752 7404 15804 7410
rect 15752 7346 15804 7352
rect 15764 7002 15792 7346
rect 15752 6996 15804 7002
rect 15580 6956 15700 6984
rect 15568 6860 15620 6866
rect 15568 6802 15620 6808
rect 15476 6384 15528 6390
rect 15476 6326 15528 6332
rect 15580 5710 15608 6802
rect 15672 6118 15700 6956
rect 15752 6938 15804 6944
rect 15764 6798 15792 6938
rect 15752 6792 15804 6798
rect 15752 6734 15804 6740
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15660 6112 15712 6118
rect 15660 6054 15712 6060
rect 15764 5914 15792 6598
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 15568 5704 15620 5710
rect 15568 5646 15620 5652
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 15384 2576 15436 2582
rect 15384 2518 15436 2524
rect 15488 2514 15516 5510
rect 15580 4010 15608 5646
rect 15750 4720 15806 4729
rect 15750 4655 15806 4664
rect 15764 4486 15792 4655
rect 15752 4480 15804 4486
rect 15752 4422 15804 4428
rect 15568 4004 15620 4010
rect 15568 3946 15620 3952
rect 15764 3602 15792 4422
rect 15752 3596 15804 3602
rect 15752 3538 15804 3544
rect 15856 2922 15884 10118
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 16040 9654 16068 9998
rect 16028 9648 16080 9654
rect 16028 9590 16080 9596
rect 16028 8968 16080 8974
rect 16028 8910 16080 8916
rect 15936 8560 15988 8566
rect 15936 8502 15988 8508
rect 15948 5710 15976 8502
rect 16040 8022 16068 8910
rect 16120 8288 16172 8294
rect 16120 8230 16172 8236
rect 16028 8016 16080 8022
rect 16028 7958 16080 7964
rect 16026 7576 16082 7585
rect 16026 7511 16082 7520
rect 15936 5704 15988 5710
rect 15936 5646 15988 5652
rect 15936 5024 15988 5030
rect 15936 4966 15988 4972
rect 15844 2916 15896 2922
rect 15844 2858 15896 2864
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 15290 2408 15346 2417
rect 15290 2343 15346 2352
rect 15476 2100 15528 2106
rect 15476 2042 15528 2048
rect 15200 1692 15252 1698
rect 15200 1634 15252 1640
rect 15488 480 15516 2042
rect 15948 480 15976 4966
rect 16040 4690 16068 7511
rect 16028 4684 16080 4690
rect 16028 4626 16080 4632
rect 16028 3936 16080 3942
rect 16028 3878 16080 3884
rect 16040 3777 16068 3878
rect 16026 3768 16082 3777
rect 16026 3703 16082 3712
rect 16132 1834 16160 8230
rect 16224 7585 16252 13738
rect 16684 12850 16712 13874
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16776 12714 16804 18022
rect 16868 17814 16896 18770
rect 17052 18086 17080 18770
rect 17040 18080 17092 18086
rect 17040 18022 17092 18028
rect 16856 17808 16908 17814
rect 16856 17750 16908 17756
rect 16764 12708 16816 12714
rect 16764 12650 16816 12656
rect 16868 12594 16896 17750
rect 17040 17740 17092 17746
rect 17040 17682 17092 17688
rect 17052 17202 17080 17682
rect 17132 17264 17184 17270
rect 17132 17206 17184 17212
rect 17040 17196 17092 17202
rect 17040 17138 17092 17144
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 16960 16658 16988 16934
rect 16948 16652 17000 16658
rect 16948 16594 17000 16600
rect 17144 16590 17172 17206
rect 17132 16584 17184 16590
rect 17132 16526 17184 16532
rect 17144 14482 17172 16526
rect 17236 16017 17264 20334
rect 17958 20295 18014 20304
rect 18052 20324 18104 20330
rect 17972 20074 18000 20295
rect 18052 20266 18104 20272
rect 17880 20058 18000 20074
rect 17868 20052 18000 20058
rect 17920 20046 18000 20052
rect 17868 19994 17920 20000
rect 17958 19952 18014 19961
rect 17958 19887 18014 19896
rect 17774 19000 17830 19009
rect 17774 18935 17830 18944
rect 17316 18896 17368 18902
rect 17316 18838 17368 18844
rect 17328 16726 17356 18838
rect 17788 18698 17816 18935
rect 17972 18714 18000 19887
rect 18064 19281 18092 20266
rect 18156 19854 18184 20470
rect 18248 19990 18276 20470
rect 18880 20460 18932 20466
rect 18880 20402 18932 20408
rect 18788 20392 18840 20398
rect 18788 20334 18840 20340
rect 18604 20256 18656 20262
rect 18604 20198 18656 20204
rect 18236 19984 18288 19990
rect 18236 19926 18288 19932
rect 18144 19848 18196 19854
rect 18144 19790 18196 19796
rect 18156 19378 18184 19790
rect 18282 19612 18578 19632
rect 18338 19610 18362 19612
rect 18418 19610 18442 19612
rect 18498 19610 18522 19612
rect 18360 19558 18362 19610
rect 18424 19558 18436 19610
rect 18498 19558 18500 19610
rect 18338 19556 18362 19558
rect 18418 19556 18442 19558
rect 18498 19556 18522 19558
rect 18282 19536 18578 19556
rect 18144 19372 18196 19378
rect 18144 19314 18196 19320
rect 18050 19272 18106 19281
rect 18616 19242 18644 20198
rect 18694 19408 18750 19417
rect 18694 19343 18750 19352
rect 18050 19207 18106 19216
rect 18604 19236 18656 19242
rect 18604 19178 18656 19184
rect 18052 19168 18104 19174
rect 18052 19110 18104 19116
rect 18064 18970 18092 19110
rect 18052 18964 18104 18970
rect 18052 18906 18104 18912
rect 17776 18692 17828 18698
rect 17776 18634 17828 18640
rect 17880 18686 18000 18714
rect 18144 18692 18196 18698
rect 17880 18630 17908 18686
rect 18144 18634 18196 18640
rect 17868 18624 17920 18630
rect 17868 18566 17920 18572
rect 18052 18624 18104 18630
rect 18052 18566 18104 18572
rect 18064 18465 18092 18566
rect 18050 18456 18106 18465
rect 18050 18391 18106 18400
rect 18052 18352 18104 18358
rect 18052 18294 18104 18300
rect 17592 18080 17644 18086
rect 18064 18057 18092 18294
rect 17592 18022 17644 18028
rect 18050 18048 18106 18057
rect 17500 17604 17552 17610
rect 17500 17546 17552 17552
rect 17408 17536 17460 17542
rect 17408 17478 17460 17484
rect 17420 16998 17448 17478
rect 17408 16992 17460 16998
rect 17408 16934 17460 16940
rect 17316 16720 17368 16726
rect 17316 16662 17368 16668
rect 17408 16720 17460 16726
rect 17408 16662 17460 16668
rect 17222 16008 17278 16017
rect 17222 15943 17278 15952
rect 17132 14476 17184 14482
rect 17132 14418 17184 14424
rect 17144 12850 17172 14418
rect 17236 13433 17264 15943
rect 17222 13424 17278 13433
rect 17222 13359 17278 13368
rect 17328 12986 17356 16662
rect 17420 15434 17448 16662
rect 17512 15706 17540 17546
rect 17500 15700 17552 15706
rect 17500 15642 17552 15648
rect 17408 15428 17460 15434
rect 17408 15370 17460 15376
rect 17316 12980 17368 12986
rect 17316 12922 17368 12928
rect 17132 12844 17184 12850
rect 17132 12786 17184 12792
rect 16776 12566 16896 12594
rect 16580 12436 16632 12442
rect 16580 12378 16632 12384
rect 16304 12096 16356 12102
rect 16304 12038 16356 12044
rect 16210 7576 16266 7585
rect 16210 7511 16266 7520
rect 16316 7426 16344 12038
rect 16592 11898 16620 12378
rect 16580 11892 16632 11898
rect 16580 11834 16632 11840
rect 16488 11688 16540 11694
rect 16488 11630 16540 11636
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16224 7398 16344 7426
rect 16224 1970 16252 7398
rect 16408 5522 16436 11494
rect 16316 5494 16436 5522
rect 16316 4146 16344 5494
rect 16396 5364 16448 5370
rect 16396 5306 16448 5312
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 16316 3738 16344 3878
rect 16304 3732 16356 3738
rect 16304 3674 16356 3680
rect 16212 1964 16264 1970
rect 16212 1906 16264 1912
rect 16120 1828 16172 1834
rect 16120 1770 16172 1776
rect 16408 1034 16436 5306
rect 16500 3534 16528 11630
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16684 8945 16712 11494
rect 16776 10266 16804 12566
rect 17144 12306 17172 12786
rect 17316 12640 17368 12646
rect 17316 12582 17368 12588
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 17224 12300 17276 12306
rect 17224 12242 17276 12248
rect 16946 11656 17002 11665
rect 16946 11591 16948 11600
rect 17000 11591 17002 11600
rect 16948 11562 17000 11568
rect 17236 11354 17264 12242
rect 17328 12209 17356 12582
rect 17314 12200 17370 12209
rect 17314 12135 17370 12144
rect 17224 11348 17276 11354
rect 17224 11290 17276 11296
rect 17132 11212 17184 11218
rect 17132 11154 17184 11160
rect 16856 10532 16908 10538
rect 16856 10474 16908 10480
rect 16764 10260 16816 10266
rect 16764 10202 16816 10208
rect 16776 10130 16804 10202
rect 16764 10124 16816 10130
rect 16764 10066 16816 10072
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 16776 9518 16804 9862
rect 16764 9512 16816 9518
rect 16764 9454 16816 9460
rect 16764 9172 16816 9178
rect 16764 9114 16816 9120
rect 16670 8936 16726 8945
rect 16670 8871 16726 8880
rect 16580 8356 16632 8362
rect 16580 8298 16632 8304
rect 16592 7954 16620 8298
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 16580 5092 16632 5098
rect 16580 5034 16632 5040
rect 16592 3670 16620 5034
rect 16672 5024 16724 5030
rect 16672 4966 16724 4972
rect 16684 4010 16712 4966
rect 16776 4434 16804 9114
rect 16868 5370 16896 10474
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 16960 5914 16988 9318
rect 17040 9036 17092 9042
rect 17040 8978 17092 8984
rect 17052 8498 17080 8978
rect 17040 8492 17092 8498
rect 17040 8434 17092 8440
rect 17040 7472 17092 7478
rect 17040 7414 17092 7420
rect 17052 7313 17080 7414
rect 17038 7304 17094 7313
rect 17038 7239 17094 7248
rect 17040 6996 17092 7002
rect 17040 6938 17092 6944
rect 16948 5908 17000 5914
rect 16948 5850 17000 5856
rect 17052 5778 17080 6938
rect 17144 6322 17172 11154
rect 17236 10674 17264 11290
rect 17224 10668 17276 10674
rect 17224 10610 17276 10616
rect 17420 10554 17448 15370
rect 17500 14884 17552 14890
rect 17500 14826 17552 14832
rect 17512 14074 17540 14826
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 17500 13320 17552 13326
rect 17500 13262 17552 13268
rect 17512 12646 17540 13262
rect 17604 12782 17632 18022
rect 18050 17983 18106 17992
rect 17696 17598 17908 17626
rect 17696 16454 17724 17598
rect 17880 17542 17908 17598
rect 17868 17536 17920 17542
rect 17868 17478 17920 17484
rect 17868 17128 17920 17134
rect 17868 17070 17920 17076
rect 17880 16726 17908 17070
rect 17868 16720 17920 16726
rect 17868 16662 17920 16668
rect 17684 16448 17736 16454
rect 17684 16390 17736 16396
rect 17776 16176 17828 16182
rect 17776 16118 17828 16124
rect 17788 13326 17816 16118
rect 18156 15688 18184 18634
rect 18282 18524 18578 18544
rect 18338 18522 18362 18524
rect 18418 18522 18442 18524
rect 18498 18522 18522 18524
rect 18360 18470 18362 18522
rect 18424 18470 18436 18522
rect 18498 18470 18500 18522
rect 18338 18468 18362 18470
rect 18418 18468 18442 18470
rect 18498 18468 18522 18470
rect 18282 18448 18578 18468
rect 18604 18420 18656 18426
rect 18604 18362 18656 18368
rect 18234 18320 18290 18329
rect 18234 18255 18290 18264
rect 18248 18154 18276 18255
rect 18236 18148 18288 18154
rect 18236 18090 18288 18096
rect 18512 18080 18564 18086
rect 18616 18057 18644 18362
rect 18512 18022 18564 18028
rect 18602 18048 18658 18057
rect 18524 17921 18552 18022
rect 18602 17983 18658 17992
rect 18510 17912 18566 17921
rect 18708 17882 18736 19343
rect 18800 18222 18828 20334
rect 18892 19854 18920 20402
rect 18880 19848 18932 19854
rect 18880 19790 18932 19796
rect 18984 19394 19012 22607
rect 20074 22520 20130 23000
rect 19154 22264 19210 22273
rect 19154 22199 19210 22208
rect 19168 20058 19196 22199
rect 19246 21312 19302 21321
rect 19246 21247 19302 21256
rect 19156 20052 19208 20058
rect 19156 19994 19208 20000
rect 18892 19366 19012 19394
rect 18788 18216 18840 18222
rect 18788 18158 18840 18164
rect 18510 17847 18566 17856
rect 18696 17876 18748 17882
rect 18696 17818 18748 17824
rect 18282 17436 18578 17456
rect 18338 17434 18362 17436
rect 18418 17434 18442 17436
rect 18498 17434 18522 17436
rect 18360 17382 18362 17434
rect 18424 17382 18436 17434
rect 18498 17382 18500 17434
rect 18338 17380 18362 17382
rect 18418 17380 18442 17382
rect 18498 17380 18522 17382
rect 18282 17360 18578 17380
rect 18604 16992 18656 16998
rect 18604 16934 18656 16940
rect 18616 16794 18644 16934
rect 18604 16788 18656 16794
rect 18604 16730 18656 16736
rect 18788 16516 18840 16522
rect 18788 16458 18840 16464
rect 18282 16348 18578 16368
rect 18338 16346 18362 16348
rect 18418 16346 18442 16348
rect 18498 16346 18522 16348
rect 18360 16294 18362 16346
rect 18424 16294 18436 16346
rect 18498 16294 18500 16346
rect 18338 16292 18362 16294
rect 18418 16292 18442 16294
rect 18498 16292 18522 16294
rect 18282 16272 18578 16292
rect 18694 16280 18750 16289
rect 18694 16215 18750 16224
rect 18604 15904 18656 15910
rect 18604 15846 18656 15852
rect 17972 15660 18184 15688
rect 17972 13870 18000 15660
rect 18050 15600 18106 15609
rect 18050 15535 18052 15544
rect 18104 15535 18106 15544
rect 18052 15506 18104 15512
rect 18144 15496 18196 15502
rect 18144 15438 18196 15444
rect 18326 15464 18382 15473
rect 18052 15360 18104 15366
rect 18052 15302 18104 15308
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 18064 13546 18092 15302
rect 18156 14074 18184 15438
rect 18326 15399 18328 15408
rect 18380 15399 18382 15408
rect 18328 15370 18380 15376
rect 18282 15260 18578 15280
rect 18338 15258 18362 15260
rect 18418 15258 18442 15260
rect 18498 15258 18522 15260
rect 18360 15206 18362 15258
rect 18424 15206 18436 15258
rect 18498 15206 18500 15258
rect 18338 15204 18362 15206
rect 18418 15204 18442 15206
rect 18498 15204 18522 15206
rect 18282 15184 18578 15204
rect 18616 14385 18644 15846
rect 18708 15162 18736 16215
rect 18696 15156 18748 15162
rect 18696 15098 18748 15104
rect 18696 14816 18748 14822
rect 18696 14758 18748 14764
rect 18602 14376 18658 14385
rect 18602 14311 18658 14320
rect 18604 14272 18656 14278
rect 18604 14214 18656 14220
rect 18282 14172 18578 14192
rect 18338 14170 18362 14172
rect 18418 14170 18442 14172
rect 18498 14170 18522 14172
rect 18360 14118 18362 14170
rect 18424 14118 18436 14170
rect 18498 14118 18500 14170
rect 18338 14116 18362 14118
rect 18418 14116 18442 14118
rect 18498 14116 18522 14118
rect 18282 14096 18578 14116
rect 18144 14068 18196 14074
rect 18144 14010 18196 14016
rect 18616 13977 18644 14214
rect 18602 13968 18658 13977
rect 18708 13938 18736 14758
rect 18602 13903 18658 13912
rect 18696 13932 18748 13938
rect 18696 13874 18748 13880
rect 18800 13802 18828 16458
rect 18892 16153 18920 19366
rect 18972 19236 19024 19242
rect 18972 19178 19024 19184
rect 18984 18902 19012 19178
rect 19064 19168 19116 19174
rect 19064 19110 19116 19116
rect 18972 18896 19024 18902
rect 18972 18838 19024 18844
rect 19076 18086 19104 19110
rect 19064 18080 19116 18086
rect 19064 18022 19116 18028
rect 18970 16688 19026 16697
rect 19168 16658 19196 19994
rect 19260 18970 19288 21247
rect 20088 20074 20116 22520
rect 20166 21720 20222 21729
rect 20166 21655 20222 21664
rect 20180 20602 20208 21655
rect 20168 20596 20220 20602
rect 20168 20538 20220 20544
rect 19536 20046 20116 20074
rect 19340 19916 19392 19922
rect 19340 19858 19392 19864
rect 19352 19514 19380 19858
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 19248 18964 19300 18970
rect 19248 18906 19300 18912
rect 19432 18828 19484 18834
rect 19432 18770 19484 18776
rect 19340 18760 19392 18766
rect 19340 18702 19392 18708
rect 19352 18290 19380 18702
rect 19340 18284 19392 18290
rect 19340 18226 19392 18232
rect 19248 18080 19300 18086
rect 19248 18022 19300 18028
rect 18970 16623 19026 16632
rect 19156 16652 19208 16658
rect 18878 16144 18934 16153
rect 18878 16079 18934 16088
rect 18880 15904 18932 15910
rect 18880 15846 18932 15852
rect 18892 14521 18920 15846
rect 18878 14512 18934 14521
rect 18878 14447 18934 14456
rect 18788 13796 18840 13802
rect 18788 13738 18840 13744
rect 18064 13518 18184 13546
rect 17868 13456 17920 13462
rect 17868 13398 17920 13404
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 17592 12776 17644 12782
rect 17592 12718 17644 12724
rect 17500 12640 17552 12646
rect 17500 12582 17552 12588
rect 17328 10526 17448 10554
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 17132 6316 17184 6322
rect 17132 6258 17184 6264
rect 17040 5772 17092 5778
rect 17040 5714 17092 5720
rect 16856 5364 16908 5370
rect 16856 5306 16908 5312
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 16868 4826 16896 4966
rect 16856 4820 16908 4826
rect 16856 4762 16908 4768
rect 16960 4758 16988 5170
rect 17052 5166 17080 5714
rect 17132 5704 17184 5710
rect 17132 5646 17184 5652
rect 17040 5160 17092 5166
rect 17040 5102 17092 5108
rect 16948 4752 17000 4758
rect 16948 4694 17000 4700
rect 17052 4622 17080 5102
rect 17040 4616 17092 4622
rect 17040 4558 17092 4564
rect 17144 4554 17172 5646
rect 17132 4548 17184 4554
rect 17132 4490 17184 4496
rect 16776 4406 16988 4434
rect 16672 4004 16724 4010
rect 16672 3946 16724 3952
rect 16580 3664 16632 3670
rect 16580 3606 16632 3612
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 16408 1006 16528 1034
rect 16500 480 16528 1006
rect 16960 480 16988 4406
rect 17144 4282 17172 4490
rect 17132 4276 17184 4282
rect 17132 4218 17184 4224
rect 17236 2582 17264 10406
rect 17328 6769 17356 10526
rect 17604 10418 17632 12718
rect 17684 12708 17736 12714
rect 17684 12650 17736 12656
rect 17420 10390 17632 10418
rect 17314 6760 17370 6769
rect 17314 6695 17370 6704
rect 17316 6656 17368 6662
rect 17316 6598 17368 6604
rect 17328 6322 17356 6598
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 17328 5778 17356 6258
rect 17420 6254 17448 10390
rect 17592 10260 17644 10266
rect 17592 10202 17644 10208
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17408 6248 17460 6254
rect 17408 6190 17460 6196
rect 17512 6066 17540 9318
rect 17604 8294 17632 10202
rect 17592 8288 17644 8294
rect 17592 8230 17644 8236
rect 17420 6038 17540 6066
rect 17316 5772 17368 5778
rect 17316 5714 17368 5720
rect 17316 5364 17368 5370
rect 17316 5306 17368 5312
rect 17328 2961 17356 5306
rect 17314 2952 17370 2961
rect 17314 2887 17370 2896
rect 17224 2576 17276 2582
rect 17224 2518 17276 2524
rect 17224 2440 17276 2446
rect 17224 2382 17276 2388
rect 17236 1562 17264 2382
rect 17224 1556 17276 1562
rect 17224 1498 17276 1504
rect 17420 480 17448 6038
rect 17500 5772 17552 5778
rect 17500 5714 17552 5720
rect 17512 1766 17540 5714
rect 17696 2009 17724 12650
rect 17776 12640 17828 12646
rect 17776 12582 17828 12588
rect 17788 12322 17816 12582
rect 17880 12442 17908 13398
rect 18052 13388 18104 13394
rect 18052 13330 18104 13336
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 17868 12436 17920 12442
rect 17972 12424 18000 13262
rect 18064 12617 18092 13330
rect 18156 12646 18184 13518
rect 18788 13252 18840 13258
rect 18788 13194 18840 13200
rect 18696 13184 18748 13190
rect 18696 13126 18748 13132
rect 18282 13084 18578 13104
rect 18338 13082 18362 13084
rect 18418 13082 18442 13084
rect 18498 13082 18522 13084
rect 18360 13030 18362 13082
rect 18424 13030 18436 13082
rect 18498 13030 18500 13082
rect 18338 13028 18362 13030
rect 18418 13028 18442 13030
rect 18498 13028 18522 13030
rect 18282 13008 18578 13028
rect 18604 12980 18656 12986
rect 18604 12922 18656 12928
rect 18144 12640 18196 12646
rect 18050 12608 18106 12617
rect 18144 12582 18196 12588
rect 18050 12543 18106 12552
rect 17972 12396 18184 12424
rect 17868 12378 17920 12384
rect 17788 12294 18000 12322
rect 17972 11762 18000 12294
rect 18052 12096 18104 12102
rect 18052 12038 18104 12044
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 18064 11626 18092 12038
rect 18052 11620 18104 11626
rect 18052 11562 18104 11568
rect 18156 11506 18184 12396
rect 18282 11996 18578 12016
rect 18338 11994 18362 11996
rect 18418 11994 18442 11996
rect 18498 11994 18522 11996
rect 18360 11942 18362 11994
rect 18424 11942 18436 11994
rect 18498 11942 18500 11994
rect 18338 11940 18362 11942
rect 18418 11940 18442 11942
rect 18498 11940 18522 11942
rect 18282 11920 18578 11940
rect 18064 11478 18184 11506
rect 17776 11008 17828 11014
rect 17776 10950 17828 10956
rect 17788 10606 17816 10950
rect 17776 10600 17828 10606
rect 17776 10542 17828 10548
rect 18064 10470 18092 11478
rect 18142 11384 18198 11393
rect 18142 11319 18144 11328
rect 18196 11319 18198 11328
rect 18144 11290 18196 11296
rect 18144 11076 18196 11082
rect 18144 11018 18196 11024
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 17866 10296 17922 10305
rect 18156 10266 18184 11018
rect 18282 10908 18578 10928
rect 18338 10906 18362 10908
rect 18418 10906 18442 10908
rect 18498 10906 18522 10908
rect 18360 10854 18362 10906
rect 18424 10854 18436 10906
rect 18498 10854 18500 10906
rect 18338 10852 18362 10854
rect 18418 10852 18442 10854
rect 18498 10852 18522 10854
rect 18282 10832 18578 10852
rect 18236 10736 18288 10742
rect 18236 10678 18288 10684
rect 17866 10231 17922 10240
rect 18144 10260 18196 10266
rect 17776 10124 17828 10130
rect 17776 10066 17828 10072
rect 17788 9178 17816 10066
rect 17880 9926 17908 10231
rect 18144 10202 18196 10208
rect 18050 10160 18106 10169
rect 18248 10146 18276 10678
rect 18050 10095 18106 10104
rect 18156 10118 18276 10146
rect 17958 10024 18014 10033
rect 17958 9959 17960 9968
rect 18012 9959 18014 9968
rect 17960 9930 18012 9936
rect 17868 9920 17920 9926
rect 17868 9862 17920 9868
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17774 8528 17830 8537
rect 17774 8463 17830 8472
rect 17788 6984 17816 8463
rect 17880 8362 17908 9862
rect 17960 9512 18012 9518
rect 17960 9454 18012 9460
rect 17868 8356 17920 8362
rect 17868 8298 17920 8304
rect 17972 7154 18000 9454
rect 18064 9353 18092 10095
rect 18156 9704 18184 10118
rect 18282 9820 18578 9840
rect 18338 9818 18362 9820
rect 18418 9818 18442 9820
rect 18498 9818 18522 9820
rect 18360 9766 18362 9818
rect 18424 9766 18436 9818
rect 18498 9766 18500 9818
rect 18338 9764 18362 9766
rect 18418 9764 18442 9766
rect 18498 9764 18522 9766
rect 18282 9744 18578 9764
rect 18156 9676 18552 9704
rect 18524 9625 18552 9676
rect 18510 9616 18566 9625
rect 18510 9551 18566 9560
rect 18234 9480 18290 9489
rect 18234 9415 18290 9424
rect 18050 9344 18106 9353
rect 18050 9279 18106 9288
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 18156 9081 18184 9114
rect 18142 9072 18198 9081
rect 18052 9036 18104 9042
rect 18142 9007 18198 9016
rect 18052 8978 18104 8984
rect 18064 8634 18092 8978
rect 18142 8936 18198 8945
rect 18248 8906 18276 9415
rect 18142 8871 18198 8880
rect 18236 8900 18288 8906
rect 18156 8838 18184 8871
rect 18236 8842 18288 8848
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 18282 8732 18578 8752
rect 18338 8730 18362 8732
rect 18418 8730 18442 8732
rect 18498 8730 18522 8732
rect 18360 8678 18362 8730
rect 18424 8678 18436 8730
rect 18498 8678 18500 8730
rect 18338 8676 18362 8678
rect 18418 8676 18442 8678
rect 18498 8676 18522 8678
rect 18282 8656 18578 8676
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 18144 8288 18196 8294
rect 18144 8230 18196 8236
rect 18156 7410 18184 8230
rect 18282 7644 18578 7664
rect 18338 7642 18362 7644
rect 18418 7642 18442 7644
rect 18498 7642 18522 7644
rect 18360 7590 18362 7642
rect 18424 7590 18436 7642
rect 18498 7590 18500 7642
rect 18338 7588 18362 7590
rect 18418 7588 18442 7590
rect 18498 7588 18522 7590
rect 18282 7568 18578 7588
rect 18144 7404 18196 7410
rect 18144 7346 18196 7352
rect 17972 7126 18092 7154
rect 17958 7032 18014 7041
rect 17788 6956 17908 6984
rect 17958 6967 18014 6976
rect 17880 6390 17908 6956
rect 17972 6934 18000 6967
rect 17960 6928 18012 6934
rect 17960 6870 18012 6876
rect 17960 6792 18012 6798
rect 17960 6734 18012 6740
rect 17972 6458 18000 6734
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 17868 6384 17920 6390
rect 17868 6326 17920 6332
rect 17776 6248 17828 6254
rect 17776 6190 17828 6196
rect 17788 4486 17816 6190
rect 17958 6080 18014 6089
rect 17958 6015 18014 6024
rect 17972 5846 18000 6015
rect 17960 5840 18012 5846
rect 17960 5782 18012 5788
rect 17776 4480 17828 4486
rect 17776 4422 17828 4428
rect 17788 2961 17816 4422
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 17774 2952 17830 2961
rect 17774 2887 17830 2896
rect 17682 2000 17738 2009
rect 17682 1935 17738 1944
rect 17500 1760 17552 1766
rect 17500 1702 17552 1708
rect 17880 480 17908 4082
rect 17960 4072 18012 4078
rect 17960 4014 18012 4020
rect 17972 3369 18000 4014
rect 17958 3360 18014 3369
rect 17958 3295 18014 3304
rect 18064 3126 18092 7126
rect 18144 6792 18196 6798
rect 18144 6734 18196 6740
rect 18156 6254 18184 6734
rect 18282 6556 18578 6576
rect 18338 6554 18362 6556
rect 18418 6554 18442 6556
rect 18498 6554 18522 6556
rect 18360 6502 18362 6554
rect 18424 6502 18436 6554
rect 18498 6502 18500 6554
rect 18338 6500 18362 6502
rect 18418 6500 18442 6502
rect 18498 6500 18522 6502
rect 18282 6480 18578 6500
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 18282 5468 18578 5488
rect 18338 5466 18362 5468
rect 18418 5466 18442 5468
rect 18498 5466 18522 5468
rect 18360 5414 18362 5466
rect 18424 5414 18436 5466
rect 18498 5414 18500 5466
rect 18338 5412 18362 5414
rect 18418 5412 18442 5414
rect 18498 5412 18522 5414
rect 18282 5392 18578 5412
rect 18144 5160 18196 5166
rect 18144 5102 18196 5108
rect 18156 4026 18184 5102
rect 18282 4380 18578 4400
rect 18338 4378 18362 4380
rect 18418 4378 18442 4380
rect 18498 4378 18522 4380
rect 18360 4326 18362 4378
rect 18424 4326 18436 4378
rect 18498 4326 18500 4378
rect 18338 4324 18362 4326
rect 18418 4324 18442 4326
rect 18498 4324 18522 4326
rect 18282 4304 18578 4324
rect 18156 3998 18276 4026
rect 18248 3534 18276 3998
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 18282 3292 18578 3312
rect 18338 3290 18362 3292
rect 18418 3290 18442 3292
rect 18498 3290 18522 3292
rect 18360 3238 18362 3290
rect 18424 3238 18436 3290
rect 18498 3238 18500 3290
rect 18338 3236 18362 3238
rect 18418 3236 18442 3238
rect 18498 3236 18522 3238
rect 18282 3216 18578 3236
rect 18052 3120 18104 3126
rect 18052 3062 18104 3068
rect 18282 2204 18578 2224
rect 18338 2202 18362 2204
rect 18418 2202 18442 2204
rect 18498 2202 18522 2204
rect 18360 2150 18362 2202
rect 18424 2150 18436 2202
rect 18498 2150 18500 2202
rect 18338 2148 18362 2150
rect 18418 2148 18442 2150
rect 18498 2148 18522 2150
rect 18282 2128 18578 2148
rect 18616 1601 18644 12922
rect 18708 2514 18736 13126
rect 18800 12646 18828 13194
rect 18788 12640 18840 12646
rect 18788 12582 18840 12588
rect 18800 10742 18828 12582
rect 18984 12458 19012 16623
rect 19156 16594 19208 16600
rect 19168 16402 19196 16594
rect 19260 16522 19288 18022
rect 19352 17678 19380 18226
rect 19340 17672 19392 17678
rect 19340 17614 19392 17620
rect 19248 16516 19300 16522
rect 19248 16458 19300 16464
rect 19168 16374 19288 16402
rect 19260 14958 19288 16374
rect 19444 16096 19472 18770
rect 19352 16068 19472 16096
rect 19352 15434 19380 16068
rect 19432 15972 19484 15978
rect 19432 15914 19484 15920
rect 19340 15428 19392 15434
rect 19340 15370 19392 15376
rect 19248 14952 19300 14958
rect 19248 14894 19300 14900
rect 19248 14816 19300 14822
rect 19248 14758 19300 14764
rect 19260 14618 19288 14758
rect 19248 14612 19300 14618
rect 19248 14554 19300 14560
rect 19260 13870 19288 14554
rect 19352 14482 19380 15370
rect 19444 14550 19472 15914
rect 19432 14544 19484 14550
rect 19432 14486 19484 14492
rect 19340 14476 19392 14482
rect 19340 14418 19392 14424
rect 19432 14408 19484 14414
rect 19432 14350 19484 14356
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 19248 13864 19300 13870
rect 19248 13806 19300 13812
rect 19156 13524 19208 13530
rect 19156 13466 19208 13472
rect 19064 12708 19116 12714
rect 19064 12650 19116 12656
rect 18892 12430 19012 12458
rect 18892 10810 18920 12430
rect 18972 12368 19024 12374
rect 18972 12310 19024 12316
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 18788 10736 18840 10742
rect 18788 10678 18840 10684
rect 18878 10704 18934 10713
rect 18878 10639 18934 10648
rect 18786 10568 18842 10577
rect 18786 10503 18842 10512
rect 18800 9081 18828 10503
rect 18786 9072 18842 9081
rect 18786 9007 18842 9016
rect 18788 8968 18840 8974
rect 18788 8910 18840 8916
rect 18800 8634 18828 8910
rect 18788 8628 18840 8634
rect 18788 8570 18840 8576
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 18800 8090 18828 8434
rect 18892 8129 18920 10639
rect 18984 8922 19012 12310
rect 19076 12102 19104 12650
rect 19064 12096 19116 12102
rect 19064 12038 19116 12044
rect 19076 11762 19104 12038
rect 19064 11756 19116 11762
rect 19064 11698 19116 11704
rect 19168 10606 19196 13466
rect 19248 13388 19300 13394
rect 19248 13330 19300 13336
rect 19260 11898 19288 13330
rect 19248 11892 19300 11898
rect 19248 11834 19300 11840
rect 19246 10704 19302 10713
rect 19352 10674 19380 14282
rect 19444 11694 19472 14350
rect 19432 11688 19484 11694
rect 19432 11630 19484 11636
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 19246 10639 19302 10648
rect 19340 10668 19392 10674
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 19260 10266 19288 10639
rect 19340 10610 19392 10616
rect 19340 10532 19392 10538
rect 19340 10474 19392 10480
rect 19248 10260 19300 10266
rect 19248 10202 19300 10208
rect 19156 10192 19208 10198
rect 19352 10146 19380 10474
rect 19208 10140 19380 10146
rect 19156 10134 19380 10140
rect 19168 10118 19380 10134
rect 19168 9518 19196 10118
rect 19156 9512 19208 9518
rect 19156 9454 19208 9460
rect 19154 9344 19210 9353
rect 19154 9279 19210 9288
rect 19168 9178 19196 9279
rect 19156 9172 19208 9178
rect 19156 9114 19208 9120
rect 18984 8894 19288 8922
rect 19064 8832 19116 8838
rect 19064 8774 19116 8780
rect 18972 8356 19024 8362
rect 18972 8298 19024 8304
rect 18878 8120 18934 8129
rect 18788 8084 18840 8090
rect 18878 8055 18934 8064
rect 18788 8026 18840 8032
rect 18880 8016 18932 8022
rect 18880 7958 18932 7964
rect 18786 7576 18842 7585
rect 18786 7511 18788 7520
rect 18840 7511 18842 7520
rect 18788 7482 18840 7488
rect 18892 6730 18920 7958
rect 18880 6724 18932 6730
rect 18880 6666 18932 6672
rect 18892 5914 18920 6666
rect 18880 5908 18932 5914
rect 18880 5850 18932 5856
rect 18984 5234 19012 8298
rect 18972 5228 19024 5234
rect 18972 5170 19024 5176
rect 18788 4684 18840 4690
rect 18788 4626 18840 4632
rect 18696 2508 18748 2514
rect 18696 2450 18748 2456
rect 18602 1592 18658 1601
rect 18602 1527 18658 1536
rect 18328 1420 18380 1426
rect 18328 1362 18380 1368
rect 18340 480 18368 1362
rect 18800 1057 18828 4626
rect 18972 4480 19024 4486
rect 18972 4422 19024 4428
rect 18984 4146 19012 4422
rect 18972 4140 19024 4146
rect 18972 4082 19024 4088
rect 18984 3670 19012 4082
rect 19076 3670 19104 8774
rect 19156 7948 19208 7954
rect 19156 7890 19208 7896
rect 19168 7410 19196 7890
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 19156 6656 19208 6662
rect 19156 6598 19208 6604
rect 18972 3664 19024 3670
rect 18972 3606 19024 3612
rect 19064 3664 19116 3670
rect 19064 3606 19116 3612
rect 19062 3224 19118 3233
rect 19062 3159 19118 3168
rect 19076 1426 19104 3159
rect 19168 2990 19196 6598
rect 19156 2984 19208 2990
rect 19156 2926 19208 2932
rect 19064 1420 19116 1426
rect 19064 1362 19116 1368
rect 18880 1352 18932 1358
rect 18880 1294 18932 1300
rect 18786 1048 18842 1057
rect 18786 983 18842 992
rect 18892 480 18920 1294
rect 6276 332 6328 338
rect 6276 274 6328 280
rect 6366 0 6422 480
rect 6826 0 6882 480
rect 7378 0 7434 480
rect 7838 0 7894 480
rect 8298 0 8354 480
rect 8758 0 8814 480
rect 9218 0 9274 480
rect 9770 0 9826 480
rect 10230 0 10286 480
rect 10690 0 10746 480
rect 11150 0 11206 480
rect 11702 0 11758 480
rect 12162 0 12218 480
rect 12622 0 12678 480
rect 13082 0 13138 480
rect 13542 0 13598 480
rect 14094 0 14150 480
rect 14554 0 14610 480
rect 15014 0 15070 480
rect 15474 0 15530 480
rect 15934 0 15990 480
rect 16486 0 16542 480
rect 16946 0 17002 480
rect 17406 0 17462 480
rect 17866 0 17922 480
rect 18326 0 18382 480
rect 18878 0 18934 480
rect 19260 241 19288 8894
rect 19444 6322 19472 11494
rect 19536 6882 19564 20046
rect 20076 19916 20128 19922
rect 20076 19858 20128 19864
rect 19984 18692 20036 18698
rect 19984 18634 20036 18640
rect 19996 18154 20024 18634
rect 20088 18170 20116 19858
rect 20168 19848 20220 19854
rect 20168 19790 20220 19796
rect 20180 19378 20208 19790
rect 20168 19372 20220 19378
rect 20168 19314 20220 19320
rect 20088 18154 20208 18170
rect 19984 18148 20036 18154
rect 20088 18148 20220 18154
rect 20088 18142 20168 18148
rect 19984 18090 20036 18096
rect 20168 18090 20220 18096
rect 20444 18148 20496 18154
rect 20444 18090 20496 18096
rect 19800 17740 19852 17746
rect 19800 17682 19852 17688
rect 19708 17060 19760 17066
rect 19708 17002 19760 17008
rect 19616 16720 19668 16726
rect 19616 16662 19668 16668
rect 19628 14618 19656 16662
rect 19720 16658 19748 17002
rect 19708 16652 19760 16658
rect 19708 16594 19760 16600
rect 19812 15570 19840 17682
rect 19984 16788 20036 16794
rect 19984 16730 20036 16736
rect 19890 15736 19946 15745
rect 19890 15671 19892 15680
rect 19944 15671 19946 15680
rect 19892 15642 19944 15648
rect 19800 15564 19852 15570
rect 19800 15506 19852 15512
rect 19616 14612 19668 14618
rect 19616 14554 19668 14560
rect 19708 12300 19760 12306
rect 19708 12242 19760 12248
rect 19720 11286 19748 12242
rect 19708 11280 19760 11286
rect 19708 11222 19760 11228
rect 19616 10124 19668 10130
rect 19616 10066 19668 10072
rect 19628 9722 19656 10066
rect 19616 9716 19668 9722
rect 19616 9658 19668 9664
rect 19708 9444 19760 9450
rect 19708 9386 19760 9392
rect 19720 7342 19748 9386
rect 19812 7546 19840 15506
rect 19996 14929 20024 16730
rect 19982 14920 20038 14929
rect 19982 14855 20038 14864
rect 19984 13864 20036 13870
rect 19984 13806 20036 13812
rect 20352 13864 20404 13870
rect 20352 13806 20404 13812
rect 19890 13016 19946 13025
rect 19890 12951 19946 12960
rect 19904 12442 19932 12951
rect 19892 12436 19944 12442
rect 19892 12378 19944 12384
rect 19996 12374 20024 13806
rect 19984 12368 20036 12374
rect 19984 12310 20036 12316
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 19892 8900 19944 8906
rect 19892 8842 19944 8848
rect 19800 7540 19852 7546
rect 19800 7482 19852 7488
rect 19708 7336 19760 7342
rect 19708 7278 19760 7284
rect 19536 6854 19748 6882
rect 19524 6724 19576 6730
rect 19524 6666 19576 6672
rect 19432 6316 19484 6322
rect 19432 6258 19484 6264
rect 19430 5264 19486 5273
rect 19430 5199 19486 5208
rect 19444 2990 19472 5199
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 19340 2848 19392 2854
rect 19340 2790 19392 2796
rect 19352 480 19380 2790
rect 19536 1494 19564 6666
rect 19614 5128 19670 5137
rect 19614 5063 19670 5072
rect 19628 4826 19656 5063
rect 19720 5030 19748 6854
rect 19904 5846 19932 8842
rect 20076 8288 20128 8294
rect 20076 8230 20128 8236
rect 19892 5840 19944 5846
rect 19892 5782 19944 5788
rect 19708 5024 19760 5030
rect 19708 4966 19760 4972
rect 19616 4820 19668 4826
rect 19616 4762 19668 4768
rect 19798 3632 19854 3641
rect 19798 3567 19854 3576
rect 19524 1488 19576 1494
rect 19524 1430 19576 1436
rect 19812 480 19840 3567
rect 20088 3505 20116 8230
rect 20074 3496 20130 3505
rect 20074 3431 20130 3440
rect 20180 3380 20208 9658
rect 20258 4040 20314 4049
rect 20258 3975 20314 3984
rect 20088 3352 20208 3380
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 19996 1902 20024 2450
rect 19984 1896 20036 1902
rect 19984 1838 20036 1844
rect 20088 649 20116 3352
rect 20168 2916 20220 2922
rect 20168 2858 20220 2864
rect 20180 2650 20208 2858
rect 20168 2644 20220 2650
rect 20168 2586 20220 2592
rect 20074 640 20130 649
rect 20074 575 20130 584
rect 20272 480 20300 3975
rect 20364 3777 20392 13806
rect 20456 9994 20484 18090
rect 20718 17640 20774 17649
rect 20718 17575 20774 17584
rect 20732 16250 20760 17575
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 20718 15328 20774 15337
rect 20718 15263 20774 15272
rect 20732 15162 20760 15263
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20720 13728 20772 13734
rect 20720 13670 20772 13676
rect 20732 13569 20760 13670
rect 20718 13560 20774 13569
rect 20718 13495 20774 13504
rect 20812 10464 20864 10470
rect 20812 10406 20864 10412
rect 20628 10056 20680 10062
rect 20628 9998 20680 10004
rect 20444 9988 20496 9994
rect 20444 9930 20496 9936
rect 20456 9722 20484 9930
rect 20536 9920 20588 9926
rect 20536 9862 20588 9868
rect 20444 9716 20496 9722
rect 20444 9658 20496 9664
rect 20548 8498 20576 9862
rect 20536 8492 20588 8498
rect 20536 8434 20588 8440
rect 20536 8356 20588 8362
rect 20536 8298 20588 8304
rect 20548 7274 20576 8298
rect 20640 7546 20668 9998
rect 20824 9518 20852 10406
rect 20812 9512 20864 9518
rect 20812 9454 20864 9460
rect 20628 7540 20680 7546
rect 20628 7482 20680 7488
rect 20536 7268 20588 7274
rect 20536 7210 20588 7216
rect 20548 5370 20576 7210
rect 20536 5364 20588 5370
rect 20536 5306 20588 5312
rect 20640 5166 20668 7482
rect 20628 5160 20680 5166
rect 20628 5102 20680 5108
rect 20534 4312 20590 4321
rect 20534 4247 20590 4256
rect 20548 4078 20576 4247
rect 20536 4072 20588 4078
rect 20536 4014 20588 4020
rect 21732 3936 21784 3942
rect 20534 3904 20590 3913
rect 21732 3878 21784 3884
rect 20534 3839 20590 3848
rect 20350 3768 20406 3777
rect 20350 3703 20406 3712
rect 20548 2990 20576 3839
rect 20720 3188 20772 3194
rect 20720 3130 20772 3136
rect 20536 2984 20588 2990
rect 20536 2926 20588 2932
rect 20732 480 20760 3130
rect 21272 3120 21324 3126
rect 21272 3062 21324 3068
rect 21284 480 21312 3062
rect 21744 480 21772 3878
rect 22652 2916 22704 2922
rect 22652 2858 22704 2864
rect 22192 2848 22244 2854
rect 22192 2790 22244 2796
rect 22204 480 22232 2790
rect 22664 480 22692 2858
rect 19246 232 19302 241
rect 19246 167 19302 176
rect 19338 0 19394 480
rect 19798 0 19854 480
rect 20258 0 20314 480
rect 20718 0 20774 480
rect 21270 0 21326 480
rect 21730 0 21786 480
rect 22190 0 22246 480
rect 22650 0 22706 480
<< via2 >>
rect 3882 22616 3938 22672
rect 3514 22208 3570 22264
rect 3146 21256 3202 21312
rect 18970 22616 19026 22672
rect 4250 21800 4306 21856
rect 4066 20868 4122 20904
rect 4066 20848 4068 20868
rect 4068 20848 4120 20868
rect 4120 20848 4122 20868
rect 3974 20440 4030 20496
rect 2870 18536 2926 18592
rect 1950 17720 2006 17776
rect 1030 15000 1086 15056
rect 1674 14592 1730 14648
rect 3054 18128 3110 18184
rect 2962 16768 3018 16824
rect 2686 16360 2742 16416
rect 2134 13232 2190 13288
rect 2778 13640 2834 13696
rect 3146 14048 3202 14104
rect 2962 10240 3018 10296
rect 3330 19488 3386 19544
rect 3330 15816 3386 15872
rect 3514 15408 3570 15464
rect 3238 10648 3294 10704
rect 2962 9696 3018 9752
rect 2042 6840 2098 6896
rect 1674 3440 1730 3496
rect 1766 2624 1822 2680
rect 1306 584 1362 640
rect 2226 6024 2282 6080
rect 2226 2916 2282 2952
rect 2226 2896 2228 2916
rect 2228 2896 2280 2916
rect 2280 2896 2282 2916
rect 2778 7112 2834 7168
rect 2870 6704 2926 6760
rect 2594 6332 2596 6352
rect 2596 6332 2648 6352
rect 2648 6332 2650 6352
rect 2594 6296 2650 6332
rect 2502 6024 2558 6080
rect 2502 5636 2558 5672
rect 2502 5616 2504 5636
rect 2504 5616 2556 5636
rect 2556 5616 2558 5636
rect 2410 4936 2466 4992
rect 2134 2352 2190 2408
rect 3330 9696 3386 9752
rect 4066 19896 4122 19952
rect 4066 19080 4122 19136
rect 4158 17176 4214 17232
rect 4421 20698 4477 20700
rect 4501 20698 4557 20700
rect 4581 20698 4637 20700
rect 4661 20698 4717 20700
rect 4421 20646 4447 20698
rect 4447 20646 4477 20698
rect 4501 20646 4511 20698
rect 4511 20646 4557 20698
rect 4581 20646 4627 20698
rect 4627 20646 4637 20698
rect 4661 20646 4691 20698
rect 4691 20646 4717 20698
rect 4421 20644 4477 20646
rect 4501 20644 4557 20646
rect 4581 20644 4637 20646
rect 4661 20644 4717 20646
rect 4421 19610 4477 19612
rect 4501 19610 4557 19612
rect 4581 19610 4637 19612
rect 4661 19610 4717 19612
rect 4421 19558 4447 19610
rect 4447 19558 4477 19610
rect 4501 19558 4511 19610
rect 4511 19558 4557 19610
rect 4581 19558 4627 19610
rect 4627 19558 4637 19610
rect 4661 19558 4691 19610
rect 4691 19558 4717 19610
rect 4421 19556 4477 19558
rect 4501 19556 4557 19558
rect 4581 19556 4637 19558
rect 4661 19556 4717 19558
rect 4421 18522 4477 18524
rect 4501 18522 4557 18524
rect 4581 18522 4637 18524
rect 4661 18522 4717 18524
rect 4421 18470 4447 18522
rect 4447 18470 4477 18522
rect 4501 18470 4511 18522
rect 4511 18470 4557 18522
rect 4581 18470 4627 18522
rect 4627 18470 4637 18522
rect 4661 18470 4691 18522
rect 4691 18470 4717 18522
rect 4421 18468 4477 18470
rect 4501 18468 4557 18470
rect 4581 18468 4637 18470
rect 4661 18468 4717 18470
rect 4421 17434 4477 17436
rect 4501 17434 4557 17436
rect 4581 17434 4637 17436
rect 4661 17434 4717 17436
rect 4421 17382 4447 17434
rect 4447 17382 4477 17434
rect 4501 17382 4511 17434
rect 4511 17382 4557 17434
rect 4581 17382 4627 17434
rect 4627 17382 4637 17434
rect 4661 17382 4691 17434
rect 4691 17382 4717 17434
rect 4421 17380 4477 17382
rect 4501 17380 4557 17382
rect 4581 17380 4637 17382
rect 4661 17380 4717 17382
rect 4421 16346 4477 16348
rect 4501 16346 4557 16348
rect 4581 16346 4637 16348
rect 4661 16346 4717 16348
rect 4421 16294 4447 16346
rect 4447 16294 4477 16346
rect 4501 16294 4511 16346
rect 4511 16294 4557 16346
rect 4581 16294 4627 16346
rect 4627 16294 4637 16346
rect 4661 16294 4691 16346
rect 4691 16294 4717 16346
rect 4421 16292 4477 16294
rect 4501 16292 4557 16294
rect 4581 16292 4637 16294
rect 4661 16292 4717 16294
rect 3974 13504 4030 13560
rect 3882 11872 3938 11928
rect 3790 11328 3846 11384
rect 3790 9560 3846 9616
rect 3790 8200 3846 8256
rect 3698 7248 3754 7304
rect 3238 5208 3294 5264
rect 3146 3984 3202 4040
rect 3330 3576 3386 3632
rect 3054 3304 3110 3360
rect 3054 3168 3110 3224
rect 2778 3068 2780 3088
rect 2780 3068 2832 3088
rect 2832 3068 2834 3088
rect 2778 3032 2834 3068
rect 2226 1400 2282 1456
rect 3882 5480 3938 5536
rect 3790 5072 3846 5128
rect 3606 4664 3662 4720
rect 3698 3576 3754 3632
rect 3514 1944 3570 2000
rect 3882 4528 3938 4584
rect 4066 12708 4122 12744
rect 4066 12688 4068 12708
rect 4068 12688 4120 12708
rect 4120 12688 4122 12708
rect 4066 12280 4122 12336
rect 4250 13504 4306 13560
rect 4421 15258 4477 15260
rect 4501 15258 4557 15260
rect 4581 15258 4637 15260
rect 4661 15258 4717 15260
rect 4421 15206 4447 15258
rect 4447 15206 4477 15258
rect 4501 15206 4511 15258
rect 4511 15206 4557 15258
rect 4581 15206 4627 15258
rect 4627 15206 4637 15258
rect 4661 15206 4691 15258
rect 4691 15206 4717 15258
rect 4421 15204 4477 15206
rect 4501 15204 4557 15206
rect 4581 15204 4637 15206
rect 4661 15204 4717 15206
rect 4421 14170 4477 14172
rect 4501 14170 4557 14172
rect 4581 14170 4637 14172
rect 4661 14170 4717 14172
rect 4421 14118 4447 14170
rect 4447 14118 4477 14170
rect 4501 14118 4511 14170
rect 4511 14118 4557 14170
rect 4581 14118 4627 14170
rect 4627 14118 4637 14170
rect 4661 14118 4691 14170
rect 4691 14118 4717 14170
rect 4421 14116 4477 14118
rect 4501 14116 4557 14118
rect 4581 14116 4637 14118
rect 4661 14116 4717 14118
rect 4434 13912 4490 13968
rect 4421 13082 4477 13084
rect 4501 13082 4557 13084
rect 4581 13082 4637 13084
rect 4661 13082 4717 13084
rect 4421 13030 4447 13082
rect 4447 13030 4477 13082
rect 4501 13030 4511 13082
rect 4511 13030 4557 13082
rect 4581 13030 4627 13082
rect 4627 13030 4637 13082
rect 4661 13030 4691 13082
rect 4691 13030 4717 13082
rect 4421 13028 4477 13030
rect 4501 13028 4557 13030
rect 4581 13028 4637 13030
rect 4661 13028 4717 13030
rect 4421 11994 4477 11996
rect 4501 11994 4557 11996
rect 4581 11994 4637 11996
rect 4661 11994 4717 11996
rect 4421 11942 4447 11994
rect 4447 11942 4477 11994
rect 4501 11942 4511 11994
rect 4511 11942 4557 11994
rect 4581 11942 4627 11994
rect 4627 11942 4637 11994
rect 4661 11942 4691 11994
rect 4691 11942 4717 11994
rect 4421 11940 4477 11942
rect 4501 11940 4557 11942
rect 4581 11940 4637 11942
rect 4661 11940 4717 11942
rect 4066 10532 4122 10568
rect 4066 10512 4068 10532
rect 4068 10512 4120 10532
rect 4120 10512 4122 10532
rect 4421 10906 4477 10908
rect 4501 10906 4557 10908
rect 4581 10906 4637 10908
rect 4661 10906 4717 10908
rect 4421 10854 4447 10906
rect 4447 10854 4477 10906
rect 4501 10854 4511 10906
rect 4511 10854 4557 10906
rect 4581 10854 4627 10906
rect 4627 10854 4637 10906
rect 4661 10854 4691 10906
rect 4691 10854 4717 10906
rect 4421 10852 4477 10854
rect 4501 10852 4557 10854
rect 4581 10852 4637 10854
rect 4661 10852 4717 10854
rect 4342 10512 4398 10568
rect 4066 9172 4122 9208
rect 4066 9152 4068 9172
rect 4068 9152 4120 9172
rect 4120 9152 4122 9172
rect 4066 8608 4122 8664
rect 4066 7792 4122 7848
rect 4421 9818 4477 9820
rect 4501 9818 4557 9820
rect 4581 9818 4637 9820
rect 4661 9818 4717 9820
rect 4421 9766 4447 9818
rect 4447 9766 4477 9818
rect 4501 9766 4511 9818
rect 4511 9766 4557 9818
rect 4581 9766 4627 9818
rect 4627 9766 4637 9818
rect 4661 9766 4691 9818
rect 4691 9766 4717 9818
rect 4421 9764 4477 9766
rect 4501 9764 4557 9766
rect 4581 9764 4637 9766
rect 4661 9764 4717 9766
rect 4421 8730 4477 8732
rect 4501 8730 4557 8732
rect 4581 8730 4637 8732
rect 4661 8730 4717 8732
rect 4421 8678 4447 8730
rect 4447 8678 4477 8730
rect 4501 8678 4511 8730
rect 4511 8678 4557 8730
rect 4581 8678 4627 8730
rect 4627 8678 4637 8730
rect 4661 8678 4691 8730
rect 4691 8678 4717 8730
rect 4421 8676 4477 8678
rect 4501 8676 4557 8678
rect 4581 8676 4637 8678
rect 4661 8676 4717 8678
rect 4421 7642 4477 7644
rect 4501 7642 4557 7644
rect 4581 7642 4637 7644
rect 4661 7642 4717 7644
rect 4421 7590 4447 7642
rect 4447 7590 4477 7642
rect 4501 7590 4511 7642
rect 4511 7590 4557 7642
rect 4581 7590 4627 7642
rect 4627 7590 4637 7642
rect 4661 7590 4691 7642
rect 4691 7590 4717 7642
rect 4421 7588 4477 7590
rect 4501 7588 4557 7590
rect 4581 7588 4637 7590
rect 4661 7588 4717 7590
rect 4421 6554 4477 6556
rect 4501 6554 4557 6556
rect 4581 6554 4637 6556
rect 4661 6554 4717 6556
rect 4421 6502 4447 6554
rect 4447 6502 4477 6554
rect 4501 6502 4511 6554
rect 4511 6502 4557 6554
rect 4581 6502 4627 6554
rect 4627 6502 4637 6554
rect 4661 6502 4691 6554
rect 4691 6502 4717 6554
rect 4421 6500 4477 6502
rect 4501 6500 4557 6502
rect 4581 6500 4637 6502
rect 4661 6500 4717 6502
rect 4618 6296 4674 6352
rect 4066 5092 4122 5128
rect 4066 5072 4068 5092
rect 4068 5072 4120 5092
rect 4120 5072 4122 5092
rect 3974 4256 4030 4312
rect 4066 3848 4122 3904
rect 4421 5466 4477 5468
rect 4501 5466 4557 5468
rect 4581 5466 4637 5468
rect 4661 5466 4717 5468
rect 4421 5414 4447 5466
rect 4447 5414 4477 5466
rect 4501 5414 4511 5466
rect 4511 5414 4557 5466
rect 4581 5414 4627 5466
rect 4627 5414 4637 5466
rect 4661 5414 4691 5466
rect 4691 5414 4717 5466
rect 4421 5412 4477 5414
rect 4501 5412 4557 5414
rect 4581 5412 4637 5414
rect 4661 5412 4717 5414
rect 4421 4378 4477 4380
rect 4501 4378 4557 4380
rect 4581 4378 4637 4380
rect 4661 4378 4717 4380
rect 4421 4326 4447 4378
rect 4447 4326 4477 4378
rect 4501 4326 4511 4378
rect 4511 4326 4557 4378
rect 4581 4326 4627 4378
rect 4627 4326 4637 4378
rect 4661 4326 4691 4378
rect 4691 4326 4717 4378
rect 4421 4324 4477 4326
rect 4501 4324 4557 4326
rect 4581 4324 4637 4326
rect 4661 4324 4717 4326
rect 4434 4020 4436 4040
rect 4436 4020 4488 4040
rect 4488 4020 4490 4040
rect 4434 3984 4490 4020
rect 4066 2760 4122 2816
rect 4421 3290 4477 3292
rect 4501 3290 4557 3292
rect 4581 3290 4637 3292
rect 4661 3290 4717 3292
rect 4421 3238 4447 3290
rect 4447 3238 4477 3290
rect 4501 3238 4511 3290
rect 4511 3238 4557 3290
rect 4581 3238 4627 3290
rect 4627 3238 4637 3290
rect 4661 3238 4691 3290
rect 4691 3238 4717 3290
rect 4421 3236 4477 3238
rect 4501 3236 4557 3238
rect 4581 3236 4637 3238
rect 4661 3236 4717 3238
rect 5078 8336 5134 8392
rect 5262 5752 5318 5808
rect 5906 9968 5962 10024
rect 5814 5616 5870 5672
rect 5078 3848 5134 3904
rect 4421 2202 4477 2204
rect 4501 2202 4557 2204
rect 4581 2202 4637 2204
rect 4661 2202 4717 2204
rect 4421 2150 4447 2202
rect 4447 2150 4477 2202
rect 4501 2150 4511 2202
rect 4511 2150 4557 2202
rect 4581 2150 4627 2202
rect 4627 2150 4637 2202
rect 4661 2150 4691 2202
rect 4691 2150 4717 2202
rect 4421 2148 4477 2150
rect 4501 2148 4557 2150
rect 4581 2148 4637 2150
rect 4661 2148 4717 2150
rect 5170 3440 5226 3496
rect 5722 4936 5778 4992
rect 5446 2760 5502 2816
rect 6826 15544 6882 15600
rect 5630 2352 5686 2408
rect 6274 5888 6330 5944
rect 6550 9968 6606 10024
rect 3606 176 3662 232
rect 7102 10240 7158 10296
rect 7286 10140 7288 10160
rect 7288 10140 7340 10160
rect 7340 10140 7342 10160
rect 7286 10104 7342 10140
rect 6366 3440 6422 3496
rect 6642 5636 6698 5672
rect 6642 5616 6644 5636
rect 6644 5616 6696 5636
rect 6696 5616 6698 5636
rect 7194 6976 7250 7032
rect 7010 4528 7066 4584
rect 6642 992 6698 1048
rect 7286 6024 7342 6080
rect 7378 5888 7434 5944
rect 7378 4120 7434 4176
rect 7378 3304 7434 3360
rect 7378 2896 7434 2952
rect 7886 20154 7942 20156
rect 7966 20154 8022 20156
rect 8046 20154 8102 20156
rect 8126 20154 8182 20156
rect 7886 20102 7912 20154
rect 7912 20102 7942 20154
rect 7966 20102 7976 20154
rect 7976 20102 8022 20154
rect 8046 20102 8092 20154
rect 8092 20102 8102 20154
rect 8126 20102 8156 20154
rect 8156 20102 8182 20154
rect 7886 20100 7942 20102
rect 7966 20100 8022 20102
rect 8046 20100 8102 20102
rect 8126 20100 8182 20102
rect 7886 19066 7942 19068
rect 7966 19066 8022 19068
rect 8046 19066 8102 19068
rect 8126 19066 8182 19068
rect 7886 19014 7912 19066
rect 7912 19014 7942 19066
rect 7966 19014 7976 19066
rect 7976 19014 8022 19066
rect 8046 19014 8092 19066
rect 8092 19014 8102 19066
rect 8126 19014 8156 19066
rect 8156 19014 8182 19066
rect 7886 19012 7942 19014
rect 7966 19012 8022 19014
rect 8046 19012 8102 19014
rect 8126 19012 8182 19014
rect 7886 17978 7942 17980
rect 7966 17978 8022 17980
rect 8046 17978 8102 17980
rect 8126 17978 8182 17980
rect 7886 17926 7912 17978
rect 7912 17926 7942 17978
rect 7966 17926 7976 17978
rect 7976 17926 8022 17978
rect 8046 17926 8092 17978
rect 8092 17926 8102 17978
rect 8126 17926 8156 17978
rect 8156 17926 8182 17978
rect 7886 17924 7942 17926
rect 7966 17924 8022 17926
rect 8046 17924 8102 17926
rect 8126 17924 8182 17926
rect 7886 16890 7942 16892
rect 7966 16890 8022 16892
rect 8046 16890 8102 16892
rect 8126 16890 8182 16892
rect 7886 16838 7912 16890
rect 7912 16838 7942 16890
rect 7966 16838 7976 16890
rect 7976 16838 8022 16890
rect 8046 16838 8092 16890
rect 8092 16838 8102 16890
rect 8126 16838 8156 16890
rect 8156 16838 8182 16890
rect 7886 16836 7942 16838
rect 7966 16836 8022 16838
rect 8046 16836 8102 16838
rect 8126 16836 8182 16838
rect 7886 15802 7942 15804
rect 7966 15802 8022 15804
rect 8046 15802 8102 15804
rect 8126 15802 8182 15804
rect 7886 15750 7912 15802
rect 7912 15750 7942 15802
rect 7966 15750 7976 15802
rect 7976 15750 8022 15802
rect 8046 15750 8092 15802
rect 8092 15750 8102 15802
rect 8126 15750 8156 15802
rect 8156 15750 8182 15802
rect 7886 15748 7942 15750
rect 7966 15748 8022 15750
rect 8046 15748 8102 15750
rect 8126 15748 8182 15750
rect 7886 14714 7942 14716
rect 7966 14714 8022 14716
rect 8046 14714 8102 14716
rect 8126 14714 8182 14716
rect 7886 14662 7912 14714
rect 7912 14662 7942 14714
rect 7966 14662 7976 14714
rect 7976 14662 8022 14714
rect 8046 14662 8092 14714
rect 8092 14662 8102 14714
rect 8126 14662 8156 14714
rect 8156 14662 8182 14714
rect 7886 14660 7942 14662
rect 7966 14660 8022 14662
rect 8046 14660 8102 14662
rect 8126 14660 8182 14662
rect 7886 13626 7942 13628
rect 7966 13626 8022 13628
rect 8046 13626 8102 13628
rect 8126 13626 8182 13628
rect 7886 13574 7912 13626
rect 7912 13574 7942 13626
rect 7966 13574 7976 13626
rect 7976 13574 8022 13626
rect 8046 13574 8092 13626
rect 8092 13574 8102 13626
rect 8126 13574 8156 13626
rect 8156 13574 8182 13626
rect 7886 13572 7942 13574
rect 7966 13572 8022 13574
rect 8046 13572 8102 13574
rect 8126 13572 8182 13574
rect 7886 12538 7942 12540
rect 7966 12538 8022 12540
rect 8046 12538 8102 12540
rect 8126 12538 8182 12540
rect 7886 12486 7912 12538
rect 7912 12486 7942 12538
rect 7966 12486 7976 12538
rect 7976 12486 8022 12538
rect 8046 12486 8092 12538
rect 8092 12486 8102 12538
rect 8126 12486 8156 12538
rect 8156 12486 8182 12538
rect 7886 12484 7942 12486
rect 7966 12484 8022 12486
rect 8046 12484 8102 12486
rect 8126 12484 8182 12486
rect 7562 10512 7618 10568
rect 7886 11450 7942 11452
rect 7966 11450 8022 11452
rect 8046 11450 8102 11452
rect 8126 11450 8182 11452
rect 7886 11398 7912 11450
rect 7912 11398 7942 11450
rect 7966 11398 7976 11450
rect 7976 11398 8022 11450
rect 8046 11398 8092 11450
rect 8092 11398 8102 11450
rect 8126 11398 8156 11450
rect 8156 11398 8182 11450
rect 7886 11396 7942 11398
rect 7966 11396 8022 11398
rect 8046 11396 8102 11398
rect 8126 11396 8182 11398
rect 7838 11056 7894 11112
rect 7886 10362 7942 10364
rect 7966 10362 8022 10364
rect 8046 10362 8102 10364
rect 8126 10362 8182 10364
rect 7886 10310 7912 10362
rect 7912 10310 7942 10362
rect 7966 10310 7976 10362
rect 7976 10310 8022 10362
rect 8046 10310 8092 10362
rect 8092 10310 8102 10362
rect 8126 10310 8156 10362
rect 8156 10310 8182 10362
rect 7886 10308 7942 10310
rect 7966 10308 8022 10310
rect 8046 10308 8102 10310
rect 8126 10308 8182 10310
rect 7886 9274 7942 9276
rect 7966 9274 8022 9276
rect 8046 9274 8102 9276
rect 8126 9274 8182 9276
rect 7886 9222 7912 9274
rect 7912 9222 7942 9274
rect 7966 9222 7976 9274
rect 7976 9222 8022 9274
rect 8046 9222 8092 9274
rect 8092 9222 8102 9274
rect 8126 9222 8156 9274
rect 8156 9222 8182 9274
rect 7886 9220 7942 9222
rect 7966 9220 8022 9222
rect 8046 9220 8102 9222
rect 8126 9220 8182 9222
rect 7562 7148 7564 7168
rect 7564 7148 7616 7168
rect 7616 7148 7618 7168
rect 7562 7112 7618 7148
rect 7470 2624 7526 2680
rect 7886 8186 7942 8188
rect 7966 8186 8022 8188
rect 8046 8186 8102 8188
rect 8126 8186 8182 8188
rect 7886 8134 7912 8186
rect 7912 8134 7942 8186
rect 7966 8134 7976 8186
rect 7976 8134 8022 8186
rect 8046 8134 8092 8186
rect 8092 8134 8102 8186
rect 8126 8134 8156 8186
rect 8156 8134 8182 8186
rect 7886 8132 7942 8134
rect 7966 8132 8022 8134
rect 8046 8132 8102 8134
rect 8126 8132 8182 8134
rect 7886 7098 7942 7100
rect 7966 7098 8022 7100
rect 8046 7098 8102 7100
rect 8126 7098 8182 7100
rect 7886 7046 7912 7098
rect 7912 7046 7942 7098
rect 7966 7046 7976 7098
rect 7976 7046 8022 7098
rect 8046 7046 8092 7098
rect 8092 7046 8102 7098
rect 8126 7046 8156 7098
rect 8156 7046 8182 7098
rect 7886 7044 7942 7046
rect 7966 7044 8022 7046
rect 8046 7044 8102 7046
rect 8126 7044 8182 7046
rect 7886 6010 7942 6012
rect 7966 6010 8022 6012
rect 8046 6010 8102 6012
rect 8126 6010 8182 6012
rect 7886 5958 7912 6010
rect 7912 5958 7942 6010
rect 7966 5958 7976 6010
rect 7976 5958 8022 6010
rect 8046 5958 8092 6010
rect 8092 5958 8102 6010
rect 8126 5958 8156 6010
rect 8156 5958 8182 6010
rect 7886 5956 7942 5958
rect 7966 5956 8022 5958
rect 8046 5956 8102 5958
rect 8126 5956 8182 5958
rect 7886 4922 7942 4924
rect 7966 4922 8022 4924
rect 8046 4922 8102 4924
rect 8126 4922 8182 4924
rect 7886 4870 7912 4922
rect 7912 4870 7942 4922
rect 7966 4870 7976 4922
rect 7976 4870 8022 4922
rect 8046 4870 8092 4922
rect 8092 4870 8102 4922
rect 8126 4870 8156 4922
rect 8156 4870 8182 4922
rect 7886 4868 7942 4870
rect 7966 4868 8022 4870
rect 8046 4868 8102 4870
rect 8126 4868 8182 4870
rect 7930 4664 7986 4720
rect 8114 4664 8170 4720
rect 7886 3834 7942 3836
rect 7966 3834 8022 3836
rect 8046 3834 8102 3836
rect 8126 3834 8182 3836
rect 7886 3782 7912 3834
rect 7912 3782 7942 3834
rect 7966 3782 7976 3834
rect 7976 3782 8022 3834
rect 8046 3782 8092 3834
rect 8092 3782 8102 3834
rect 8126 3782 8156 3834
rect 8156 3782 8182 3834
rect 7886 3780 7942 3782
rect 7966 3780 8022 3782
rect 8046 3780 8102 3782
rect 8126 3780 8182 3782
rect 7746 3068 7748 3088
rect 7748 3068 7800 3088
rect 7800 3068 7802 3088
rect 7746 3032 7802 3068
rect 7746 2916 7802 2952
rect 7746 2896 7748 2916
rect 7748 2896 7800 2916
rect 7800 2896 7802 2916
rect 7886 2746 7942 2748
rect 7966 2746 8022 2748
rect 8046 2746 8102 2748
rect 8126 2746 8182 2748
rect 7886 2694 7912 2746
rect 7912 2694 7942 2746
rect 7966 2694 7976 2746
rect 7976 2694 8022 2746
rect 8046 2694 8092 2746
rect 8092 2694 8102 2746
rect 8126 2694 8156 2746
rect 8156 2694 8182 2746
rect 7886 2692 7942 2694
rect 7966 2692 8022 2694
rect 8046 2692 8102 2694
rect 8126 2692 8182 2694
rect 8758 13912 8814 13968
rect 8574 10648 8630 10704
rect 8574 8336 8630 8392
rect 8390 5772 8446 5808
rect 8390 5752 8392 5772
rect 8392 5752 8444 5772
rect 8444 5752 8446 5772
rect 8482 2352 8538 2408
rect 8850 10512 8906 10568
rect 8850 6704 8906 6760
rect 8850 5616 8906 5672
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11378 20698
rect 11378 20646 11408 20698
rect 11432 20646 11442 20698
rect 11442 20646 11488 20698
rect 11512 20646 11558 20698
rect 11558 20646 11568 20698
rect 11592 20646 11622 20698
rect 11622 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11378 19610
rect 11378 19558 11408 19610
rect 11432 19558 11442 19610
rect 11442 19558 11488 19610
rect 11512 19558 11558 19610
rect 11558 19558 11568 19610
rect 11592 19558 11622 19610
rect 11622 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 10230 19116 10232 19136
rect 10232 19116 10284 19136
rect 10284 19116 10286 19136
rect 10230 19080 10286 19116
rect 8942 2760 8998 2816
rect 9862 16088 9918 16144
rect 9678 9016 9734 9072
rect 9586 7384 9642 7440
rect 9586 7248 9642 7304
rect 9586 5616 9642 5672
rect 9494 5208 9550 5264
rect 9678 5208 9734 5264
rect 9310 3168 9366 3224
rect 9310 2896 9366 2952
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11378 18522
rect 11378 18470 11408 18522
rect 11432 18470 11442 18522
rect 11442 18470 11488 18522
rect 11512 18470 11558 18522
rect 11558 18470 11568 18522
rect 11592 18470 11622 18522
rect 11622 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 10322 9460 10324 9480
rect 10324 9460 10376 9480
rect 10376 9460 10378 9480
rect 10322 9424 10378 9460
rect 9862 5480 9918 5536
rect 9954 4936 10010 4992
rect 9862 4664 9918 4720
rect 9862 3848 9918 3904
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11378 17434
rect 11378 17382 11408 17434
rect 11432 17382 11442 17434
rect 11442 17382 11488 17434
rect 11512 17382 11558 17434
rect 11558 17382 11568 17434
rect 11592 17382 11622 17434
rect 11622 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11378 16346
rect 11378 16294 11408 16346
rect 11432 16294 11442 16346
rect 11442 16294 11488 16346
rect 11512 16294 11558 16346
rect 11558 16294 11568 16346
rect 11592 16294 11622 16346
rect 11622 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 10966 15408 11022 15464
rect 11518 15972 11574 16008
rect 11518 15952 11520 15972
rect 11520 15952 11572 15972
rect 11572 15952 11574 15972
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11378 15258
rect 11378 15206 11408 15258
rect 11432 15206 11442 15258
rect 11442 15206 11488 15258
rect 11512 15206 11558 15258
rect 11558 15206 11568 15258
rect 11592 15206 11622 15258
rect 11622 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11378 14170
rect 11378 14118 11408 14170
rect 11432 14118 11442 14170
rect 11442 14118 11488 14170
rect 11512 14118 11558 14170
rect 11558 14118 11568 14170
rect 11592 14118 11622 14170
rect 11622 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11378 13082
rect 11378 13030 11408 13082
rect 11432 13030 11442 13082
rect 11442 13030 11488 13082
rect 11512 13030 11558 13082
rect 11558 13030 11568 13082
rect 11592 13030 11622 13082
rect 11622 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11242 12552 11298 12608
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11378 11994
rect 11378 11942 11408 11994
rect 11432 11942 11442 11994
rect 11442 11942 11488 11994
rect 11512 11942 11558 11994
rect 11558 11942 11568 11994
rect 11592 11942 11622 11994
rect 11622 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 12254 17176 12310 17232
rect 11886 15272 11942 15328
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11378 10906
rect 11378 10854 11408 10906
rect 11432 10854 11442 10906
rect 11442 10854 11488 10906
rect 11512 10854 11558 10906
rect 11558 10854 11568 10906
rect 11592 10854 11622 10906
rect 11622 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 10782 9016 10838 9072
rect 10230 4392 10286 4448
rect 10230 4120 10286 4176
rect 10322 3848 10378 3904
rect 11426 10512 11482 10568
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11378 9818
rect 11378 9766 11408 9818
rect 11432 9766 11442 9818
rect 11442 9766 11488 9818
rect 11512 9766 11558 9818
rect 11558 9766 11568 9818
rect 11592 9766 11622 9818
rect 11622 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 10966 8880 11022 8936
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11378 8730
rect 11378 8678 11408 8730
rect 11432 8678 11442 8730
rect 11442 8678 11488 8730
rect 11512 8678 11558 8730
rect 11558 8678 11568 8730
rect 11592 8678 11622 8730
rect 11622 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11378 7642
rect 11378 7590 11408 7642
rect 11432 7590 11442 7642
rect 11442 7590 11488 7642
rect 11512 7590 11558 7642
rect 11558 7590 11568 7642
rect 11592 7590 11622 7642
rect 11622 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 10414 3168 10470 3224
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11378 6554
rect 11378 6502 11408 6554
rect 11432 6502 11442 6554
rect 11442 6502 11488 6554
rect 11512 6502 11558 6554
rect 11558 6502 11568 6554
rect 11592 6502 11622 6554
rect 11622 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11610 6296 11666 6352
rect 11242 5616 11298 5672
rect 11794 9152 11850 9208
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11378 5466
rect 11378 5414 11408 5466
rect 11432 5414 11442 5466
rect 11442 5414 11488 5466
rect 11512 5414 11558 5466
rect 11558 5414 11568 5466
rect 11592 5414 11622 5466
rect 11622 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11058 5208 11114 5264
rect 11150 4392 11206 4448
rect 10966 3168 11022 3224
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11378 4378
rect 11378 4326 11408 4378
rect 11432 4326 11442 4378
rect 11442 4326 11488 4378
rect 11512 4326 11558 4378
rect 11558 4326 11568 4378
rect 11592 4326 11622 4378
rect 11622 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 12530 14456 12586 14512
rect 12438 13776 12494 13832
rect 12990 19080 13046 19136
rect 18050 20848 18106 20904
rect 18282 20698 18338 20700
rect 18362 20698 18418 20700
rect 18442 20698 18498 20700
rect 18522 20698 18578 20700
rect 18282 20646 18308 20698
rect 18308 20646 18338 20698
rect 18362 20646 18372 20698
rect 18372 20646 18418 20698
rect 18442 20646 18488 20698
rect 18488 20646 18498 20698
rect 18522 20646 18552 20698
rect 18552 20646 18578 20698
rect 18282 20644 18338 20646
rect 18362 20644 18418 20646
rect 18442 20644 18498 20646
rect 18522 20644 18578 20646
rect 14817 20154 14873 20156
rect 14897 20154 14953 20156
rect 14977 20154 15033 20156
rect 15057 20154 15113 20156
rect 14817 20102 14843 20154
rect 14843 20102 14873 20154
rect 14897 20102 14907 20154
rect 14907 20102 14953 20154
rect 14977 20102 15023 20154
rect 15023 20102 15033 20154
rect 15057 20102 15087 20154
rect 15087 20102 15113 20154
rect 14817 20100 14873 20102
rect 14897 20100 14953 20102
rect 14977 20100 15033 20102
rect 15057 20100 15113 20102
rect 14817 19066 14873 19068
rect 14897 19066 14953 19068
rect 14977 19066 15033 19068
rect 15057 19066 15113 19068
rect 14817 19014 14843 19066
rect 14843 19014 14873 19066
rect 14897 19014 14907 19066
rect 14907 19014 14953 19066
rect 14977 19014 15023 19066
rect 15023 19014 15033 19066
rect 15057 19014 15087 19066
rect 15087 19014 15113 19066
rect 14817 19012 14873 19014
rect 14897 19012 14953 19014
rect 14977 19012 15033 19014
rect 15057 19012 15113 19014
rect 12806 13776 12862 13832
rect 12346 12144 12402 12200
rect 12714 12688 12770 12744
rect 11978 7792 12034 7848
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11378 3290
rect 11378 3238 11408 3290
rect 11432 3238 11442 3290
rect 11442 3238 11488 3290
rect 11512 3238 11558 3290
rect 11558 3238 11568 3290
rect 11592 3238 11622 3290
rect 11622 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11378 2202
rect 11378 2150 11408 2202
rect 11432 2150 11442 2202
rect 11442 2150 11488 2202
rect 11512 2150 11558 2202
rect 11558 2150 11568 2202
rect 11592 2150 11622 2202
rect 11622 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 11794 3576 11850 3632
rect 11794 3304 11850 3360
rect 12162 9696 12218 9752
rect 12162 7268 12218 7304
rect 12162 7248 12164 7268
rect 12164 7248 12216 7268
rect 12216 7248 12218 7268
rect 12254 7112 12310 7168
rect 12162 6876 12164 6896
rect 12164 6876 12216 6896
rect 12216 6876 12218 6896
rect 12162 6840 12218 6876
rect 12162 6704 12218 6760
rect 12622 9832 12678 9888
rect 12530 7928 12586 7984
rect 12530 6876 12532 6896
rect 12532 6876 12584 6896
rect 12584 6876 12586 6896
rect 12530 6840 12586 6876
rect 12898 12688 12954 12744
rect 12806 11872 12862 11928
rect 12990 7792 13046 7848
rect 12990 4936 13046 4992
rect 13542 15272 13598 15328
rect 13450 12416 13506 12472
rect 13818 12588 13820 12608
rect 13820 12588 13872 12608
rect 13872 12588 13874 12608
rect 13818 12552 13874 12588
rect 13726 12416 13782 12472
rect 14817 17978 14873 17980
rect 14897 17978 14953 17980
rect 14977 17978 15033 17980
rect 15057 17978 15113 17980
rect 14817 17926 14843 17978
rect 14843 17926 14873 17978
rect 14897 17926 14907 17978
rect 14907 17926 14953 17978
rect 14977 17926 15023 17978
rect 15023 17926 15033 17978
rect 15057 17926 15087 17978
rect 15087 17926 15113 17978
rect 14817 17924 14873 17926
rect 14897 17924 14953 17926
rect 14977 17924 15033 17926
rect 15057 17924 15113 17926
rect 13634 8356 13690 8392
rect 13634 8336 13636 8356
rect 13636 8336 13688 8356
rect 13688 8336 13690 8356
rect 13450 4800 13506 4856
rect 13266 4664 13322 4720
rect 12898 4392 12954 4448
rect 13542 4664 13598 4720
rect 14002 10140 14004 10160
rect 14004 10140 14056 10160
rect 14056 10140 14058 10160
rect 14002 10104 14058 10140
rect 14817 16890 14873 16892
rect 14897 16890 14953 16892
rect 14977 16890 15033 16892
rect 15057 16890 15113 16892
rect 14817 16838 14843 16890
rect 14843 16838 14873 16890
rect 14897 16838 14907 16890
rect 14907 16838 14953 16890
rect 14977 16838 15023 16890
rect 15023 16838 15033 16890
rect 15057 16838 15087 16890
rect 15087 16838 15113 16890
rect 14817 16836 14873 16838
rect 14897 16836 14953 16838
rect 14977 16836 15033 16838
rect 15057 16836 15113 16838
rect 14817 15802 14873 15804
rect 14897 15802 14953 15804
rect 14977 15802 15033 15804
rect 15057 15802 15113 15804
rect 14817 15750 14843 15802
rect 14843 15750 14873 15802
rect 14897 15750 14907 15802
rect 14907 15750 14953 15802
rect 14977 15750 15023 15802
rect 15023 15750 15033 15802
rect 15057 15750 15087 15802
rect 15087 15750 15113 15802
rect 14817 15748 14873 15750
rect 14897 15748 14953 15750
rect 14977 15748 15033 15750
rect 15057 15748 15113 15750
rect 14817 14714 14873 14716
rect 14897 14714 14953 14716
rect 14977 14714 15033 14716
rect 15057 14714 15113 14716
rect 14817 14662 14843 14714
rect 14843 14662 14873 14714
rect 14897 14662 14907 14714
rect 14907 14662 14953 14714
rect 14977 14662 15023 14714
rect 15023 14662 15033 14714
rect 15057 14662 15087 14714
rect 15087 14662 15113 14714
rect 14817 14660 14873 14662
rect 14897 14660 14953 14662
rect 14977 14660 15033 14662
rect 15057 14660 15113 14662
rect 14817 13626 14873 13628
rect 14897 13626 14953 13628
rect 14977 13626 15033 13628
rect 15057 13626 15113 13628
rect 14817 13574 14843 13626
rect 14843 13574 14873 13626
rect 14897 13574 14907 13626
rect 14907 13574 14953 13626
rect 14977 13574 15023 13626
rect 15023 13574 15033 13626
rect 15057 13574 15087 13626
rect 15087 13574 15113 13626
rect 14817 13572 14873 13574
rect 14897 13572 14953 13574
rect 14977 13572 15033 13574
rect 15057 13572 15113 13574
rect 14817 12538 14873 12540
rect 14897 12538 14953 12540
rect 14977 12538 15033 12540
rect 15057 12538 15113 12540
rect 14817 12486 14843 12538
rect 14843 12486 14873 12538
rect 14897 12486 14907 12538
rect 14907 12486 14953 12538
rect 14977 12486 15023 12538
rect 15023 12486 15033 12538
rect 15057 12486 15087 12538
rect 15087 12486 15113 12538
rect 14817 12484 14873 12486
rect 14897 12484 14953 12486
rect 14977 12484 15033 12486
rect 15057 12484 15113 12486
rect 14817 11450 14873 11452
rect 14897 11450 14953 11452
rect 14977 11450 15033 11452
rect 15057 11450 15113 11452
rect 14817 11398 14843 11450
rect 14843 11398 14873 11450
rect 14897 11398 14907 11450
rect 14907 11398 14953 11450
rect 14977 11398 15023 11450
rect 15023 11398 15033 11450
rect 15057 11398 15087 11450
rect 15087 11398 15113 11450
rect 14817 11396 14873 11398
rect 14897 11396 14953 11398
rect 14977 11396 15033 11398
rect 15057 11396 15113 11398
rect 15198 11192 15254 11248
rect 14646 9696 14702 9752
rect 14370 9016 14426 9072
rect 13910 7112 13966 7168
rect 14094 3440 14150 3496
rect 14278 3984 14334 4040
rect 14278 3440 14334 3496
rect 14817 10362 14873 10364
rect 14897 10362 14953 10364
rect 14977 10362 15033 10364
rect 15057 10362 15113 10364
rect 14817 10310 14843 10362
rect 14843 10310 14873 10362
rect 14897 10310 14907 10362
rect 14907 10310 14953 10362
rect 14977 10310 15023 10362
rect 15023 10310 15033 10362
rect 15057 10310 15087 10362
rect 15087 10310 15113 10362
rect 14817 10308 14873 10310
rect 14897 10308 14953 10310
rect 14977 10308 15033 10310
rect 15057 10308 15113 10310
rect 15106 9968 15162 10024
rect 14817 9274 14873 9276
rect 14897 9274 14953 9276
rect 14977 9274 15033 9276
rect 15057 9274 15113 9276
rect 14817 9222 14843 9274
rect 14843 9222 14873 9274
rect 14897 9222 14907 9274
rect 14907 9222 14953 9274
rect 14977 9222 15023 9274
rect 15023 9222 15033 9274
rect 15057 9222 15087 9274
rect 15087 9222 15113 9274
rect 14817 9220 14873 9222
rect 14897 9220 14953 9222
rect 14977 9220 15033 9222
rect 15057 9220 15113 9222
rect 14646 8472 14702 8528
rect 14554 4120 14610 4176
rect 14817 8186 14873 8188
rect 14897 8186 14953 8188
rect 14977 8186 15033 8188
rect 15057 8186 15113 8188
rect 14817 8134 14843 8186
rect 14843 8134 14873 8186
rect 14897 8134 14907 8186
rect 14907 8134 14953 8186
rect 14977 8134 15023 8186
rect 15023 8134 15033 8186
rect 15057 8134 15087 8186
rect 15087 8134 15113 8186
rect 14817 8132 14873 8134
rect 14897 8132 14953 8134
rect 14977 8132 15033 8134
rect 15057 8132 15113 8134
rect 14817 7098 14873 7100
rect 14897 7098 14953 7100
rect 14977 7098 15033 7100
rect 15057 7098 15113 7100
rect 14817 7046 14843 7098
rect 14843 7046 14873 7098
rect 14897 7046 14907 7098
rect 14907 7046 14953 7098
rect 14977 7046 15023 7098
rect 15023 7046 15033 7098
rect 15057 7046 15087 7098
rect 15087 7046 15113 7098
rect 14817 7044 14873 7046
rect 14897 7044 14953 7046
rect 14977 7044 15033 7046
rect 15057 7044 15113 7046
rect 14817 6010 14873 6012
rect 14897 6010 14953 6012
rect 14977 6010 15033 6012
rect 15057 6010 15113 6012
rect 14817 5958 14843 6010
rect 14843 5958 14873 6010
rect 14897 5958 14907 6010
rect 14907 5958 14953 6010
rect 14977 5958 15023 6010
rect 15023 5958 15033 6010
rect 15057 5958 15087 6010
rect 15087 5958 15113 6010
rect 14817 5956 14873 5958
rect 14897 5956 14953 5958
rect 14977 5956 15033 5958
rect 15057 5956 15113 5958
rect 14817 4922 14873 4924
rect 14897 4922 14953 4924
rect 14977 4922 15033 4924
rect 15057 4922 15113 4924
rect 14817 4870 14843 4922
rect 14843 4870 14873 4922
rect 14897 4870 14907 4922
rect 14907 4870 14953 4922
rect 14977 4870 15023 4922
rect 15023 4870 15033 4922
rect 15057 4870 15087 4922
rect 15087 4870 15113 4922
rect 14817 4868 14873 4870
rect 14897 4868 14953 4870
rect 14977 4868 15033 4870
rect 15057 4868 15113 4870
rect 14817 3834 14873 3836
rect 14897 3834 14953 3836
rect 14977 3834 15033 3836
rect 15057 3834 15113 3836
rect 14817 3782 14843 3834
rect 14843 3782 14873 3834
rect 14897 3782 14907 3834
rect 14907 3782 14953 3834
rect 14977 3782 15023 3834
rect 15023 3782 15033 3834
rect 15057 3782 15087 3834
rect 15087 3782 15113 3834
rect 14817 3780 14873 3782
rect 14897 3780 14953 3782
rect 14977 3780 15033 3782
rect 15057 3780 15113 3782
rect 14817 2746 14873 2748
rect 14897 2746 14953 2748
rect 14977 2746 15033 2748
rect 15057 2746 15113 2748
rect 14817 2694 14843 2746
rect 14843 2694 14873 2746
rect 14897 2694 14907 2746
rect 14907 2694 14953 2746
rect 14977 2694 15023 2746
rect 15023 2694 15033 2746
rect 15057 2694 15087 2746
rect 15087 2694 15113 2746
rect 14817 2692 14873 2694
rect 14897 2692 14953 2694
rect 14977 2692 15033 2694
rect 15057 2692 15113 2694
rect 15934 16668 15936 16688
rect 15936 16668 15988 16688
rect 15988 16668 15990 16688
rect 15934 16632 15990 16668
rect 15750 4664 15806 4720
rect 16026 7520 16082 7576
rect 15290 2352 15346 2408
rect 16026 3712 16082 3768
rect 17958 20304 18014 20360
rect 17958 19896 18014 19952
rect 17774 18944 17830 19000
rect 18282 19610 18338 19612
rect 18362 19610 18418 19612
rect 18442 19610 18498 19612
rect 18522 19610 18578 19612
rect 18282 19558 18308 19610
rect 18308 19558 18338 19610
rect 18362 19558 18372 19610
rect 18372 19558 18418 19610
rect 18442 19558 18488 19610
rect 18488 19558 18498 19610
rect 18522 19558 18552 19610
rect 18552 19558 18578 19610
rect 18282 19556 18338 19558
rect 18362 19556 18418 19558
rect 18442 19556 18498 19558
rect 18522 19556 18578 19558
rect 18050 19216 18106 19272
rect 18694 19352 18750 19408
rect 18050 18400 18106 18456
rect 17222 15952 17278 16008
rect 17222 13368 17278 13424
rect 16210 7520 16266 7576
rect 16946 11620 17002 11656
rect 16946 11600 16948 11620
rect 16948 11600 17000 11620
rect 17000 11600 17002 11620
rect 17314 12144 17370 12200
rect 16670 8880 16726 8936
rect 17038 7248 17094 7304
rect 18050 17992 18106 18048
rect 18282 18522 18338 18524
rect 18362 18522 18418 18524
rect 18442 18522 18498 18524
rect 18522 18522 18578 18524
rect 18282 18470 18308 18522
rect 18308 18470 18338 18522
rect 18362 18470 18372 18522
rect 18372 18470 18418 18522
rect 18442 18470 18488 18522
rect 18488 18470 18498 18522
rect 18522 18470 18552 18522
rect 18552 18470 18578 18522
rect 18282 18468 18338 18470
rect 18362 18468 18418 18470
rect 18442 18468 18498 18470
rect 18522 18468 18578 18470
rect 18234 18264 18290 18320
rect 18602 17992 18658 18048
rect 18510 17856 18566 17912
rect 19154 22208 19210 22264
rect 19246 21256 19302 21312
rect 18282 17434 18338 17436
rect 18362 17434 18418 17436
rect 18442 17434 18498 17436
rect 18522 17434 18578 17436
rect 18282 17382 18308 17434
rect 18308 17382 18338 17434
rect 18362 17382 18372 17434
rect 18372 17382 18418 17434
rect 18442 17382 18488 17434
rect 18488 17382 18498 17434
rect 18522 17382 18552 17434
rect 18552 17382 18578 17434
rect 18282 17380 18338 17382
rect 18362 17380 18418 17382
rect 18442 17380 18498 17382
rect 18522 17380 18578 17382
rect 18282 16346 18338 16348
rect 18362 16346 18418 16348
rect 18442 16346 18498 16348
rect 18522 16346 18578 16348
rect 18282 16294 18308 16346
rect 18308 16294 18338 16346
rect 18362 16294 18372 16346
rect 18372 16294 18418 16346
rect 18442 16294 18488 16346
rect 18488 16294 18498 16346
rect 18522 16294 18552 16346
rect 18552 16294 18578 16346
rect 18282 16292 18338 16294
rect 18362 16292 18418 16294
rect 18442 16292 18498 16294
rect 18522 16292 18578 16294
rect 18694 16224 18750 16280
rect 18050 15564 18106 15600
rect 18050 15544 18052 15564
rect 18052 15544 18104 15564
rect 18104 15544 18106 15564
rect 18326 15428 18382 15464
rect 18326 15408 18328 15428
rect 18328 15408 18380 15428
rect 18380 15408 18382 15428
rect 18282 15258 18338 15260
rect 18362 15258 18418 15260
rect 18442 15258 18498 15260
rect 18522 15258 18578 15260
rect 18282 15206 18308 15258
rect 18308 15206 18338 15258
rect 18362 15206 18372 15258
rect 18372 15206 18418 15258
rect 18442 15206 18488 15258
rect 18488 15206 18498 15258
rect 18522 15206 18552 15258
rect 18552 15206 18578 15258
rect 18282 15204 18338 15206
rect 18362 15204 18418 15206
rect 18442 15204 18498 15206
rect 18522 15204 18578 15206
rect 18602 14320 18658 14376
rect 18282 14170 18338 14172
rect 18362 14170 18418 14172
rect 18442 14170 18498 14172
rect 18522 14170 18578 14172
rect 18282 14118 18308 14170
rect 18308 14118 18338 14170
rect 18362 14118 18372 14170
rect 18372 14118 18418 14170
rect 18442 14118 18488 14170
rect 18488 14118 18498 14170
rect 18522 14118 18552 14170
rect 18552 14118 18578 14170
rect 18282 14116 18338 14118
rect 18362 14116 18418 14118
rect 18442 14116 18498 14118
rect 18522 14116 18578 14118
rect 18602 13912 18658 13968
rect 18970 16632 19026 16688
rect 20166 21664 20222 21720
rect 18878 16088 18934 16144
rect 18878 14456 18934 14512
rect 17314 6704 17370 6760
rect 17314 2896 17370 2952
rect 18282 13082 18338 13084
rect 18362 13082 18418 13084
rect 18442 13082 18498 13084
rect 18522 13082 18578 13084
rect 18282 13030 18308 13082
rect 18308 13030 18338 13082
rect 18362 13030 18372 13082
rect 18372 13030 18418 13082
rect 18442 13030 18488 13082
rect 18488 13030 18498 13082
rect 18522 13030 18552 13082
rect 18552 13030 18578 13082
rect 18282 13028 18338 13030
rect 18362 13028 18418 13030
rect 18442 13028 18498 13030
rect 18522 13028 18578 13030
rect 18050 12552 18106 12608
rect 18282 11994 18338 11996
rect 18362 11994 18418 11996
rect 18442 11994 18498 11996
rect 18522 11994 18578 11996
rect 18282 11942 18308 11994
rect 18308 11942 18338 11994
rect 18362 11942 18372 11994
rect 18372 11942 18418 11994
rect 18442 11942 18488 11994
rect 18488 11942 18498 11994
rect 18522 11942 18552 11994
rect 18552 11942 18578 11994
rect 18282 11940 18338 11942
rect 18362 11940 18418 11942
rect 18442 11940 18498 11942
rect 18522 11940 18578 11942
rect 18142 11348 18198 11384
rect 18142 11328 18144 11348
rect 18144 11328 18196 11348
rect 18196 11328 18198 11348
rect 17866 10240 17922 10296
rect 18282 10906 18338 10908
rect 18362 10906 18418 10908
rect 18442 10906 18498 10908
rect 18522 10906 18578 10908
rect 18282 10854 18308 10906
rect 18308 10854 18338 10906
rect 18362 10854 18372 10906
rect 18372 10854 18418 10906
rect 18442 10854 18488 10906
rect 18488 10854 18498 10906
rect 18522 10854 18552 10906
rect 18552 10854 18578 10906
rect 18282 10852 18338 10854
rect 18362 10852 18418 10854
rect 18442 10852 18498 10854
rect 18522 10852 18578 10854
rect 18050 10104 18106 10160
rect 17958 9988 18014 10024
rect 17958 9968 17960 9988
rect 17960 9968 18012 9988
rect 18012 9968 18014 9988
rect 17774 8472 17830 8528
rect 18282 9818 18338 9820
rect 18362 9818 18418 9820
rect 18442 9818 18498 9820
rect 18522 9818 18578 9820
rect 18282 9766 18308 9818
rect 18308 9766 18338 9818
rect 18362 9766 18372 9818
rect 18372 9766 18418 9818
rect 18442 9766 18488 9818
rect 18488 9766 18498 9818
rect 18522 9766 18552 9818
rect 18552 9766 18578 9818
rect 18282 9764 18338 9766
rect 18362 9764 18418 9766
rect 18442 9764 18498 9766
rect 18522 9764 18578 9766
rect 18510 9560 18566 9616
rect 18234 9424 18290 9480
rect 18050 9288 18106 9344
rect 18142 9016 18198 9072
rect 18142 8880 18198 8936
rect 18282 8730 18338 8732
rect 18362 8730 18418 8732
rect 18442 8730 18498 8732
rect 18522 8730 18578 8732
rect 18282 8678 18308 8730
rect 18308 8678 18338 8730
rect 18362 8678 18372 8730
rect 18372 8678 18418 8730
rect 18442 8678 18488 8730
rect 18488 8678 18498 8730
rect 18522 8678 18552 8730
rect 18552 8678 18578 8730
rect 18282 8676 18338 8678
rect 18362 8676 18418 8678
rect 18442 8676 18498 8678
rect 18522 8676 18578 8678
rect 18282 7642 18338 7644
rect 18362 7642 18418 7644
rect 18442 7642 18498 7644
rect 18522 7642 18578 7644
rect 18282 7590 18308 7642
rect 18308 7590 18338 7642
rect 18362 7590 18372 7642
rect 18372 7590 18418 7642
rect 18442 7590 18488 7642
rect 18488 7590 18498 7642
rect 18522 7590 18552 7642
rect 18552 7590 18578 7642
rect 18282 7588 18338 7590
rect 18362 7588 18418 7590
rect 18442 7588 18498 7590
rect 18522 7588 18578 7590
rect 17958 6976 18014 7032
rect 17958 6024 18014 6080
rect 17774 2896 17830 2952
rect 17682 1944 17738 2000
rect 17958 3304 18014 3360
rect 18282 6554 18338 6556
rect 18362 6554 18418 6556
rect 18442 6554 18498 6556
rect 18522 6554 18578 6556
rect 18282 6502 18308 6554
rect 18308 6502 18338 6554
rect 18362 6502 18372 6554
rect 18372 6502 18418 6554
rect 18442 6502 18488 6554
rect 18488 6502 18498 6554
rect 18522 6502 18552 6554
rect 18552 6502 18578 6554
rect 18282 6500 18338 6502
rect 18362 6500 18418 6502
rect 18442 6500 18498 6502
rect 18522 6500 18578 6502
rect 18282 5466 18338 5468
rect 18362 5466 18418 5468
rect 18442 5466 18498 5468
rect 18522 5466 18578 5468
rect 18282 5414 18308 5466
rect 18308 5414 18338 5466
rect 18362 5414 18372 5466
rect 18372 5414 18418 5466
rect 18442 5414 18488 5466
rect 18488 5414 18498 5466
rect 18522 5414 18552 5466
rect 18552 5414 18578 5466
rect 18282 5412 18338 5414
rect 18362 5412 18418 5414
rect 18442 5412 18498 5414
rect 18522 5412 18578 5414
rect 18282 4378 18338 4380
rect 18362 4378 18418 4380
rect 18442 4378 18498 4380
rect 18522 4378 18578 4380
rect 18282 4326 18308 4378
rect 18308 4326 18338 4378
rect 18362 4326 18372 4378
rect 18372 4326 18418 4378
rect 18442 4326 18488 4378
rect 18488 4326 18498 4378
rect 18522 4326 18552 4378
rect 18552 4326 18578 4378
rect 18282 4324 18338 4326
rect 18362 4324 18418 4326
rect 18442 4324 18498 4326
rect 18522 4324 18578 4326
rect 18282 3290 18338 3292
rect 18362 3290 18418 3292
rect 18442 3290 18498 3292
rect 18522 3290 18578 3292
rect 18282 3238 18308 3290
rect 18308 3238 18338 3290
rect 18362 3238 18372 3290
rect 18372 3238 18418 3290
rect 18442 3238 18488 3290
rect 18488 3238 18498 3290
rect 18522 3238 18552 3290
rect 18552 3238 18578 3290
rect 18282 3236 18338 3238
rect 18362 3236 18418 3238
rect 18442 3236 18498 3238
rect 18522 3236 18578 3238
rect 18282 2202 18338 2204
rect 18362 2202 18418 2204
rect 18442 2202 18498 2204
rect 18522 2202 18578 2204
rect 18282 2150 18308 2202
rect 18308 2150 18338 2202
rect 18362 2150 18372 2202
rect 18372 2150 18418 2202
rect 18442 2150 18488 2202
rect 18488 2150 18498 2202
rect 18522 2150 18552 2202
rect 18552 2150 18578 2202
rect 18282 2148 18338 2150
rect 18362 2148 18418 2150
rect 18442 2148 18498 2150
rect 18522 2148 18578 2150
rect 18878 10648 18934 10704
rect 18786 10512 18842 10568
rect 18786 9016 18842 9072
rect 19246 10648 19302 10704
rect 19154 9288 19210 9344
rect 18878 8064 18934 8120
rect 18786 7540 18842 7576
rect 18786 7520 18788 7540
rect 18788 7520 18840 7540
rect 18840 7520 18842 7540
rect 18602 1536 18658 1592
rect 19062 3168 19118 3224
rect 18786 992 18842 1048
rect 19890 15700 19946 15736
rect 19890 15680 19892 15700
rect 19892 15680 19944 15700
rect 19944 15680 19946 15700
rect 19982 14864 20038 14920
rect 19890 12960 19946 13016
rect 19430 5208 19486 5264
rect 19614 5072 19670 5128
rect 19798 3576 19854 3632
rect 20074 3440 20130 3496
rect 20258 3984 20314 4040
rect 20074 584 20130 640
rect 20718 17584 20774 17640
rect 20718 15272 20774 15328
rect 20718 13504 20774 13560
rect 20534 4256 20590 4312
rect 20534 3848 20590 3904
rect 20350 3712 20406 3768
rect 19246 176 19302 232
<< metal3 >>
rect 0 22674 480 22704
rect 3877 22674 3943 22677
rect 0 22672 3943 22674
rect 0 22616 3882 22672
rect 3938 22616 3943 22672
rect 0 22614 3943 22616
rect 0 22584 480 22614
rect 3877 22611 3943 22614
rect 18965 22674 19031 22677
rect 22520 22674 23000 22704
rect 18965 22672 23000 22674
rect 18965 22616 18970 22672
rect 19026 22616 23000 22672
rect 18965 22614 23000 22616
rect 18965 22611 19031 22614
rect 22520 22584 23000 22614
rect 0 22266 480 22296
rect 3509 22266 3575 22269
rect 0 22264 3575 22266
rect 0 22208 3514 22264
rect 3570 22208 3575 22264
rect 0 22206 3575 22208
rect 0 22176 480 22206
rect 3509 22203 3575 22206
rect 19149 22266 19215 22269
rect 22520 22266 23000 22296
rect 19149 22264 23000 22266
rect 19149 22208 19154 22264
rect 19210 22208 23000 22264
rect 19149 22206 23000 22208
rect 19149 22203 19215 22206
rect 22520 22176 23000 22206
rect 0 21858 480 21888
rect 4245 21858 4311 21861
rect 0 21856 4311 21858
rect 0 21800 4250 21856
rect 4306 21800 4311 21856
rect 0 21798 4311 21800
rect 0 21768 480 21798
rect 4245 21795 4311 21798
rect 20161 21722 20227 21725
rect 22520 21722 23000 21752
rect 20161 21720 23000 21722
rect 20161 21664 20166 21720
rect 20222 21664 23000 21720
rect 20161 21662 23000 21664
rect 20161 21659 20227 21662
rect 22520 21632 23000 21662
rect 0 21314 480 21344
rect 3141 21314 3207 21317
rect 0 21312 3207 21314
rect 0 21256 3146 21312
rect 3202 21256 3207 21312
rect 0 21254 3207 21256
rect 0 21224 480 21254
rect 3141 21251 3207 21254
rect 19241 21314 19307 21317
rect 22520 21314 23000 21344
rect 19241 21312 23000 21314
rect 19241 21256 19246 21312
rect 19302 21256 23000 21312
rect 19241 21254 23000 21256
rect 19241 21251 19307 21254
rect 22520 21224 23000 21254
rect 0 20906 480 20936
rect 4061 20906 4127 20909
rect 0 20904 4127 20906
rect 0 20848 4066 20904
rect 4122 20848 4127 20904
rect 0 20846 4127 20848
rect 0 20816 480 20846
rect 4061 20843 4127 20846
rect 18045 20906 18111 20909
rect 22520 20906 23000 20936
rect 18045 20904 23000 20906
rect 18045 20848 18050 20904
rect 18106 20848 23000 20904
rect 18045 20846 23000 20848
rect 18045 20843 18111 20846
rect 22520 20816 23000 20846
rect 4409 20704 4729 20705
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 20639 4729 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 18270 20704 18590 20705
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 18270 20639 18590 20640
rect 0 20498 480 20528
rect 3969 20498 4035 20501
rect 0 20496 4035 20498
rect 0 20440 3974 20496
rect 4030 20440 4035 20496
rect 0 20438 4035 20440
rect 0 20408 480 20438
rect 3969 20435 4035 20438
rect 17953 20362 18019 20365
rect 22520 20362 23000 20392
rect 17953 20360 23000 20362
rect 17953 20304 17958 20360
rect 18014 20304 23000 20360
rect 17953 20302 23000 20304
rect 17953 20299 18019 20302
rect 22520 20272 23000 20302
rect 7874 20160 8194 20161
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8194 20160
rect 7874 20095 8194 20096
rect 14805 20160 15125 20161
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 20095 15125 20096
rect 0 19954 480 19984
rect 4061 19954 4127 19957
rect 0 19952 4127 19954
rect 0 19896 4066 19952
rect 4122 19896 4127 19952
rect 0 19894 4127 19896
rect 0 19864 480 19894
rect 4061 19891 4127 19894
rect 17953 19954 18019 19957
rect 22520 19954 23000 19984
rect 17953 19952 23000 19954
rect 17953 19896 17958 19952
rect 18014 19896 23000 19952
rect 17953 19894 23000 19896
rect 17953 19891 18019 19894
rect 22520 19864 23000 19894
rect 4409 19616 4729 19617
rect 0 19546 480 19576
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 19551 4729 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 18270 19616 18590 19617
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 19551 18590 19552
rect 3325 19546 3391 19549
rect 0 19544 3391 19546
rect 0 19488 3330 19544
rect 3386 19488 3391 19544
rect 0 19486 3391 19488
rect 0 19456 480 19486
rect 3325 19483 3391 19486
rect 18689 19410 18755 19413
rect 22520 19410 23000 19440
rect 18689 19408 23000 19410
rect 18689 19352 18694 19408
rect 18750 19352 23000 19408
rect 18689 19350 23000 19352
rect 18689 19347 18755 19350
rect 22520 19320 23000 19350
rect 18045 19274 18111 19277
rect 18822 19274 18828 19276
rect 18045 19272 18828 19274
rect 18045 19216 18050 19272
rect 18106 19216 18828 19272
rect 18045 19214 18828 19216
rect 18045 19211 18111 19214
rect 18822 19212 18828 19214
rect 18892 19212 18898 19276
rect 0 19138 480 19168
rect 4061 19138 4127 19141
rect 0 19136 4127 19138
rect 0 19080 4066 19136
rect 4122 19080 4127 19136
rect 0 19078 4127 19080
rect 0 19048 480 19078
rect 4061 19075 4127 19078
rect 10225 19138 10291 19141
rect 12985 19138 13051 19141
rect 10225 19136 13051 19138
rect 10225 19080 10230 19136
rect 10286 19080 12990 19136
rect 13046 19080 13051 19136
rect 10225 19078 13051 19080
rect 10225 19075 10291 19078
rect 12985 19075 13051 19078
rect 7874 19072 8194 19073
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8194 19072
rect 7874 19007 8194 19008
rect 14805 19072 15125 19073
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 19007 15125 19008
rect 17769 19002 17835 19005
rect 22520 19002 23000 19032
rect 17769 19000 23000 19002
rect 17769 18944 17774 19000
rect 17830 18944 23000 19000
rect 17769 18942 23000 18944
rect 17769 18939 17835 18942
rect 22520 18912 23000 18942
rect 0 18594 480 18624
rect 2865 18594 2931 18597
rect 22520 18594 23000 18624
rect 0 18592 2931 18594
rect 0 18536 2870 18592
rect 2926 18536 2931 18592
rect 0 18534 2931 18536
rect 0 18504 480 18534
rect 2865 18531 2931 18534
rect 19014 18534 23000 18594
rect 4409 18528 4729 18529
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 18463 4729 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 18270 18528 18590 18529
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18270 18463 18590 18464
rect 18045 18460 18111 18461
rect 18045 18458 18092 18460
rect 18000 18456 18092 18458
rect 18000 18400 18050 18456
rect 18000 18398 18092 18400
rect 18045 18396 18092 18398
rect 18156 18396 18162 18460
rect 18045 18395 18111 18396
rect 18229 18322 18295 18325
rect 19014 18322 19074 18534
rect 22520 18504 23000 18534
rect 18229 18320 19074 18322
rect 18229 18264 18234 18320
rect 18290 18264 19074 18320
rect 18229 18262 19074 18264
rect 18229 18259 18295 18262
rect 0 18186 480 18216
rect 3049 18186 3115 18189
rect 0 18184 3115 18186
rect 0 18128 3054 18184
rect 3110 18128 3115 18184
rect 0 18126 3115 18128
rect 0 18096 480 18126
rect 3049 18123 3115 18126
rect 17902 17988 17908 18052
rect 17972 18050 17978 18052
rect 18045 18050 18111 18053
rect 17972 18048 18111 18050
rect 17972 17992 18050 18048
rect 18106 17992 18111 18048
rect 17972 17990 18111 17992
rect 17972 17988 17978 17990
rect 18045 17987 18111 17990
rect 18597 18050 18663 18053
rect 22520 18050 23000 18080
rect 18597 18048 23000 18050
rect 18597 17992 18602 18048
rect 18658 17992 23000 18048
rect 18597 17990 23000 17992
rect 18597 17987 18663 17990
rect 7874 17984 8194 17985
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8194 17984
rect 7874 17919 8194 17920
rect 14805 17984 15125 17985
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 22520 17960 23000 17990
rect 14805 17919 15125 17920
rect 17534 17852 17540 17916
rect 17604 17914 17610 17916
rect 18505 17914 18571 17917
rect 17604 17912 18571 17914
rect 17604 17856 18510 17912
rect 18566 17856 18571 17912
rect 17604 17854 18571 17856
rect 17604 17852 17610 17854
rect 18505 17851 18571 17854
rect 0 17778 480 17808
rect 1945 17778 2011 17781
rect 0 17776 2011 17778
rect 0 17720 1950 17776
rect 2006 17720 2011 17776
rect 0 17718 2011 17720
rect 0 17688 480 17718
rect 1945 17715 2011 17718
rect 20713 17642 20779 17645
rect 22520 17642 23000 17672
rect 20713 17640 23000 17642
rect 20713 17584 20718 17640
rect 20774 17584 23000 17640
rect 20713 17582 23000 17584
rect 20713 17579 20779 17582
rect 22520 17552 23000 17582
rect 4409 17440 4729 17441
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 17375 4729 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 18270 17440 18590 17441
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 18270 17375 18590 17376
rect 0 17234 480 17264
rect 4153 17234 4219 17237
rect 0 17232 4219 17234
rect 0 17176 4158 17232
rect 4214 17176 4219 17232
rect 0 17174 4219 17176
rect 0 17144 480 17174
rect 4153 17171 4219 17174
rect 12249 17234 12315 17237
rect 22520 17234 23000 17264
rect 12249 17232 23000 17234
rect 12249 17176 12254 17232
rect 12310 17176 23000 17232
rect 12249 17174 23000 17176
rect 12249 17171 12315 17174
rect 22520 17144 23000 17174
rect 7874 16896 8194 16897
rect 0 16826 480 16856
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8194 16896
rect 7874 16831 8194 16832
rect 14805 16896 15125 16897
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 16831 15125 16832
rect 2957 16826 3023 16829
rect 0 16824 3023 16826
rect 0 16768 2962 16824
rect 3018 16768 3023 16824
rect 0 16766 3023 16768
rect 0 16736 480 16766
rect 2957 16763 3023 16766
rect 15929 16690 15995 16693
rect 18822 16690 18828 16692
rect 15929 16688 18828 16690
rect 15929 16632 15934 16688
rect 15990 16632 18828 16688
rect 15929 16630 18828 16632
rect 15929 16627 15995 16630
rect 18822 16628 18828 16630
rect 18892 16628 18898 16692
rect 18965 16690 19031 16693
rect 22520 16690 23000 16720
rect 18965 16688 23000 16690
rect 18965 16632 18970 16688
rect 19026 16632 23000 16688
rect 18965 16630 23000 16632
rect 18965 16627 19031 16630
rect 22520 16600 23000 16630
rect 0 16418 480 16448
rect 2681 16418 2747 16421
rect 0 16416 2747 16418
rect 0 16360 2686 16416
rect 2742 16360 2747 16416
rect 0 16358 2747 16360
rect 0 16328 480 16358
rect 2681 16355 2747 16358
rect 4409 16352 4729 16353
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 16287 4729 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 18270 16352 18590 16353
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 16287 18590 16288
rect 18689 16282 18755 16285
rect 22520 16282 23000 16312
rect 18689 16280 23000 16282
rect 18689 16224 18694 16280
rect 18750 16224 23000 16280
rect 18689 16222 23000 16224
rect 18689 16219 18755 16222
rect 22520 16192 23000 16222
rect 9857 16146 9923 16149
rect 18873 16146 18939 16149
rect 9857 16144 18939 16146
rect 9857 16088 9862 16144
rect 9918 16088 18878 16144
rect 18934 16088 18939 16144
rect 9857 16086 18939 16088
rect 9857 16083 9923 16086
rect 18873 16083 18939 16086
rect 11513 16010 11579 16013
rect 17217 16010 17283 16013
rect 11513 16008 17283 16010
rect 11513 15952 11518 16008
rect 11574 15952 17222 16008
rect 17278 15952 17283 16008
rect 11513 15950 17283 15952
rect 11513 15947 11579 15950
rect 17217 15947 17283 15950
rect 0 15874 480 15904
rect 3325 15874 3391 15877
rect 0 15872 3391 15874
rect 0 15816 3330 15872
rect 3386 15816 3391 15872
rect 0 15814 3391 15816
rect 0 15784 480 15814
rect 3325 15811 3391 15814
rect 7874 15808 8194 15809
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8194 15808
rect 7874 15743 8194 15744
rect 14805 15808 15125 15809
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 15743 15125 15744
rect 19885 15738 19951 15741
rect 22520 15738 23000 15768
rect 19885 15736 23000 15738
rect 19885 15680 19890 15736
rect 19946 15680 23000 15736
rect 19885 15678 23000 15680
rect 19885 15675 19951 15678
rect 22520 15648 23000 15678
rect 6821 15602 6887 15605
rect 18045 15602 18111 15605
rect 6821 15600 18111 15602
rect 6821 15544 6826 15600
rect 6882 15544 18050 15600
rect 18106 15544 18111 15600
rect 6821 15542 18111 15544
rect 6821 15539 6887 15542
rect 18045 15539 18111 15542
rect 0 15466 480 15496
rect 3509 15466 3575 15469
rect 0 15464 3575 15466
rect 0 15408 3514 15464
rect 3570 15408 3575 15464
rect 0 15406 3575 15408
rect 0 15376 480 15406
rect 3509 15403 3575 15406
rect 10961 15466 11027 15469
rect 18321 15466 18387 15469
rect 10961 15464 18387 15466
rect 10961 15408 10966 15464
rect 11022 15408 18326 15464
rect 18382 15408 18387 15464
rect 10961 15406 18387 15408
rect 10961 15403 11027 15406
rect 18321 15403 18387 15406
rect 11881 15330 11947 15333
rect 13537 15330 13603 15333
rect 11881 15328 13603 15330
rect 11881 15272 11886 15328
rect 11942 15272 13542 15328
rect 13598 15272 13603 15328
rect 11881 15270 13603 15272
rect 11881 15267 11947 15270
rect 13537 15267 13603 15270
rect 20713 15330 20779 15333
rect 22520 15330 23000 15360
rect 20713 15328 23000 15330
rect 20713 15272 20718 15328
rect 20774 15272 23000 15328
rect 20713 15270 23000 15272
rect 20713 15267 20779 15270
rect 4409 15264 4729 15265
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 15199 4729 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 18270 15264 18590 15265
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 22520 15240 23000 15270
rect 18270 15199 18590 15200
rect 0 15058 480 15088
rect 1025 15058 1091 15061
rect 0 15056 1091 15058
rect 0 15000 1030 15056
rect 1086 15000 1091 15056
rect 0 14998 1091 15000
rect 0 14968 480 14998
rect 1025 14995 1091 14998
rect 19977 14922 20043 14925
rect 22520 14922 23000 14952
rect 19977 14920 23000 14922
rect 19977 14864 19982 14920
rect 20038 14864 23000 14920
rect 19977 14862 23000 14864
rect 19977 14859 20043 14862
rect 22520 14832 23000 14862
rect 7874 14720 8194 14721
rect 0 14650 480 14680
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8194 14720
rect 7874 14655 8194 14656
rect 14805 14720 15125 14721
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 14655 15125 14656
rect 1669 14650 1735 14653
rect 0 14648 1735 14650
rect 0 14592 1674 14648
rect 1730 14592 1735 14648
rect 0 14590 1735 14592
rect 0 14560 480 14590
rect 1669 14587 1735 14590
rect 12525 14514 12591 14517
rect 18873 14514 18939 14517
rect 12525 14512 18939 14514
rect 12525 14456 12530 14512
rect 12586 14456 18878 14512
rect 18934 14456 18939 14512
rect 12525 14454 18939 14456
rect 12525 14451 12591 14454
rect 18873 14451 18939 14454
rect 18597 14378 18663 14381
rect 22520 14378 23000 14408
rect 18597 14376 23000 14378
rect 18597 14320 18602 14376
rect 18658 14320 23000 14376
rect 18597 14318 23000 14320
rect 18597 14315 18663 14318
rect 22520 14288 23000 14318
rect 4409 14176 4729 14177
rect 0 14106 480 14136
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 14111 4729 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 18270 14176 18590 14177
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 18270 14111 18590 14112
rect 3141 14106 3207 14109
rect 0 14104 3207 14106
rect 0 14048 3146 14104
rect 3202 14048 3207 14104
rect 0 14046 3207 14048
rect 0 14016 480 14046
rect 3141 14043 3207 14046
rect 4429 13970 4495 13973
rect 8753 13970 8819 13973
rect 4429 13968 8819 13970
rect 4429 13912 4434 13968
rect 4490 13912 8758 13968
rect 8814 13912 8819 13968
rect 4429 13910 8819 13912
rect 4429 13907 4495 13910
rect 8753 13907 8819 13910
rect 18597 13970 18663 13973
rect 22520 13970 23000 14000
rect 18597 13968 23000 13970
rect 18597 13912 18602 13968
rect 18658 13912 23000 13968
rect 18597 13910 23000 13912
rect 18597 13907 18663 13910
rect 22520 13880 23000 13910
rect 12433 13834 12499 13837
rect 12801 13834 12867 13837
rect 12433 13832 12867 13834
rect 12433 13776 12438 13832
rect 12494 13776 12806 13832
rect 12862 13776 12867 13832
rect 12433 13774 12867 13776
rect 12433 13771 12499 13774
rect 12801 13771 12867 13774
rect 0 13698 480 13728
rect 2773 13698 2839 13701
rect 0 13696 2839 13698
rect 0 13640 2778 13696
rect 2834 13640 2839 13696
rect 0 13638 2839 13640
rect 0 13608 480 13638
rect 2773 13635 2839 13638
rect 7874 13632 8194 13633
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8194 13632
rect 7874 13567 8194 13568
rect 14805 13632 15125 13633
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 13567 15125 13568
rect 3969 13562 4035 13565
rect 4245 13562 4311 13565
rect 3969 13560 4311 13562
rect 3969 13504 3974 13560
rect 4030 13504 4250 13560
rect 4306 13504 4311 13560
rect 3969 13502 4311 13504
rect 3969 13499 4035 13502
rect 4245 13499 4311 13502
rect 20713 13562 20779 13565
rect 22520 13562 23000 13592
rect 20713 13560 23000 13562
rect 20713 13504 20718 13560
rect 20774 13504 23000 13560
rect 20713 13502 23000 13504
rect 20713 13499 20779 13502
rect 22520 13472 23000 13502
rect 17217 13426 17283 13429
rect 17718 13426 17724 13428
rect 17217 13424 17724 13426
rect 17217 13368 17222 13424
rect 17278 13368 17724 13424
rect 17217 13366 17724 13368
rect 17217 13363 17283 13366
rect 17718 13364 17724 13366
rect 17788 13364 17794 13428
rect 0 13290 480 13320
rect 2129 13290 2195 13293
rect 0 13288 2195 13290
rect 0 13232 2134 13288
rect 2190 13232 2195 13288
rect 0 13230 2195 13232
rect 0 13200 480 13230
rect 2129 13227 2195 13230
rect 4409 13088 4729 13089
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 13023 4729 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 18270 13088 18590 13089
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 13023 18590 13024
rect 19885 13018 19951 13021
rect 22520 13018 23000 13048
rect 19885 13016 23000 13018
rect 19885 12960 19890 13016
rect 19946 12960 23000 13016
rect 19885 12958 23000 12960
rect 19885 12955 19951 12958
rect 22520 12928 23000 12958
rect 0 12746 480 12776
rect 4061 12746 4127 12749
rect 0 12744 4127 12746
rect 0 12688 4066 12744
rect 4122 12688 4127 12744
rect 0 12686 4127 12688
rect 0 12656 480 12686
rect 4061 12683 4127 12686
rect 12709 12746 12775 12749
rect 12893 12746 12959 12749
rect 12709 12744 12959 12746
rect 12709 12688 12714 12744
rect 12770 12688 12898 12744
rect 12954 12688 12959 12744
rect 12709 12686 12959 12688
rect 12709 12683 12775 12686
rect 12893 12683 12959 12686
rect 11237 12610 11303 12613
rect 13813 12610 13879 12613
rect 11237 12608 13879 12610
rect 11237 12552 11242 12608
rect 11298 12552 13818 12608
rect 13874 12552 13879 12608
rect 11237 12550 13879 12552
rect 11237 12547 11303 12550
rect 13813 12547 13879 12550
rect 18045 12610 18111 12613
rect 22520 12610 23000 12640
rect 18045 12608 23000 12610
rect 18045 12552 18050 12608
rect 18106 12552 23000 12608
rect 18045 12550 23000 12552
rect 18045 12547 18111 12550
rect 7874 12544 8194 12545
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8194 12544
rect 7874 12479 8194 12480
rect 14805 12544 15125 12545
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 22520 12520 23000 12550
rect 14805 12479 15125 12480
rect 13445 12474 13511 12477
rect 13721 12474 13787 12477
rect 13445 12472 13787 12474
rect 13445 12416 13450 12472
rect 13506 12416 13726 12472
rect 13782 12416 13787 12472
rect 13445 12414 13787 12416
rect 13445 12411 13511 12414
rect 13721 12411 13787 12414
rect 0 12338 480 12368
rect 4061 12338 4127 12341
rect 0 12336 4127 12338
rect 0 12280 4066 12336
rect 4122 12280 4127 12336
rect 0 12278 4127 12280
rect 0 12248 480 12278
rect 4061 12275 4127 12278
rect 12341 12202 12407 12205
rect 17309 12202 17375 12205
rect 12341 12200 12818 12202
rect 12341 12144 12346 12200
rect 12402 12144 12818 12200
rect 12341 12142 12818 12144
rect 12341 12139 12407 12142
rect 4409 12000 4729 12001
rect 0 11930 480 11960
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 11935 4729 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 12758 11933 12818 12142
rect 17309 12200 19994 12202
rect 17309 12144 17314 12200
rect 17370 12144 19994 12200
rect 17309 12142 19994 12144
rect 17309 12139 17375 12142
rect 19934 12066 19994 12142
rect 22520 12066 23000 12096
rect 19934 12006 23000 12066
rect 18270 12000 18590 12001
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 22520 11976 23000 12006
rect 18270 11935 18590 11936
rect 3877 11930 3943 11933
rect 0 11928 3943 11930
rect 0 11872 3882 11928
rect 3938 11872 3943 11928
rect 0 11870 3943 11872
rect 12758 11928 12867 11933
rect 12758 11872 12806 11928
rect 12862 11872 12867 11928
rect 12758 11870 12867 11872
rect 0 11840 480 11870
rect 3877 11867 3943 11870
rect 12801 11867 12867 11870
rect 16941 11658 17007 11661
rect 22520 11658 23000 11688
rect 16941 11656 23000 11658
rect 16941 11600 16946 11656
rect 17002 11600 23000 11656
rect 16941 11598 23000 11600
rect 16941 11595 17007 11598
rect 22520 11568 23000 11598
rect 7874 11456 8194 11457
rect 0 11386 480 11416
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8194 11456
rect 7874 11391 8194 11392
rect 14805 11456 15125 11457
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 11391 15125 11392
rect 3785 11386 3851 11389
rect 0 11384 3851 11386
rect 0 11328 3790 11384
rect 3846 11328 3851 11384
rect 0 11326 3851 11328
rect 0 11296 480 11326
rect 3785 11323 3851 11326
rect 17718 11324 17724 11388
rect 17788 11386 17794 11388
rect 18137 11386 18203 11389
rect 17788 11384 18203 11386
rect 17788 11328 18142 11384
rect 18198 11328 18203 11384
rect 17788 11326 18203 11328
rect 17788 11324 17794 11326
rect 18137 11323 18203 11326
rect 15193 11250 15259 11253
rect 22520 11250 23000 11280
rect 15193 11248 23000 11250
rect 15193 11192 15198 11248
rect 15254 11192 23000 11248
rect 15193 11190 23000 11192
rect 15193 11187 15259 11190
rect 22520 11160 23000 11190
rect 7833 11114 7899 11117
rect 4156 11112 7899 11114
rect 4156 11056 7838 11112
rect 7894 11056 7899 11112
rect 4156 11054 7899 11056
rect 0 10978 480 11008
rect 4156 10978 4216 11054
rect 7833 11051 7899 11054
rect 0 10918 4216 10978
rect 0 10888 480 10918
rect 4409 10912 4729 10913
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 10847 4729 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 18270 10912 18590 10913
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 18270 10847 18590 10848
rect 3233 10706 3299 10709
rect 8569 10706 8635 10709
rect 18873 10708 18939 10709
rect 18822 10706 18828 10708
rect 3233 10704 8635 10706
rect 3233 10648 3238 10704
rect 3294 10648 8574 10704
rect 8630 10648 8635 10704
rect 3233 10646 8635 10648
rect 18782 10646 18828 10706
rect 18892 10704 18939 10708
rect 18934 10648 18939 10704
rect 3233 10643 3299 10646
rect 8569 10643 8635 10646
rect 18822 10644 18828 10646
rect 18892 10644 18939 10648
rect 18873 10643 18939 10644
rect 19241 10706 19307 10709
rect 22520 10706 23000 10736
rect 19241 10704 23000 10706
rect 19241 10648 19246 10704
rect 19302 10648 23000 10704
rect 19241 10646 23000 10648
rect 19241 10643 19307 10646
rect 22520 10616 23000 10646
rect 0 10570 480 10600
rect 4061 10570 4127 10573
rect 0 10568 4127 10570
rect 0 10512 4066 10568
rect 4122 10512 4127 10568
rect 0 10510 4127 10512
rect 0 10480 480 10510
rect 4061 10507 4127 10510
rect 4337 10570 4403 10573
rect 7557 10570 7623 10573
rect 8845 10570 8911 10573
rect 4337 10568 8911 10570
rect 4337 10512 4342 10568
rect 4398 10512 7562 10568
rect 7618 10512 8850 10568
rect 8906 10512 8911 10568
rect 4337 10510 8911 10512
rect 4337 10507 4403 10510
rect 7557 10507 7623 10510
rect 8845 10507 8911 10510
rect 11421 10570 11487 10573
rect 18781 10570 18847 10573
rect 11421 10568 18847 10570
rect 11421 10512 11426 10568
rect 11482 10512 18786 10568
rect 18842 10512 18847 10568
rect 11421 10510 18847 10512
rect 11421 10507 11487 10510
rect 18781 10507 18847 10510
rect 7874 10368 8194 10369
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8194 10368
rect 7874 10303 8194 10304
rect 14805 10368 15125 10369
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 10303 15125 10304
rect 2957 10298 3023 10301
rect 7097 10298 7163 10301
rect 2957 10296 7163 10298
rect 2957 10240 2962 10296
rect 3018 10240 7102 10296
rect 7158 10240 7163 10296
rect 2957 10238 7163 10240
rect 2957 10235 3023 10238
rect 7097 10235 7163 10238
rect 17861 10298 17927 10301
rect 22520 10298 23000 10328
rect 17861 10296 23000 10298
rect 17861 10240 17866 10296
rect 17922 10240 23000 10296
rect 17861 10238 23000 10240
rect 17861 10235 17927 10238
rect 22520 10208 23000 10238
rect 7281 10162 7347 10165
rect 4846 10160 7347 10162
rect 4846 10104 7286 10160
rect 7342 10104 7347 10160
rect 4846 10102 7347 10104
rect 0 10026 480 10056
rect 4846 10026 4906 10102
rect 7281 10099 7347 10102
rect 13997 10162 14063 10165
rect 17534 10162 17540 10164
rect 13997 10160 17540 10162
rect 13997 10104 14002 10160
rect 14058 10104 17540 10160
rect 13997 10102 17540 10104
rect 13997 10099 14063 10102
rect 17534 10100 17540 10102
rect 17604 10162 17610 10164
rect 18045 10162 18111 10165
rect 17604 10160 18111 10162
rect 17604 10104 18050 10160
rect 18106 10104 18111 10160
rect 17604 10102 18111 10104
rect 17604 10100 17610 10102
rect 18045 10099 18111 10102
rect 0 9966 4906 10026
rect 5901 10026 5967 10029
rect 6545 10026 6611 10029
rect 5901 10024 6611 10026
rect 5901 9968 5906 10024
rect 5962 9968 6550 10024
rect 6606 9968 6611 10024
rect 5901 9966 6611 9968
rect 0 9936 480 9966
rect 5901 9963 5967 9966
rect 6545 9963 6611 9966
rect 15101 10026 15167 10029
rect 17953 10026 18019 10029
rect 15101 10024 18019 10026
rect 15101 9968 15106 10024
rect 15162 9968 17958 10024
rect 18014 9968 18019 10024
rect 18232 9992 18752 10026
rect 15101 9966 18019 9968
rect 15101 9963 15167 9966
rect 17953 9963 18019 9966
rect 18094 9966 18752 9992
rect 18094 9932 18292 9966
rect 12617 9890 12683 9893
rect 18094 9890 18154 9932
rect 12617 9888 18154 9890
rect 12617 9832 12622 9888
rect 12678 9832 18154 9888
rect 12617 9830 18154 9832
rect 12617 9827 12683 9830
rect 4409 9824 4729 9825
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 9759 4729 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 18270 9824 18590 9825
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 9759 18590 9760
rect 2957 9754 3023 9757
rect 3325 9754 3391 9757
rect 2957 9752 3391 9754
rect 2957 9696 2962 9752
rect 3018 9696 3330 9752
rect 3386 9696 3391 9752
rect 2957 9694 3391 9696
rect 2957 9691 3023 9694
rect 3325 9691 3391 9694
rect 12157 9754 12223 9757
rect 14641 9754 14707 9757
rect 12157 9752 14707 9754
rect 12157 9696 12162 9752
rect 12218 9696 14646 9752
rect 14702 9696 14707 9752
rect 12157 9694 14707 9696
rect 18692 9754 18752 9966
rect 22520 9754 23000 9784
rect 18692 9694 23000 9754
rect 12157 9691 12223 9694
rect 14641 9691 14707 9694
rect 22520 9664 23000 9694
rect 0 9618 480 9648
rect 3785 9618 3851 9621
rect 0 9616 3851 9618
rect 0 9560 3790 9616
rect 3846 9560 3851 9616
rect 0 9558 3851 9560
rect 0 9528 480 9558
rect 3785 9555 3851 9558
rect 11094 9556 11100 9620
rect 11164 9618 11170 9620
rect 18505 9618 18571 9621
rect 11164 9616 18571 9618
rect 11164 9560 18510 9616
rect 18566 9560 18571 9616
rect 11164 9558 18571 9560
rect 11164 9556 11170 9558
rect 18505 9555 18571 9558
rect 10317 9482 10383 9485
rect 18229 9482 18295 9485
rect 10317 9480 18295 9482
rect 10317 9424 10322 9480
rect 10378 9424 18234 9480
rect 18290 9424 18295 9480
rect 10317 9422 18295 9424
rect 10317 9419 10383 9422
rect 18229 9419 18295 9422
rect 18045 9346 18111 9349
rect 19006 9346 19012 9348
rect 18045 9344 19012 9346
rect 18045 9288 18050 9344
rect 18106 9288 19012 9344
rect 18045 9286 19012 9288
rect 18045 9283 18111 9286
rect 19006 9284 19012 9286
rect 19076 9284 19082 9348
rect 19149 9346 19215 9349
rect 22520 9346 23000 9376
rect 19149 9344 23000 9346
rect 19149 9288 19154 9344
rect 19210 9288 23000 9344
rect 19149 9286 23000 9288
rect 19149 9283 19215 9286
rect 7874 9280 8194 9281
rect 0 9210 480 9240
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8194 9280
rect 7874 9215 8194 9216
rect 14805 9280 15125 9281
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 22520 9256 23000 9286
rect 14805 9215 15125 9216
rect 4061 9210 4127 9213
rect 11789 9212 11855 9213
rect 11789 9210 11836 9212
rect 0 9208 4127 9210
rect 0 9152 4066 9208
rect 4122 9152 4127 9208
rect 0 9150 4127 9152
rect 11744 9208 11836 9210
rect 11744 9152 11794 9208
rect 11744 9150 11836 9152
rect 0 9120 480 9150
rect 4061 9147 4127 9150
rect 11789 9148 11836 9150
rect 11900 9148 11906 9212
rect 11789 9147 11855 9148
rect 9673 9074 9739 9077
rect 10777 9074 10843 9077
rect 14365 9074 14431 9077
rect 18137 9074 18203 9077
rect 18781 9076 18847 9077
rect 18781 9074 18828 9076
rect 9673 9072 18203 9074
rect 9673 9016 9678 9072
rect 9734 9016 10782 9072
rect 10838 9016 14370 9072
rect 14426 9016 18142 9072
rect 18198 9016 18203 9072
rect 9673 9014 18203 9016
rect 18736 9072 18828 9074
rect 18736 9016 18786 9072
rect 18736 9014 18828 9016
rect 9673 9011 9739 9014
rect 10777 9011 10843 9014
rect 14365 9011 14431 9014
rect 18137 9011 18203 9014
rect 18781 9012 18828 9014
rect 18892 9012 18898 9076
rect 18781 9011 18847 9012
rect 10961 8938 11027 8941
rect 16665 8938 16731 8941
rect 10961 8936 16731 8938
rect 10961 8880 10966 8936
rect 11022 8880 16670 8936
rect 16726 8880 16731 8936
rect 10961 8878 16731 8880
rect 10961 8875 11027 8878
rect 16665 8875 16731 8878
rect 18137 8938 18203 8941
rect 22520 8938 23000 8968
rect 18137 8936 23000 8938
rect 18137 8880 18142 8936
rect 18198 8880 23000 8936
rect 18137 8878 23000 8880
rect 18137 8875 18203 8878
rect 22520 8848 23000 8878
rect 4409 8736 4729 8737
rect 0 8666 480 8696
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 8671 4729 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 18270 8736 18590 8737
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 8671 18590 8672
rect 4061 8666 4127 8669
rect 0 8664 4127 8666
rect 0 8608 4066 8664
rect 4122 8608 4127 8664
rect 0 8606 4127 8608
rect 0 8576 480 8606
rect 4061 8603 4127 8606
rect 14641 8530 14707 8533
rect 17769 8530 17835 8533
rect 14641 8528 17835 8530
rect 14641 8472 14646 8528
rect 14702 8472 17774 8528
rect 17830 8472 17835 8528
rect 14641 8470 17835 8472
rect 14641 8467 14707 8470
rect 17769 8467 17835 8470
rect 5073 8394 5139 8397
rect 8569 8394 8635 8397
rect 5073 8392 8635 8394
rect 5073 8336 5078 8392
rect 5134 8336 8574 8392
rect 8630 8336 8635 8392
rect 5073 8334 8635 8336
rect 5073 8331 5139 8334
rect 8569 8331 8635 8334
rect 13629 8394 13695 8397
rect 22520 8394 23000 8424
rect 13629 8392 23000 8394
rect 13629 8336 13634 8392
rect 13690 8336 23000 8392
rect 13629 8334 23000 8336
rect 13629 8331 13695 8334
rect 22520 8304 23000 8334
rect 0 8258 480 8288
rect 3785 8258 3851 8261
rect 0 8256 3851 8258
rect 0 8200 3790 8256
rect 3846 8200 3851 8256
rect 0 8198 3851 8200
rect 0 8168 480 8198
rect 3785 8195 3851 8198
rect 7874 8192 8194 8193
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8194 8192
rect 7874 8127 8194 8128
rect 14805 8192 15125 8193
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 8127 15125 8128
rect 18873 8122 18939 8125
rect 19006 8122 19012 8124
rect 18873 8120 19012 8122
rect 18873 8064 18878 8120
rect 18934 8064 19012 8120
rect 18873 8062 19012 8064
rect 18873 8059 18939 8062
rect 19006 8060 19012 8062
rect 19076 8060 19082 8124
rect 12525 7986 12591 7989
rect 22520 7986 23000 8016
rect 12525 7984 23000 7986
rect 12525 7928 12530 7984
rect 12586 7928 23000 7984
rect 12525 7926 23000 7928
rect 12525 7923 12591 7926
rect 22520 7896 23000 7926
rect 0 7850 480 7880
rect 4061 7850 4127 7853
rect 0 7848 4127 7850
rect 0 7792 4066 7848
rect 4122 7792 4127 7848
rect 0 7790 4127 7792
rect 0 7760 480 7790
rect 4061 7787 4127 7790
rect 11973 7850 12039 7853
rect 12985 7850 13051 7853
rect 11973 7848 13051 7850
rect 11973 7792 11978 7848
rect 12034 7792 12990 7848
rect 13046 7792 13051 7848
rect 11973 7790 13051 7792
rect 11973 7787 12039 7790
rect 12985 7787 13051 7790
rect 4409 7648 4729 7649
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 7583 4729 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 18270 7648 18590 7649
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 18270 7583 18590 7584
rect 16021 7578 16087 7581
rect 16205 7578 16271 7581
rect 16021 7576 16271 7578
rect 16021 7520 16026 7576
rect 16082 7520 16210 7576
rect 16266 7520 16271 7576
rect 16021 7518 16271 7520
rect 16021 7515 16087 7518
rect 16205 7515 16271 7518
rect 18781 7578 18847 7581
rect 22520 7578 23000 7608
rect 18781 7576 23000 7578
rect 18781 7520 18786 7576
rect 18842 7520 23000 7576
rect 18781 7518 23000 7520
rect 18781 7515 18847 7518
rect 22520 7488 23000 7518
rect 0 7442 480 7472
rect 9581 7442 9647 7445
rect 0 7440 9647 7442
rect 0 7384 9586 7440
rect 9642 7384 9647 7440
rect 0 7382 9647 7384
rect 0 7352 480 7382
rect 9581 7379 9647 7382
rect 3693 7306 3759 7309
rect 9581 7306 9647 7309
rect 3693 7304 9647 7306
rect 3693 7248 3698 7304
rect 3754 7248 9586 7304
rect 9642 7248 9647 7304
rect 3693 7246 9647 7248
rect 3693 7243 3759 7246
rect 9581 7243 9647 7246
rect 12157 7306 12223 7309
rect 17033 7306 17099 7309
rect 12157 7304 17099 7306
rect 12157 7248 12162 7304
rect 12218 7248 17038 7304
rect 17094 7248 17099 7304
rect 12157 7246 17099 7248
rect 12157 7243 12223 7246
rect 17033 7243 17099 7246
rect 2773 7170 2839 7173
rect 7557 7170 7623 7173
rect 2773 7168 7623 7170
rect 2773 7112 2778 7168
rect 2834 7112 7562 7168
rect 7618 7112 7623 7168
rect 2773 7110 7623 7112
rect 2773 7107 2839 7110
rect 7557 7107 7623 7110
rect 12249 7170 12315 7173
rect 13905 7170 13971 7173
rect 12249 7168 13971 7170
rect 12249 7112 12254 7168
rect 12310 7112 13910 7168
rect 13966 7112 13971 7168
rect 12249 7110 13971 7112
rect 12249 7107 12315 7110
rect 13905 7107 13971 7110
rect 7874 7104 8194 7105
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8194 7104
rect 7874 7039 8194 7040
rect 14805 7104 15125 7105
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 7039 15125 7040
rect 7189 7034 7255 7037
rect 2638 7032 7255 7034
rect 2638 6976 7194 7032
rect 7250 6976 7255 7032
rect 2638 6974 7255 6976
rect 0 6898 480 6928
rect 2037 6898 2103 6901
rect 0 6896 2103 6898
rect 0 6840 2042 6896
rect 2098 6840 2103 6896
rect 0 6838 2103 6840
rect 0 6808 480 6838
rect 2037 6835 2103 6838
rect 0 6490 480 6520
rect 2638 6490 2698 6974
rect 7189 6971 7255 6974
rect 17953 7034 18019 7037
rect 22520 7034 23000 7064
rect 17953 7032 23000 7034
rect 17953 6976 17958 7032
rect 18014 6976 23000 7032
rect 17953 6974 23000 6976
rect 17953 6971 18019 6974
rect 22520 6944 23000 6974
rect 12157 6898 12223 6901
rect 12525 6898 12591 6901
rect 12157 6896 12591 6898
rect 12157 6840 12162 6896
rect 12218 6840 12530 6896
rect 12586 6840 12591 6896
rect 12157 6838 12591 6840
rect 12157 6835 12223 6838
rect 12525 6835 12591 6838
rect 2865 6762 2931 6765
rect 2998 6762 3004 6764
rect 2865 6760 3004 6762
rect 2865 6704 2870 6760
rect 2926 6704 3004 6760
rect 2865 6702 3004 6704
rect 2865 6699 2931 6702
rect 2998 6700 3004 6702
rect 3068 6762 3074 6764
rect 8845 6762 8911 6765
rect 3068 6760 8911 6762
rect 3068 6704 8850 6760
rect 8906 6704 8911 6760
rect 3068 6702 8911 6704
rect 3068 6700 3074 6702
rect 8845 6699 8911 6702
rect 12157 6762 12223 6765
rect 17309 6762 17375 6765
rect 12157 6760 17375 6762
rect 12157 6704 12162 6760
rect 12218 6704 17314 6760
rect 17370 6704 17375 6760
rect 12157 6702 17375 6704
rect 12157 6699 12223 6702
rect 17309 6699 17375 6702
rect 22520 6626 23000 6656
rect 18784 6566 23000 6626
rect 4409 6560 4729 6561
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 6495 4729 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 18270 6560 18590 6561
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 6495 18590 6496
rect 0 6430 2698 6490
rect 0 6400 480 6430
rect 2589 6354 2655 6357
rect 4613 6354 4679 6357
rect 2589 6352 4679 6354
rect 2589 6296 2594 6352
rect 2650 6296 4618 6352
rect 4674 6296 4679 6352
rect 2589 6294 4679 6296
rect 2589 6291 2655 6294
rect 4613 6291 4679 6294
rect 11605 6354 11671 6357
rect 18784 6354 18844 6566
rect 22520 6536 23000 6566
rect 11605 6352 18844 6354
rect 11605 6296 11610 6352
rect 11666 6296 18844 6352
rect 11605 6294 18844 6296
rect 11605 6291 11671 6294
rect 0 6082 480 6112
rect 2221 6082 2287 6085
rect 0 6080 2287 6082
rect 0 6024 2226 6080
rect 2282 6024 2287 6080
rect 0 6022 2287 6024
rect 0 5992 480 6022
rect 2221 6019 2287 6022
rect 2497 6082 2563 6085
rect 7281 6082 7347 6085
rect 2497 6080 7347 6082
rect 2497 6024 2502 6080
rect 2558 6024 7286 6080
rect 7342 6024 7347 6080
rect 2497 6022 7347 6024
rect 2497 6019 2563 6022
rect 7281 6019 7347 6022
rect 17953 6082 18019 6085
rect 22520 6082 23000 6112
rect 17953 6080 23000 6082
rect 17953 6024 17958 6080
rect 18014 6024 23000 6080
rect 17953 6022 23000 6024
rect 17953 6019 18019 6022
rect 7874 6016 8194 6017
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8194 6016
rect 7874 5951 8194 5952
rect 14805 6016 15125 6017
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 22520 5992 23000 6022
rect 14805 5951 15125 5952
rect 6269 5946 6335 5949
rect 7373 5946 7439 5949
rect 6269 5944 7439 5946
rect 6269 5888 6274 5944
rect 6330 5888 7378 5944
rect 7434 5888 7439 5944
rect 6269 5886 7439 5888
rect 6269 5883 6335 5886
rect 7373 5883 7439 5886
rect 5257 5810 5323 5813
rect 8385 5810 8451 5813
rect 5257 5808 8451 5810
rect 5257 5752 5262 5808
rect 5318 5752 8390 5808
rect 8446 5752 8451 5808
rect 5257 5750 8451 5752
rect 5257 5747 5323 5750
rect 8385 5747 8451 5750
rect 2497 5674 2563 5677
rect 5809 5674 5875 5677
rect 6637 5674 6703 5677
rect 2497 5672 6703 5674
rect 2497 5616 2502 5672
rect 2558 5616 5814 5672
rect 5870 5616 6642 5672
rect 6698 5616 6703 5672
rect 2497 5614 6703 5616
rect 2497 5611 2563 5614
rect 5809 5611 5875 5614
rect 6637 5611 6703 5614
rect 8845 5674 8911 5677
rect 9581 5674 9647 5677
rect 8845 5672 9647 5674
rect 8845 5616 8850 5672
rect 8906 5616 9586 5672
rect 9642 5616 9647 5672
rect 8845 5614 9647 5616
rect 8845 5611 8911 5614
rect 9581 5611 9647 5614
rect 11237 5674 11303 5677
rect 22520 5674 23000 5704
rect 11237 5672 23000 5674
rect 11237 5616 11242 5672
rect 11298 5616 23000 5672
rect 11237 5614 23000 5616
rect 11237 5611 11303 5614
rect 22520 5584 23000 5614
rect 0 5538 480 5568
rect 3877 5538 3943 5541
rect 9857 5540 9923 5541
rect 9806 5538 9812 5540
rect 0 5536 3943 5538
rect 0 5480 3882 5536
rect 3938 5480 3943 5536
rect 0 5478 3943 5480
rect 9766 5478 9812 5538
rect 9876 5536 9923 5540
rect 9918 5480 9923 5536
rect 0 5448 480 5478
rect 3877 5475 3943 5478
rect 9806 5476 9812 5478
rect 9876 5476 9923 5480
rect 9857 5475 9923 5476
rect 4409 5472 4729 5473
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 5407 4729 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 18270 5472 18590 5473
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 5407 18590 5408
rect 3233 5266 3299 5269
rect 9489 5266 9555 5269
rect 3233 5264 9555 5266
rect 3233 5208 3238 5264
rect 3294 5208 9494 5264
rect 9550 5208 9555 5264
rect 3233 5206 9555 5208
rect 3233 5203 3299 5206
rect 9489 5203 9555 5206
rect 9673 5266 9739 5269
rect 11053 5266 11119 5269
rect 9673 5264 11119 5266
rect 9673 5208 9678 5264
rect 9734 5208 11058 5264
rect 11114 5208 11119 5264
rect 9673 5206 11119 5208
rect 9673 5203 9739 5206
rect 11053 5203 11119 5206
rect 19425 5266 19491 5269
rect 22520 5266 23000 5296
rect 19425 5264 23000 5266
rect 19425 5208 19430 5264
rect 19486 5208 23000 5264
rect 19425 5206 23000 5208
rect 19425 5203 19491 5206
rect 22520 5176 23000 5206
rect 0 5130 480 5160
rect 3785 5130 3851 5133
rect 0 5128 3851 5130
rect 0 5072 3790 5128
rect 3846 5072 3851 5128
rect 0 5070 3851 5072
rect 0 5040 480 5070
rect 3785 5067 3851 5070
rect 4061 5130 4127 5133
rect 19609 5130 19675 5133
rect 4061 5128 19675 5130
rect 4061 5072 4066 5128
rect 4122 5072 19614 5128
rect 19670 5072 19675 5128
rect 4061 5070 19675 5072
rect 4061 5067 4127 5070
rect 19609 5067 19675 5070
rect 2405 4994 2471 4997
rect 5717 4994 5783 4997
rect 2405 4992 5783 4994
rect 2405 4936 2410 4992
rect 2466 4936 5722 4992
rect 5778 4936 5783 4992
rect 2405 4934 5783 4936
rect 2405 4931 2471 4934
rect 5717 4931 5783 4934
rect 9949 4994 10015 4997
rect 12985 4994 13051 4997
rect 9949 4992 13051 4994
rect 9949 4936 9954 4992
rect 10010 4936 12990 4992
rect 13046 4936 13051 4992
rect 9949 4934 13051 4936
rect 9949 4931 10015 4934
rect 12985 4931 13051 4934
rect 7874 4928 8194 4929
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8194 4928
rect 7874 4863 8194 4864
rect 14805 4928 15125 4929
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 4863 15125 4864
rect 13445 4858 13511 4861
rect 3374 4798 7436 4858
rect 0 4722 480 4752
rect 3374 4722 3434 4798
rect 0 4662 3434 4722
rect 3601 4722 3667 4725
rect 7376 4722 7436 4798
rect 10320 4856 13511 4858
rect 10320 4800 13450 4856
rect 13506 4800 13511 4856
rect 10320 4798 13511 4800
rect 7925 4722 7991 4725
rect 3601 4720 7252 4722
rect 3601 4664 3606 4720
rect 3662 4664 7252 4720
rect 3601 4662 7252 4664
rect 7376 4720 7991 4722
rect 7376 4664 7930 4720
rect 7986 4664 7991 4720
rect 7376 4662 7991 4664
rect 0 4632 480 4662
rect 3601 4659 3667 4662
rect 3877 4586 3943 4589
rect 7005 4586 7071 4589
rect 3877 4584 7071 4586
rect 3877 4528 3882 4584
rect 3938 4528 7010 4584
rect 7066 4528 7071 4584
rect 3877 4526 7071 4528
rect 7192 4586 7252 4662
rect 7925 4659 7991 4662
rect 8109 4722 8175 4725
rect 9857 4722 9923 4725
rect 10320 4722 10380 4798
rect 13445 4795 13511 4798
rect 8109 4720 8540 4722
rect 8109 4664 8114 4720
rect 8170 4688 8540 4720
rect 9857 4720 10380 4722
rect 8170 4664 8586 4688
rect 8109 4662 8586 4664
rect 8109 4659 8175 4662
rect 8480 4628 8586 4662
rect 9857 4664 9862 4720
rect 9918 4664 10380 4720
rect 9857 4662 10380 4664
rect 13261 4722 13327 4725
rect 13537 4722 13603 4725
rect 13261 4720 13603 4722
rect 13261 4664 13266 4720
rect 13322 4664 13542 4720
rect 13598 4664 13603 4720
rect 13261 4662 13603 4664
rect 9857 4659 9923 4662
rect 13261 4659 13327 4662
rect 13537 4659 13603 4662
rect 15745 4722 15811 4725
rect 22520 4722 23000 4752
rect 15745 4720 23000 4722
rect 15745 4664 15750 4720
rect 15806 4664 23000 4720
rect 15745 4662 23000 4664
rect 15745 4659 15811 4662
rect 22520 4632 23000 4662
rect 8526 4586 8586 4628
rect 7192 4552 7666 4586
rect 7974 4554 8402 4586
rect 7974 4552 8340 4554
rect 7192 4526 8340 4552
rect 3877 4523 3943 4526
rect 7005 4523 7071 4526
rect 7606 4492 8034 4526
rect 8334 4490 8340 4526
rect 8404 4490 8410 4554
rect 8526 4552 9644 4586
rect 9814 4552 11852 4586
rect 8526 4526 11852 4552
rect 9584 4492 9874 4526
rect 10225 4450 10291 4453
rect 11145 4450 11211 4453
rect 10225 4448 11211 4450
rect 10225 4392 10230 4448
rect 10286 4392 11150 4448
rect 11206 4392 11211 4448
rect 10225 4390 11211 4392
rect 11792 4452 11852 4526
rect 11792 4390 11836 4452
rect 10225 4387 10291 4390
rect 11145 4387 11211 4390
rect 11830 4388 11836 4390
rect 11900 4450 11906 4452
rect 12893 4450 12959 4453
rect 11900 4448 12959 4450
rect 11900 4392 12898 4448
rect 12954 4392 12959 4448
rect 11900 4390 12959 4392
rect 11900 4388 11906 4390
rect 12893 4387 12959 4390
rect 4409 4384 4729 4385
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 4319 4729 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 18270 4384 18590 4385
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 18270 4319 18590 4320
rect 3969 4314 4035 4317
rect 3788 4312 4035 4314
rect 3788 4256 3974 4312
rect 4030 4256 4035 4312
rect 3788 4254 4035 4256
rect 0 4178 480 4208
rect 3788 4178 3848 4254
rect 3969 4251 4035 4254
rect 20529 4314 20595 4317
rect 22520 4314 23000 4344
rect 20529 4312 23000 4314
rect 20529 4256 20534 4312
rect 20590 4256 23000 4312
rect 20529 4254 23000 4256
rect 20529 4251 20595 4254
rect 22520 4224 23000 4254
rect 7373 4178 7439 4181
rect 0 4118 3848 4178
rect 3926 4176 7439 4178
rect 3926 4120 7378 4176
rect 7434 4120 7439 4176
rect 3926 4118 7439 4120
rect 0 4088 480 4118
rect 3141 4042 3207 4045
rect 3926 4042 3986 4118
rect 7373 4115 7439 4118
rect 10225 4178 10291 4181
rect 14549 4178 14615 4181
rect 10225 4176 14615 4178
rect 10225 4120 10230 4176
rect 10286 4120 14554 4176
rect 14610 4120 14615 4176
rect 10225 4118 14615 4120
rect 10225 4115 10291 4118
rect 14549 4115 14615 4118
rect 3141 4040 3986 4042
rect 3141 3984 3146 4040
rect 3202 3984 3986 4040
rect 3141 3982 3986 3984
rect 4429 4042 4495 4045
rect 14273 4042 14339 4045
rect 20253 4042 20319 4045
rect 4429 4040 14339 4042
rect 4429 3984 4434 4040
rect 4490 3984 14278 4040
rect 14334 3984 14339 4040
rect 4429 3982 14339 3984
rect 3141 3979 3207 3982
rect 4429 3979 4495 3982
rect 14273 3979 14339 3982
rect 14598 4040 20319 4042
rect 14598 3984 20258 4040
rect 20314 3984 20319 4040
rect 14598 3982 20319 3984
rect 4061 3906 4127 3909
rect 5073 3906 5139 3909
rect 9857 3908 9923 3909
rect 4061 3904 5139 3906
rect 4061 3848 4066 3904
rect 4122 3848 5078 3904
rect 5134 3848 5139 3904
rect 4061 3846 5139 3848
rect 4061 3843 4127 3846
rect 5073 3843 5139 3846
rect 9806 3844 9812 3908
rect 9876 3906 9923 3908
rect 10317 3906 10383 3909
rect 14598 3906 14658 3982
rect 20253 3979 20319 3982
rect 9876 3904 9968 3906
rect 9918 3848 9968 3904
rect 9876 3846 9968 3848
rect 10317 3904 14658 3906
rect 10317 3848 10322 3904
rect 10378 3848 14658 3904
rect 10317 3846 14658 3848
rect 20529 3906 20595 3909
rect 22520 3906 23000 3936
rect 20529 3904 23000 3906
rect 20529 3848 20534 3904
rect 20590 3848 23000 3904
rect 20529 3846 23000 3848
rect 9876 3844 9923 3846
rect 9857 3843 9923 3844
rect 10317 3843 10383 3846
rect 20529 3843 20595 3846
rect 7874 3840 8194 3841
rect 0 3770 480 3800
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8194 3840
rect 7874 3775 8194 3776
rect 14805 3840 15125 3841
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 22520 3816 23000 3846
rect 14805 3775 15125 3776
rect 0 3710 3066 3770
rect 0 3680 480 3710
rect 3006 3634 3066 3710
rect 8334 3708 8340 3772
rect 8404 3770 8410 3772
rect 16021 3770 16087 3773
rect 20345 3770 20411 3773
rect 8404 3710 12082 3770
rect 8404 3708 8410 3710
rect 3325 3634 3391 3637
rect 3006 3632 3391 3634
rect 3006 3576 3330 3632
rect 3386 3576 3391 3632
rect 3006 3574 3391 3576
rect 3325 3571 3391 3574
rect 3693 3634 3759 3637
rect 11789 3634 11855 3637
rect 3693 3632 11855 3634
rect 3693 3576 3698 3632
rect 3754 3576 11794 3632
rect 11850 3576 11855 3632
rect 3693 3574 11855 3576
rect 12022 3634 12082 3710
rect 16021 3768 20411 3770
rect 16021 3712 16026 3768
rect 16082 3712 20350 3768
rect 20406 3712 20411 3768
rect 16021 3710 20411 3712
rect 16021 3707 16087 3710
rect 20345 3707 20411 3710
rect 19793 3634 19859 3637
rect 12022 3632 19859 3634
rect 12022 3576 19798 3632
rect 19854 3576 19859 3632
rect 12022 3574 19859 3576
rect 3693 3571 3759 3574
rect 11789 3571 11855 3574
rect 19793 3571 19859 3574
rect 1669 3498 1735 3501
rect 5165 3498 5231 3501
rect 1669 3496 5231 3498
rect 1669 3440 1674 3496
rect 1730 3440 5170 3496
rect 5226 3440 5231 3496
rect 1669 3438 5231 3440
rect 1669 3435 1735 3438
rect 5165 3435 5231 3438
rect 6361 3498 6427 3501
rect 14089 3498 14155 3501
rect 6361 3496 14155 3498
rect 6361 3440 6366 3496
rect 6422 3440 14094 3496
rect 14150 3440 14155 3496
rect 6361 3438 14155 3440
rect 6361 3435 6427 3438
rect 14089 3435 14155 3438
rect 14273 3498 14339 3501
rect 20069 3498 20135 3501
rect 14273 3496 20135 3498
rect 14273 3440 14278 3496
rect 14334 3440 20074 3496
rect 20130 3440 20135 3496
rect 14273 3438 20135 3440
rect 14273 3435 14339 3438
rect 20069 3435 20135 3438
rect 0 3362 480 3392
rect 3049 3362 3115 3365
rect 0 3360 3115 3362
rect 0 3304 3054 3360
rect 3110 3304 3115 3360
rect 0 3302 3115 3304
rect 0 3272 480 3302
rect 3049 3299 3115 3302
rect 7373 3362 7439 3365
rect 11094 3362 11100 3364
rect 7373 3360 11100 3362
rect 7373 3304 7378 3360
rect 7434 3304 11100 3360
rect 7373 3302 11100 3304
rect 7373 3299 7439 3302
rect 11094 3300 11100 3302
rect 11164 3300 11170 3364
rect 11789 3362 11855 3365
rect 17953 3362 18019 3365
rect 11789 3360 18019 3362
rect 11789 3304 11794 3360
rect 11850 3304 17958 3360
rect 18014 3304 18019 3360
rect 11789 3302 18019 3304
rect 11789 3299 11855 3302
rect 17953 3299 18019 3302
rect 19006 3300 19012 3364
rect 19076 3362 19082 3364
rect 22520 3362 23000 3392
rect 19076 3302 23000 3362
rect 19076 3300 19082 3302
rect 4409 3296 4729 3297
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 3231 4729 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 18270 3296 18590 3297
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 22520 3272 23000 3302
rect 18270 3231 18590 3232
rect 3049 3228 3115 3229
rect 2998 3226 3004 3228
rect 2958 3166 3004 3226
rect 3068 3224 3115 3228
rect 9305 3226 9371 3229
rect 3110 3168 3115 3224
rect 2998 3164 3004 3166
rect 3068 3164 3115 3168
rect 3049 3163 3115 3164
rect 7054 3224 9371 3226
rect 7054 3168 9310 3224
rect 9366 3168 9371 3224
rect 7054 3166 9371 3168
rect 2773 3090 2839 3093
rect 7054 3090 7114 3166
rect 9305 3163 9371 3166
rect 10409 3226 10475 3229
rect 10961 3226 11027 3229
rect 10409 3224 11027 3226
rect 10409 3168 10414 3224
rect 10470 3168 10966 3224
rect 11022 3168 11027 3224
rect 10409 3166 11027 3168
rect 10409 3163 10475 3166
rect 10961 3163 11027 3166
rect 18822 3164 18828 3228
rect 18892 3226 18898 3228
rect 19057 3226 19123 3229
rect 18892 3224 19123 3226
rect 18892 3168 19062 3224
rect 19118 3168 19123 3224
rect 18892 3166 19123 3168
rect 18892 3164 18898 3166
rect 19057 3163 19123 3166
rect 2773 3088 7114 3090
rect 2773 3032 2778 3088
rect 2834 3032 7114 3088
rect 2773 3030 7114 3032
rect 7741 3090 7807 3093
rect 18086 3090 18092 3092
rect 7741 3088 18092 3090
rect 7741 3032 7746 3088
rect 7802 3032 18092 3088
rect 7741 3030 18092 3032
rect 2773 3027 2839 3030
rect 7741 3027 7807 3030
rect 18086 3028 18092 3030
rect 18156 3028 18162 3092
rect 2221 2954 2287 2957
rect 7373 2954 7439 2957
rect 2221 2952 7439 2954
rect 2221 2896 2226 2952
rect 2282 2896 7378 2952
rect 7434 2896 7439 2952
rect 2221 2894 7439 2896
rect 2221 2891 2287 2894
rect 7373 2891 7439 2894
rect 7741 2954 7807 2957
rect 9305 2954 9371 2957
rect 17309 2954 17375 2957
rect 7741 2952 9138 2954
rect 7741 2896 7746 2952
rect 7802 2896 9138 2952
rect 7741 2894 9138 2896
rect 7741 2891 7807 2894
rect 0 2818 480 2848
rect 4061 2818 4127 2821
rect 0 2816 4127 2818
rect 0 2760 4066 2816
rect 4122 2760 4127 2816
rect 0 2758 4127 2760
rect 0 2728 480 2758
rect 4061 2755 4127 2758
rect 5441 2818 5507 2821
rect 8937 2818 9003 2821
rect 5441 2816 7666 2818
rect 5441 2760 5446 2816
rect 5502 2760 7666 2816
rect 5441 2758 7666 2760
rect 5441 2755 5507 2758
rect 1761 2682 1827 2685
rect 7465 2682 7531 2685
rect 1761 2680 7531 2682
rect 1761 2624 1766 2680
rect 1822 2624 7470 2680
rect 7526 2624 7531 2680
rect 1761 2622 7531 2624
rect 1761 2619 1827 2622
rect 7465 2619 7531 2622
rect 7606 2546 7666 2758
rect 8342 2816 9003 2818
rect 8342 2760 8942 2816
rect 8998 2760 9003 2816
rect 8342 2758 9003 2760
rect 9078 2818 9138 2894
rect 9305 2952 17375 2954
rect 9305 2896 9310 2952
rect 9366 2896 17314 2952
rect 17370 2896 17375 2952
rect 9305 2894 17375 2896
rect 9305 2891 9371 2894
rect 17309 2891 17375 2894
rect 17769 2954 17835 2957
rect 22520 2954 23000 2984
rect 17769 2952 23000 2954
rect 17769 2896 17774 2952
rect 17830 2896 23000 2952
rect 17769 2894 23000 2896
rect 17769 2891 17835 2894
rect 22520 2864 23000 2894
rect 17902 2818 17908 2820
rect 9078 2758 14658 2818
rect 7874 2752 8194 2753
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8194 2752
rect 7874 2687 8194 2688
rect 8342 2546 8402 2758
rect 8937 2755 9003 2758
rect 7606 2486 8402 2546
rect 14598 2546 14658 2758
rect 15334 2758 17908 2818
rect 14805 2752 15125 2753
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2687 15125 2688
rect 15334 2546 15394 2758
rect 17902 2756 17908 2758
rect 17972 2756 17978 2820
rect 14598 2486 15394 2546
rect 0 2410 480 2440
rect 2129 2410 2195 2413
rect 0 2408 2195 2410
rect 0 2352 2134 2408
rect 2190 2352 2195 2408
rect 0 2350 2195 2352
rect 0 2320 480 2350
rect 2129 2347 2195 2350
rect 5625 2410 5691 2413
rect 8477 2410 8543 2413
rect 15285 2410 15351 2413
rect 5625 2408 15351 2410
rect 5625 2352 5630 2408
rect 5686 2352 8482 2408
rect 8538 2352 15290 2408
rect 15346 2352 15351 2408
rect 5625 2350 15351 2352
rect 5625 2347 5691 2350
rect 8477 2347 8543 2350
rect 15285 2347 15351 2350
rect 19190 2348 19196 2412
rect 19260 2410 19266 2412
rect 22520 2410 23000 2440
rect 19260 2350 23000 2410
rect 19260 2348 19266 2350
rect 22520 2320 23000 2350
rect 4409 2208 4729 2209
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2143 4729 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 18270 2208 18590 2209
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2143 18590 2144
rect 0 2002 480 2032
rect 3509 2002 3575 2005
rect 0 2000 3575 2002
rect 0 1944 3514 2000
rect 3570 1944 3575 2000
rect 0 1942 3575 1944
rect 0 1912 480 1942
rect 3509 1939 3575 1942
rect 17677 2002 17743 2005
rect 22520 2002 23000 2032
rect 17677 2000 23000 2002
rect 17677 1944 17682 2000
rect 17738 1944 23000 2000
rect 17677 1942 23000 1944
rect 17677 1939 17743 1942
rect 22520 1912 23000 1942
rect 18597 1594 18663 1597
rect 22520 1594 23000 1624
rect 18597 1592 23000 1594
rect 18597 1536 18602 1592
rect 18658 1536 23000 1592
rect 18597 1534 23000 1536
rect 18597 1531 18663 1534
rect 22520 1504 23000 1534
rect 0 1458 480 1488
rect 2221 1458 2287 1461
rect 0 1456 2287 1458
rect 0 1400 2226 1456
rect 2282 1400 2287 1456
rect 0 1398 2287 1400
rect 0 1368 480 1398
rect 2221 1395 2287 1398
rect 0 1050 480 1080
rect 6637 1050 6703 1053
rect 0 1048 6703 1050
rect 0 992 6642 1048
rect 6698 992 6703 1048
rect 0 990 6703 992
rect 0 960 480 990
rect 6637 987 6703 990
rect 18781 1050 18847 1053
rect 22520 1050 23000 1080
rect 18781 1048 23000 1050
rect 18781 992 18786 1048
rect 18842 992 23000 1048
rect 18781 990 23000 992
rect 18781 987 18847 990
rect 22520 960 23000 990
rect 0 642 480 672
rect 1301 642 1367 645
rect 0 640 1367 642
rect 0 584 1306 640
rect 1362 584 1367 640
rect 0 582 1367 584
rect 0 552 480 582
rect 1301 579 1367 582
rect 20069 642 20135 645
rect 22520 642 23000 672
rect 20069 640 23000 642
rect 20069 584 20074 640
rect 20130 584 23000 640
rect 20069 582 23000 584
rect 20069 579 20135 582
rect 22520 552 23000 582
rect 0 234 480 264
rect 3601 234 3667 237
rect 0 232 3667 234
rect 0 176 3606 232
rect 3662 176 3667 232
rect 0 174 3667 176
rect 0 144 480 174
rect 3601 171 3667 174
rect 19241 234 19307 237
rect 22520 234 23000 264
rect 19241 232 23000 234
rect 19241 176 19246 232
rect 19302 176 23000 232
rect 19241 174 23000 176
rect 19241 171 19307 174
rect 22520 144 23000 174
<< via3 >>
rect 4417 20700 4481 20704
rect 4417 20644 4421 20700
rect 4421 20644 4477 20700
rect 4477 20644 4481 20700
rect 4417 20640 4481 20644
rect 4497 20700 4561 20704
rect 4497 20644 4501 20700
rect 4501 20644 4557 20700
rect 4557 20644 4561 20700
rect 4497 20640 4561 20644
rect 4577 20700 4641 20704
rect 4577 20644 4581 20700
rect 4581 20644 4637 20700
rect 4637 20644 4641 20700
rect 4577 20640 4641 20644
rect 4657 20700 4721 20704
rect 4657 20644 4661 20700
rect 4661 20644 4717 20700
rect 4717 20644 4721 20700
rect 4657 20640 4721 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 18278 20700 18342 20704
rect 18278 20644 18282 20700
rect 18282 20644 18338 20700
rect 18338 20644 18342 20700
rect 18278 20640 18342 20644
rect 18358 20700 18422 20704
rect 18358 20644 18362 20700
rect 18362 20644 18418 20700
rect 18418 20644 18422 20700
rect 18358 20640 18422 20644
rect 18438 20700 18502 20704
rect 18438 20644 18442 20700
rect 18442 20644 18498 20700
rect 18498 20644 18502 20700
rect 18438 20640 18502 20644
rect 18518 20700 18582 20704
rect 18518 20644 18522 20700
rect 18522 20644 18578 20700
rect 18578 20644 18582 20700
rect 18518 20640 18582 20644
rect 7882 20156 7946 20160
rect 7882 20100 7886 20156
rect 7886 20100 7942 20156
rect 7942 20100 7946 20156
rect 7882 20096 7946 20100
rect 7962 20156 8026 20160
rect 7962 20100 7966 20156
rect 7966 20100 8022 20156
rect 8022 20100 8026 20156
rect 7962 20096 8026 20100
rect 8042 20156 8106 20160
rect 8042 20100 8046 20156
rect 8046 20100 8102 20156
rect 8102 20100 8106 20156
rect 8042 20096 8106 20100
rect 8122 20156 8186 20160
rect 8122 20100 8126 20156
rect 8126 20100 8182 20156
rect 8182 20100 8186 20156
rect 8122 20096 8186 20100
rect 14813 20156 14877 20160
rect 14813 20100 14817 20156
rect 14817 20100 14873 20156
rect 14873 20100 14877 20156
rect 14813 20096 14877 20100
rect 14893 20156 14957 20160
rect 14893 20100 14897 20156
rect 14897 20100 14953 20156
rect 14953 20100 14957 20156
rect 14893 20096 14957 20100
rect 14973 20156 15037 20160
rect 14973 20100 14977 20156
rect 14977 20100 15033 20156
rect 15033 20100 15037 20156
rect 14973 20096 15037 20100
rect 15053 20156 15117 20160
rect 15053 20100 15057 20156
rect 15057 20100 15113 20156
rect 15113 20100 15117 20156
rect 15053 20096 15117 20100
rect 4417 19612 4481 19616
rect 4417 19556 4421 19612
rect 4421 19556 4477 19612
rect 4477 19556 4481 19612
rect 4417 19552 4481 19556
rect 4497 19612 4561 19616
rect 4497 19556 4501 19612
rect 4501 19556 4557 19612
rect 4557 19556 4561 19612
rect 4497 19552 4561 19556
rect 4577 19612 4641 19616
rect 4577 19556 4581 19612
rect 4581 19556 4637 19612
rect 4637 19556 4641 19612
rect 4577 19552 4641 19556
rect 4657 19612 4721 19616
rect 4657 19556 4661 19612
rect 4661 19556 4717 19612
rect 4717 19556 4721 19612
rect 4657 19552 4721 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 18278 19612 18342 19616
rect 18278 19556 18282 19612
rect 18282 19556 18338 19612
rect 18338 19556 18342 19612
rect 18278 19552 18342 19556
rect 18358 19612 18422 19616
rect 18358 19556 18362 19612
rect 18362 19556 18418 19612
rect 18418 19556 18422 19612
rect 18358 19552 18422 19556
rect 18438 19612 18502 19616
rect 18438 19556 18442 19612
rect 18442 19556 18498 19612
rect 18498 19556 18502 19612
rect 18438 19552 18502 19556
rect 18518 19612 18582 19616
rect 18518 19556 18522 19612
rect 18522 19556 18578 19612
rect 18578 19556 18582 19612
rect 18518 19552 18582 19556
rect 18828 19212 18892 19276
rect 7882 19068 7946 19072
rect 7882 19012 7886 19068
rect 7886 19012 7942 19068
rect 7942 19012 7946 19068
rect 7882 19008 7946 19012
rect 7962 19068 8026 19072
rect 7962 19012 7966 19068
rect 7966 19012 8022 19068
rect 8022 19012 8026 19068
rect 7962 19008 8026 19012
rect 8042 19068 8106 19072
rect 8042 19012 8046 19068
rect 8046 19012 8102 19068
rect 8102 19012 8106 19068
rect 8042 19008 8106 19012
rect 8122 19068 8186 19072
rect 8122 19012 8126 19068
rect 8126 19012 8182 19068
rect 8182 19012 8186 19068
rect 8122 19008 8186 19012
rect 14813 19068 14877 19072
rect 14813 19012 14817 19068
rect 14817 19012 14873 19068
rect 14873 19012 14877 19068
rect 14813 19008 14877 19012
rect 14893 19068 14957 19072
rect 14893 19012 14897 19068
rect 14897 19012 14953 19068
rect 14953 19012 14957 19068
rect 14893 19008 14957 19012
rect 14973 19068 15037 19072
rect 14973 19012 14977 19068
rect 14977 19012 15033 19068
rect 15033 19012 15037 19068
rect 14973 19008 15037 19012
rect 15053 19068 15117 19072
rect 15053 19012 15057 19068
rect 15057 19012 15113 19068
rect 15113 19012 15117 19068
rect 15053 19008 15117 19012
rect 4417 18524 4481 18528
rect 4417 18468 4421 18524
rect 4421 18468 4477 18524
rect 4477 18468 4481 18524
rect 4417 18464 4481 18468
rect 4497 18524 4561 18528
rect 4497 18468 4501 18524
rect 4501 18468 4557 18524
rect 4557 18468 4561 18524
rect 4497 18464 4561 18468
rect 4577 18524 4641 18528
rect 4577 18468 4581 18524
rect 4581 18468 4637 18524
rect 4637 18468 4641 18524
rect 4577 18464 4641 18468
rect 4657 18524 4721 18528
rect 4657 18468 4661 18524
rect 4661 18468 4717 18524
rect 4717 18468 4721 18524
rect 4657 18464 4721 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 18278 18524 18342 18528
rect 18278 18468 18282 18524
rect 18282 18468 18338 18524
rect 18338 18468 18342 18524
rect 18278 18464 18342 18468
rect 18358 18524 18422 18528
rect 18358 18468 18362 18524
rect 18362 18468 18418 18524
rect 18418 18468 18422 18524
rect 18358 18464 18422 18468
rect 18438 18524 18502 18528
rect 18438 18468 18442 18524
rect 18442 18468 18498 18524
rect 18498 18468 18502 18524
rect 18438 18464 18502 18468
rect 18518 18524 18582 18528
rect 18518 18468 18522 18524
rect 18522 18468 18578 18524
rect 18578 18468 18582 18524
rect 18518 18464 18582 18468
rect 18092 18456 18156 18460
rect 18092 18400 18106 18456
rect 18106 18400 18156 18456
rect 18092 18396 18156 18400
rect 17908 17988 17972 18052
rect 7882 17980 7946 17984
rect 7882 17924 7886 17980
rect 7886 17924 7942 17980
rect 7942 17924 7946 17980
rect 7882 17920 7946 17924
rect 7962 17980 8026 17984
rect 7962 17924 7966 17980
rect 7966 17924 8022 17980
rect 8022 17924 8026 17980
rect 7962 17920 8026 17924
rect 8042 17980 8106 17984
rect 8042 17924 8046 17980
rect 8046 17924 8102 17980
rect 8102 17924 8106 17980
rect 8042 17920 8106 17924
rect 8122 17980 8186 17984
rect 8122 17924 8126 17980
rect 8126 17924 8182 17980
rect 8182 17924 8186 17980
rect 8122 17920 8186 17924
rect 14813 17980 14877 17984
rect 14813 17924 14817 17980
rect 14817 17924 14873 17980
rect 14873 17924 14877 17980
rect 14813 17920 14877 17924
rect 14893 17980 14957 17984
rect 14893 17924 14897 17980
rect 14897 17924 14953 17980
rect 14953 17924 14957 17980
rect 14893 17920 14957 17924
rect 14973 17980 15037 17984
rect 14973 17924 14977 17980
rect 14977 17924 15033 17980
rect 15033 17924 15037 17980
rect 14973 17920 15037 17924
rect 15053 17980 15117 17984
rect 15053 17924 15057 17980
rect 15057 17924 15113 17980
rect 15113 17924 15117 17980
rect 15053 17920 15117 17924
rect 17540 17852 17604 17916
rect 4417 17436 4481 17440
rect 4417 17380 4421 17436
rect 4421 17380 4477 17436
rect 4477 17380 4481 17436
rect 4417 17376 4481 17380
rect 4497 17436 4561 17440
rect 4497 17380 4501 17436
rect 4501 17380 4557 17436
rect 4557 17380 4561 17436
rect 4497 17376 4561 17380
rect 4577 17436 4641 17440
rect 4577 17380 4581 17436
rect 4581 17380 4637 17436
rect 4637 17380 4641 17436
rect 4577 17376 4641 17380
rect 4657 17436 4721 17440
rect 4657 17380 4661 17436
rect 4661 17380 4717 17436
rect 4717 17380 4721 17436
rect 4657 17376 4721 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 18278 17436 18342 17440
rect 18278 17380 18282 17436
rect 18282 17380 18338 17436
rect 18338 17380 18342 17436
rect 18278 17376 18342 17380
rect 18358 17436 18422 17440
rect 18358 17380 18362 17436
rect 18362 17380 18418 17436
rect 18418 17380 18422 17436
rect 18358 17376 18422 17380
rect 18438 17436 18502 17440
rect 18438 17380 18442 17436
rect 18442 17380 18498 17436
rect 18498 17380 18502 17436
rect 18438 17376 18502 17380
rect 18518 17436 18582 17440
rect 18518 17380 18522 17436
rect 18522 17380 18578 17436
rect 18578 17380 18582 17436
rect 18518 17376 18582 17380
rect 7882 16892 7946 16896
rect 7882 16836 7886 16892
rect 7886 16836 7942 16892
rect 7942 16836 7946 16892
rect 7882 16832 7946 16836
rect 7962 16892 8026 16896
rect 7962 16836 7966 16892
rect 7966 16836 8022 16892
rect 8022 16836 8026 16892
rect 7962 16832 8026 16836
rect 8042 16892 8106 16896
rect 8042 16836 8046 16892
rect 8046 16836 8102 16892
rect 8102 16836 8106 16892
rect 8042 16832 8106 16836
rect 8122 16892 8186 16896
rect 8122 16836 8126 16892
rect 8126 16836 8182 16892
rect 8182 16836 8186 16892
rect 8122 16832 8186 16836
rect 14813 16892 14877 16896
rect 14813 16836 14817 16892
rect 14817 16836 14873 16892
rect 14873 16836 14877 16892
rect 14813 16832 14877 16836
rect 14893 16892 14957 16896
rect 14893 16836 14897 16892
rect 14897 16836 14953 16892
rect 14953 16836 14957 16892
rect 14893 16832 14957 16836
rect 14973 16892 15037 16896
rect 14973 16836 14977 16892
rect 14977 16836 15033 16892
rect 15033 16836 15037 16892
rect 14973 16832 15037 16836
rect 15053 16892 15117 16896
rect 15053 16836 15057 16892
rect 15057 16836 15113 16892
rect 15113 16836 15117 16892
rect 15053 16832 15117 16836
rect 18828 16628 18892 16692
rect 4417 16348 4481 16352
rect 4417 16292 4421 16348
rect 4421 16292 4477 16348
rect 4477 16292 4481 16348
rect 4417 16288 4481 16292
rect 4497 16348 4561 16352
rect 4497 16292 4501 16348
rect 4501 16292 4557 16348
rect 4557 16292 4561 16348
rect 4497 16288 4561 16292
rect 4577 16348 4641 16352
rect 4577 16292 4581 16348
rect 4581 16292 4637 16348
rect 4637 16292 4641 16348
rect 4577 16288 4641 16292
rect 4657 16348 4721 16352
rect 4657 16292 4661 16348
rect 4661 16292 4717 16348
rect 4717 16292 4721 16348
rect 4657 16288 4721 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 18278 16348 18342 16352
rect 18278 16292 18282 16348
rect 18282 16292 18338 16348
rect 18338 16292 18342 16348
rect 18278 16288 18342 16292
rect 18358 16348 18422 16352
rect 18358 16292 18362 16348
rect 18362 16292 18418 16348
rect 18418 16292 18422 16348
rect 18358 16288 18422 16292
rect 18438 16348 18502 16352
rect 18438 16292 18442 16348
rect 18442 16292 18498 16348
rect 18498 16292 18502 16348
rect 18438 16288 18502 16292
rect 18518 16348 18582 16352
rect 18518 16292 18522 16348
rect 18522 16292 18578 16348
rect 18578 16292 18582 16348
rect 18518 16288 18582 16292
rect 7882 15804 7946 15808
rect 7882 15748 7886 15804
rect 7886 15748 7942 15804
rect 7942 15748 7946 15804
rect 7882 15744 7946 15748
rect 7962 15804 8026 15808
rect 7962 15748 7966 15804
rect 7966 15748 8022 15804
rect 8022 15748 8026 15804
rect 7962 15744 8026 15748
rect 8042 15804 8106 15808
rect 8042 15748 8046 15804
rect 8046 15748 8102 15804
rect 8102 15748 8106 15804
rect 8042 15744 8106 15748
rect 8122 15804 8186 15808
rect 8122 15748 8126 15804
rect 8126 15748 8182 15804
rect 8182 15748 8186 15804
rect 8122 15744 8186 15748
rect 14813 15804 14877 15808
rect 14813 15748 14817 15804
rect 14817 15748 14873 15804
rect 14873 15748 14877 15804
rect 14813 15744 14877 15748
rect 14893 15804 14957 15808
rect 14893 15748 14897 15804
rect 14897 15748 14953 15804
rect 14953 15748 14957 15804
rect 14893 15744 14957 15748
rect 14973 15804 15037 15808
rect 14973 15748 14977 15804
rect 14977 15748 15033 15804
rect 15033 15748 15037 15804
rect 14973 15744 15037 15748
rect 15053 15804 15117 15808
rect 15053 15748 15057 15804
rect 15057 15748 15113 15804
rect 15113 15748 15117 15804
rect 15053 15744 15117 15748
rect 4417 15260 4481 15264
rect 4417 15204 4421 15260
rect 4421 15204 4477 15260
rect 4477 15204 4481 15260
rect 4417 15200 4481 15204
rect 4497 15260 4561 15264
rect 4497 15204 4501 15260
rect 4501 15204 4557 15260
rect 4557 15204 4561 15260
rect 4497 15200 4561 15204
rect 4577 15260 4641 15264
rect 4577 15204 4581 15260
rect 4581 15204 4637 15260
rect 4637 15204 4641 15260
rect 4577 15200 4641 15204
rect 4657 15260 4721 15264
rect 4657 15204 4661 15260
rect 4661 15204 4717 15260
rect 4717 15204 4721 15260
rect 4657 15200 4721 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 18278 15260 18342 15264
rect 18278 15204 18282 15260
rect 18282 15204 18338 15260
rect 18338 15204 18342 15260
rect 18278 15200 18342 15204
rect 18358 15260 18422 15264
rect 18358 15204 18362 15260
rect 18362 15204 18418 15260
rect 18418 15204 18422 15260
rect 18358 15200 18422 15204
rect 18438 15260 18502 15264
rect 18438 15204 18442 15260
rect 18442 15204 18498 15260
rect 18498 15204 18502 15260
rect 18438 15200 18502 15204
rect 18518 15260 18582 15264
rect 18518 15204 18522 15260
rect 18522 15204 18578 15260
rect 18578 15204 18582 15260
rect 18518 15200 18582 15204
rect 7882 14716 7946 14720
rect 7882 14660 7886 14716
rect 7886 14660 7942 14716
rect 7942 14660 7946 14716
rect 7882 14656 7946 14660
rect 7962 14716 8026 14720
rect 7962 14660 7966 14716
rect 7966 14660 8022 14716
rect 8022 14660 8026 14716
rect 7962 14656 8026 14660
rect 8042 14716 8106 14720
rect 8042 14660 8046 14716
rect 8046 14660 8102 14716
rect 8102 14660 8106 14716
rect 8042 14656 8106 14660
rect 8122 14716 8186 14720
rect 8122 14660 8126 14716
rect 8126 14660 8182 14716
rect 8182 14660 8186 14716
rect 8122 14656 8186 14660
rect 14813 14716 14877 14720
rect 14813 14660 14817 14716
rect 14817 14660 14873 14716
rect 14873 14660 14877 14716
rect 14813 14656 14877 14660
rect 14893 14716 14957 14720
rect 14893 14660 14897 14716
rect 14897 14660 14953 14716
rect 14953 14660 14957 14716
rect 14893 14656 14957 14660
rect 14973 14716 15037 14720
rect 14973 14660 14977 14716
rect 14977 14660 15033 14716
rect 15033 14660 15037 14716
rect 14973 14656 15037 14660
rect 15053 14716 15117 14720
rect 15053 14660 15057 14716
rect 15057 14660 15113 14716
rect 15113 14660 15117 14716
rect 15053 14656 15117 14660
rect 4417 14172 4481 14176
rect 4417 14116 4421 14172
rect 4421 14116 4477 14172
rect 4477 14116 4481 14172
rect 4417 14112 4481 14116
rect 4497 14172 4561 14176
rect 4497 14116 4501 14172
rect 4501 14116 4557 14172
rect 4557 14116 4561 14172
rect 4497 14112 4561 14116
rect 4577 14172 4641 14176
rect 4577 14116 4581 14172
rect 4581 14116 4637 14172
rect 4637 14116 4641 14172
rect 4577 14112 4641 14116
rect 4657 14172 4721 14176
rect 4657 14116 4661 14172
rect 4661 14116 4717 14172
rect 4717 14116 4721 14172
rect 4657 14112 4721 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 18278 14172 18342 14176
rect 18278 14116 18282 14172
rect 18282 14116 18338 14172
rect 18338 14116 18342 14172
rect 18278 14112 18342 14116
rect 18358 14172 18422 14176
rect 18358 14116 18362 14172
rect 18362 14116 18418 14172
rect 18418 14116 18422 14172
rect 18358 14112 18422 14116
rect 18438 14172 18502 14176
rect 18438 14116 18442 14172
rect 18442 14116 18498 14172
rect 18498 14116 18502 14172
rect 18438 14112 18502 14116
rect 18518 14172 18582 14176
rect 18518 14116 18522 14172
rect 18522 14116 18578 14172
rect 18578 14116 18582 14172
rect 18518 14112 18582 14116
rect 7882 13628 7946 13632
rect 7882 13572 7886 13628
rect 7886 13572 7942 13628
rect 7942 13572 7946 13628
rect 7882 13568 7946 13572
rect 7962 13628 8026 13632
rect 7962 13572 7966 13628
rect 7966 13572 8022 13628
rect 8022 13572 8026 13628
rect 7962 13568 8026 13572
rect 8042 13628 8106 13632
rect 8042 13572 8046 13628
rect 8046 13572 8102 13628
rect 8102 13572 8106 13628
rect 8042 13568 8106 13572
rect 8122 13628 8186 13632
rect 8122 13572 8126 13628
rect 8126 13572 8182 13628
rect 8182 13572 8186 13628
rect 8122 13568 8186 13572
rect 14813 13628 14877 13632
rect 14813 13572 14817 13628
rect 14817 13572 14873 13628
rect 14873 13572 14877 13628
rect 14813 13568 14877 13572
rect 14893 13628 14957 13632
rect 14893 13572 14897 13628
rect 14897 13572 14953 13628
rect 14953 13572 14957 13628
rect 14893 13568 14957 13572
rect 14973 13628 15037 13632
rect 14973 13572 14977 13628
rect 14977 13572 15033 13628
rect 15033 13572 15037 13628
rect 14973 13568 15037 13572
rect 15053 13628 15117 13632
rect 15053 13572 15057 13628
rect 15057 13572 15113 13628
rect 15113 13572 15117 13628
rect 15053 13568 15117 13572
rect 17724 13364 17788 13428
rect 4417 13084 4481 13088
rect 4417 13028 4421 13084
rect 4421 13028 4477 13084
rect 4477 13028 4481 13084
rect 4417 13024 4481 13028
rect 4497 13084 4561 13088
rect 4497 13028 4501 13084
rect 4501 13028 4557 13084
rect 4557 13028 4561 13084
rect 4497 13024 4561 13028
rect 4577 13084 4641 13088
rect 4577 13028 4581 13084
rect 4581 13028 4637 13084
rect 4637 13028 4641 13084
rect 4577 13024 4641 13028
rect 4657 13084 4721 13088
rect 4657 13028 4661 13084
rect 4661 13028 4717 13084
rect 4717 13028 4721 13084
rect 4657 13024 4721 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 18278 13084 18342 13088
rect 18278 13028 18282 13084
rect 18282 13028 18338 13084
rect 18338 13028 18342 13084
rect 18278 13024 18342 13028
rect 18358 13084 18422 13088
rect 18358 13028 18362 13084
rect 18362 13028 18418 13084
rect 18418 13028 18422 13084
rect 18358 13024 18422 13028
rect 18438 13084 18502 13088
rect 18438 13028 18442 13084
rect 18442 13028 18498 13084
rect 18498 13028 18502 13084
rect 18438 13024 18502 13028
rect 18518 13084 18582 13088
rect 18518 13028 18522 13084
rect 18522 13028 18578 13084
rect 18578 13028 18582 13084
rect 18518 13024 18582 13028
rect 7882 12540 7946 12544
rect 7882 12484 7886 12540
rect 7886 12484 7942 12540
rect 7942 12484 7946 12540
rect 7882 12480 7946 12484
rect 7962 12540 8026 12544
rect 7962 12484 7966 12540
rect 7966 12484 8022 12540
rect 8022 12484 8026 12540
rect 7962 12480 8026 12484
rect 8042 12540 8106 12544
rect 8042 12484 8046 12540
rect 8046 12484 8102 12540
rect 8102 12484 8106 12540
rect 8042 12480 8106 12484
rect 8122 12540 8186 12544
rect 8122 12484 8126 12540
rect 8126 12484 8182 12540
rect 8182 12484 8186 12540
rect 8122 12480 8186 12484
rect 14813 12540 14877 12544
rect 14813 12484 14817 12540
rect 14817 12484 14873 12540
rect 14873 12484 14877 12540
rect 14813 12480 14877 12484
rect 14893 12540 14957 12544
rect 14893 12484 14897 12540
rect 14897 12484 14953 12540
rect 14953 12484 14957 12540
rect 14893 12480 14957 12484
rect 14973 12540 15037 12544
rect 14973 12484 14977 12540
rect 14977 12484 15033 12540
rect 15033 12484 15037 12540
rect 14973 12480 15037 12484
rect 15053 12540 15117 12544
rect 15053 12484 15057 12540
rect 15057 12484 15113 12540
rect 15113 12484 15117 12540
rect 15053 12480 15117 12484
rect 4417 11996 4481 12000
rect 4417 11940 4421 11996
rect 4421 11940 4477 11996
rect 4477 11940 4481 11996
rect 4417 11936 4481 11940
rect 4497 11996 4561 12000
rect 4497 11940 4501 11996
rect 4501 11940 4557 11996
rect 4557 11940 4561 11996
rect 4497 11936 4561 11940
rect 4577 11996 4641 12000
rect 4577 11940 4581 11996
rect 4581 11940 4637 11996
rect 4637 11940 4641 11996
rect 4577 11936 4641 11940
rect 4657 11996 4721 12000
rect 4657 11940 4661 11996
rect 4661 11940 4717 11996
rect 4717 11940 4721 11996
rect 4657 11936 4721 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 18278 11996 18342 12000
rect 18278 11940 18282 11996
rect 18282 11940 18338 11996
rect 18338 11940 18342 11996
rect 18278 11936 18342 11940
rect 18358 11996 18422 12000
rect 18358 11940 18362 11996
rect 18362 11940 18418 11996
rect 18418 11940 18422 11996
rect 18358 11936 18422 11940
rect 18438 11996 18502 12000
rect 18438 11940 18442 11996
rect 18442 11940 18498 11996
rect 18498 11940 18502 11996
rect 18438 11936 18502 11940
rect 18518 11996 18582 12000
rect 18518 11940 18522 11996
rect 18522 11940 18578 11996
rect 18578 11940 18582 11996
rect 18518 11936 18582 11940
rect 7882 11452 7946 11456
rect 7882 11396 7886 11452
rect 7886 11396 7942 11452
rect 7942 11396 7946 11452
rect 7882 11392 7946 11396
rect 7962 11452 8026 11456
rect 7962 11396 7966 11452
rect 7966 11396 8022 11452
rect 8022 11396 8026 11452
rect 7962 11392 8026 11396
rect 8042 11452 8106 11456
rect 8042 11396 8046 11452
rect 8046 11396 8102 11452
rect 8102 11396 8106 11452
rect 8042 11392 8106 11396
rect 8122 11452 8186 11456
rect 8122 11396 8126 11452
rect 8126 11396 8182 11452
rect 8182 11396 8186 11452
rect 8122 11392 8186 11396
rect 14813 11452 14877 11456
rect 14813 11396 14817 11452
rect 14817 11396 14873 11452
rect 14873 11396 14877 11452
rect 14813 11392 14877 11396
rect 14893 11452 14957 11456
rect 14893 11396 14897 11452
rect 14897 11396 14953 11452
rect 14953 11396 14957 11452
rect 14893 11392 14957 11396
rect 14973 11452 15037 11456
rect 14973 11396 14977 11452
rect 14977 11396 15033 11452
rect 15033 11396 15037 11452
rect 14973 11392 15037 11396
rect 15053 11452 15117 11456
rect 15053 11396 15057 11452
rect 15057 11396 15113 11452
rect 15113 11396 15117 11452
rect 15053 11392 15117 11396
rect 17724 11324 17788 11388
rect 4417 10908 4481 10912
rect 4417 10852 4421 10908
rect 4421 10852 4477 10908
rect 4477 10852 4481 10908
rect 4417 10848 4481 10852
rect 4497 10908 4561 10912
rect 4497 10852 4501 10908
rect 4501 10852 4557 10908
rect 4557 10852 4561 10908
rect 4497 10848 4561 10852
rect 4577 10908 4641 10912
rect 4577 10852 4581 10908
rect 4581 10852 4637 10908
rect 4637 10852 4641 10908
rect 4577 10848 4641 10852
rect 4657 10908 4721 10912
rect 4657 10852 4661 10908
rect 4661 10852 4717 10908
rect 4717 10852 4721 10908
rect 4657 10848 4721 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 18278 10908 18342 10912
rect 18278 10852 18282 10908
rect 18282 10852 18338 10908
rect 18338 10852 18342 10908
rect 18278 10848 18342 10852
rect 18358 10908 18422 10912
rect 18358 10852 18362 10908
rect 18362 10852 18418 10908
rect 18418 10852 18422 10908
rect 18358 10848 18422 10852
rect 18438 10908 18502 10912
rect 18438 10852 18442 10908
rect 18442 10852 18498 10908
rect 18498 10852 18502 10908
rect 18438 10848 18502 10852
rect 18518 10908 18582 10912
rect 18518 10852 18522 10908
rect 18522 10852 18578 10908
rect 18578 10852 18582 10908
rect 18518 10848 18582 10852
rect 18828 10704 18892 10708
rect 18828 10648 18878 10704
rect 18878 10648 18892 10704
rect 18828 10644 18892 10648
rect 7882 10364 7946 10368
rect 7882 10308 7886 10364
rect 7886 10308 7942 10364
rect 7942 10308 7946 10364
rect 7882 10304 7946 10308
rect 7962 10364 8026 10368
rect 7962 10308 7966 10364
rect 7966 10308 8022 10364
rect 8022 10308 8026 10364
rect 7962 10304 8026 10308
rect 8042 10364 8106 10368
rect 8042 10308 8046 10364
rect 8046 10308 8102 10364
rect 8102 10308 8106 10364
rect 8042 10304 8106 10308
rect 8122 10364 8186 10368
rect 8122 10308 8126 10364
rect 8126 10308 8182 10364
rect 8182 10308 8186 10364
rect 8122 10304 8186 10308
rect 14813 10364 14877 10368
rect 14813 10308 14817 10364
rect 14817 10308 14873 10364
rect 14873 10308 14877 10364
rect 14813 10304 14877 10308
rect 14893 10364 14957 10368
rect 14893 10308 14897 10364
rect 14897 10308 14953 10364
rect 14953 10308 14957 10364
rect 14893 10304 14957 10308
rect 14973 10364 15037 10368
rect 14973 10308 14977 10364
rect 14977 10308 15033 10364
rect 15033 10308 15037 10364
rect 14973 10304 15037 10308
rect 15053 10364 15117 10368
rect 15053 10308 15057 10364
rect 15057 10308 15113 10364
rect 15113 10308 15117 10364
rect 15053 10304 15117 10308
rect 17540 10100 17604 10164
rect 4417 9820 4481 9824
rect 4417 9764 4421 9820
rect 4421 9764 4477 9820
rect 4477 9764 4481 9820
rect 4417 9760 4481 9764
rect 4497 9820 4561 9824
rect 4497 9764 4501 9820
rect 4501 9764 4557 9820
rect 4557 9764 4561 9820
rect 4497 9760 4561 9764
rect 4577 9820 4641 9824
rect 4577 9764 4581 9820
rect 4581 9764 4637 9820
rect 4637 9764 4641 9820
rect 4577 9760 4641 9764
rect 4657 9820 4721 9824
rect 4657 9764 4661 9820
rect 4661 9764 4717 9820
rect 4717 9764 4721 9820
rect 4657 9760 4721 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 18278 9820 18342 9824
rect 18278 9764 18282 9820
rect 18282 9764 18338 9820
rect 18338 9764 18342 9820
rect 18278 9760 18342 9764
rect 18358 9820 18422 9824
rect 18358 9764 18362 9820
rect 18362 9764 18418 9820
rect 18418 9764 18422 9820
rect 18358 9760 18422 9764
rect 18438 9820 18502 9824
rect 18438 9764 18442 9820
rect 18442 9764 18498 9820
rect 18498 9764 18502 9820
rect 18438 9760 18502 9764
rect 18518 9820 18582 9824
rect 18518 9764 18522 9820
rect 18522 9764 18578 9820
rect 18578 9764 18582 9820
rect 18518 9760 18582 9764
rect 11100 9556 11164 9620
rect 19012 9284 19076 9348
rect 7882 9276 7946 9280
rect 7882 9220 7886 9276
rect 7886 9220 7942 9276
rect 7942 9220 7946 9276
rect 7882 9216 7946 9220
rect 7962 9276 8026 9280
rect 7962 9220 7966 9276
rect 7966 9220 8022 9276
rect 8022 9220 8026 9276
rect 7962 9216 8026 9220
rect 8042 9276 8106 9280
rect 8042 9220 8046 9276
rect 8046 9220 8102 9276
rect 8102 9220 8106 9276
rect 8042 9216 8106 9220
rect 8122 9276 8186 9280
rect 8122 9220 8126 9276
rect 8126 9220 8182 9276
rect 8182 9220 8186 9276
rect 8122 9216 8186 9220
rect 14813 9276 14877 9280
rect 14813 9220 14817 9276
rect 14817 9220 14873 9276
rect 14873 9220 14877 9276
rect 14813 9216 14877 9220
rect 14893 9276 14957 9280
rect 14893 9220 14897 9276
rect 14897 9220 14953 9276
rect 14953 9220 14957 9276
rect 14893 9216 14957 9220
rect 14973 9276 15037 9280
rect 14973 9220 14977 9276
rect 14977 9220 15033 9276
rect 15033 9220 15037 9276
rect 14973 9216 15037 9220
rect 15053 9276 15117 9280
rect 15053 9220 15057 9276
rect 15057 9220 15113 9276
rect 15113 9220 15117 9276
rect 15053 9216 15117 9220
rect 11836 9208 11900 9212
rect 11836 9152 11850 9208
rect 11850 9152 11900 9208
rect 11836 9148 11900 9152
rect 18828 9072 18892 9076
rect 18828 9016 18842 9072
rect 18842 9016 18892 9072
rect 18828 9012 18892 9016
rect 4417 8732 4481 8736
rect 4417 8676 4421 8732
rect 4421 8676 4477 8732
rect 4477 8676 4481 8732
rect 4417 8672 4481 8676
rect 4497 8732 4561 8736
rect 4497 8676 4501 8732
rect 4501 8676 4557 8732
rect 4557 8676 4561 8732
rect 4497 8672 4561 8676
rect 4577 8732 4641 8736
rect 4577 8676 4581 8732
rect 4581 8676 4637 8732
rect 4637 8676 4641 8732
rect 4577 8672 4641 8676
rect 4657 8732 4721 8736
rect 4657 8676 4661 8732
rect 4661 8676 4717 8732
rect 4717 8676 4721 8732
rect 4657 8672 4721 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 18278 8732 18342 8736
rect 18278 8676 18282 8732
rect 18282 8676 18338 8732
rect 18338 8676 18342 8732
rect 18278 8672 18342 8676
rect 18358 8732 18422 8736
rect 18358 8676 18362 8732
rect 18362 8676 18418 8732
rect 18418 8676 18422 8732
rect 18358 8672 18422 8676
rect 18438 8732 18502 8736
rect 18438 8676 18442 8732
rect 18442 8676 18498 8732
rect 18498 8676 18502 8732
rect 18438 8672 18502 8676
rect 18518 8732 18582 8736
rect 18518 8676 18522 8732
rect 18522 8676 18578 8732
rect 18578 8676 18582 8732
rect 18518 8672 18582 8676
rect 7882 8188 7946 8192
rect 7882 8132 7886 8188
rect 7886 8132 7942 8188
rect 7942 8132 7946 8188
rect 7882 8128 7946 8132
rect 7962 8188 8026 8192
rect 7962 8132 7966 8188
rect 7966 8132 8022 8188
rect 8022 8132 8026 8188
rect 7962 8128 8026 8132
rect 8042 8188 8106 8192
rect 8042 8132 8046 8188
rect 8046 8132 8102 8188
rect 8102 8132 8106 8188
rect 8042 8128 8106 8132
rect 8122 8188 8186 8192
rect 8122 8132 8126 8188
rect 8126 8132 8182 8188
rect 8182 8132 8186 8188
rect 8122 8128 8186 8132
rect 14813 8188 14877 8192
rect 14813 8132 14817 8188
rect 14817 8132 14873 8188
rect 14873 8132 14877 8188
rect 14813 8128 14877 8132
rect 14893 8188 14957 8192
rect 14893 8132 14897 8188
rect 14897 8132 14953 8188
rect 14953 8132 14957 8188
rect 14893 8128 14957 8132
rect 14973 8188 15037 8192
rect 14973 8132 14977 8188
rect 14977 8132 15033 8188
rect 15033 8132 15037 8188
rect 14973 8128 15037 8132
rect 15053 8188 15117 8192
rect 15053 8132 15057 8188
rect 15057 8132 15113 8188
rect 15113 8132 15117 8188
rect 15053 8128 15117 8132
rect 19012 8060 19076 8124
rect 4417 7644 4481 7648
rect 4417 7588 4421 7644
rect 4421 7588 4477 7644
rect 4477 7588 4481 7644
rect 4417 7584 4481 7588
rect 4497 7644 4561 7648
rect 4497 7588 4501 7644
rect 4501 7588 4557 7644
rect 4557 7588 4561 7644
rect 4497 7584 4561 7588
rect 4577 7644 4641 7648
rect 4577 7588 4581 7644
rect 4581 7588 4637 7644
rect 4637 7588 4641 7644
rect 4577 7584 4641 7588
rect 4657 7644 4721 7648
rect 4657 7588 4661 7644
rect 4661 7588 4717 7644
rect 4717 7588 4721 7644
rect 4657 7584 4721 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 18278 7644 18342 7648
rect 18278 7588 18282 7644
rect 18282 7588 18338 7644
rect 18338 7588 18342 7644
rect 18278 7584 18342 7588
rect 18358 7644 18422 7648
rect 18358 7588 18362 7644
rect 18362 7588 18418 7644
rect 18418 7588 18422 7644
rect 18358 7584 18422 7588
rect 18438 7644 18502 7648
rect 18438 7588 18442 7644
rect 18442 7588 18498 7644
rect 18498 7588 18502 7644
rect 18438 7584 18502 7588
rect 18518 7644 18582 7648
rect 18518 7588 18522 7644
rect 18522 7588 18578 7644
rect 18578 7588 18582 7644
rect 18518 7584 18582 7588
rect 7882 7100 7946 7104
rect 7882 7044 7886 7100
rect 7886 7044 7942 7100
rect 7942 7044 7946 7100
rect 7882 7040 7946 7044
rect 7962 7100 8026 7104
rect 7962 7044 7966 7100
rect 7966 7044 8022 7100
rect 8022 7044 8026 7100
rect 7962 7040 8026 7044
rect 8042 7100 8106 7104
rect 8042 7044 8046 7100
rect 8046 7044 8102 7100
rect 8102 7044 8106 7100
rect 8042 7040 8106 7044
rect 8122 7100 8186 7104
rect 8122 7044 8126 7100
rect 8126 7044 8182 7100
rect 8182 7044 8186 7100
rect 8122 7040 8186 7044
rect 14813 7100 14877 7104
rect 14813 7044 14817 7100
rect 14817 7044 14873 7100
rect 14873 7044 14877 7100
rect 14813 7040 14877 7044
rect 14893 7100 14957 7104
rect 14893 7044 14897 7100
rect 14897 7044 14953 7100
rect 14953 7044 14957 7100
rect 14893 7040 14957 7044
rect 14973 7100 15037 7104
rect 14973 7044 14977 7100
rect 14977 7044 15033 7100
rect 15033 7044 15037 7100
rect 14973 7040 15037 7044
rect 15053 7100 15117 7104
rect 15053 7044 15057 7100
rect 15057 7044 15113 7100
rect 15113 7044 15117 7100
rect 15053 7040 15117 7044
rect 3004 6700 3068 6764
rect 4417 6556 4481 6560
rect 4417 6500 4421 6556
rect 4421 6500 4477 6556
rect 4477 6500 4481 6556
rect 4417 6496 4481 6500
rect 4497 6556 4561 6560
rect 4497 6500 4501 6556
rect 4501 6500 4557 6556
rect 4557 6500 4561 6556
rect 4497 6496 4561 6500
rect 4577 6556 4641 6560
rect 4577 6500 4581 6556
rect 4581 6500 4637 6556
rect 4637 6500 4641 6556
rect 4577 6496 4641 6500
rect 4657 6556 4721 6560
rect 4657 6500 4661 6556
rect 4661 6500 4717 6556
rect 4717 6500 4721 6556
rect 4657 6496 4721 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 18278 6556 18342 6560
rect 18278 6500 18282 6556
rect 18282 6500 18338 6556
rect 18338 6500 18342 6556
rect 18278 6496 18342 6500
rect 18358 6556 18422 6560
rect 18358 6500 18362 6556
rect 18362 6500 18418 6556
rect 18418 6500 18422 6556
rect 18358 6496 18422 6500
rect 18438 6556 18502 6560
rect 18438 6500 18442 6556
rect 18442 6500 18498 6556
rect 18498 6500 18502 6556
rect 18438 6496 18502 6500
rect 18518 6556 18582 6560
rect 18518 6500 18522 6556
rect 18522 6500 18578 6556
rect 18578 6500 18582 6556
rect 18518 6496 18582 6500
rect 7882 6012 7946 6016
rect 7882 5956 7886 6012
rect 7886 5956 7942 6012
rect 7942 5956 7946 6012
rect 7882 5952 7946 5956
rect 7962 6012 8026 6016
rect 7962 5956 7966 6012
rect 7966 5956 8022 6012
rect 8022 5956 8026 6012
rect 7962 5952 8026 5956
rect 8042 6012 8106 6016
rect 8042 5956 8046 6012
rect 8046 5956 8102 6012
rect 8102 5956 8106 6012
rect 8042 5952 8106 5956
rect 8122 6012 8186 6016
rect 8122 5956 8126 6012
rect 8126 5956 8182 6012
rect 8182 5956 8186 6012
rect 8122 5952 8186 5956
rect 14813 6012 14877 6016
rect 14813 5956 14817 6012
rect 14817 5956 14873 6012
rect 14873 5956 14877 6012
rect 14813 5952 14877 5956
rect 14893 6012 14957 6016
rect 14893 5956 14897 6012
rect 14897 5956 14953 6012
rect 14953 5956 14957 6012
rect 14893 5952 14957 5956
rect 14973 6012 15037 6016
rect 14973 5956 14977 6012
rect 14977 5956 15033 6012
rect 15033 5956 15037 6012
rect 14973 5952 15037 5956
rect 15053 6012 15117 6016
rect 15053 5956 15057 6012
rect 15057 5956 15113 6012
rect 15113 5956 15117 6012
rect 15053 5952 15117 5956
rect 9812 5536 9876 5540
rect 9812 5480 9862 5536
rect 9862 5480 9876 5536
rect 9812 5476 9876 5480
rect 4417 5468 4481 5472
rect 4417 5412 4421 5468
rect 4421 5412 4477 5468
rect 4477 5412 4481 5468
rect 4417 5408 4481 5412
rect 4497 5468 4561 5472
rect 4497 5412 4501 5468
rect 4501 5412 4557 5468
rect 4557 5412 4561 5468
rect 4497 5408 4561 5412
rect 4577 5468 4641 5472
rect 4577 5412 4581 5468
rect 4581 5412 4637 5468
rect 4637 5412 4641 5468
rect 4577 5408 4641 5412
rect 4657 5468 4721 5472
rect 4657 5412 4661 5468
rect 4661 5412 4717 5468
rect 4717 5412 4721 5468
rect 4657 5408 4721 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 18278 5468 18342 5472
rect 18278 5412 18282 5468
rect 18282 5412 18338 5468
rect 18338 5412 18342 5468
rect 18278 5408 18342 5412
rect 18358 5468 18422 5472
rect 18358 5412 18362 5468
rect 18362 5412 18418 5468
rect 18418 5412 18422 5468
rect 18358 5408 18422 5412
rect 18438 5468 18502 5472
rect 18438 5412 18442 5468
rect 18442 5412 18498 5468
rect 18498 5412 18502 5468
rect 18438 5408 18502 5412
rect 18518 5468 18582 5472
rect 18518 5412 18522 5468
rect 18522 5412 18578 5468
rect 18578 5412 18582 5468
rect 18518 5408 18582 5412
rect 7882 4924 7946 4928
rect 7882 4868 7886 4924
rect 7886 4868 7942 4924
rect 7942 4868 7946 4924
rect 7882 4864 7946 4868
rect 7962 4924 8026 4928
rect 7962 4868 7966 4924
rect 7966 4868 8022 4924
rect 8022 4868 8026 4924
rect 7962 4864 8026 4868
rect 8042 4924 8106 4928
rect 8042 4868 8046 4924
rect 8046 4868 8102 4924
rect 8102 4868 8106 4924
rect 8042 4864 8106 4868
rect 8122 4924 8186 4928
rect 8122 4868 8126 4924
rect 8126 4868 8182 4924
rect 8182 4868 8186 4924
rect 8122 4864 8186 4868
rect 14813 4924 14877 4928
rect 14813 4868 14817 4924
rect 14817 4868 14873 4924
rect 14873 4868 14877 4924
rect 14813 4864 14877 4868
rect 14893 4924 14957 4928
rect 14893 4868 14897 4924
rect 14897 4868 14953 4924
rect 14953 4868 14957 4924
rect 14893 4864 14957 4868
rect 14973 4924 15037 4928
rect 14973 4868 14977 4924
rect 14977 4868 15033 4924
rect 15033 4868 15037 4924
rect 14973 4864 15037 4868
rect 15053 4924 15117 4928
rect 15053 4868 15057 4924
rect 15057 4868 15113 4924
rect 15113 4868 15117 4924
rect 15053 4864 15117 4868
rect 8340 4490 8404 4554
rect 11836 4388 11900 4452
rect 4417 4380 4481 4384
rect 4417 4324 4421 4380
rect 4421 4324 4477 4380
rect 4477 4324 4481 4380
rect 4417 4320 4481 4324
rect 4497 4380 4561 4384
rect 4497 4324 4501 4380
rect 4501 4324 4557 4380
rect 4557 4324 4561 4380
rect 4497 4320 4561 4324
rect 4577 4380 4641 4384
rect 4577 4324 4581 4380
rect 4581 4324 4637 4380
rect 4637 4324 4641 4380
rect 4577 4320 4641 4324
rect 4657 4380 4721 4384
rect 4657 4324 4661 4380
rect 4661 4324 4717 4380
rect 4717 4324 4721 4380
rect 4657 4320 4721 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 18278 4380 18342 4384
rect 18278 4324 18282 4380
rect 18282 4324 18338 4380
rect 18338 4324 18342 4380
rect 18278 4320 18342 4324
rect 18358 4380 18422 4384
rect 18358 4324 18362 4380
rect 18362 4324 18418 4380
rect 18418 4324 18422 4380
rect 18358 4320 18422 4324
rect 18438 4380 18502 4384
rect 18438 4324 18442 4380
rect 18442 4324 18498 4380
rect 18498 4324 18502 4380
rect 18438 4320 18502 4324
rect 18518 4380 18582 4384
rect 18518 4324 18522 4380
rect 18522 4324 18578 4380
rect 18578 4324 18582 4380
rect 18518 4320 18582 4324
rect 9812 3904 9876 3908
rect 9812 3848 9862 3904
rect 9862 3848 9876 3904
rect 9812 3844 9876 3848
rect 7882 3836 7946 3840
rect 7882 3780 7886 3836
rect 7886 3780 7942 3836
rect 7942 3780 7946 3836
rect 7882 3776 7946 3780
rect 7962 3836 8026 3840
rect 7962 3780 7966 3836
rect 7966 3780 8022 3836
rect 8022 3780 8026 3836
rect 7962 3776 8026 3780
rect 8042 3836 8106 3840
rect 8042 3780 8046 3836
rect 8046 3780 8102 3836
rect 8102 3780 8106 3836
rect 8042 3776 8106 3780
rect 8122 3836 8186 3840
rect 8122 3780 8126 3836
rect 8126 3780 8182 3836
rect 8182 3780 8186 3836
rect 8122 3776 8186 3780
rect 14813 3836 14877 3840
rect 14813 3780 14817 3836
rect 14817 3780 14873 3836
rect 14873 3780 14877 3836
rect 14813 3776 14877 3780
rect 14893 3836 14957 3840
rect 14893 3780 14897 3836
rect 14897 3780 14953 3836
rect 14953 3780 14957 3836
rect 14893 3776 14957 3780
rect 14973 3836 15037 3840
rect 14973 3780 14977 3836
rect 14977 3780 15033 3836
rect 15033 3780 15037 3836
rect 14973 3776 15037 3780
rect 15053 3836 15117 3840
rect 15053 3780 15057 3836
rect 15057 3780 15113 3836
rect 15113 3780 15117 3836
rect 15053 3776 15117 3780
rect 8340 3708 8404 3772
rect 11100 3300 11164 3364
rect 19012 3300 19076 3364
rect 4417 3292 4481 3296
rect 4417 3236 4421 3292
rect 4421 3236 4477 3292
rect 4477 3236 4481 3292
rect 4417 3232 4481 3236
rect 4497 3292 4561 3296
rect 4497 3236 4501 3292
rect 4501 3236 4557 3292
rect 4557 3236 4561 3292
rect 4497 3232 4561 3236
rect 4577 3292 4641 3296
rect 4577 3236 4581 3292
rect 4581 3236 4637 3292
rect 4637 3236 4641 3292
rect 4577 3232 4641 3236
rect 4657 3292 4721 3296
rect 4657 3236 4661 3292
rect 4661 3236 4717 3292
rect 4717 3236 4721 3292
rect 4657 3232 4721 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 18278 3292 18342 3296
rect 18278 3236 18282 3292
rect 18282 3236 18338 3292
rect 18338 3236 18342 3292
rect 18278 3232 18342 3236
rect 18358 3292 18422 3296
rect 18358 3236 18362 3292
rect 18362 3236 18418 3292
rect 18418 3236 18422 3292
rect 18358 3232 18422 3236
rect 18438 3292 18502 3296
rect 18438 3236 18442 3292
rect 18442 3236 18498 3292
rect 18498 3236 18502 3292
rect 18438 3232 18502 3236
rect 18518 3292 18582 3296
rect 18518 3236 18522 3292
rect 18522 3236 18578 3292
rect 18578 3236 18582 3292
rect 18518 3232 18582 3236
rect 3004 3224 3068 3228
rect 3004 3168 3054 3224
rect 3054 3168 3068 3224
rect 3004 3164 3068 3168
rect 18828 3164 18892 3228
rect 18092 3028 18156 3092
rect 7882 2748 7946 2752
rect 7882 2692 7886 2748
rect 7886 2692 7942 2748
rect 7942 2692 7946 2748
rect 7882 2688 7946 2692
rect 7962 2748 8026 2752
rect 7962 2692 7966 2748
rect 7966 2692 8022 2748
rect 8022 2692 8026 2748
rect 7962 2688 8026 2692
rect 8042 2748 8106 2752
rect 8042 2692 8046 2748
rect 8046 2692 8102 2748
rect 8102 2692 8106 2748
rect 8042 2688 8106 2692
rect 8122 2748 8186 2752
rect 8122 2692 8126 2748
rect 8126 2692 8182 2748
rect 8182 2692 8186 2748
rect 8122 2688 8186 2692
rect 14813 2748 14877 2752
rect 14813 2692 14817 2748
rect 14817 2692 14873 2748
rect 14873 2692 14877 2748
rect 14813 2688 14877 2692
rect 14893 2748 14957 2752
rect 14893 2692 14897 2748
rect 14897 2692 14953 2748
rect 14953 2692 14957 2748
rect 14893 2688 14957 2692
rect 14973 2748 15037 2752
rect 14973 2692 14977 2748
rect 14977 2692 15033 2748
rect 15033 2692 15037 2748
rect 14973 2688 15037 2692
rect 15053 2748 15117 2752
rect 15053 2692 15057 2748
rect 15057 2692 15113 2748
rect 15113 2692 15117 2748
rect 15053 2688 15117 2692
rect 17908 2756 17972 2820
rect 19196 2348 19260 2412
rect 4417 2204 4481 2208
rect 4417 2148 4421 2204
rect 4421 2148 4477 2204
rect 4477 2148 4481 2204
rect 4417 2144 4481 2148
rect 4497 2204 4561 2208
rect 4497 2148 4501 2204
rect 4501 2148 4557 2204
rect 4557 2148 4561 2204
rect 4497 2144 4561 2148
rect 4577 2204 4641 2208
rect 4577 2148 4581 2204
rect 4581 2148 4637 2204
rect 4637 2148 4641 2204
rect 4577 2144 4641 2148
rect 4657 2204 4721 2208
rect 4657 2148 4661 2204
rect 4661 2148 4717 2204
rect 4717 2148 4721 2204
rect 4657 2144 4721 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 18278 2204 18342 2208
rect 18278 2148 18282 2204
rect 18282 2148 18338 2204
rect 18338 2148 18342 2204
rect 18278 2144 18342 2148
rect 18358 2204 18422 2208
rect 18358 2148 18362 2204
rect 18362 2148 18418 2204
rect 18418 2148 18422 2204
rect 18358 2144 18422 2148
rect 18438 2204 18502 2208
rect 18438 2148 18442 2204
rect 18442 2148 18498 2204
rect 18498 2148 18502 2204
rect 18438 2144 18502 2148
rect 18518 2204 18582 2208
rect 18518 2148 18522 2204
rect 18522 2148 18578 2204
rect 18578 2148 18582 2204
rect 18518 2144 18582 2148
<< metal4 >>
rect 4409 20704 4729 20720
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 19616 4729 20640
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 18528 4729 19552
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 17440 4729 18464
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 16352 4729 17376
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 15264 4729 16288
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 14176 4729 15200
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 13088 4729 14112
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 12000 4729 13024
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 10912 4729 11936
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 9824 4729 10848
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 8736 4729 9760
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 7648 4729 8672
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 3003 6764 3069 6765
rect 3003 6700 3004 6764
rect 3068 6700 3069 6764
rect 3003 6699 3069 6700
rect 3006 3229 3066 6699
rect 4409 6560 4729 7584
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 5472 4729 6496
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 4384 4729 5408
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 3296 4729 4320
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 3003 3228 3069 3229
rect 3003 3164 3004 3228
rect 3068 3164 3069 3228
rect 3003 3163 3069 3164
rect 4409 2208 4729 3232
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2128 4729 2144
rect 7874 20160 8195 20720
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8195 20160
rect 7874 19072 8195 20096
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8195 19072
rect 7874 17984 8195 19008
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8195 17984
rect 7874 16896 8195 17920
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8195 16896
rect 7874 15808 8195 16832
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8195 15808
rect 7874 14720 8195 15744
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8195 14720
rect 7874 13632 8195 14656
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8195 13632
rect 7874 12544 8195 13568
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8195 12544
rect 7874 11456 8195 12480
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8195 11456
rect 7874 10368 8195 11392
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8195 10368
rect 7874 9280 8195 10304
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11099 9620 11165 9621
rect 11099 9556 11100 9620
rect 11164 9556 11165 9620
rect 11099 9555 11165 9556
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8195 9280
rect 7874 8192 8195 9216
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8195 8192
rect 7874 7104 8195 8128
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8195 7104
rect 7874 6016 8195 7040
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8195 6016
rect 7874 4928 8195 5952
rect 9811 5540 9877 5541
rect 9811 5476 9812 5540
rect 9876 5476 9877 5540
rect 9811 5475 9877 5476
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8195 4928
rect 7874 3840 8195 4864
rect 8339 4554 8405 4555
rect 8339 4490 8340 4554
rect 8404 4490 8405 4554
rect 8339 4489 8405 4490
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8195 3840
rect 7874 2752 8195 3776
rect 8342 3773 8402 4489
rect 9814 3909 9874 5475
rect 9811 3908 9877 3909
rect 9811 3844 9812 3908
rect 9876 3844 9877 3908
rect 9811 3843 9877 3844
rect 8339 3772 8405 3773
rect 8339 3708 8340 3772
rect 8404 3708 8405 3772
rect 8339 3707 8405 3708
rect 11102 3365 11162 9555
rect 11340 8736 11660 9760
rect 14805 20160 15125 20720
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 19072 15125 20096
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 17984 15125 19008
rect 18270 20704 18590 20720
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 18270 19616 18590 20640
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 18528 18590 19552
rect 18827 19276 18893 19277
rect 18827 19212 18828 19276
rect 18892 19212 18893 19276
rect 18827 19211 18893 19212
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18091 18460 18157 18461
rect 18091 18396 18092 18460
rect 18156 18396 18157 18460
rect 18091 18395 18157 18396
rect 17907 18052 17973 18053
rect 17907 17988 17908 18052
rect 17972 17988 17973 18052
rect 17907 17987 17973 17988
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 16896 15125 17920
rect 17539 17916 17605 17917
rect 17539 17852 17540 17916
rect 17604 17852 17605 17916
rect 17539 17851 17605 17852
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 15808 15125 16832
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 14720 15125 15744
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 13632 15125 14656
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 12544 15125 13568
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 11456 15125 12480
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 10368 15125 11392
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 9280 15125 10304
rect 17542 10165 17602 17851
rect 17723 13428 17789 13429
rect 17723 13364 17724 13428
rect 17788 13364 17789 13428
rect 17723 13363 17789 13364
rect 17726 11389 17786 13363
rect 17723 11388 17789 11389
rect 17723 11324 17724 11388
rect 17788 11324 17789 11388
rect 17723 11323 17789 11324
rect 17539 10164 17605 10165
rect 17539 10100 17540 10164
rect 17604 10100 17605 10164
rect 17539 10099 17605 10100
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 11835 9212 11901 9213
rect 11835 9148 11836 9212
rect 11900 9148 11901 9212
rect 11835 9147 11901 9148
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11838 4453 11898 9147
rect 14805 8192 15125 9216
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 7104 15125 8128
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 6016 15125 7040
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 4928 15125 5952
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 11835 4452 11901 4453
rect 11835 4388 11836 4452
rect 11900 4388 11901 4452
rect 11835 4387 11901 4388
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11099 3364 11165 3365
rect 11099 3300 11100 3364
rect 11164 3300 11165 3364
rect 11099 3299 11165 3300
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8195 2752
rect 7874 2128 8195 2688
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 14805 3840 15125 4864
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 2752 15125 3776
rect 17910 2821 17970 17987
rect 18094 3093 18154 18395
rect 18270 17440 18590 18464
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 18270 16352 18590 17376
rect 18830 16693 18890 19211
rect 18827 16692 18893 16693
rect 18827 16628 18828 16692
rect 18892 16628 18893 16692
rect 18827 16627 18893 16628
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 15264 18590 16288
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 14176 18590 15200
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 18270 13088 18590 14112
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 12000 18590 13024
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 18270 10912 18590 11936
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 18270 9824 18590 10848
rect 18830 10709 18890 16627
rect 18827 10708 18893 10709
rect 18827 10644 18828 10708
rect 18892 10644 18893 10708
rect 18827 10643 18893 10644
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 8736 18590 9760
rect 19011 9348 19077 9349
rect 19011 9284 19012 9348
rect 19076 9284 19077 9348
rect 19011 9283 19077 9284
rect 19014 9210 19074 9283
rect 19014 9150 19258 9210
rect 18827 9076 18893 9077
rect 18827 9012 18828 9076
rect 18892 9012 18893 9076
rect 18827 9011 18893 9012
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 7648 18590 8672
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 18270 6560 18590 7584
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 5472 18590 6496
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 4384 18590 5408
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 18270 3296 18590 4320
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 18091 3092 18157 3093
rect 18091 3028 18092 3092
rect 18156 3028 18157 3092
rect 18091 3027 18157 3028
rect 17907 2820 17973 2821
rect 17907 2756 17908 2820
rect 17972 2756 17973 2820
rect 17907 2755 17973 2756
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2128 15125 2688
rect 18270 2208 18590 3232
rect 18830 3229 18890 9011
rect 19011 8124 19077 8125
rect 19011 8060 19012 8124
rect 19076 8060 19077 8124
rect 19011 8059 19077 8060
rect 19014 3365 19074 8059
rect 19011 3364 19077 3365
rect 19011 3300 19012 3364
rect 19076 3300 19077 3364
rect 19011 3299 19077 3300
rect 18827 3228 18893 3229
rect 18827 3164 18828 3228
rect 18892 3164 18893 3228
rect 18827 3163 18893 3164
rect 19198 2413 19258 9150
rect 19195 2412 19261 2413
rect 19195 2348 19196 2412
rect 19260 2348 19261 2412
rect 19195 2347 19261 2348
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2128 18590 2144
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2852 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2852 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 3772 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28
timestamp 1604681595
transform 1 0 3680 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_28 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3680 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _114_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6348 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5520 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5244 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6072 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1604681595
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_60
timestamp 1604681595
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1604681595
transform 1 0 8556 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 7820 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 7728 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_79 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8372 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9292 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1604681595
transform 1 0 8924 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103
timestamp 1604681595
transform 1 0 10580 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_87 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 9108 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1604681595
transform 1 0 11316 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1604681595
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_123 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 1604681595
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_117
timestamp 1604681595
transform 1 0 11868 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_116
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_1_105 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 10764 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1604681595
transform 1 0 14168 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 14352 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12788 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_0_134
timestamp 1604681595
transform 1 0 13432 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_136
timestamp 1604681595
transform 1 0 13616 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15916 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_146
timestamp 1604681595
transform 1 0 14536 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154
timestamp 1604681595
transform 1 0 15272 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_162
timestamp 1604681595
transform 1 0 16008 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_153
timestamp 1604681595
transform 1 0 15180 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_177
timestamp 1604681595
transform 1 0 17388 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_170
timestamp 1604681595
transform 1 0 16744 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16836 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_179
timestamp 1604681595
transform 1 0 17572 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_185
timestamp 1604681595
transform 1 0 18124 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_167
timestamp 1604681595
transform 1 0 16468 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1604681595
transform 1 0 19964 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1604681595
transform 1 0 19412 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18676 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1604681595
transform 1 0 19228 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_190
timestamp 1604681595
transform 1 0 18584 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_198
timestamp 1604681595
transform 1 0 19320 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_203
timestamp 1604681595
transform 1 0 19780 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1604681595
transform 1 0 20516 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 21896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 21896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_209
timestamp 1604681595
transform 1 0 20332 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_222
timestamp 1604681595
transform 1 0 21528 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_215
timestamp 1604681595
transform 1 0 20884 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 1564 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 3036 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_30
timestamp 1604681595
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6624 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 5520 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_2_57
timestamp 1604681595
transform 1 0 6348 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _028_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8556 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_69
timestamp 1604681595
transform 1 0 7452 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10212 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_84
timestamp 1604681595
transform 1 0 8832 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_93 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1604681595
transform 1 0 11776 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_108
timestamp 1604681595
transform 1 0 11040 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_125
timestamp 1604681595
transform 1 0 12604 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13524 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_133
timestamp 1604681595
transform 1 0 13340 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_144
timestamp 1604681595
transform 1 0 14352 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_152
timestamp 1604681595
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_163
timestamp 1604681595
transform 1 0 16100 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 17112 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_2_171
timestamp 1604681595
transform 1 0 16836 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_180
timestamp 1604681595
transform 1 0 17664 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18584 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_188
timestamp 1604681595
transform 1 0 18400 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_206
timestamp 1604681595
transform 1 0 20056 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 21896 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_215
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 2944 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 1472 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4416 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_42
timestamp 1604681595
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_53
timestamp 1604681595
transform 1 0 5980 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 7452 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_68
timestamp 1604681595
transform 1 0 7360 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_75
timestamp 1604681595
transform 1 0 8004 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1604681595
transform 1 0 9476 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10580 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_87
timestamp 1604681595
transform 1 0 9108 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_95
timestamp 1604681595
transform 1 0 9844 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_112
timestamp 1604681595
transform 1 0 11408 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1604681595
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13432 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_126
timestamp 1604681595
transform 1 0 12696 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_143
timestamp 1604681595
transform 1 0 14260 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1604681595
transform 1 0 16284 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 14996 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_157
timestamp 1604681595
transform 1 0 15548 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_168
timestamp 1604681595
transform 1 0 16560 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_180
timestamp 1604681595
transform 1 0 17664 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_184
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18492 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_188
timestamp 1604681595
transform 1 0 18400 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_198
timestamp 1604681595
transform 1 0 19320 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1604681595
transform 1 0 20516 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_210
timestamp 1604681595
transform 1 0 20424 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_215
timestamp 1604681595
transform 1 0 20884 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2852 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1604681595
transform 1 0 3680 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4876 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1604681595
transform 1 0 5704 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1604681595
transform 1 0 5980 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7360 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_4_65
timestamp 1604681595
transform 1 0 7084 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_84
timestamp 1604681595
transform 1 0 8832 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_102
timestamp 1604681595
transform 1 0 10488 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11408 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_110
timestamp 1604681595
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_118
timestamp 1604681595
transform 1 0 11960 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12696 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_4_142
timestamp 1604681595
transform 1 0 14168 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16008 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_150
timestamp 1604681595
transform 1 0 14904 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_154
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 17572 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_4_171
timestamp 1604681595
transform 1 0 16836 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1604681595
transform 1 0 19780 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1604681595
transform 1 0 19596 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_195
timestamp 1604681595
transform 1 0 19044 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_206
timestamp 1604681595
transform 1 0 20056 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 21896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_215
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_19
timestamp 1604681595
transform 1 0 2852 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1604681595
transform 1 0 3680 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1604681595
transform 1 0 3496 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_25
timestamp 1604681595
transform 1 0 3404 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_37
timestamp 1604681595
transform 1 0 4508 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1604681595
transform 1 0 5060 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_52
timestamp 1604681595
transform 1 0 5888 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_60
timestamp 1604681595
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1604681595
transform 1 0 7820 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_65
timestamp 1604681595
transform 1 0 7084 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_76
timestamp 1604681595
transform 1 0 8096 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1604681595
transform 1 0 8832 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9844 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_87
timestamp 1604681595
transform 1 0 9108 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_104
timestamp 1604681595
transform 1 0 10672 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12512 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_116
timestamp 1604681595
transform 1 0 11776 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1604681595
transform 1 0 14168 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_130
timestamp 1604681595
transform 1 0 13064 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1604681595
transform 1 0 15272 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_146
timestamp 1604681595
transform 1 0 14536 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_158
timestamp 1604681595
transform 1 0 15640 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_175
timestamp 1604681595
transform 1 0 17204 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_184
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1604681595
transform 1 0 18400 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 19412 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_5_191
timestamp 1604681595
transform 1 0 18676 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 21896 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_215
timestamp 1604681595
transform 1 0 20884 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1604681595
transform 1 0 2392 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1604681595
transform 1 0 1564 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1604681595
transform 1 0 2208 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_18
timestamp 1604681595
transform 1 0 2760 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1604681595
transform 1 0 3404 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4508 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_23
timestamp 1604681595
transform 1 0 3220 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_35
timestamp 1604681595
transform 1 0 4324 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_24
timestamp 1604681595
transform 1 0 3312 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_29
timestamp 1604681595
transform 1 0 3772 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 5336 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_43
timestamp 1604681595
transform 1 0 5060 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_62
timestamp 1604681595
transform 1 0 6808 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_53
timestamp 1604681595
transform 1 0 5980 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6992 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7544 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_6_79
timestamp 1604681595
transform 1 0 8372 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_80
timestamp 1604681595
transform 1 0 8464 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9384 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10028 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1604681595
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_88
timestamp 1604681595
transform 1 0 9200 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11960 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_106
timestamp 1604681595
transform 1 0 10856 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_106
timestamp 1604681595
transform 1 0 10856 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1604681595
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1604681595
transform 1 0 14168 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_134
timestamp 1604681595
transform 1 0 13432 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_145
timestamp 1604681595
transform 1 0 14444 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_139
timestamp 1604681595
transform 1 0 13892 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_1_
timestamp 1604681595
transform 1 0 14904 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_163
timestamp 1604681595
transform 1 0 16100 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_147
timestamp 1604681595
transform 1 0 14628 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1604681595
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1604681595
transform 1 0 16928 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 17204 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_171
timestamp 1604681595
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_175
timestamp 1604681595
transform 1 0 17204 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1604681595
transform 1 0 19596 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19412 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_191
timestamp 1604681595
transform 1 0 18676 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_205
timestamp 1604681595
transform 1 0 19964 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_193
timestamp 1604681595
transform 1 0 18860 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_204
timestamp 1604681595
transform 1 0 19872 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1604681595
transform 1 0 20608 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 21896 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 21896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp 1604681595
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_215
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_215
timestamp 1604681595
transform 1 0 20884 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1604681595
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_11
timestamp 1604681595
transform 1 0 2116 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_3_
timestamp 1604681595
transform 1 0 4692 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_23
timestamp 1604681595
transform 1 0 3220 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_38
timestamp 1604681595
transform 1 0 4600 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6256 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_48
timestamp 1604681595
transform 1 0 5520 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7820 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_65
timestamp 1604681595
transform 1 0 7084 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_82
timestamp 1604681595
transform 1 0 8648 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1604681595
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_102
timestamp 1604681595
transform 1 0 10488 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l3_in_0_
timestamp 1604681595
transform 1 0 11960 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_114
timestamp 1604681595
transform 1 0 11592 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_127
timestamp 1604681595
transform 1 0 12788 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_135
timestamp 1604681595
transform 1 0 13524 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_145
timestamp 1604681595
transform 1 0 14444 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15824 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1604681595
transform 1 0 18124 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_176
timestamp 1604681595
transform 1 0 17296 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_184
timestamp 1604681595
transform 1 0 18032 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19136 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_188
timestamp 1604681595
transform 1 0 18400 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_205
timestamp 1604681595
transform 1 0 19964 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 21896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1604681595
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1604681595
transform 1 0 2208 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 2576 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4784 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_32
timestamp 1604681595
transform 1 0 4048 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_2_
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_49
timestamp 1604681595
transform 1 0 5612 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 8372 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_9_71
timestamp 1604681595
transform 1 0 7636 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10580 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_95
timestamp 1604681595
transform 1 0 9844 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_112
timestamp 1604681595
transform 1 0 11408 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1604681595
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13984 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_132
timestamp 1604681595
transform 1 0 13248 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15732 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_9_149
timestamp 1604681595
transform 1 0 14812 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_157
timestamp 1604681595
transform 1 0 15548 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1604681595
transform 1 0 18124 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_175
timestamp 1604681595
transform 1 0 17204 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_184
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19412 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_9_188
timestamp 1604681595
transform 1 0 18400 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_196
timestamp 1604681595
transform 1 0 19136 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 21896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_215
timestamp 1604681595
transform 1 0 20884 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1604681595
transform 1 0 1840 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 2116 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_7
timestamp 1604681595
transform 1 0 1748 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_20
timestamp 1604681595
transform 1 0 2944 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4784 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_28
timestamp 1604681595
transform 1 0 3680 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_56
timestamp 1604681595
transform 1 0 6256 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 7084 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8648 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_64
timestamp 1604681595
transform 1 0 6992 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_74
timestamp 1604681595
transform 1 0 7912 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_85
timestamp 1604681595
transform 1 0 8924 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1604681595
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_102
timestamp 1604681595
transform 1 0 10488 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11500 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_10_110
timestamp 1604681595
transform 1 0 11224 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13892 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_129
timestamp 1604681595
transform 1 0 12972 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_137
timestamp 1604681595
transform 1 0 13708 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_145
timestamp 1604681595
transform 1 0 14444 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 17940 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 17480 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_170
timestamp 1604681595
transform 1 0 16744 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_181
timestamp 1604681595
transform 1 0 17756 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_199
timestamp 1604681595
transform 1 0 19412 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 21896 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_211
timestamp 1604681595
transform 1 0 20516 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2116 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_20
timestamp 1604681595
transform 1 0 2944 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4416 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_32
timestamp 1604681595
transform 1 0 4048 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1604681595
transform 1 0 5980 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_45
timestamp 1604681595
transform 1 0 5244 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_56
timestamp 1604681595
transform 1 0 6256 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_60
timestamp 1604681595
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6992 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_11_73
timestamp 1604681595
transform 1 0 7820 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9200 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_11_85
timestamp 1604681595
transform 1 0 8924 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_104
timestamp 1604681595
transform 1 0 10672 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_116
timestamp 1604681595
transform 1 0 11776 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 14168 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_11_132
timestamp 1604681595
transform 1 0 13248 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_140
timestamp 1604681595
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_158
timestamp 1604681595
transform 1 0 15640 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_175
timestamp 1604681595
transform 1 0 17204 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20056 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1604681595
transform 1 0 18860 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_205
timestamp 1604681595
transform 1 0 19964 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 21896 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_215
timestamp 1604681595
transform 1 0 20884 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 1748 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_23
timestamp 1604681595
transform 1 0 3220 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6716 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 6440 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_48
timestamp 1604681595
transform 1 0 5520 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_56
timestamp 1604681595
transform 1 0 6256 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1604681595
transform 1 0 8464 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_70
timestamp 1604681595
transform 1 0 7544 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_78
timestamp 1604681595
transform 1 0 8280 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10488 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_84
timestamp 1604681595
transform 1 0 8832 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_101
timestamp 1604681595
transform 1 0 10396 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_118
timestamp 1604681595
transform 1 0 11960 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 12972 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 12696 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_145
timestamp 1604681595
transform 1 0 14444 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16376 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_158
timestamp 1604681595
transform 1 0 15640 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_182
timestamp 1604681595
transform 1 0 17848 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18584 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_12_199
timestamp 1604681595
transform 1 0 19412 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 21896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_211
timestamp 1604681595
transform 1 0 20516 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_9
timestamp 1604681595
transform 1 0 1932 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 1604681595
transform 1 0 1748 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 1840 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 2024 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_13_17
timestamp 1604681595
transform 1 0 2668 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_19
timestamp 1604681595
transform 1 0 2852 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 4508 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 3588 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_25
timestamp 1604681595
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_36
timestamp 1604681595
transform 1 0 4416 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_36
timestamp 1604681595
transform 1 0 4416 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1604681595
transform 1 0 6716 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1604681595
transform 1 0 5152 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_53
timestamp 1604681595
transform 1 0 5980 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_53
timestamp 1604681595
transform 1 0 5980 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1604681595
transform 1 0 8280 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1604681595
transform 1 0 8648 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_71
timestamp 1604681595
transform 1 0 7636 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_79
timestamp 1604681595
transform 1 0 8372 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_70
timestamp 1604681595
transform 1 0 7544 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_82
timestamp 1604681595
transform 1 0 8648 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 9752 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_86
timestamp 1604681595
transform 1 0 9016 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_103
timestamp 1604681595
transform 1 0 10580 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1604681595
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1604681595
transform 1 0 11316 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12052 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_114
timestamp 1604681595
transform 1 0 11592 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_109
timestamp 1604681595
transform 1 0 11132 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_117
timestamp 1604681595
transform 1 0 11868 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_13_139
timestamp 1604681595
transform 1 0 13892 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_128
timestamp 1604681595
transform 1 0 12880 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_145
timestamp 1604681595
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 14812 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15364 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_147
timestamp 1604681595
transform 1 0 14628 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_158
timestamp 1604681595
transform 1 0 15640 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_154
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_164
timestamp 1604681595
transform 1 0 16192 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 16928 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_175
timestamp 1604681595
transform 1 0 17204 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 19228 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_13_188
timestamp 1604681595
transform 1 0 18400 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_196
timestamp 1604681595
transform 1 0 19136 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_188
timestamp 1604681595
transform 1 0 18400 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_196
timestamp 1604681595
transform 1 0 19136 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_206
timestamp 1604681595
transform 1 0 20056 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 21896 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 21896 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_213
timestamp 1604681595
transform 1 0 20700 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_221
timestamp 1604681595
transform 1 0 21436 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 2852 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1564 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_11
timestamp 1604681595
transform 1 0 2116 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_35
timestamp 1604681595
transform 1 0 4324 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_43
timestamp 1604681595
transform 1 0 5060 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_53
timestamp 1604681595
transform 1 0 5980 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_78
timestamp 1604681595
transform 1 0 8280 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1604681595
transform 1 0 10304 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9476 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1604681595
transform 1 0 9016 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_89
timestamp 1604681595
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_104
timestamp 1604681595
transform 1 0 10672 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1604681595
transform 1 0 11224 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_114
timestamp 1604681595
transform 1 0 11592 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_123
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13248 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_131
timestamp 1604681595
transform 1 0 13156 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_141
timestamp 1604681595
transform 1 0 14076 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14812 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_15_158
timestamp 1604681595
transform 1 0 15640 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1604681595
transform 1 0 18308 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_175
timestamp 1604681595
transform 1 0 17204 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_184
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 19412 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_15_191
timestamp 1604681595
transform 1 0 18676 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_215
timestamp 1604681595
transform 1 0 20884 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_6
timestamp 1604681595
transform 1 0 1656 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_23
timestamp 1604681595
transform 1 0 3220 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_38
timestamp 1604681595
transform 1 0 4600 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1604681595
transform 1 0 5336 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_16_55
timestamp 1604681595
transform 1 0 6164 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7360 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_16_67
timestamp 1604681595
transform 1 0 7268 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 10396 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_16_84
timestamp 1604681595
transform 1 0 8832 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 12236 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13708 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15548 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_146
timestamp 1604681595
transform 1 0 14536 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1604681595
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_154
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_1_
timestamp 1604681595
transform 1 0 17756 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_173
timestamp 1604681595
transform 1 0 17020 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19504 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_190
timestamp 1604681595
transform 1 0 18584 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_198
timestamp 1604681595
transform 1 0 19320 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_206
timestamp 1604681595
transform 1 0 20056 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 21896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 1840 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_7
timestamp 1604681595
transform 1 0 1748 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_17
timestamp 1604681595
transform 1 0 2668 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 3404 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_34
timestamp 1604681595
transform 1 0 4232 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4968 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1604681595
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1604681595
transform 1 0 7360 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_17_77
timestamp 1604681595
transform 1 0 8188 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9660 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_89
timestamp 1604681595
transform 1 0 9292 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1604681595
transform 1 0 12052 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_109
timestamp 1604681595
transform 1 0 11132 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_117
timestamp 1604681595
transform 1 0 11868 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12972 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_17_145
timestamp 1604681595
transform 1 0 14444 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1604681595
transform 1 0 15272 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_153
timestamp 1604681595
transform 1 0 15180 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_158
timestamp 1604681595
transform 1 0 15640 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_175
timestamp 1604681595
transform 1 0 17204 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_187
timestamp 1604681595
transform 1 0 18308 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_1_
timestamp 1604681595
transform 1 0 19044 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_204
timestamp 1604681595
transform 1 0 19872 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1604681595
transform 1 0 20608 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 21896 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_215
timestamp 1604681595
transform 1 0 20884 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 2208 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_11
timestamp 1604681595
transform 1 0 2116 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_21
timestamp 1604681595
transform 1 0 3036 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1604681595
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_35
timestamp 1604681595
transform 1 0 4324 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_3_
timestamp 1604681595
transform 1 0 6808 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5060 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_52
timestamp 1604681595
transform 1 0 5888 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_60
timestamp 1604681595
transform 1 0 6624 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1604681595
transform 1 0 8464 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_71
timestamp 1604681595
transform 1 0 7636 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_79
timestamp 1604681595
transform 1 0 8372 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_84
timestamp 1604681595
transform 1 0 8832 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_102
timestamp 1604681595
transform 1 0 10488 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1604681595
transform 1 0 11868 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_18_114
timestamp 1604681595
transform 1 0 11592 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13432 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_126
timestamp 1604681595
transform 1 0 12696 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_143
timestamp 1604681595
transform 1 0 14260 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1604681595
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_163
timestamp 1604681595
transform 1 0 16100 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 17112 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_18_171
timestamp 1604681595
transform 1 0 16836 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1604681595
transform 1 0 19688 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_190
timestamp 1604681595
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_206
timestamp 1604681595
transform 1 0 20056 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 21896 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_215
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 2300 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_11
timestamp 1604681595
transform 1 0 2116 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_6
timestamp 1604681595
transform 1 0 1656 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1604681595
transform 1 0 3864 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_22
timestamp 1604681595
transform 1 0 3128 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_34
timestamp 1604681595
transform 1 0 4232 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_23
timestamp 1604681595
transform 1 0 3220 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_38
timestamp 1604681595
transform 1 0 4600 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5520 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1604681595
transform 1 0 4968 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1604681595
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_46
timestamp 1604681595
transform 1 0 5336 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_57
timestamp 1604681595
transform 1 0 6348 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7084 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 8372 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 8648 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_71
timestamp 1604681595
transform 1 0 7636 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_82
timestamp 1604681595
transform 1 0 8648 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_74
timestamp 1604681595
transform 1 0 7912 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9200 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_97
timestamp 1604681595
transform 1 0 10028 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1604681595
transform 1 0 8924 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1604681595
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_102
timestamp 1604681595
transform 1 0 10488 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1604681595
transform 1 0 11224 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 12236 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_114
timestamp 1604681595
transform 1 0 11592 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_113
timestamp 1604681595
transform 1 0 11500 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13892 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_3_
timestamp 1604681595
transform 1 0 14352 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 13984 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_132
timestamp 1604681595
transform 1 0 13248 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_143
timestamp 1604681595
transform 1 0 14260 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_130
timestamp 1604681595
transform 1 0 13064 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_138
timestamp 1604681595
transform 1 0 13800 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_145
timestamp 1604681595
transform 1 0 14444 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15916 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_153
timestamp 1604681595
transform 1 0 15180 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_163
timestamp 1604681595
transform 1 0 16100 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 17296 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_170
timestamp 1604681595
transform 1 0 16744 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_182
timestamp 1604681595
transform 1 0 17848 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_175
timestamp 1604681595
transform 1 0 17204 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_185
timestamp 1604681595
transform 1 0 18124 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18768 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18860 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1604681595
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_202
timestamp 1604681595
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 21896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 21896 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_220
timestamp 1604681595
transform 1 0 21344 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1604681595
transform 1 0 1472 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 2576 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_8
timestamp 1604681595
transform 1 0 1840 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4784 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_32
timestamp 1604681595
transform 1 0 4048 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 6348 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_49
timestamp 1604681595
transform 1 0 5612 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_60
timestamp 1604681595
transform 1 0 6624 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1604681595
transform 1 0 8372 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_71
timestamp 1604681595
transform 1 0 7636 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 10120 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_21_88
timestamp 1604681595
transform 1 0 9200 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_96
timestamp 1604681595
transform 1 0 9936 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_114
timestamp 1604681595
transform 1 0 11592 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13984 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_132
timestamp 1604681595
transform 1 0 13248 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15916 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1604681595
transform 1 0 14812 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18216 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_170
timestamp 1604681595
transform 1 0 16744 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_182
timestamp 1604681595
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_195
timestamp 1604681595
transform 1 0 19044 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_207
timestamp 1604681595
transform 1 0 20148 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1604681595
transform 1 0 20516 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 21896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_215
timestamp 1604681595
transform 1 0 20884 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_6_
timestamp 1604681595
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_6
timestamp 1604681595
transform 1 0 1656 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_23
timestamp 1604681595
transform 1 0 3220 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_41
timestamp 1604681595
transform 1 0 4876 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5796 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_49
timestamp 1604681595
transform 1 0 5612 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_3_
timestamp 1604681595
transform 1 0 8004 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_22_67
timestamp 1604681595
transform 1 0 7268 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_84
timestamp 1604681595
transform 1 0 8832 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_97
timestamp 1604681595
transform 1 0 10028 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 11040 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_22_105
timestamp 1604681595
transform 1 0 10764 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_124
timestamp 1604681595
transform 1 0 12512 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 13248 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_22_141
timestamp 1604681595
transform 1 0 14076 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 14812 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_152
timestamp 1604681595
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_170
timestamp 1604681595
transform 1 0 16744 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_182
timestamp 1604681595
transform 1 0 17848 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1604681595
transform 1 0 18400 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19504 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_192
timestamp 1604681595
transform 1 0 18768 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_206
timestamp 1604681595
transform 1 0 20056 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 21896 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_5_
timestamp 1604681595
transform 1 0 1932 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_18
timestamp 1604681595
transform 1 0 2760 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 3496 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1604681595
transform 1 0 5704 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_42
timestamp 1604681595
transform 1 0 4968 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_53
timestamp 1604681595
transform 1 0 5980 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_78
timestamp 1604681595
transform 1 0 8280 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9016 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_23_102
timestamp 1604681595
transform 1 0 10488 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1604681595
transform 1 0 11224 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_114
timestamp 1604681595
transform 1 0 11592 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_123
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13064 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_23_129
timestamp 1604681595
transform 1 0 12972 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15272 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_23_146
timestamp 1604681595
transform 1 0 14536 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_170
timestamp 1604681595
transform 1 0 16744 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_182
timestamp 1604681595
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18860 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_192
timestamp 1604681595
transform 1 0 18768 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_202
timestamp 1604681595
transform 1 0 19688 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1604681595
transform 1 0 20516 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 21896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_210
timestamp 1604681595
transform 1 0 20424 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_215
timestamp 1604681595
transform 1 0 20884 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1604681595
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_6
timestamp 1604681595
transform 1 0 1656 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4232 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_23
timestamp 1604681595
transform 1 0 3220 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_32
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6440 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_24_50
timestamp 1604681595
transform 1 0 5704 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_24_67
timestamp 1604681595
transform 1 0 7268 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_84
timestamp 1604681595
transform 1 0 8832 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_102
timestamp 1604681595
transform 1 0 10488 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1604681595
transform 1 0 11500 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_24_110
timestamp 1604681595
transform 1 0 11224 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_122
timestamp 1604681595
transform 1 0 12328 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1604681595
transform 1 0 13064 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_24_139
timestamp 1604681595
transform 1 0 13892 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 16100 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_151
timestamp 1604681595
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_162
timestamp 1604681595
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 17664 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_24_172
timestamp 1604681595
transform 1 0 16928 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1604681595
transform 1 0 19688 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_189
timestamp 1604681595
transform 1 0 18492 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_201
timestamp 1604681595
transform 1 0 19596 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_206
timestamp 1604681595
transform 1 0 20056 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 21896 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_4_
timestamp 1604681595
transform 1 0 1472 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_13
timestamp 1604681595
transform 1 0 2300 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4600 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1604681595
transform 1 0 3036 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_25_30
timestamp 1604681595
transform 1 0 3864 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_47
timestamp 1604681595
transform 1 0 5428 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8372 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_25_71
timestamp 1604681595
transform 1 0 7636 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_95
timestamp 1604681595
transform 1 0 9844 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_103
timestamp 1604681595
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1604681595
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_114
timestamp 1604681595
transform 1 0 11592 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_123
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 12880 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_25_127
timestamp 1604681595
transform 1 0 12788 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_144
timestamp 1604681595
transform 1 0 14352 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15088 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1604681595
transform 1 0 18124 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_168
timestamp 1604681595
transform 1 0 16560 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_180
timestamp 1604681595
transform 1 0 17664 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_184
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19228 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_189
timestamp 1604681595
transform 1 0 18492 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_203
timestamp 1604681595
transform 1 0 19780 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1604681595
transform 1 0 20516 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 21896 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_215
timestamp 1604681595
transform 1 0 20884 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1932 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_6
timestamp 1604681595
transform 1 0 1656 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_15
timestamp 1604681595
transform 1 0 2484 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 3496 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4140 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_23
timestamp 1604681595
transform 1 0 3220 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_32
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_23
timestamp 1604681595
transform 1 0 3220 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1604681595
transform 1 0 5704 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5704 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_42
timestamp 1604681595
transform 1 0 4968 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_42
timestamp 1604681595
transform 1 0 4968 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_53
timestamp 1604681595
transform 1 0 5980 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8372 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_26_66
timestamp 1604681595
transform 1 0 7176 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_74
timestamp 1604681595
transform 1 0 7912 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_71
timestamp 1604681595
transform 1 0 7636 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10488 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_84
timestamp 1604681595
transform 1 0 8832 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_97
timestamp 1604681595
transform 1 0 10028 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_88
timestamp 1604681595
transform 1 0 9200 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_100
timestamp 1604681595
transform 1 0 10304 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 10948 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_105
timestamp 1604681595
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_123
timestamp 1604681595
transform 1 0 12420 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_111
timestamp 1604681595
transform 1 0 11316 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_119
timestamp 1604681595
transform 1 0 12052 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13708 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 13156 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_134
timestamp 1604681595
transform 1 0 13432 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_145
timestamp 1604681595
transform 1 0 14444 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_129
timestamp 1604681595
transform 1 0 12972 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1604681595
transform 1 0 15272 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15548 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_154
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_166
timestamp 1604681595
transform 1 0 16376 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_146
timestamp 1604681595
transform 1 0 14536 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_158
timestamp 1604681595
transform 1 0 15640 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 17388 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18124 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_174
timestamp 1604681595
transform 1 0 17112 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_175
timestamp 1604681595
transform 1 0 17204 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1604681595
transform 1 0 19688 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_193
timestamp 1604681595
transform 1 0 18860 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_201
timestamp 1604681595
transform 1 0 19596 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_206
timestamp 1604681595
transform 1 0 20056 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_201
timestamp 1604681595
transform 1 0 19596 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20332 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 21896 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 21896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_215
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_215
timestamp 1604681595
transform 1 0 20884 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2024 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_9
timestamp 1604681595
transform 1 0 1932 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_16
timestamp 1604681595
transform 1 0 2576 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4876 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_28
timestamp 1604681595
transform 1 0 3680 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_40
timestamp 1604681595
transform 1 0 4784 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_57
timestamp 1604681595
transform 1 0 6348 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1604681595
transform 1 0 7084 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_28_74
timestamp 1604681595
transform 1 0 7912 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_3_
timestamp 1604681595
transform 1 0 10488 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_86
timestamp 1604681595
transform 1 0 9016 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_93
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_101
timestamp 1604681595
transform 1 0 10396 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12052 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_28_111
timestamp 1604681595
transform 1 0 11316 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_5_
timestamp 1604681595
transform 1 0 13616 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_28_128
timestamp 1604681595
transform 1 0 12880 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_145
timestamp 1604681595
transform 1 0 14444 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1604681595
transform 1 0 15364 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_154
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_159
timestamp 1604681595
transform 1 0 15732 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16468 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_28_183
timestamp 1604681595
transform 1 0 17940 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_6_
timestamp 1604681595
transform 1 0 18952 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_28_191
timestamp 1604681595
transform 1 0 18676 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_203
timestamp 1604681595
transform 1 0 19780 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 21896 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_211
timestamp 1604681595
transform 1 0 20516 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1604681595
transform 1 0 1564 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 2668 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_9
timestamp 1604681595
transform 1 0 1932 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_33
timestamp 1604681595
transform 1 0 4140 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5428 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_45
timestamp 1604681595
transform 1 0 5244 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_53
timestamp 1604681595
transform 1 0 5980 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 8372 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_29_71
timestamp 1604681595
transform 1 0 7636 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10580 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_29_95
timestamp 1604681595
transform 1 0 9844 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_112
timestamp 1604681595
transform 1 0 11408 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1604681595
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_4_
timestamp 1604681595
transform 1 0 14352 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_29_132
timestamp 1604681595
transform 1 0 13248 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15916 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_29_153
timestamp 1604681595
transform 1 0 15180 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_170
timestamp 1604681595
transform 1 0 16744 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_182
timestamp 1604681595
transform 1 0 17848 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 19596 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_29_193
timestamp 1604681595
transform 1 0 18860 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_210
timestamp 1604681595
transform 1 0 20424 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_222
timestamp 1604681595
transform 1 0 21528 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1604681595
transform 1 0 2852 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1604681595
transform 1 0 1748 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_11
timestamp 1604681595
transform 1 0 2116 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_23
timestamp 1604681595
transform 1 0 3220 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_36
timestamp 1604681595
transform 1 0 4416 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5612 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_30_48
timestamp 1604681595
transform 1 0 5520 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7820 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_30_65
timestamp 1604681595
transform 1 0 7084 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_82
timestamp 1604681595
transform 1 0 8648 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1604681595
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11868 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_30_109
timestamp 1604681595
transform 1 0 11132 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1604681595
transform 1 0 14076 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_133
timestamp 1604681595
transform 1 0 13340 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_145
timestamp 1604681595
transform 1 0 14444 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_163
timestamp 1604681595
transform 1 0 16100 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1604681595
transform 1 0 16928 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18032 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_30_171
timestamp 1604681595
transform 1 0 16836 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_176
timestamp 1604681595
transform 1 0 17296 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1604681595
transform 1 0 19688 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_193
timestamp 1604681595
transform 1 0 18860 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_201
timestamp 1604681595
transform 1 0 19596 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_206
timestamp 1604681595
transform 1 0 20056 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 21896 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1604681595
transform 1 0 2852 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1604681595
transform 1 0 1748 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_11
timestamp 1604681595
transform 1 0 2116 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4784 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_23
timestamp 1604681595
transform 1 0 3220 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_35
timestamp 1604681595
transform 1 0 4324 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_39
timestamp 1604681595
transform 1 0 4692 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_46
timestamp 1604681595
transform 1 0 5336 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_58
timestamp 1604681595
transform 1 0 6440 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 8648 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_31_71
timestamp 1604681595
transform 1 0 7636 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_79
timestamp 1604681595
transform 1 0 8372 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1604681595
transform 1 0 10212 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_31_91
timestamp 1604681595
transform 1 0 9476 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1604681595
transform 1 0 12512 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_108
timestamp 1604681595
transform 1 0 11040 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_120
timestamp 1604681595
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 13616 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_31_128
timestamp 1604681595
transform 1 0 12880 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 15824 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_31_152
timestamp 1604681595
transform 1 0 15088 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_169
timestamp 1604681595
transform 1 0 16652 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_181
timestamp 1604681595
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 19596 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_31_193
timestamp 1604681595
transform 1 0 18860 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 21896 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_210
timestamp 1604681595
transform 1 0 20424 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_222
timestamp 1604681595
transform 1 0 21528 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1604681595
transform 1 0 2852 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1604681595
transform 1 0 1748 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_11
timestamp 1604681595
transform 1 0 2116 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_23
timestamp 1604681595
transform 1 0 3220 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_36
timestamp 1604681595
transform 1 0 4416 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6716 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1604681595
transform 1 0 5152 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_32_53
timestamp 1604681595
transform 1 0 5980 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_77
timestamp 1604681595
transform 1 0 8188 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_89
timestamp 1604681595
transform 1 0 9292 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 12236 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_32_109
timestamp 1604681595
transform 1 0 11132 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_137
timestamp 1604681595
transform 1 0 13708 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_149
timestamp 1604681595
transform 1 0 14812 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 17480 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_32_170
timestamp 1604681595
transform 1 0 16744 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_187
timestamp 1604681595
transform 1 0 18308 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19044 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_32_204
timestamp 1604681595
transform 1 0 19872 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 21896 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_212
timestamp 1604681595
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1604681595
transform 1 0 2852 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1604681595
transform 1 0 1748 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_11
timestamp 1604681595
transform 1 0 2116 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1604681595
transform 1 0 4048 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 3956 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_23
timestamp 1604681595
transform 1 0 3220 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_36
timestamp 1604681595
transform 1 0 4416 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1604681595
transform 1 0 5152 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_48
timestamp 1604681595
transform 1 0 5520 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_60
timestamp 1604681595
transform 1 0 6624 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1604681595
transform 1 0 8004 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1604681595
transform 1 0 6900 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_67
timestamp 1604681595
transform 1 0 7268 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_79
timestamp 1604681595
transform 1 0 8372 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1604681595
transform 1 0 9844 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9660 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_91
timestamp 1604681595
transform 1 0 9476 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_94
timestamp 1604681595
transform 1 0 9752 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_99
timestamp 1604681595
transform 1 0 10212 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 10948 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 12512 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_116
timestamp 1604681595
transform 1 0 11776 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_125
timestamp 1604681595
transform 1 0 12604 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 13064 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_33_129
timestamp 1604681595
transform 1 0 12972 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_139
timestamp 1604681595
transform 1 0 13892 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 15456 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 15364 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_151
timestamp 1604681595
transform 1 0 14996 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_165
timestamp 1604681595
transform 1 0 16284 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604681595
transform 1 0 17112 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18308 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 18216 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_173
timestamp 1604681595
transform 1 0 17020 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_178
timestamp 1604681595
transform 1 0 17480 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1604681595
transform 1 0 19964 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_196
timestamp 1604681595
transform 1 0 19136 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_204
timestamp 1604681595
transform 1 0 19872 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 21896 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 21068 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_209
timestamp 1604681595
transform 1 0 20332 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_218
timestamp 1604681595
transform 1 0 21160 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_222
timestamp 1604681595
transform 1 0 21528 0 1 20128
box -38 -48 130 592
<< labels >>
rlabel metal3 s 0 22176 480 22296 6 SC_IN_BOT
port 0 nsew default input
rlabel metal3 s 22520 22584 23000 22704 6 SC_IN_TOP
port 1 nsew default input
rlabel metal3 s 0 22584 480 22704 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 20074 22520 20130 23000 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal2 s 202 0 258 480 6 bottom_left_grid_pin_42_
port 4 nsew default input
rlabel metal2 s 662 0 718 480 6 bottom_left_grid_pin_43_
port 5 nsew default input
rlabel metal2 s 1122 0 1178 480 6 bottom_left_grid_pin_44_
port 6 nsew default input
rlabel metal2 s 1582 0 1638 480 6 bottom_left_grid_pin_45_
port 7 nsew default input
rlabel metal2 s 2042 0 2098 480 6 bottom_left_grid_pin_46_
port 8 nsew default input
rlabel metal2 s 2594 0 2650 480 6 bottom_left_grid_pin_47_
port 9 nsew default input
rlabel metal2 s 3054 0 3110 480 6 bottom_left_grid_pin_48_
port 10 nsew default input
rlabel metal2 s 3514 0 3570 480 6 bottom_left_grid_pin_49_
port 11 nsew default input
rlabel metal2 s 8574 22520 8630 23000 6 ccff_head
port 12 nsew default input
rlabel metal2 s 14370 22520 14426 23000 6 ccff_tail
port 13 nsew default tristate
rlabel metal3 s 0 3680 480 3800 6 chanx_left_in[0]
port 14 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_left_in[10]
port 15 nsew default input
rlabel metal3 s 0 8576 480 8696 6 chanx_left_in[11]
port 16 nsew default input
rlabel metal3 s 0 9120 480 9240 6 chanx_left_in[12]
port 17 nsew default input
rlabel metal3 s 0 9528 480 9648 6 chanx_left_in[13]
port 18 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[14]
port 19 nsew default input
rlabel metal3 s 0 10480 480 10600 6 chanx_left_in[15]
port 20 nsew default input
rlabel metal3 s 0 10888 480 11008 6 chanx_left_in[16]
port 21 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[17]
port 22 nsew default input
rlabel metal3 s 0 11840 480 11960 6 chanx_left_in[18]
port 23 nsew default input
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[19]
port 24 nsew default input
rlabel metal3 s 0 4088 480 4208 6 chanx_left_in[1]
port 25 nsew default input
rlabel metal3 s 0 4632 480 4752 6 chanx_left_in[2]
port 26 nsew default input
rlabel metal3 s 0 5040 480 5160 6 chanx_left_in[3]
port 27 nsew default input
rlabel metal3 s 0 5448 480 5568 6 chanx_left_in[4]
port 28 nsew default input
rlabel metal3 s 0 5992 480 6112 6 chanx_left_in[5]
port 29 nsew default input
rlabel metal3 s 0 6400 480 6520 6 chanx_left_in[6]
port 30 nsew default input
rlabel metal3 s 0 6808 480 6928 6 chanx_left_in[7]
port 31 nsew default input
rlabel metal3 s 0 7352 480 7472 6 chanx_left_in[8]
port 32 nsew default input
rlabel metal3 s 0 7760 480 7880 6 chanx_left_in[9]
port 33 nsew default input
rlabel metal3 s 0 12656 480 12776 6 chanx_left_out[0]
port 34 nsew default tristate
rlabel metal3 s 0 17144 480 17264 6 chanx_left_out[10]
port 35 nsew default tristate
rlabel metal3 s 0 17688 480 17808 6 chanx_left_out[11]
port 36 nsew default tristate
rlabel metal3 s 0 18096 480 18216 6 chanx_left_out[12]
port 37 nsew default tristate
rlabel metal3 s 0 18504 480 18624 6 chanx_left_out[13]
port 38 nsew default tristate
rlabel metal3 s 0 19048 480 19168 6 chanx_left_out[14]
port 39 nsew default tristate
rlabel metal3 s 0 19456 480 19576 6 chanx_left_out[15]
port 40 nsew default tristate
rlabel metal3 s 0 19864 480 19984 6 chanx_left_out[16]
port 41 nsew default tristate
rlabel metal3 s 0 20408 480 20528 6 chanx_left_out[17]
port 42 nsew default tristate
rlabel metal3 s 0 20816 480 20936 6 chanx_left_out[18]
port 43 nsew default tristate
rlabel metal3 s 0 21224 480 21344 6 chanx_left_out[19]
port 44 nsew default tristate
rlabel metal3 s 0 13200 480 13320 6 chanx_left_out[1]
port 45 nsew default tristate
rlabel metal3 s 0 13608 480 13728 6 chanx_left_out[2]
port 46 nsew default tristate
rlabel metal3 s 0 14016 480 14136 6 chanx_left_out[3]
port 47 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[4]
port 48 nsew default tristate
rlabel metal3 s 0 14968 480 15088 6 chanx_left_out[5]
port 49 nsew default tristate
rlabel metal3 s 0 15376 480 15496 6 chanx_left_out[6]
port 50 nsew default tristate
rlabel metal3 s 0 15784 480 15904 6 chanx_left_out[7]
port 51 nsew default tristate
rlabel metal3 s 0 16328 480 16448 6 chanx_left_out[8]
port 52 nsew default tristate
rlabel metal3 s 0 16736 480 16856 6 chanx_left_out[9]
port 53 nsew default tristate
rlabel metal3 s 22520 3816 23000 3936 6 chanx_right_in[0]
port 54 nsew default input
rlabel metal3 s 22520 8304 23000 8424 6 chanx_right_in[10]
port 55 nsew default input
rlabel metal3 s 22520 8848 23000 8968 6 chanx_right_in[11]
port 56 nsew default input
rlabel metal3 s 22520 9256 23000 9376 6 chanx_right_in[12]
port 57 nsew default input
rlabel metal3 s 22520 9664 23000 9784 6 chanx_right_in[13]
port 58 nsew default input
rlabel metal3 s 22520 10208 23000 10328 6 chanx_right_in[14]
port 59 nsew default input
rlabel metal3 s 22520 10616 23000 10736 6 chanx_right_in[15]
port 60 nsew default input
rlabel metal3 s 22520 11160 23000 11280 6 chanx_right_in[16]
port 61 nsew default input
rlabel metal3 s 22520 11568 23000 11688 6 chanx_right_in[17]
port 62 nsew default input
rlabel metal3 s 22520 11976 23000 12096 6 chanx_right_in[18]
port 63 nsew default input
rlabel metal3 s 22520 12520 23000 12640 6 chanx_right_in[19]
port 64 nsew default input
rlabel metal3 s 22520 4224 23000 4344 6 chanx_right_in[1]
port 65 nsew default input
rlabel metal3 s 22520 4632 23000 4752 6 chanx_right_in[2]
port 66 nsew default input
rlabel metal3 s 22520 5176 23000 5296 6 chanx_right_in[3]
port 67 nsew default input
rlabel metal3 s 22520 5584 23000 5704 6 chanx_right_in[4]
port 68 nsew default input
rlabel metal3 s 22520 5992 23000 6112 6 chanx_right_in[5]
port 69 nsew default input
rlabel metal3 s 22520 6536 23000 6656 6 chanx_right_in[6]
port 70 nsew default input
rlabel metal3 s 22520 6944 23000 7064 6 chanx_right_in[7]
port 71 nsew default input
rlabel metal3 s 22520 7488 23000 7608 6 chanx_right_in[8]
port 72 nsew default input
rlabel metal3 s 22520 7896 23000 8016 6 chanx_right_in[9]
port 73 nsew default input
rlabel metal3 s 22520 12928 23000 13048 6 chanx_right_out[0]
port 74 nsew default tristate
rlabel metal3 s 22520 17552 23000 17672 6 chanx_right_out[10]
port 75 nsew default tristate
rlabel metal3 s 22520 17960 23000 18080 6 chanx_right_out[11]
port 76 nsew default tristate
rlabel metal3 s 22520 18504 23000 18624 6 chanx_right_out[12]
port 77 nsew default tristate
rlabel metal3 s 22520 18912 23000 19032 6 chanx_right_out[13]
port 78 nsew default tristate
rlabel metal3 s 22520 19320 23000 19440 6 chanx_right_out[14]
port 79 nsew default tristate
rlabel metal3 s 22520 19864 23000 19984 6 chanx_right_out[15]
port 80 nsew default tristate
rlabel metal3 s 22520 20272 23000 20392 6 chanx_right_out[16]
port 81 nsew default tristate
rlabel metal3 s 22520 20816 23000 20936 6 chanx_right_out[17]
port 82 nsew default tristate
rlabel metal3 s 22520 21224 23000 21344 6 chanx_right_out[18]
port 83 nsew default tristate
rlabel metal3 s 22520 21632 23000 21752 6 chanx_right_out[19]
port 84 nsew default tristate
rlabel metal3 s 22520 13472 23000 13592 6 chanx_right_out[1]
port 85 nsew default tristate
rlabel metal3 s 22520 13880 23000 14000 6 chanx_right_out[2]
port 86 nsew default tristate
rlabel metal3 s 22520 14288 23000 14408 6 chanx_right_out[3]
port 87 nsew default tristate
rlabel metal3 s 22520 14832 23000 14952 6 chanx_right_out[4]
port 88 nsew default tristate
rlabel metal3 s 22520 15240 23000 15360 6 chanx_right_out[5]
port 89 nsew default tristate
rlabel metal3 s 22520 15648 23000 15768 6 chanx_right_out[6]
port 90 nsew default tristate
rlabel metal3 s 22520 16192 23000 16312 6 chanx_right_out[7]
port 91 nsew default tristate
rlabel metal3 s 22520 16600 23000 16720 6 chanx_right_out[8]
port 92 nsew default tristate
rlabel metal3 s 22520 17144 23000 17264 6 chanx_right_out[9]
port 93 nsew default tristate
rlabel metal2 s 3974 0 4030 480 6 chany_bottom_in[0]
port 94 nsew default input
rlabel metal2 s 8758 0 8814 480 6 chany_bottom_in[10]
port 95 nsew default input
rlabel metal2 s 9218 0 9274 480 6 chany_bottom_in[11]
port 96 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chany_bottom_in[12]
port 97 nsew default input
rlabel metal2 s 10230 0 10286 480 6 chany_bottom_in[13]
port 98 nsew default input
rlabel metal2 s 10690 0 10746 480 6 chany_bottom_in[14]
port 99 nsew default input
rlabel metal2 s 11150 0 11206 480 6 chany_bottom_in[15]
port 100 nsew default input
rlabel metal2 s 11702 0 11758 480 6 chany_bottom_in[16]
port 101 nsew default input
rlabel metal2 s 12162 0 12218 480 6 chany_bottom_in[17]
port 102 nsew default input
rlabel metal2 s 12622 0 12678 480 6 chany_bottom_in[18]
port 103 nsew default input
rlabel metal2 s 13082 0 13138 480 6 chany_bottom_in[19]
port 104 nsew default input
rlabel metal2 s 4434 0 4490 480 6 chany_bottom_in[1]
port 105 nsew default input
rlabel metal2 s 4986 0 5042 480 6 chany_bottom_in[2]
port 106 nsew default input
rlabel metal2 s 5446 0 5502 480 6 chany_bottom_in[3]
port 107 nsew default input
rlabel metal2 s 5906 0 5962 480 6 chany_bottom_in[4]
port 108 nsew default input
rlabel metal2 s 6366 0 6422 480 6 chany_bottom_in[5]
port 109 nsew default input
rlabel metal2 s 6826 0 6882 480 6 chany_bottom_in[6]
port 110 nsew default input
rlabel metal2 s 7378 0 7434 480 6 chany_bottom_in[7]
port 111 nsew default input
rlabel metal2 s 7838 0 7894 480 6 chany_bottom_in[8]
port 112 nsew default input
rlabel metal2 s 8298 0 8354 480 6 chany_bottom_in[9]
port 113 nsew default input
rlabel metal2 s 13542 0 13598 480 6 chany_bottom_out[0]
port 114 nsew default tristate
rlabel metal2 s 18326 0 18382 480 6 chany_bottom_out[10]
port 115 nsew default tristate
rlabel metal2 s 18878 0 18934 480 6 chany_bottom_out[11]
port 116 nsew default tristate
rlabel metal2 s 19338 0 19394 480 6 chany_bottom_out[12]
port 117 nsew default tristate
rlabel metal2 s 19798 0 19854 480 6 chany_bottom_out[13]
port 118 nsew default tristate
rlabel metal2 s 20258 0 20314 480 6 chany_bottom_out[14]
port 119 nsew default tristate
rlabel metal2 s 20718 0 20774 480 6 chany_bottom_out[15]
port 120 nsew default tristate
rlabel metal2 s 21270 0 21326 480 6 chany_bottom_out[16]
port 121 nsew default tristate
rlabel metal2 s 21730 0 21786 480 6 chany_bottom_out[17]
port 122 nsew default tristate
rlabel metal2 s 22190 0 22246 480 6 chany_bottom_out[18]
port 123 nsew default tristate
rlabel metal2 s 22650 0 22706 480 6 chany_bottom_out[19]
port 124 nsew default tristate
rlabel metal2 s 14094 0 14150 480 6 chany_bottom_out[1]
port 125 nsew default tristate
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_out[2]
port 126 nsew default tristate
rlabel metal2 s 15014 0 15070 480 6 chany_bottom_out[3]
port 127 nsew default tristate
rlabel metal2 s 15474 0 15530 480 6 chany_bottom_out[4]
port 128 nsew default tristate
rlabel metal2 s 15934 0 15990 480 6 chany_bottom_out[5]
port 129 nsew default tristate
rlabel metal2 s 16486 0 16542 480 6 chany_bottom_out[6]
port 130 nsew default tristate
rlabel metal2 s 16946 0 17002 480 6 chany_bottom_out[7]
port 131 nsew default tristate
rlabel metal2 s 17406 0 17462 480 6 chany_bottom_out[8]
port 132 nsew default tristate
rlabel metal2 s 17866 0 17922 480 6 chany_bottom_out[9]
port 133 nsew default tristate
rlabel metal3 s 0 144 480 264 6 left_bottom_grid_pin_34_
port 134 nsew default input
rlabel metal3 s 0 552 480 672 6 left_bottom_grid_pin_35_
port 135 nsew default input
rlabel metal3 s 0 960 480 1080 6 left_bottom_grid_pin_36_
port 136 nsew default input
rlabel metal3 s 0 1368 480 1488 6 left_bottom_grid_pin_37_
port 137 nsew default input
rlabel metal3 s 0 1912 480 2032 6 left_bottom_grid_pin_38_
port 138 nsew default input
rlabel metal3 s 0 2320 480 2440 6 left_bottom_grid_pin_39_
port 139 nsew default input
rlabel metal3 s 0 2728 480 2848 6 left_bottom_grid_pin_40_
port 140 nsew default input
rlabel metal3 s 0 3272 480 3392 6 left_bottom_grid_pin_41_
port 141 nsew default input
rlabel metal3 s 0 21768 480 21888 6 left_top_grid_pin_1_
port 142 nsew default input
rlabel metal2 s 2870 22520 2926 23000 6 prog_clk
port 143 nsew default input
rlabel metal3 s 22520 144 23000 264 6 right_bottom_grid_pin_34_
port 144 nsew default input
rlabel metal3 s 22520 552 23000 672 6 right_bottom_grid_pin_35_
port 145 nsew default input
rlabel metal3 s 22520 960 23000 1080 6 right_bottom_grid_pin_36_
port 146 nsew default input
rlabel metal3 s 22520 1504 23000 1624 6 right_bottom_grid_pin_37_
port 147 nsew default input
rlabel metal3 s 22520 1912 23000 2032 6 right_bottom_grid_pin_38_
port 148 nsew default input
rlabel metal3 s 22520 2320 23000 2440 6 right_bottom_grid_pin_39_
port 149 nsew default input
rlabel metal3 s 22520 2864 23000 2984 6 right_bottom_grid_pin_40_
port 150 nsew default input
rlabel metal3 s 22520 3272 23000 3392 6 right_bottom_grid_pin_41_
port 151 nsew default input
rlabel metal3 s 22520 22176 23000 22296 6 right_top_grid_pin_1_
port 152 nsew default input
rlabel metal4 s 4409 2128 4729 20720 6 VPWR
port 153 nsew default input
rlabel metal4 s 7875 2128 8195 20720 6 VGND
port 154 nsew default input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
