magic
tech sky130A
magscale 1 2
timestamp 1606225624
<< locali >>
rect 6193 14263 6227 14501
rect 7205 14263 7239 14365
rect 8769 13243 8803 13481
rect 6561 12631 6595 12937
rect 6653 12767 6687 12937
rect 6653 12733 6745 12767
rect 10425 12631 10459 12937
rect 6561 12597 6653 12631
rect 3801 12087 3835 12257
rect 11621 12087 11655 12189
rect 8309 11611 8343 11713
rect 12207 11169 12299 11203
rect 12265 10999 12299 11169
rect 13185 10999 13219 11101
rect 3249 10455 3283 10625
rect 8401 10455 8435 10693
rect 9321 10455 9355 10625
rect 14289 10455 14323 10761
rect 9815 9605 9873 9639
rect 11897 9503 11931 9673
rect 3249 7395 3283 7497
rect 12173 7259 12207 7497
rect 13277 7327 13311 7497
rect 14381 7191 14415 7497
rect 5365 6851 5399 6953
rect 9505 6851 9539 6953
rect 4997 6171 5031 6341
rect 10149 6103 10183 6409
rect 12173 6239 12207 6341
rect 13277 6239 13311 6341
rect 11713 6205 11805 6239
rect 11713 6103 11747 6205
rect 3801 5559 3835 5865
rect 9137 5627 9171 5865
rect 11621 5559 11655 5865
rect 11563 5525 11655 5559
rect 12541 5559 12575 5865
rect 8309 5015 8343 5253
rect 9965 5015 9999 5253
rect 8309 4471 8343 4573
rect 5583 4233 5675 4267
rect 5549 3927 5583 4097
rect 5641 3927 5675 4233
rect 9321 3995 9355 4233
rect 10425 3927 10459 4097
rect 12541 3485 12633 3519
rect 11621 3383 11655 3485
rect 12541 3451 12575 3485
rect 8769 2975 8803 3077
rect 2881 2295 2915 2533
rect 5641 2431 5675 2601
rect 9539 2533 9597 2567
rect 13645 2499 13679 2601
rect 8125 935 8159 1649
<< viali >>
rect 4445 15657 4479 15691
rect 9321 15657 9355 15691
rect 9965 15657 9999 15691
rect 10517 15657 10551 15691
rect 6285 15589 6319 15623
rect 3249 15521 3283 15555
rect 4261 15521 4295 15555
rect 4813 15521 4847 15555
rect 6193 15521 6227 15555
rect 7481 15521 7515 15555
rect 8493 15521 8527 15555
rect 8585 15521 8619 15555
rect 9137 15521 9171 15555
rect 9781 15521 9815 15555
rect 10333 15521 10367 15555
rect 6469 15453 6503 15487
rect 7573 15453 7607 15487
rect 7665 15453 7699 15487
rect 8677 15453 8711 15487
rect 4997 15385 5031 15419
rect 3433 15317 3467 15351
rect 5825 15317 5859 15351
rect 7113 15317 7147 15351
rect 8125 15317 8159 15351
rect 5365 15113 5399 15147
rect 9689 15113 9723 15147
rect 2973 15045 3007 15079
rect 3525 15045 3559 15079
rect 4813 15045 4847 15079
rect 7389 15045 7423 15079
rect 6193 14977 6227 15011
rect 6377 14977 6411 15011
rect 8217 14977 8251 15011
rect 9229 14977 9263 15011
rect 10149 14977 10183 15011
rect 10333 14977 10367 15011
rect 2237 14909 2271 14943
rect 2789 14909 2823 14943
rect 3341 14909 3375 14943
rect 3893 14909 3927 14943
rect 4169 14909 4203 14943
rect 4629 14909 4663 14943
rect 5181 14909 5215 14943
rect 6837 14909 6871 14943
rect 7573 14909 7607 14943
rect 8125 14909 8159 14943
rect 10701 14909 10735 14943
rect 9137 14841 9171 14875
rect 2421 14773 2455 14807
rect 5733 14773 5767 14807
rect 6101 14773 6135 14807
rect 7021 14773 7055 14807
rect 7665 14773 7699 14807
rect 8033 14773 8067 14807
rect 8677 14773 8711 14807
rect 9045 14773 9079 14807
rect 10057 14773 10091 14807
rect 10885 14773 10919 14807
rect 11253 14773 11287 14807
rect 2605 14569 2639 14603
rect 5733 14569 5767 14603
rect 5825 14569 5859 14603
rect 8861 14569 8895 14603
rect 9689 14569 9723 14603
rect 6193 14501 6227 14535
rect 6745 14501 6779 14535
rect 6837 14501 6871 14535
rect 8769 14501 8803 14535
rect 10057 14501 10091 14535
rect 11069 14501 11103 14535
rect 1869 14433 1903 14467
rect 2421 14433 2455 14467
rect 2973 14433 3007 14467
rect 4721 14433 4755 14467
rect 3157 14365 3191 14399
rect 4813 14365 4847 14399
rect 4997 14365 5031 14399
rect 6009 14365 6043 14399
rect 2053 14297 2087 14331
rect 7757 14433 7791 14467
rect 7849 14433 7883 14467
rect 11161 14433 11195 14467
rect 11713 14433 11747 14467
rect 12449 14433 12483 14467
rect 6929 14365 6963 14399
rect 7205 14365 7239 14399
rect 8033 14365 8067 14399
rect 9045 14365 9079 14399
rect 10149 14365 10183 14399
rect 10333 14365 10367 14399
rect 11253 14365 11287 14399
rect 7389 14297 7423 14331
rect 10701 14297 10735 14331
rect 4353 14229 4387 14263
rect 5365 14229 5399 14263
rect 6193 14229 6227 14263
rect 6377 14229 6411 14263
rect 7205 14229 7239 14263
rect 8401 14229 8435 14263
rect 11897 14229 11931 14263
rect 12265 14229 12299 14263
rect 5733 14025 5767 14059
rect 6837 14025 6871 14059
rect 7849 14025 7883 14059
rect 9873 14025 9907 14059
rect 12633 14025 12667 14059
rect 1777 13957 1811 13991
rect 8861 13957 8895 13991
rect 10885 13957 10919 13991
rect 3065 13889 3099 13923
rect 4261 13889 4295 13923
rect 5273 13889 5307 13923
rect 6285 13889 6319 13923
rect 7297 13889 7331 13923
rect 7481 13889 7515 13923
rect 8309 13889 8343 13923
rect 8401 13889 8435 13923
rect 9505 13889 9539 13923
rect 10425 13889 10459 13923
rect 11529 13889 11563 13923
rect 1593 13821 1627 13855
rect 2145 13821 2179 13855
rect 2421 13821 2455 13855
rect 2881 13821 2915 13855
rect 5181 13821 5215 13855
rect 6193 13821 6227 13855
rect 9229 13821 9263 13855
rect 10333 13821 10367 13855
rect 11345 13821 11379 13855
rect 12449 13821 12483 13855
rect 4077 13753 4111 13787
rect 6101 13753 6135 13787
rect 7205 13753 7239 13787
rect 8217 13753 8251 13787
rect 10241 13753 10275 13787
rect 3709 13685 3743 13719
rect 4169 13685 4203 13719
rect 4721 13685 4755 13719
rect 5089 13685 5123 13719
rect 9321 13685 9355 13719
rect 11253 13685 11287 13719
rect 11897 13685 11931 13719
rect 3433 13481 3467 13515
rect 4629 13481 4663 13515
rect 5273 13481 5307 13515
rect 5641 13481 5675 13515
rect 8769 13481 8803 13515
rect 10149 13481 10183 13515
rect 11069 13481 11103 13515
rect 11713 13481 11747 13515
rect 12173 13481 12207 13515
rect 8309 13413 8343 13447
rect 1501 13345 1535 13379
rect 2237 13345 2271 13379
rect 2513 13345 2547 13379
rect 3341 13345 3375 13379
rect 6285 13345 6319 13379
rect 6552 13345 6586 13379
rect 8401 13345 8435 13379
rect 1685 13277 1719 13311
rect 3617 13277 3651 13311
rect 4721 13277 4755 13311
rect 4905 13277 4939 13311
rect 5733 13277 5767 13311
rect 5825 13277 5859 13311
rect 8585 13277 8619 13311
rect 10057 13413 10091 13447
rect 14013 13413 14047 13447
rect 8953 13345 8987 13379
rect 12081 13345 12115 13379
rect 13093 13345 13127 13379
rect 13737 13345 13771 13379
rect 10333 13277 10367 13311
rect 11161 13277 11195 13311
rect 11345 13277 11379 13311
rect 12265 13277 12299 13311
rect 13185 13277 13219 13311
rect 13369 13277 13403 13311
rect 7941 13209 7975 13243
rect 8769 13209 8803 13243
rect 9137 13209 9171 13243
rect 9689 13209 9723 13243
rect 12725 13209 12759 13243
rect 2973 13141 3007 13175
rect 4261 13141 4295 13175
rect 7665 13141 7699 13175
rect 10701 13141 10735 13175
rect 6561 12937 6595 12971
rect 2329 12801 2363 12835
rect 3157 12801 3191 12835
rect 3249 12801 3283 12835
rect 4169 12801 4203 12835
rect 4353 12801 4387 12835
rect 5273 12801 5307 12835
rect 6377 12801 6411 12835
rect 4077 12733 4111 12767
rect 5089 12733 5123 12767
rect 6193 12733 6227 12767
rect 3065 12665 3099 12699
rect 6101 12665 6135 12699
rect 6653 12937 6687 12971
rect 8217 12937 8251 12971
rect 9505 12937 9539 12971
rect 10425 12937 10459 12971
rect 11713 12937 11747 12971
rect 13461 12937 13495 12971
rect 8493 12869 8527 12903
rect 8953 12801 8987 12835
rect 9045 12801 9079 12835
rect 10057 12801 10091 12835
rect 6745 12733 6779 12767
rect 6837 12733 6871 12767
rect 7093 12733 7127 12767
rect 9873 12733 9907 12767
rect 8861 12665 8895 12699
rect 10517 12869 10551 12903
rect 12449 12869 12483 12903
rect 10977 12801 11011 12835
rect 11161 12801 11195 12835
rect 13093 12801 13127 12835
rect 14013 12801 14047 12835
rect 10885 12733 10919 12767
rect 11529 12733 11563 12767
rect 12265 12733 12299 12767
rect 12909 12733 12943 12767
rect 13829 12733 13863 12767
rect 1685 12597 1719 12631
rect 2053 12597 2087 12631
rect 2145 12597 2179 12631
rect 2697 12597 2731 12631
rect 3709 12597 3743 12631
rect 4721 12597 4755 12631
rect 5181 12597 5215 12631
rect 5733 12597 5767 12631
rect 6653 12597 6687 12631
rect 9965 12597 9999 12631
rect 10425 12597 10459 12631
rect 12081 12597 12115 12631
rect 12817 12597 12851 12631
rect 13921 12597 13955 12631
rect 1961 12393 1995 12427
rect 2973 12393 3007 12427
rect 3433 12393 3467 12427
rect 4077 12393 4111 12427
rect 4537 12393 4571 12427
rect 9689 12393 9723 12427
rect 12081 12393 12115 12427
rect 13185 12393 13219 12427
rect 13737 12393 13771 12427
rect 14197 12393 14231 12427
rect 4445 12325 4479 12359
rect 5356 12325 5390 12359
rect 6990 12325 7024 12359
rect 10057 12325 10091 12359
rect 1869 12257 1903 12291
rect 2329 12257 2363 12291
rect 3341 12257 3375 12291
rect 3801 12257 3835 12291
rect 5089 12257 5123 12291
rect 6745 12257 6779 12291
rect 8769 12257 8803 12291
rect 10149 12257 10183 12291
rect 11069 12257 11103 12291
rect 12173 12257 12207 12291
rect 13093 12257 13127 12291
rect 14105 12257 14139 12291
rect 2421 12189 2455 12223
rect 2605 12189 2639 12223
rect 3617 12189 3651 12223
rect 4721 12189 4755 12223
rect 8861 12189 8895 12223
rect 9045 12189 9079 12223
rect 10333 12189 10367 12223
rect 11161 12189 11195 12223
rect 11345 12189 11379 12223
rect 11621 12189 11655 12223
rect 12357 12189 12391 12223
rect 13277 12189 13311 12223
rect 14289 12189 14323 12223
rect 14749 12189 14783 12223
rect 10701 12121 10735 12155
rect 1685 12053 1719 12087
rect 3801 12053 3835 12087
rect 6469 12053 6503 12087
rect 8125 12053 8159 12087
rect 8401 12053 8435 12087
rect 11621 12053 11655 12087
rect 11713 12053 11747 12087
rect 12725 12053 12759 12087
rect 2053 11849 2087 11883
rect 9873 11849 9907 11883
rect 11529 11849 11563 11883
rect 14473 11849 14507 11883
rect 6469 11781 6503 11815
rect 2697 11713 2731 11747
rect 3709 11713 3743 11747
rect 4537 11713 4571 11747
rect 4721 11713 4755 11747
rect 6837 11713 6871 11747
rect 8309 11713 8343 11747
rect 13001 11713 13035 11747
rect 14013 11713 14047 11747
rect 15025 11713 15059 11747
rect 1961 11645 1995 11679
rect 5089 11645 5123 11679
rect 8493 11645 8527 11679
rect 8749 11645 8783 11679
rect 10149 11645 10183 11679
rect 13829 11645 13863 11679
rect 13921 11645 13955 11679
rect 14933 11645 14967 11679
rect 2421 11577 2455 11611
rect 3433 11577 3467 11611
rect 4445 11577 4479 11611
rect 5356 11577 5390 11611
rect 7082 11577 7116 11611
rect 8309 11577 8343 11611
rect 10416 11577 10450 11611
rect 12817 11577 12851 11611
rect 1777 11509 1811 11543
rect 2513 11509 2547 11543
rect 3065 11509 3099 11543
rect 3525 11509 3559 11543
rect 4077 11509 4111 11543
rect 8217 11509 8251 11543
rect 11805 11509 11839 11543
rect 12449 11509 12483 11543
rect 12909 11509 12943 11543
rect 13461 11509 13495 11543
rect 14841 11509 14875 11543
rect 1961 11305 1995 11339
rect 2329 11305 2363 11339
rect 3341 11305 3375 11339
rect 5733 11305 5767 11339
rect 7389 11305 7423 11339
rect 9045 11305 9079 11339
rect 9321 11305 9355 11339
rect 11345 11305 11379 11339
rect 12357 11305 12391 11339
rect 12817 11305 12851 11339
rect 13369 11305 13403 11339
rect 13737 11305 13771 11339
rect 3433 11237 3467 11271
rect 6276 11237 6310 11271
rect 11713 11237 11747 11271
rect 12725 11237 12759 11271
rect 14381 11237 14415 11271
rect 4620 11169 4654 11203
rect 6009 11169 6043 11203
rect 7921 11169 7955 11203
rect 9505 11169 9539 11203
rect 9956 11169 9990 11203
rect 11805 11169 11839 11203
rect 12173 11169 12207 11203
rect 13829 11169 13863 11203
rect 15025 11169 15059 11203
rect 1501 11101 1535 11135
rect 2421 11101 2455 11135
rect 2513 11101 2547 11135
rect 3617 11101 3651 11135
rect 4353 11101 4387 11135
rect 7665 11101 7699 11135
rect 9689 11101 9723 11135
rect 11897 11101 11931 11135
rect 1869 11033 1903 11067
rect 2973 11033 3007 11067
rect 13001 11101 13035 11135
rect 13185 11101 13219 11135
rect 13921 11101 13955 11135
rect 11069 10965 11103 10999
rect 12265 10965 12299 10999
rect 14841 11033 14875 11067
rect 13185 10965 13219 10999
rect 14289 10761 14323 10795
rect 4813 10693 4847 10727
rect 6469 10693 6503 10727
rect 8401 10693 8435 10727
rect 8493 10693 8527 10727
rect 11161 10693 11195 10727
rect 12449 10693 12483 10727
rect 13461 10693 13495 10727
rect 1869 10625 1903 10659
rect 2053 10625 2087 10659
rect 2881 10625 2915 10659
rect 3065 10625 3099 10659
rect 3249 10625 3283 10659
rect 6837 10625 6871 10659
rect 1777 10557 1811 10591
rect 3433 10557 3467 10591
rect 5089 10557 5123 10591
rect 5356 10557 5390 10591
rect 3700 10489 3734 10523
rect 7104 10489 7138 10523
rect 9045 10625 9079 10659
rect 9321 10625 9355 10659
rect 9505 10625 9539 10659
rect 11713 10625 11747 10659
rect 13001 10625 13035 10659
rect 13921 10625 13955 10659
rect 14013 10625 14047 10659
rect 11529 10557 11563 10591
rect 12817 10557 12851 10591
rect 9772 10489 9806 10523
rect 13829 10489 13863 10523
rect 15025 10625 15059 10659
rect 14933 10489 14967 10523
rect 1409 10421 1443 10455
rect 2421 10421 2455 10455
rect 2789 10421 2823 10455
rect 3249 10421 3283 10455
rect 8217 10421 8251 10455
rect 8401 10421 8435 10455
rect 8861 10421 8895 10455
rect 8953 10421 8987 10455
rect 9321 10421 9355 10455
rect 10885 10421 10919 10455
rect 11621 10421 11655 10455
rect 12909 10421 12943 10455
rect 14289 10421 14323 10455
rect 14473 10421 14507 10455
rect 14841 10421 14875 10455
rect 5549 10217 5583 10251
rect 7481 10217 7515 10251
rect 9321 10217 9355 10251
rect 12725 10217 12759 10251
rect 13461 10217 13495 10251
rect 14013 10217 14047 10251
rect 1869 10149 1903 10183
rect 2596 10149 2630 10183
rect 4436 10149 4470 10183
rect 8208 10149 8242 10183
rect 1593 10081 1627 10115
rect 4169 10081 4203 10115
rect 6081 10081 6115 10115
rect 7941 10081 7975 10115
rect 9689 10081 9723 10115
rect 9956 10081 9990 10115
rect 11601 10081 11635 10115
rect 13369 10081 13403 10115
rect 14381 10081 14415 10115
rect 2329 10013 2363 10047
rect 5825 10013 5859 10047
rect 11345 10013 11379 10047
rect 13553 10013 13587 10047
rect 14473 10013 14507 10047
rect 14565 10013 14599 10047
rect 3709 9877 3743 9911
rect 7205 9877 7239 9911
rect 11069 9877 11103 9911
rect 13001 9877 13035 9911
rect 11897 9673 11931 9707
rect 7021 9605 7055 9639
rect 9781 9605 9815 9639
rect 9873 9605 9907 9639
rect 1777 9537 1811 9571
rect 5089 9537 5123 9571
rect 7665 9537 7699 9571
rect 14105 9605 14139 9639
rect 12449 9537 12483 9571
rect 14657 9537 14691 9571
rect 15117 9537 15151 9571
rect 3433 9469 3467 9503
rect 7389 9469 7423 9503
rect 8217 9469 8251 9503
rect 8309 9469 8343 9503
rect 9965 9469 9999 9503
rect 11897 9469 11931 9503
rect 12265 9469 12299 9503
rect 2044 9401 2078 9435
rect 3700 9401 3734 9435
rect 5356 9401 5390 9435
rect 8576 9401 8610 9435
rect 10232 9401 10266 9435
rect 11621 9401 11655 9435
rect 12694 9401 12728 9435
rect 14473 9401 14507 9435
rect 3157 9333 3191 9367
rect 4813 9333 4847 9367
rect 6469 9333 6503 9367
rect 7481 9333 7515 9367
rect 8033 9333 8067 9367
rect 9689 9333 9723 9367
rect 11345 9333 11379 9367
rect 12081 9333 12115 9367
rect 13829 9333 13863 9367
rect 14565 9333 14599 9367
rect 3709 9129 3743 9163
rect 5641 9129 5675 9163
rect 8677 9129 8711 9163
rect 11069 9129 11103 9163
rect 14381 9129 14415 9163
rect 14657 9129 14691 9163
rect 1869 9061 1903 9095
rect 2596 9061 2630 9095
rect 4528 9061 4562 9095
rect 7389 9061 7423 9095
rect 9945 9061 9979 9095
rect 1593 8993 1627 9027
rect 4261 8993 4295 9027
rect 5733 8993 5767 9027
rect 6000 8993 6034 9027
rect 9689 8993 9723 9027
rect 11345 8993 11379 9027
rect 11612 8993 11646 9027
rect 13001 8993 13035 9027
rect 13268 8993 13302 9027
rect 2329 8925 2363 8959
rect 7113 8789 7147 8823
rect 12725 8789 12759 8823
rect 4813 8585 4847 8619
rect 7021 8585 7055 8619
rect 7389 8585 7423 8619
rect 10885 8585 10919 8619
rect 13829 8585 13863 8619
rect 6469 8517 6503 8551
rect 9321 8517 9355 8551
rect 14105 8517 14139 8551
rect 1777 8449 1811 8483
rect 7941 8449 7975 8483
rect 11437 8449 11471 8483
rect 14657 8449 14691 8483
rect 2044 8381 2078 8415
rect 3433 8381 3467 8415
rect 5089 8381 5123 8415
rect 6862 8381 6896 8415
rect 7573 8381 7607 8415
rect 8208 8381 8242 8415
rect 9413 8381 9447 8415
rect 11253 8381 11287 8415
rect 11897 8381 11931 8415
rect 12449 8381 12483 8415
rect 12705 8381 12739 8415
rect 3700 8313 3734 8347
rect 5345 8313 5379 8347
rect 9658 8313 9692 8347
rect 11345 8313 11379 8347
rect 14565 8313 14599 8347
rect 3157 8245 3191 8279
rect 10793 8245 10827 8279
rect 14473 8245 14507 8279
rect 15117 8245 15151 8279
rect 3709 8041 3743 8075
rect 6009 8041 6043 8075
rect 14381 8041 14415 8075
rect 4353 7973 4387 8007
rect 11612 7973 11646 8007
rect 13461 7973 13495 8007
rect 1593 7905 1627 7939
rect 2329 7905 2363 7939
rect 2596 7905 2630 7939
rect 4077 7905 4111 7939
rect 4896 7905 4930 7939
rect 6101 7905 6135 7939
rect 6368 7905 6402 7939
rect 7573 7905 7607 7939
rect 7829 7905 7863 7939
rect 9045 7905 9079 7939
rect 9689 7905 9723 7939
rect 9956 7905 9990 7939
rect 11345 7905 11379 7939
rect 13369 7905 13403 7939
rect 14473 7905 14507 7939
rect 1777 7837 1811 7871
rect 4629 7837 4663 7871
rect 9229 7837 9263 7871
rect 13553 7837 13587 7871
rect 14565 7837 14599 7871
rect 14013 7769 14047 7803
rect 7481 7701 7515 7735
rect 8953 7701 8987 7735
rect 11069 7701 11103 7735
rect 12725 7701 12759 7735
rect 13001 7701 13035 7735
rect 3249 7497 3283 7531
rect 8217 7497 8251 7531
rect 9873 7497 9907 7531
rect 12173 7497 12207 7531
rect 4813 7429 4847 7463
rect 11989 7429 12023 7463
rect 2053 7361 2087 7395
rect 3065 7361 3099 7395
rect 3249 7361 3283 7395
rect 5089 7361 5123 7395
rect 8493 7361 8527 7395
rect 10149 7361 10183 7395
rect 1777 7293 1811 7327
rect 3433 7293 3467 7327
rect 3700 7293 3734 7327
rect 6837 7293 6871 7327
rect 10416 7293 10450 7327
rect 11805 7293 11839 7327
rect 13277 7497 13311 7531
rect 12449 7429 12483 7463
rect 13001 7361 13035 7395
rect 14381 7497 14415 7531
rect 13921 7361 13955 7395
rect 14013 7361 14047 7395
rect 13277 7293 13311 7327
rect 2881 7225 2915 7259
rect 5356 7225 5390 7259
rect 7082 7225 7116 7259
rect 8760 7225 8794 7259
rect 12173 7225 12207 7259
rect 12817 7225 12851 7259
rect 15025 7361 15059 7395
rect 14933 7225 14967 7259
rect 1409 7157 1443 7191
rect 1869 7157 1903 7191
rect 2421 7157 2455 7191
rect 2789 7157 2823 7191
rect 6469 7157 6503 7191
rect 11529 7157 11563 7191
rect 12909 7157 12943 7191
rect 13461 7157 13495 7191
rect 13829 7157 13863 7191
rect 14381 7157 14415 7191
rect 14473 7157 14507 7191
rect 14841 7157 14875 7191
rect 4997 6953 5031 6987
rect 5365 6953 5399 6987
rect 9045 6953 9079 6987
rect 9505 6953 9539 6987
rect 11345 6953 11379 6987
rect 11713 6953 11747 6987
rect 13737 6953 13771 6987
rect 13829 6953 13863 6987
rect 14933 6953 14967 6987
rect 2574 6885 2608 6919
rect 4905 6885 4939 6919
rect 11805 6885 11839 6919
rect 12725 6885 12759 6919
rect 1593 6817 1627 6851
rect 2329 6817 2363 6851
rect 5365 6817 5399 6851
rect 5549 6817 5583 6851
rect 5816 6817 5850 6851
rect 7205 6817 7239 6851
rect 7461 6817 7495 6851
rect 9137 6817 9171 6851
rect 9505 6817 9539 6851
rect 9689 6817 9723 6851
rect 9956 6817 9990 6851
rect 12817 6817 12851 6851
rect 14381 6817 14415 6851
rect 15117 6817 15151 6851
rect 1777 6749 1811 6783
rect 4077 6749 4111 6783
rect 5181 6749 5215 6783
rect 9229 6749 9263 6783
rect 11897 6749 11931 6783
rect 12909 6749 12943 6783
rect 13921 6749 13955 6783
rect 8677 6681 8711 6715
rect 12357 6681 12391 6715
rect 13369 6681 13403 6715
rect 3709 6613 3743 6647
rect 4537 6613 4571 6647
rect 6929 6613 6963 6647
rect 8585 6613 8619 6647
rect 11069 6613 11103 6647
rect 14565 6613 14599 6647
rect 2421 6409 2455 6443
rect 9965 6409 9999 6443
rect 10149 6409 10183 6443
rect 13461 6409 13495 6443
rect 14473 6409 14507 6443
rect 4813 6341 4847 6375
rect 4997 6341 5031 6375
rect 2053 6273 2087 6307
rect 2973 6273 3007 6307
rect 3433 6273 3467 6307
rect 2881 6205 2915 6239
rect 6929 6273 6963 6307
rect 8585 6273 8619 6307
rect 5089 6205 5123 6239
rect 5345 6205 5379 6239
rect 1777 6137 1811 6171
rect 2789 6137 2823 6171
rect 3678 6137 3712 6171
rect 4997 6137 5031 6171
rect 7196 6137 7230 6171
rect 8852 6137 8886 6171
rect 11621 6341 11655 6375
rect 12173 6341 12207 6375
rect 10241 6273 10275 6307
rect 13277 6341 13311 6375
rect 13001 6273 13035 6307
rect 13921 6273 13955 6307
rect 14013 6273 14047 6307
rect 15025 6273 15059 6307
rect 10497 6205 10531 6239
rect 11805 6205 11839 6239
rect 12173 6205 12207 6239
rect 12909 6205 12943 6239
rect 13277 6205 13311 6239
rect 1409 6069 1443 6103
rect 1869 6069 1903 6103
rect 6469 6069 6503 6103
rect 8309 6069 8343 6103
rect 10149 6069 10183 6103
rect 14841 6137 14875 6171
rect 11713 6069 11747 6103
rect 11897 6069 11931 6103
rect 12449 6069 12483 6103
rect 12817 6069 12851 6103
rect 13829 6069 13863 6103
rect 14933 6069 14967 6103
rect 2421 5865 2455 5899
rect 3801 5865 3835 5899
rect 8677 5865 8711 5899
rect 9137 5865 9171 5899
rect 11161 5865 11195 5899
rect 11621 5865 11655 5899
rect 11713 5865 11747 5899
rect 12541 5865 12575 5899
rect 13093 5865 13127 5899
rect 14105 5865 14139 5899
rect 14749 5865 14783 5899
rect 1409 5729 1443 5763
rect 2329 5729 2363 5763
rect 3341 5729 3375 5763
rect 3433 5729 3467 5763
rect 2605 5661 2639 5695
rect 3617 5661 3651 5695
rect 1961 5593 1995 5627
rect 4629 5797 4663 5831
rect 4077 5729 4111 5763
rect 5253 5729 5287 5763
rect 6920 5729 6954 5763
rect 4261 5661 4295 5695
rect 4997 5661 5031 5695
rect 6653 5661 6687 5695
rect 8769 5661 8803 5695
rect 8953 5661 8987 5695
rect 10057 5797 10091 5831
rect 11069 5797 11103 5831
rect 9505 5729 9539 5763
rect 10149 5729 10183 5763
rect 10333 5661 10367 5695
rect 11345 5661 11379 5695
rect 8309 5593 8343 5627
rect 9137 5593 9171 5627
rect 12081 5797 12115 5831
rect 12173 5661 12207 5695
rect 12265 5661 12299 5695
rect 1593 5525 1627 5559
rect 2973 5525 3007 5559
rect 3801 5525 3835 5559
rect 6377 5525 6411 5559
rect 8033 5525 8067 5559
rect 9321 5525 9355 5559
rect 9689 5525 9723 5559
rect 10701 5525 10735 5559
rect 11529 5525 11563 5559
rect 13185 5661 13219 5695
rect 13277 5661 13311 5695
rect 14197 5661 14231 5695
rect 14289 5661 14323 5695
rect 12541 5525 12575 5559
rect 12725 5525 12759 5559
rect 13737 5525 13771 5559
rect 3065 5321 3099 5355
rect 4077 5321 4111 5355
rect 10149 5321 10183 5355
rect 1685 5253 1719 5287
rect 6469 5253 6503 5287
rect 8309 5253 8343 5287
rect 9873 5253 9907 5287
rect 9965 5253 9999 5287
rect 2513 5185 2547 5219
rect 2973 5185 3007 5219
rect 3525 5185 3559 5219
rect 3709 5185 3743 5219
rect 4629 5185 4663 5219
rect 6837 5185 6871 5219
rect 1501 5117 1535 5151
rect 4445 5117 4479 5151
rect 5089 5117 5123 5151
rect 2237 5049 2271 5083
rect 5334 5049 5368 5083
rect 7082 5049 7116 5083
rect 8493 5185 8527 5219
rect 8738 5049 8772 5083
rect 1869 4981 1903 5015
rect 2329 4981 2363 5015
rect 3433 4981 3467 5015
rect 4537 4981 4571 5015
rect 8217 4981 8251 5015
rect 8309 4981 8343 5015
rect 10609 5185 10643 5219
rect 10793 5185 10827 5219
rect 11713 5185 11747 5219
rect 13093 5185 13127 5219
rect 14013 5185 14047 5219
rect 15025 5185 15059 5219
rect 10517 5117 10551 5151
rect 11529 5117 11563 5151
rect 11621 5117 11655 5151
rect 12817 5049 12851 5083
rect 14841 5049 14875 5083
rect 9965 4981 9999 5015
rect 11161 4981 11195 5015
rect 12449 4981 12483 5015
rect 12909 4981 12943 5015
rect 13461 4981 13495 5015
rect 13829 4981 13863 5015
rect 13921 4981 13955 5015
rect 14473 4981 14507 5015
rect 14933 4981 14967 5015
rect 3341 4777 3375 4811
rect 4721 4777 4755 4811
rect 5089 4777 5123 4811
rect 5733 4777 5767 4811
rect 6101 4777 6135 4811
rect 10057 4777 10091 4811
rect 10149 4777 10183 4811
rect 10701 4777 10735 4811
rect 11713 4777 11747 4811
rect 14197 4777 14231 4811
rect 2421 4709 2455 4743
rect 8769 4709 8803 4743
rect 11069 4709 11103 4743
rect 11161 4709 11195 4743
rect 1409 4641 1443 4675
rect 2329 4641 2363 4675
rect 4169 4641 4203 4675
rect 5181 4641 5215 4675
rect 6745 4641 6779 4675
rect 7012 4641 7046 4675
rect 12081 4641 12115 4675
rect 12909 4641 12943 4675
rect 13553 4641 13587 4675
rect 14105 4641 14139 4675
rect 2605 4573 2639 4607
rect 3433 4573 3467 4607
rect 3525 4573 3559 4607
rect 5365 4573 5399 4607
rect 6193 4573 6227 4607
rect 6285 4573 6319 4607
rect 8309 4573 8343 4607
rect 8861 4573 8895 4607
rect 9045 4573 9079 4607
rect 10241 4573 10275 4607
rect 11345 4573 11379 4607
rect 12173 4573 12207 4607
rect 12265 4573 12299 4607
rect 13001 4573 13035 4607
rect 13093 4573 13127 4607
rect 14289 4573 14323 4607
rect 1593 4505 1627 4539
rect 2973 4505 3007 4539
rect 9689 4505 9723 4539
rect 1961 4437 1995 4471
rect 4353 4437 4387 4471
rect 8125 4437 8159 4471
rect 8309 4437 8343 4471
rect 8401 4437 8435 4471
rect 12541 4437 12575 4471
rect 13737 4437 13771 4471
rect 5549 4233 5583 4267
rect 5733 4233 5767 4267
rect 8493 4233 8527 4267
rect 9321 4233 9355 4267
rect 9505 4233 9539 4267
rect 14473 4233 14507 4267
rect 4077 4165 4111 4199
rect 2329 4097 2363 4131
rect 5181 4097 5215 4131
rect 5365 4097 5399 4131
rect 5549 4097 5583 4131
rect 2053 4029 2087 4063
rect 2697 4029 2731 4063
rect 4629 4029 4663 4063
rect 2942 3961 2976 3995
rect 1685 3893 1719 3927
rect 2145 3893 2179 3927
rect 4445 3893 4479 3927
rect 4721 3893 4755 3927
rect 5089 3893 5123 3927
rect 5549 3893 5583 3927
rect 6377 4097 6411 4131
rect 6837 4097 6871 4131
rect 9137 4097 9171 4131
rect 6193 4029 6227 4063
rect 10517 4165 10551 4199
rect 10149 4097 10183 4131
rect 10425 4097 10459 4131
rect 11161 4097 11195 4131
rect 13001 4097 13035 4131
rect 14013 4097 14047 4131
rect 15025 4097 15059 4131
rect 9873 4029 9907 4063
rect 7104 3961 7138 3995
rect 8861 3961 8895 3995
rect 9321 3961 9355 3995
rect 9965 3961 9999 3995
rect 10885 4029 10919 4063
rect 11535 4029 11569 4063
rect 13921 4029 13955 4063
rect 12817 3961 12851 3995
rect 14841 3961 14875 3995
rect 5641 3893 5675 3927
rect 6101 3893 6135 3927
rect 8217 3893 8251 3927
rect 8953 3893 8987 3927
rect 10425 3893 10459 3927
rect 10977 3893 11011 3927
rect 11713 3893 11747 3927
rect 12449 3893 12483 3927
rect 12909 3893 12943 3927
rect 13461 3893 13495 3927
rect 13829 3893 13863 3927
rect 14933 3893 14967 3927
rect 1961 3689 1995 3723
rect 2973 3689 3007 3723
rect 3433 3689 3467 3723
rect 4813 3689 4847 3723
rect 6469 3689 6503 3723
rect 7113 3689 7147 3723
rect 7757 3689 7791 3723
rect 9689 3689 9723 3723
rect 11069 3689 11103 3723
rect 11161 3689 11195 3723
rect 11713 3689 11747 3723
rect 12173 3689 12207 3723
rect 13737 3689 13771 3723
rect 14105 3689 14139 3723
rect 4721 3621 4755 3655
rect 5733 3621 5767 3655
rect 7205 3621 7239 3655
rect 10057 3621 10091 3655
rect 14197 3621 14231 3655
rect 1409 3553 1443 3587
rect 2329 3553 2363 3587
rect 3341 3553 3375 3587
rect 6653 3553 6687 3587
rect 8125 3553 8159 3587
rect 8769 3553 8803 3587
rect 12081 3553 12115 3587
rect 13093 3553 13127 3587
rect 13185 3553 13219 3587
rect 2421 3485 2455 3519
rect 2605 3485 2639 3519
rect 3617 3485 3651 3519
rect 4997 3485 5031 3519
rect 5825 3485 5859 3519
rect 6009 3485 6043 3519
rect 7297 3485 7331 3519
rect 8217 3485 8251 3519
rect 8309 3485 8343 3519
rect 10149 3485 10183 3519
rect 10333 3485 10367 3519
rect 11253 3485 11287 3519
rect 11621 3485 11655 3519
rect 12265 3485 12299 3519
rect 12633 3485 12667 3519
rect 13369 3485 13403 3519
rect 14289 3485 14323 3519
rect 6745 3417 6779 3451
rect 8953 3417 8987 3451
rect 10701 3417 10735 3451
rect 12541 3417 12575 3451
rect 12725 3417 12759 3451
rect 1593 3349 1627 3383
rect 4353 3349 4387 3383
rect 5365 3349 5399 3383
rect 11621 3349 11655 3383
rect 1685 3145 1719 3179
rect 2697 3145 2731 3179
rect 3709 3145 3743 3179
rect 4721 3145 4755 3179
rect 5733 3145 5767 3179
rect 6837 3145 6871 3179
rect 10885 3145 10919 3179
rect 12449 3145 12483 3179
rect 13645 3145 13679 3179
rect 8769 3077 8803 3111
rect 9873 3077 9907 3111
rect 14197 3077 14231 3111
rect 2237 3009 2271 3043
rect 3341 3009 3375 3043
rect 4261 3009 4295 3043
rect 5181 3009 5215 3043
rect 5365 3009 5399 3043
rect 6193 3009 6227 3043
rect 6377 3009 6411 3043
rect 7481 3009 7515 3043
rect 8493 3009 8527 3043
rect 9321 3009 9355 3043
rect 9505 3009 9539 3043
rect 10333 3009 10367 3043
rect 10517 3009 10551 3043
rect 11437 3009 11471 3043
rect 12909 3009 12943 3043
rect 13093 3009 13127 3043
rect 2145 2941 2179 2975
rect 3157 2941 3191 2975
rect 7205 2941 7239 2975
rect 8309 2941 8343 2975
rect 8769 2941 8803 2975
rect 10241 2941 10275 2975
rect 12817 2941 12851 2975
rect 13461 2941 13495 2975
rect 14013 2941 14047 2975
rect 14565 2941 14599 2975
rect 4169 2873 4203 2907
rect 5089 2873 5123 2907
rect 6101 2873 6135 2907
rect 7297 2873 7331 2907
rect 11345 2873 11379 2907
rect 2053 2805 2087 2839
rect 3065 2805 3099 2839
rect 4077 2805 4111 2839
rect 7849 2805 7883 2839
rect 8217 2805 8251 2839
rect 8861 2805 8895 2839
rect 9229 2805 9263 2839
rect 11253 2805 11287 2839
rect 11897 2805 11931 2839
rect 14749 2805 14783 2839
rect 2973 2601 3007 2635
rect 3433 2601 3467 2635
rect 4813 2601 4847 2635
rect 5181 2601 5215 2635
rect 5273 2601 5307 2635
rect 5641 2601 5675 2635
rect 5825 2601 5859 2635
rect 6285 2601 6319 2635
rect 8493 2601 8527 2635
rect 11161 2601 11195 2635
rect 12817 2601 12851 2635
rect 13645 2601 13679 2635
rect 2881 2533 2915 2567
rect 3341 2533 3375 2567
rect 1501 2465 1535 2499
rect 2237 2465 2271 2499
rect 1685 2397 1719 2431
rect 2421 2397 2455 2431
rect 4077 2465 4111 2499
rect 7573 2533 7607 2567
rect 8585 2533 8619 2567
rect 9505 2533 9539 2567
rect 9597 2533 9631 2567
rect 11253 2533 11287 2567
rect 6193 2465 6227 2499
rect 7481 2465 7515 2499
rect 9137 2465 9171 2499
rect 10149 2465 10183 2499
rect 10241 2465 10275 2499
rect 11805 2465 11839 2499
rect 12633 2465 12667 2499
rect 13185 2465 13219 2499
rect 13645 2465 13679 2499
rect 13737 2465 13771 2499
rect 14289 2465 14323 2499
rect 14841 2465 14875 2499
rect 3525 2397 3559 2431
rect 4261 2397 4295 2431
rect 5457 2397 5491 2431
rect 5641 2397 5675 2431
rect 6469 2397 6503 2431
rect 7757 2397 7791 2431
rect 8769 2397 8803 2431
rect 10425 2397 10459 2431
rect 11345 2397 11379 2431
rect 9321 2329 9355 2363
rect 13369 2329 13403 2363
rect 2881 2261 2915 2295
rect 7113 2261 7147 2295
rect 8125 2261 8159 2295
rect 9781 2261 9815 2295
rect 10793 2261 10827 2295
rect 11989 2261 12023 2295
rect 13921 2261 13955 2295
rect 14473 2261 14507 2295
rect 15025 2261 15059 2295
rect 8125 1649 8159 1683
rect 8125 901 8159 935
<< metal1 >>
rect 7466 16124 7472 16176
rect 7524 16164 7530 16176
rect 9122 16164 9128 16176
rect 7524 16136 9128 16164
rect 7524 16124 7530 16136
rect 9122 16124 9128 16136
rect 9180 16124 9186 16176
rect 8110 16056 8116 16108
rect 8168 16096 8174 16108
rect 8662 16096 8668 16108
rect 8168 16068 8668 16096
rect 8168 16056 8174 16068
rect 8662 16056 8668 16068
rect 8720 16056 8726 16108
rect 7006 15988 7012 16040
rect 7064 16028 7070 16040
rect 9398 16028 9404 16040
rect 7064 16000 9404 16028
rect 7064 15988 7070 16000
rect 9398 15988 9404 16000
rect 9456 15988 9462 16040
rect 1026 15920 1032 15972
rect 1084 15960 1090 15972
rect 3326 15960 3332 15972
rect 1084 15932 3332 15960
rect 1084 15920 1090 15932
rect 3326 15920 3332 15932
rect 3384 15920 3390 15972
rect 4246 15920 4252 15972
rect 4304 15960 4310 15972
rect 11790 15960 11796 15972
rect 4304 15932 11796 15960
rect 4304 15920 4310 15932
rect 11790 15920 11796 15932
rect 11848 15920 11854 15972
rect 3142 15852 3148 15904
rect 3200 15892 3206 15904
rect 4062 15892 4068 15904
rect 3200 15864 4068 15892
rect 3200 15852 3206 15864
rect 4062 15852 4068 15864
rect 4120 15852 4126 15904
rect 6638 15852 6644 15904
rect 6696 15892 6702 15904
rect 9858 15892 9864 15904
rect 6696 15864 9864 15892
rect 6696 15852 6702 15864
rect 9858 15852 9864 15864
rect 9916 15852 9922 15904
rect 1104 15802 15824 15824
rect 1104 15750 5912 15802
rect 5964 15750 5976 15802
rect 6028 15750 6040 15802
rect 6092 15750 6104 15802
rect 6156 15750 10843 15802
rect 10895 15750 10907 15802
rect 10959 15750 10971 15802
rect 11023 15750 11035 15802
rect 11087 15750 15824 15802
rect 1104 15728 15824 15750
rect 3602 15648 3608 15700
rect 3660 15688 3666 15700
rect 4433 15691 4491 15697
rect 4433 15688 4445 15691
rect 3660 15660 4445 15688
rect 3660 15648 3666 15660
rect 4433 15657 4445 15660
rect 4479 15657 4491 15691
rect 4433 15651 4491 15657
rect 5258 15648 5264 15700
rect 5316 15688 5322 15700
rect 5316 15660 7972 15688
rect 5316 15648 5322 15660
rect 2038 15580 2044 15632
rect 2096 15620 2102 15632
rect 6273 15623 6331 15629
rect 6273 15620 6285 15623
rect 2096 15592 6285 15620
rect 2096 15580 2102 15592
rect 6273 15589 6285 15592
rect 6319 15589 6331 15623
rect 7944 15620 7972 15660
rect 8202 15648 8208 15700
rect 8260 15688 8266 15700
rect 9309 15691 9367 15697
rect 9309 15688 9321 15691
rect 8260 15660 9321 15688
rect 8260 15648 8266 15660
rect 9309 15657 9321 15660
rect 9355 15657 9367 15691
rect 9309 15651 9367 15657
rect 9398 15648 9404 15700
rect 9456 15688 9462 15700
rect 9953 15691 10011 15697
rect 9953 15688 9965 15691
rect 9456 15660 9965 15688
rect 9456 15648 9462 15660
rect 9953 15657 9965 15660
rect 9999 15657 10011 15691
rect 9953 15651 10011 15657
rect 10505 15691 10563 15697
rect 10505 15657 10517 15691
rect 10551 15657 10563 15691
rect 10505 15651 10563 15657
rect 10520 15620 10548 15651
rect 6273 15583 6331 15589
rect 6380 15592 7696 15620
rect 7944 15592 10548 15620
rect 3237 15555 3295 15561
rect 3237 15521 3249 15555
rect 3283 15552 3295 15555
rect 3786 15552 3792 15564
rect 3283 15524 3792 15552
rect 3283 15521 3295 15524
rect 3237 15515 3295 15521
rect 3786 15512 3792 15524
rect 3844 15512 3850 15564
rect 4246 15552 4252 15564
rect 4207 15524 4252 15552
rect 4246 15512 4252 15524
rect 4304 15512 4310 15564
rect 4801 15555 4859 15561
rect 4801 15521 4813 15555
rect 4847 15552 4859 15555
rect 5810 15552 5816 15564
rect 4847 15524 5816 15552
rect 4847 15521 4859 15524
rect 4801 15515 4859 15521
rect 5810 15512 5816 15524
rect 5868 15512 5874 15564
rect 6178 15552 6184 15564
rect 6139 15524 6184 15552
rect 6178 15512 6184 15524
rect 6236 15512 6242 15564
rect 2774 15444 2780 15496
rect 2832 15484 2838 15496
rect 2832 15456 5488 15484
rect 2832 15444 2838 15456
rect 5460 15428 5488 15456
rect 5626 15444 5632 15496
rect 5684 15484 5690 15496
rect 6380 15484 6408 15592
rect 7466 15552 7472 15564
rect 7427 15524 7472 15552
rect 7466 15512 7472 15524
rect 7524 15512 7530 15564
rect 5684 15456 6408 15484
rect 6457 15487 6515 15493
rect 5684 15444 5690 15456
rect 6457 15453 6469 15487
rect 6503 15484 6515 15487
rect 6638 15484 6644 15496
rect 6503 15456 6644 15484
rect 6503 15453 6515 15456
rect 6457 15447 6515 15453
rect 6638 15444 6644 15456
rect 6696 15444 6702 15496
rect 7668 15493 7696 15592
rect 8481 15555 8539 15561
rect 8481 15521 8493 15555
rect 8527 15521 8539 15555
rect 8481 15515 8539 15521
rect 8573 15555 8631 15561
rect 8573 15521 8585 15555
rect 8619 15552 8631 15555
rect 8619 15524 8800 15552
rect 8619 15521 8631 15524
rect 8573 15515 8631 15521
rect 7561 15487 7619 15493
rect 7561 15453 7573 15487
rect 7607 15453 7619 15487
rect 7561 15447 7619 15453
rect 7653 15487 7711 15493
rect 7653 15453 7665 15487
rect 7699 15453 7711 15487
rect 7653 15447 7711 15453
rect 2682 15376 2688 15428
rect 2740 15416 2746 15428
rect 4985 15419 5043 15425
rect 4985 15416 4997 15419
rect 2740 15388 4997 15416
rect 2740 15376 2746 15388
rect 4985 15385 4997 15388
rect 5031 15385 5043 15419
rect 4985 15379 5043 15385
rect 5442 15376 5448 15428
rect 5500 15416 5506 15428
rect 7576 15416 7604 15447
rect 5500 15388 7604 15416
rect 8496 15416 8524 15515
rect 8772 15496 8800 15524
rect 9030 15512 9036 15564
rect 9088 15552 9094 15564
rect 9125 15555 9183 15561
rect 9125 15552 9137 15555
rect 9088 15524 9137 15552
rect 9088 15512 9094 15524
rect 9125 15521 9137 15524
rect 9171 15521 9183 15555
rect 9125 15515 9183 15521
rect 9769 15555 9827 15561
rect 9769 15521 9781 15555
rect 9815 15552 9827 15555
rect 10042 15552 10048 15564
rect 9815 15524 10048 15552
rect 9815 15521 9827 15524
rect 9769 15515 9827 15521
rect 10042 15512 10048 15524
rect 10100 15512 10106 15564
rect 10321 15555 10379 15561
rect 10321 15521 10333 15555
rect 10367 15552 10379 15555
rect 11146 15552 11152 15564
rect 10367 15524 11152 15552
rect 10367 15521 10379 15524
rect 10321 15515 10379 15521
rect 11146 15512 11152 15524
rect 11204 15512 11210 15564
rect 8662 15484 8668 15496
rect 8623 15456 8668 15484
rect 8662 15444 8668 15456
rect 8720 15444 8726 15496
rect 8754 15444 8760 15496
rect 8812 15484 8818 15496
rect 9950 15484 9956 15496
rect 8812 15456 9956 15484
rect 8812 15444 8818 15456
rect 9950 15444 9956 15456
rect 10008 15444 10014 15496
rect 9306 15416 9312 15428
rect 8496 15388 9312 15416
rect 5500 15376 5506 15388
rect 9306 15376 9312 15388
rect 9364 15376 9370 15428
rect 10410 15376 10416 15428
rect 10468 15416 10474 15428
rect 13906 15416 13912 15428
rect 10468 15388 13912 15416
rect 10468 15376 10474 15388
rect 13906 15376 13912 15388
rect 13964 15376 13970 15428
rect 3050 15308 3056 15360
rect 3108 15348 3114 15360
rect 3421 15351 3479 15357
rect 3421 15348 3433 15351
rect 3108 15320 3433 15348
rect 3108 15308 3114 15320
rect 3421 15317 3433 15320
rect 3467 15317 3479 15351
rect 3421 15311 3479 15317
rect 5813 15351 5871 15357
rect 5813 15317 5825 15351
rect 5859 15348 5871 15351
rect 6638 15348 6644 15360
rect 5859 15320 6644 15348
rect 5859 15317 5871 15320
rect 5813 15311 5871 15317
rect 6638 15308 6644 15320
rect 6696 15308 6702 15360
rect 7098 15348 7104 15360
rect 7059 15320 7104 15348
rect 7098 15308 7104 15320
rect 7156 15308 7162 15360
rect 7190 15308 7196 15360
rect 7248 15348 7254 15360
rect 8113 15351 8171 15357
rect 8113 15348 8125 15351
rect 7248 15320 8125 15348
rect 7248 15308 7254 15320
rect 8113 15317 8125 15320
rect 8159 15317 8171 15351
rect 8113 15311 8171 15317
rect 10318 15308 10324 15360
rect 10376 15348 10382 15360
rect 13814 15348 13820 15360
rect 10376 15320 13820 15348
rect 10376 15308 10382 15320
rect 13814 15308 13820 15320
rect 13872 15308 13878 15360
rect 1104 15258 15824 15280
rect 1104 15206 3447 15258
rect 3499 15206 3511 15258
rect 3563 15206 3575 15258
rect 3627 15206 3639 15258
rect 3691 15206 8378 15258
rect 8430 15206 8442 15258
rect 8494 15206 8506 15258
rect 8558 15206 8570 15258
rect 8622 15206 13308 15258
rect 13360 15206 13372 15258
rect 13424 15206 13436 15258
rect 13488 15206 13500 15258
rect 13552 15206 15824 15258
rect 1104 15184 15824 15206
rect 1394 15104 1400 15156
rect 1452 15144 1458 15156
rect 3050 15144 3056 15156
rect 1452 15116 3056 15144
rect 1452 15104 1458 15116
rect 3050 15104 3056 15116
rect 3108 15104 3114 15156
rect 3142 15104 3148 15156
rect 3200 15144 3206 15156
rect 5353 15147 5411 15153
rect 5353 15144 5365 15147
rect 3200 15116 5365 15144
rect 3200 15104 3206 15116
rect 5353 15113 5365 15116
rect 5399 15113 5411 15147
rect 5353 15107 5411 15113
rect 6546 15104 6552 15156
rect 6604 15144 6610 15156
rect 9677 15147 9735 15153
rect 6604 15116 8800 15144
rect 6604 15104 6610 15116
rect 566 15036 572 15088
rect 624 15076 630 15088
rect 2961 15079 3019 15085
rect 2961 15076 2973 15079
rect 624 15048 2973 15076
rect 624 15036 630 15048
rect 2961 15045 2973 15048
rect 3007 15045 3019 15079
rect 2961 15039 3019 15045
rect 3326 15036 3332 15088
rect 3384 15076 3390 15088
rect 3513 15079 3571 15085
rect 3513 15076 3525 15079
rect 3384 15048 3525 15076
rect 3384 15036 3390 15048
rect 3513 15045 3525 15048
rect 3559 15045 3571 15079
rect 3513 15039 3571 15045
rect 4801 15079 4859 15085
rect 4801 15045 4813 15079
rect 4847 15045 4859 15079
rect 4801 15039 4859 15045
rect 1854 14968 1860 15020
rect 1912 15008 1918 15020
rect 4816 15008 4844 15039
rect 5534 15036 5540 15088
rect 5592 15076 5598 15088
rect 5592 15048 6224 15076
rect 5592 15036 5598 15048
rect 6086 15008 6092 15020
rect 1912 14980 4844 15008
rect 4908 14980 6092 15008
rect 1912 14968 1918 14980
rect 2222 14940 2228 14952
rect 2183 14912 2228 14940
rect 2222 14900 2228 14912
rect 2280 14900 2286 14952
rect 2774 14940 2780 14952
rect 2735 14912 2780 14940
rect 2774 14900 2780 14912
rect 2832 14900 2838 14952
rect 3234 14900 3240 14952
rect 3292 14940 3298 14952
rect 3329 14943 3387 14949
rect 3329 14940 3341 14943
rect 3292 14912 3341 14940
rect 3292 14900 3298 14912
rect 3329 14909 3341 14912
rect 3375 14909 3387 14943
rect 3329 14903 3387 14909
rect 3694 14900 3700 14952
rect 3752 14940 3758 14952
rect 3881 14943 3939 14949
rect 3881 14940 3893 14943
rect 3752 14912 3893 14940
rect 3752 14900 3758 14912
rect 3881 14909 3893 14912
rect 3927 14909 3939 14943
rect 3881 14903 3939 14909
rect 3970 14900 3976 14952
rect 4028 14940 4034 14952
rect 4157 14943 4215 14949
rect 4157 14940 4169 14943
rect 4028 14912 4169 14940
rect 4028 14900 4034 14912
rect 4157 14909 4169 14912
rect 4203 14909 4215 14943
rect 4157 14903 4215 14909
rect 4617 14943 4675 14949
rect 4617 14909 4629 14943
rect 4663 14940 4675 14943
rect 4908 14940 4936 14980
rect 6086 14968 6092 14980
rect 6144 14968 6150 15020
rect 6196 15017 6224 15048
rect 6270 15036 6276 15088
rect 6328 15076 6334 15088
rect 6328 15048 6868 15076
rect 6328 15036 6334 15048
rect 6181 15011 6239 15017
rect 6181 14977 6193 15011
rect 6227 14977 6239 15011
rect 6362 15008 6368 15020
rect 6323 14980 6368 15008
rect 6181 14971 6239 14977
rect 6362 14968 6368 14980
rect 6420 14968 6426 15020
rect 6840 15008 6868 15048
rect 6914 15036 6920 15088
rect 6972 15076 6978 15088
rect 7377 15079 7435 15085
rect 7377 15076 7389 15079
rect 6972 15048 7389 15076
rect 6972 15036 6978 15048
rect 7377 15045 7389 15048
rect 7423 15045 7435 15079
rect 8772 15076 8800 15116
rect 9677 15113 9689 15147
rect 9723 15144 9735 15147
rect 12158 15144 12164 15156
rect 9723 15116 12164 15144
rect 9723 15113 9735 15116
rect 9677 15107 9735 15113
rect 12158 15104 12164 15116
rect 12216 15104 12222 15156
rect 14182 15076 14188 15088
rect 8772 15048 9352 15076
rect 7377 15039 7435 15045
rect 6840 14980 7236 15008
rect 4663 14912 4936 14940
rect 4663 14909 4675 14912
rect 4617 14903 4675 14909
rect 4982 14900 4988 14952
rect 5040 14940 5046 14952
rect 5169 14943 5227 14949
rect 5169 14940 5181 14943
rect 5040 14912 5181 14940
rect 5040 14900 5046 14912
rect 5169 14909 5181 14912
rect 5215 14909 5227 14943
rect 5169 14903 5227 14909
rect 5718 14900 5724 14952
rect 5776 14940 5782 14952
rect 6270 14940 6276 14952
rect 5776 14912 6276 14940
rect 5776 14900 5782 14912
rect 6270 14900 6276 14912
rect 6328 14900 6334 14952
rect 6454 14900 6460 14952
rect 6512 14940 6518 14952
rect 6825 14943 6883 14949
rect 6825 14940 6837 14943
rect 6512 14912 6837 14940
rect 6512 14900 6518 14912
rect 6825 14909 6837 14912
rect 6871 14909 6883 14943
rect 6825 14903 6883 14909
rect 4062 14832 4068 14884
rect 4120 14872 4126 14884
rect 7208 14872 7236 14980
rect 7282 14968 7288 15020
rect 7340 15008 7346 15020
rect 8205 15011 8263 15017
rect 8205 15008 8217 15011
rect 7340 14980 8217 15008
rect 7340 14968 7346 14980
rect 8205 14977 8217 14980
rect 8251 14977 8263 15011
rect 8205 14971 8263 14977
rect 8662 14968 8668 15020
rect 8720 15008 8726 15020
rect 9217 15011 9275 15017
rect 9217 15008 9229 15011
rect 8720 14980 9229 15008
rect 8720 14968 8726 14980
rect 9217 14977 9229 14980
rect 9263 14977 9275 15011
rect 9217 14971 9275 14977
rect 7374 14900 7380 14952
rect 7432 14940 7438 14952
rect 7561 14943 7619 14949
rect 7561 14940 7573 14943
rect 7432 14912 7573 14940
rect 7432 14900 7438 14912
rect 7561 14909 7573 14912
rect 7607 14909 7619 14943
rect 7561 14903 7619 14909
rect 7650 14900 7656 14952
rect 7708 14940 7714 14952
rect 7926 14940 7932 14952
rect 7708 14912 7932 14940
rect 7708 14900 7714 14912
rect 7926 14900 7932 14912
rect 7984 14900 7990 14952
rect 8018 14900 8024 14952
rect 8076 14940 8082 14952
rect 8113 14943 8171 14949
rect 8113 14940 8125 14943
rect 8076 14912 8125 14940
rect 8076 14900 8082 14912
rect 8113 14909 8125 14912
rect 8159 14909 8171 14943
rect 9324 14940 9352 15048
rect 10152 15048 14188 15076
rect 10152 15017 10180 15048
rect 14182 15036 14188 15048
rect 14240 15076 14246 15088
rect 14734 15076 14740 15088
rect 14240 15048 14740 15076
rect 14240 15036 14246 15048
rect 14734 15036 14740 15048
rect 14792 15036 14798 15088
rect 10137 15011 10195 15017
rect 10137 14977 10149 15011
rect 10183 14977 10195 15011
rect 10137 14971 10195 14977
rect 10321 15011 10379 15017
rect 10321 14977 10333 15011
rect 10367 15008 10379 15011
rect 10502 15008 10508 15020
rect 10367 14980 10508 15008
rect 10367 14977 10379 14980
rect 10321 14971 10379 14977
rect 10502 14968 10508 14980
rect 10560 14968 10566 15020
rect 9324 14912 10364 14940
rect 8113 14903 8171 14909
rect 8938 14872 8944 14884
rect 4120 14844 7052 14872
rect 7208 14844 8944 14872
rect 4120 14832 4126 14844
rect 2409 14807 2467 14813
rect 2409 14773 2421 14807
rect 2455 14804 2467 14807
rect 4798 14804 4804 14816
rect 2455 14776 4804 14804
rect 2455 14773 2467 14776
rect 2409 14767 2467 14773
rect 4798 14764 4804 14776
rect 4856 14764 4862 14816
rect 5166 14764 5172 14816
rect 5224 14804 5230 14816
rect 5721 14807 5779 14813
rect 5721 14804 5733 14807
rect 5224 14776 5733 14804
rect 5224 14764 5230 14776
rect 5721 14773 5733 14776
rect 5767 14773 5779 14807
rect 5721 14767 5779 14773
rect 5810 14764 5816 14816
rect 5868 14804 5874 14816
rect 6089 14807 6147 14813
rect 6089 14804 6101 14807
rect 5868 14776 6101 14804
rect 5868 14764 5874 14776
rect 6089 14773 6101 14776
rect 6135 14804 6147 14807
rect 6730 14804 6736 14816
rect 6135 14776 6736 14804
rect 6135 14773 6147 14776
rect 6089 14767 6147 14773
rect 6730 14764 6736 14776
rect 6788 14764 6794 14816
rect 7024 14813 7052 14844
rect 8938 14832 8944 14844
rect 8996 14832 9002 14884
rect 9125 14875 9183 14881
rect 9125 14841 9137 14875
rect 9171 14872 9183 14875
rect 10226 14872 10232 14884
rect 9171 14844 10232 14872
rect 9171 14841 9183 14844
rect 9125 14835 9183 14841
rect 10226 14832 10232 14844
rect 10284 14832 10290 14884
rect 10336 14872 10364 14912
rect 10594 14900 10600 14952
rect 10652 14940 10658 14952
rect 10689 14943 10747 14949
rect 10689 14940 10701 14943
rect 10652 14912 10701 14940
rect 10652 14900 10658 14912
rect 10689 14909 10701 14912
rect 10735 14909 10747 14943
rect 10689 14903 10747 14909
rect 10778 14900 10784 14952
rect 10836 14940 10842 14952
rect 12986 14940 12992 14952
rect 10836 14912 12992 14940
rect 10836 14900 10842 14912
rect 12986 14900 12992 14912
rect 13044 14900 13050 14952
rect 10336 14844 10916 14872
rect 7009 14807 7067 14813
rect 7009 14773 7021 14807
rect 7055 14773 7067 14807
rect 7650 14804 7656 14816
rect 7611 14776 7656 14804
rect 7009 14767 7067 14773
rect 7650 14764 7656 14776
rect 7708 14764 7714 14816
rect 8021 14807 8079 14813
rect 8021 14773 8033 14807
rect 8067 14804 8079 14807
rect 8202 14804 8208 14816
rect 8067 14776 8208 14804
rect 8067 14773 8079 14776
rect 8021 14767 8079 14773
rect 8202 14764 8208 14776
rect 8260 14764 8266 14816
rect 8662 14804 8668 14816
rect 8623 14776 8668 14804
rect 8662 14764 8668 14776
rect 8720 14764 8726 14816
rect 9030 14804 9036 14816
rect 8943 14776 9036 14804
rect 9030 14764 9036 14776
rect 9088 14804 9094 14816
rect 10888 14813 10916 14844
rect 10045 14807 10103 14813
rect 10045 14804 10057 14807
rect 9088 14776 10057 14804
rect 9088 14764 9094 14776
rect 10045 14773 10057 14776
rect 10091 14773 10103 14807
rect 10045 14767 10103 14773
rect 10873 14807 10931 14813
rect 10873 14773 10885 14807
rect 10919 14773 10931 14807
rect 11238 14804 11244 14816
rect 11199 14776 11244 14804
rect 10873 14767 10931 14773
rect 11238 14764 11244 14776
rect 11296 14764 11302 14816
rect 11330 14764 11336 14816
rect 11388 14804 11394 14816
rect 11882 14804 11888 14816
rect 11388 14776 11888 14804
rect 11388 14764 11394 14776
rect 11882 14764 11888 14776
rect 11940 14764 11946 14816
rect 1104 14714 15824 14736
rect 1104 14662 5912 14714
rect 5964 14662 5976 14714
rect 6028 14662 6040 14714
rect 6092 14662 6104 14714
rect 6156 14662 10843 14714
rect 10895 14662 10907 14714
rect 10959 14662 10971 14714
rect 11023 14662 11035 14714
rect 11087 14662 15824 14714
rect 1104 14640 15824 14662
rect 198 14560 204 14612
rect 256 14600 262 14612
rect 2593 14603 2651 14609
rect 2593 14600 2605 14603
rect 256 14572 2605 14600
rect 256 14560 262 14572
rect 2593 14569 2605 14572
rect 2639 14569 2651 14603
rect 2593 14563 2651 14569
rect 3786 14560 3792 14612
rect 3844 14600 3850 14612
rect 5718 14600 5724 14612
rect 3844 14572 5724 14600
rect 3844 14560 3850 14572
rect 5718 14560 5724 14572
rect 5776 14560 5782 14612
rect 5813 14603 5871 14609
rect 5813 14569 5825 14603
rect 5859 14600 5871 14603
rect 7098 14600 7104 14612
rect 5859 14572 7104 14600
rect 5859 14569 5871 14572
rect 5813 14563 5871 14569
rect 7098 14560 7104 14572
rect 7156 14560 7162 14612
rect 7558 14560 7564 14612
rect 7616 14600 7622 14612
rect 8478 14600 8484 14612
rect 7616 14572 8484 14600
rect 7616 14560 7622 14572
rect 8478 14560 8484 14572
rect 8536 14560 8542 14612
rect 8846 14600 8852 14612
rect 8807 14572 8852 14600
rect 8846 14560 8852 14572
rect 8904 14560 8910 14612
rect 8938 14560 8944 14612
rect 8996 14600 9002 14612
rect 9582 14600 9588 14612
rect 8996 14572 9588 14600
rect 8996 14560 9002 14572
rect 9582 14560 9588 14572
rect 9640 14560 9646 14612
rect 9677 14603 9735 14609
rect 9677 14569 9689 14603
rect 9723 14600 9735 14603
rect 12802 14600 12808 14612
rect 9723 14572 12808 14600
rect 9723 14569 9735 14572
rect 9677 14563 9735 14569
rect 12802 14560 12808 14572
rect 12860 14560 12866 14612
rect 4430 14532 4436 14544
rect 2332 14504 4436 14532
rect 1854 14464 1860 14476
rect 1815 14436 1860 14464
rect 1854 14424 1860 14436
rect 1912 14424 1918 14476
rect 2041 14331 2099 14337
rect 2041 14297 2053 14331
rect 2087 14328 2099 14331
rect 2332 14328 2360 14504
rect 4430 14492 4436 14504
rect 4488 14492 4494 14544
rect 6181 14535 6239 14541
rect 6181 14532 6193 14535
rect 4540 14504 6193 14532
rect 2409 14467 2467 14473
rect 2409 14433 2421 14467
rect 2455 14433 2467 14467
rect 2958 14464 2964 14476
rect 2919 14436 2964 14464
rect 2409 14427 2467 14433
rect 2087 14300 2360 14328
rect 2424 14328 2452 14427
rect 2958 14424 2964 14436
rect 3016 14424 3022 14476
rect 3326 14424 3332 14476
rect 3384 14464 3390 14476
rect 4540 14464 4568 14504
rect 6181 14501 6193 14504
rect 6227 14501 6239 14535
rect 6181 14495 6239 14501
rect 6546 14492 6552 14544
rect 6604 14532 6610 14544
rect 6733 14535 6791 14541
rect 6733 14532 6745 14535
rect 6604 14504 6745 14532
rect 6604 14492 6610 14504
rect 6733 14501 6745 14504
rect 6779 14501 6791 14535
rect 6733 14495 6791 14501
rect 6825 14535 6883 14541
rect 6825 14501 6837 14535
rect 6871 14532 6883 14535
rect 8570 14532 8576 14544
rect 6871 14504 8576 14532
rect 6871 14501 6883 14504
rect 6825 14495 6883 14501
rect 8570 14492 8576 14504
rect 8628 14492 8634 14544
rect 8757 14535 8815 14541
rect 8757 14501 8769 14535
rect 8803 14532 8815 14535
rect 10045 14535 10103 14541
rect 10045 14532 10057 14535
rect 8803 14504 10057 14532
rect 8803 14501 8815 14504
rect 8757 14495 8815 14501
rect 10045 14501 10057 14504
rect 10091 14532 10103 14535
rect 10594 14532 10600 14544
rect 10091 14504 10600 14532
rect 10091 14501 10103 14504
rect 10045 14495 10103 14501
rect 10594 14492 10600 14504
rect 10652 14492 10658 14544
rect 11057 14535 11115 14541
rect 11057 14501 11069 14535
rect 11103 14532 11115 14535
rect 14550 14532 14556 14544
rect 11103 14504 14556 14532
rect 11103 14501 11115 14504
rect 11057 14495 11115 14501
rect 14550 14492 14556 14504
rect 14608 14492 14614 14544
rect 4706 14464 4712 14476
rect 3384 14436 4568 14464
rect 4667 14436 4712 14464
rect 3384 14424 3390 14436
rect 4706 14424 4712 14436
rect 4764 14424 4770 14476
rect 7006 14464 7012 14476
rect 6012 14436 7012 14464
rect 3142 14396 3148 14408
rect 3103 14368 3148 14396
rect 3142 14356 3148 14368
rect 3200 14356 3206 14408
rect 4614 14356 4620 14408
rect 4672 14396 4678 14408
rect 4801 14399 4859 14405
rect 4801 14396 4813 14399
rect 4672 14368 4813 14396
rect 4672 14356 4678 14368
rect 4801 14365 4813 14368
rect 4847 14365 4859 14399
rect 4801 14359 4859 14365
rect 4985 14399 5043 14405
rect 4985 14365 4997 14399
rect 5031 14396 5043 14399
rect 5534 14396 5540 14408
rect 5031 14368 5540 14396
rect 5031 14365 5043 14368
rect 4985 14359 5043 14365
rect 5534 14356 5540 14368
rect 5592 14356 5598 14408
rect 6012 14405 6040 14436
rect 7006 14424 7012 14436
rect 7064 14424 7070 14476
rect 7742 14464 7748 14476
rect 7703 14436 7748 14464
rect 7742 14424 7748 14436
rect 7800 14424 7806 14476
rect 7837 14467 7895 14473
rect 7837 14433 7849 14467
rect 7883 14464 7895 14467
rect 9490 14464 9496 14476
rect 7883 14436 9496 14464
rect 7883 14433 7895 14436
rect 7837 14427 7895 14433
rect 9490 14424 9496 14436
rect 9548 14424 9554 14476
rect 9766 14464 9772 14476
rect 9600 14436 9772 14464
rect 5997 14399 6055 14405
rect 5997 14365 6009 14399
rect 6043 14365 6055 14399
rect 5997 14359 6055 14365
rect 6917 14399 6975 14405
rect 6917 14365 6929 14399
rect 6963 14365 6975 14399
rect 6917 14359 6975 14365
rect 7193 14399 7251 14405
rect 7193 14365 7205 14399
rect 7239 14396 7251 14399
rect 8021 14399 8079 14405
rect 8021 14396 8033 14399
rect 7239 14368 8033 14396
rect 7239 14365 7251 14368
rect 7193 14359 7251 14365
rect 8021 14365 8033 14368
rect 8067 14396 8079 14399
rect 9033 14399 9091 14405
rect 8067 14368 8524 14396
rect 8067 14365 8079 14368
rect 8021 14359 8079 14365
rect 4632 14328 4660 14356
rect 2424 14300 4660 14328
rect 2087 14297 2099 14300
rect 2041 14291 2099 14297
rect 5074 14288 5080 14340
rect 5132 14328 5138 14340
rect 6822 14328 6828 14340
rect 5132 14300 6828 14328
rect 5132 14288 5138 14300
rect 6822 14288 6828 14300
rect 6880 14288 6886 14340
rect 2774 14220 2780 14272
rect 2832 14260 2838 14272
rect 3878 14260 3884 14272
rect 2832 14232 3884 14260
rect 2832 14220 2838 14232
rect 3878 14220 3884 14232
rect 3936 14220 3942 14272
rect 4338 14260 4344 14272
rect 4299 14232 4344 14260
rect 4338 14220 4344 14232
rect 4396 14220 4402 14272
rect 5350 14260 5356 14272
rect 5311 14232 5356 14260
rect 5350 14220 5356 14232
rect 5408 14220 5414 14272
rect 5534 14220 5540 14272
rect 5592 14260 5598 14272
rect 5810 14260 5816 14272
rect 5592 14232 5816 14260
rect 5592 14220 5598 14232
rect 5810 14220 5816 14232
rect 5868 14220 5874 14272
rect 6181 14263 6239 14269
rect 6181 14229 6193 14263
rect 6227 14260 6239 14263
rect 6365 14263 6423 14269
rect 6365 14260 6377 14263
rect 6227 14232 6377 14260
rect 6227 14229 6239 14232
rect 6181 14223 6239 14229
rect 6365 14229 6377 14232
rect 6411 14229 6423 14263
rect 6932 14260 6960 14359
rect 7098 14288 7104 14340
rect 7156 14328 7162 14340
rect 7377 14331 7435 14337
rect 7377 14328 7389 14331
rect 7156 14300 7389 14328
rect 7156 14288 7162 14300
rect 7377 14297 7389 14300
rect 7423 14297 7435 14331
rect 7377 14291 7435 14297
rect 7193 14263 7251 14269
rect 7193 14260 7205 14263
rect 6932 14232 7205 14260
rect 6365 14223 6423 14229
rect 7193 14229 7205 14232
rect 7239 14229 7251 14263
rect 7193 14223 7251 14229
rect 7466 14220 7472 14272
rect 7524 14260 7530 14272
rect 8389 14263 8447 14269
rect 8389 14260 8401 14263
rect 7524 14232 8401 14260
rect 7524 14220 7530 14232
rect 8389 14229 8401 14232
rect 8435 14229 8447 14263
rect 8496 14260 8524 14368
rect 9033 14365 9045 14399
rect 9079 14396 9091 14399
rect 9079 14368 9260 14396
rect 9079 14365 9091 14368
rect 9033 14359 9091 14365
rect 8570 14288 8576 14340
rect 8628 14328 8634 14340
rect 8754 14328 8760 14340
rect 8628 14300 8760 14328
rect 8628 14288 8634 14300
rect 8754 14288 8760 14300
rect 8812 14288 8818 14340
rect 9232 14328 9260 14368
rect 9398 14356 9404 14408
rect 9456 14396 9462 14408
rect 9600 14396 9628 14436
rect 9766 14424 9772 14436
rect 9824 14424 9830 14476
rect 9858 14424 9864 14476
rect 9916 14464 9922 14476
rect 10226 14464 10232 14476
rect 9916 14436 10232 14464
rect 9916 14424 9922 14436
rect 10226 14424 10232 14436
rect 10284 14464 10290 14476
rect 10284 14436 10640 14464
rect 10284 14424 10290 14436
rect 9456 14368 9628 14396
rect 9456 14356 9462 14368
rect 9674 14356 9680 14408
rect 9732 14396 9738 14408
rect 10137 14399 10195 14405
rect 10137 14396 10149 14399
rect 9732 14368 10149 14396
rect 9732 14356 9738 14368
rect 10137 14365 10149 14368
rect 10183 14365 10195 14399
rect 10137 14359 10195 14365
rect 10321 14399 10379 14405
rect 10321 14365 10333 14399
rect 10367 14396 10379 14399
rect 10502 14396 10508 14408
rect 10367 14368 10508 14396
rect 10367 14365 10379 14368
rect 10321 14359 10379 14365
rect 10502 14356 10508 14368
rect 10560 14356 10566 14408
rect 10612 14396 10640 14436
rect 10686 14424 10692 14476
rect 10744 14464 10750 14476
rect 11149 14467 11207 14473
rect 11149 14464 11161 14467
rect 10744 14436 11161 14464
rect 10744 14424 10750 14436
rect 11149 14433 11161 14436
rect 11195 14464 11207 14467
rect 11195 14436 11652 14464
rect 11195 14433 11207 14436
rect 11149 14427 11207 14433
rect 11241 14399 11299 14405
rect 11241 14396 11253 14399
rect 10612 14368 11253 14396
rect 11241 14365 11253 14368
rect 11287 14365 11299 14399
rect 11624 14396 11652 14436
rect 11698 14424 11704 14476
rect 11756 14464 11762 14476
rect 12437 14467 12495 14473
rect 11756 14436 11801 14464
rect 11756 14424 11762 14436
rect 12437 14433 12449 14467
rect 12483 14464 12495 14467
rect 13814 14464 13820 14476
rect 12483 14436 13820 14464
rect 12483 14433 12495 14436
rect 12437 14427 12495 14433
rect 13814 14424 13820 14436
rect 13872 14424 13878 14476
rect 14458 14396 14464 14408
rect 11624 14368 14464 14396
rect 11241 14359 11299 14365
rect 14458 14356 14464 14368
rect 14516 14396 14522 14408
rect 15470 14396 15476 14408
rect 14516 14368 15476 14396
rect 14516 14356 14522 14368
rect 15470 14356 15476 14368
rect 15528 14356 15534 14408
rect 9766 14328 9772 14340
rect 9232 14300 9772 14328
rect 9766 14288 9772 14300
rect 9824 14328 9830 14340
rect 10410 14328 10416 14340
rect 9824 14300 10416 14328
rect 9824 14288 9830 14300
rect 10410 14288 10416 14300
rect 10468 14288 10474 14340
rect 10689 14331 10747 14337
rect 10689 14297 10701 14331
rect 10735 14328 10747 14331
rect 10735 14300 13400 14328
rect 10735 14297 10747 14300
rect 10689 14291 10747 14297
rect 9398 14260 9404 14272
rect 8496 14232 9404 14260
rect 8389 14223 8447 14229
rect 9398 14220 9404 14232
rect 9456 14220 9462 14272
rect 9582 14220 9588 14272
rect 9640 14260 9646 14272
rect 11885 14263 11943 14269
rect 11885 14260 11897 14263
rect 9640 14232 11897 14260
rect 9640 14220 9646 14232
rect 11885 14229 11897 14232
rect 11931 14229 11943 14263
rect 12250 14260 12256 14272
rect 12211 14232 12256 14260
rect 11885 14223 11943 14229
rect 12250 14220 12256 14232
rect 12308 14220 12314 14272
rect 13372 14260 13400 14300
rect 14182 14260 14188 14272
rect 13372 14232 14188 14260
rect 14182 14220 14188 14232
rect 14240 14220 14246 14272
rect 1104 14170 15824 14192
rect 1104 14118 3447 14170
rect 3499 14118 3511 14170
rect 3563 14118 3575 14170
rect 3627 14118 3639 14170
rect 3691 14118 8378 14170
rect 8430 14118 8442 14170
rect 8494 14118 8506 14170
rect 8558 14118 8570 14170
rect 8622 14118 13308 14170
rect 13360 14118 13372 14170
rect 13424 14118 13436 14170
rect 13488 14118 13500 14170
rect 13552 14118 15824 14170
rect 1104 14096 15824 14118
rect 2958 14016 2964 14068
rect 3016 14056 3022 14068
rect 5721 14059 5779 14065
rect 5721 14056 5733 14059
rect 3016 14028 5733 14056
rect 3016 14016 3022 14028
rect 5721 14025 5733 14028
rect 5767 14025 5779 14059
rect 6822 14056 6828 14068
rect 6783 14028 6828 14056
rect 5721 14019 5779 14025
rect 6822 14016 6828 14028
rect 6880 14016 6886 14068
rect 7006 14016 7012 14068
rect 7064 14056 7070 14068
rect 7837 14059 7895 14065
rect 7837 14056 7849 14059
rect 7064 14028 7849 14056
rect 7064 14016 7070 14028
rect 7837 14025 7849 14028
rect 7883 14025 7895 14059
rect 7837 14019 7895 14025
rect 8202 14016 8208 14068
rect 8260 14056 8266 14068
rect 9861 14059 9919 14065
rect 9861 14056 9873 14059
rect 8260 14028 9873 14056
rect 8260 14016 8266 14028
rect 9861 14025 9873 14028
rect 9907 14025 9919 14059
rect 9861 14019 9919 14025
rect 11164 14028 12020 14056
rect 1765 13991 1823 13997
rect 1765 13957 1777 13991
rect 1811 13988 1823 13991
rect 2774 13988 2780 14000
rect 1811 13960 2780 13988
rect 1811 13957 1823 13960
rect 1765 13951 1823 13957
rect 2774 13948 2780 13960
rect 2832 13948 2838 14000
rect 4062 13988 4068 14000
rect 2884 13960 4068 13988
rect 2222 13920 2228 13932
rect 1596 13892 2228 13920
rect 1596 13861 1624 13892
rect 2222 13880 2228 13892
rect 2280 13880 2286 13932
rect 1581 13855 1639 13861
rect 1581 13821 1593 13855
rect 1627 13821 1639 13855
rect 2130 13852 2136 13864
rect 2091 13824 2136 13852
rect 1581 13815 1639 13821
rect 2130 13812 2136 13824
rect 2188 13812 2194 13864
rect 2409 13855 2467 13861
rect 2409 13821 2421 13855
rect 2455 13852 2467 13855
rect 2774 13852 2780 13864
rect 2455 13824 2780 13852
rect 2455 13821 2467 13824
rect 2409 13815 2467 13821
rect 2774 13812 2780 13824
rect 2832 13812 2838 13864
rect 2884 13861 2912 13960
rect 4062 13948 4068 13960
rect 4120 13948 4126 14000
rect 5350 13948 5356 14000
rect 5408 13988 5414 14000
rect 8662 13988 8668 14000
rect 5408 13960 7328 13988
rect 5408 13948 5414 13960
rect 3050 13920 3056 13932
rect 3011 13892 3056 13920
rect 3050 13880 3056 13892
rect 3108 13880 3114 13932
rect 3786 13880 3792 13932
rect 3844 13920 3850 13932
rect 4249 13923 4307 13929
rect 4249 13920 4261 13923
rect 3844 13892 4261 13920
rect 3844 13880 3850 13892
rect 4249 13889 4261 13892
rect 4295 13889 4307 13923
rect 4249 13883 4307 13889
rect 4522 13880 4528 13932
rect 4580 13920 4586 13932
rect 5074 13920 5080 13932
rect 4580 13892 5080 13920
rect 4580 13880 4586 13892
rect 5074 13880 5080 13892
rect 5132 13880 5138 13932
rect 5258 13920 5264 13932
rect 5219 13892 5264 13920
rect 5258 13880 5264 13892
rect 5316 13880 5322 13932
rect 6270 13920 6276 13932
rect 6231 13892 6276 13920
rect 6270 13880 6276 13892
rect 6328 13880 6334 13932
rect 7300 13929 7328 13960
rect 8312 13960 8668 13988
rect 8312 13929 8340 13960
rect 8662 13948 8668 13960
rect 8720 13948 8726 14000
rect 8849 13991 8907 13997
rect 8849 13957 8861 13991
rect 8895 13988 8907 13991
rect 9582 13988 9588 14000
rect 8895 13960 9588 13988
rect 8895 13957 8907 13960
rect 8849 13951 8907 13957
rect 9582 13948 9588 13960
rect 9640 13948 9646 14000
rect 9766 13948 9772 14000
rect 9824 13988 9830 14000
rect 10873 13991 10931 13997
rect 10873 13988 10885 13991
rect 9824 13960 10885 13988
rect 9824 13948 9830 13960
rect 10873 13957 10885 13960
rect 10919 13957 10931 13991
rect 10873 13951 10931 13957
rect 7285 13923 7343 13929
rect 7285 13889 7297 13923
rect 7331 13889 7343 13923
rect 7285 13883 7343 13889
rect 7469 13923 7527 13929
rect 7469 13889 7481 13923
rect 7515 13920 7527 13923
rect 8297 13923 8355 13929
rect 7515 13892 8156 13920
rect 7515 13889 7527 13892
rect 7469 13883 7527 13889
rect 8128 13864 8156 13892
rect 8297 13889 8309 13923
rect 8343 13889 8355 13923
rect 8297 13883 8355 13889
rect 8389 13923 8447 13929
rect 8389 13889 8401 13923
rect 8435 13889 8447 13923
rect 8389 13883 8447 13889
rect 2869 13855 2927 13861
rect 2869 13821 2881 13855
rect 2915 13821 2927 13855
rect 5169 13855 5227 13861
rect 5169 13852 5181 13855
rect 2869 13815 2927 13821
rect 3804 13824 5181 13852
rect 3234 13744 3240 13796
rect 3292 13784 3298 13796
rect 3804 13784 3832 13824
rect 5169 13821 5181 13824
rect 5215 13821 5227 13855
rect 5169 13815 5227 13821
rect 5350 13812 5356 13864
rect 5408 13852 5414 13864
rect 6181 13855 6239 13861
rect 6181 13852 6193 13855
rect 5408 13824 6193 13852
rect 5408 13812 5414 13824
rect 6181 13821 6193 13824
rect 6227 13821 6239 13855
rect 7650 13852 7656 13864
rect 6181 13815 6239 13821
rect 6932 13824 7656 13852
rect 3292 13756 3832 13784
rect 4065 13787 4123 13793
rect 3292 13744 3298 13756
rect 4065 13753 4077 13787
rect 4111 13784 4123 13787
rect 5718 13784 5724 13796
rect 4111 13756 5724 13784
rect 4111 13753 4123 13756
rect 4065 13747 4123 13753
rect 5718 13744 5724 13756
rect 5776 13744 5782 13796
rect 6089 13787 6147 13793
rect 6089 13753 6101 13787
rect 6135 13784 6147 13787
rect 6932 13784 6960 13824
rect 7650 13812 7656 13824
rect 7708 13812 7714 13864
rect 8110 13812 8116 13864
rect 8168 13852 8174 13864
rect 8404 13852 8432 13883
rect 8938 13880 8944 13932
rect 8996 13920 9002 13932
rect 9398 13920 9404 13932
rect 8996 13892 9404 13920
rect 8996 13880 9002 13892
rect 9398 13880 9404 13892
rect 9456 13880 9462 13932
rect 9493 13923 9551 13929
rect 9493 13889 9505 13923
rect 9539 13889 9551 13923
rect 10410 13920 10416 13932
rect 10371 13892 10416 13920
rect 9493 13883 9551 13889
rect 8168 13824 8432 13852
rect 8168 13812 8174 13824
rect 9122 13812 9128 13864
rect 9180 13852 9186 13864
rect 9217 13855 9275 13861
rect 9217 13852 9229 13855
rect 9180 13824 9229 13852
rect 9180 13812 9186 13824
rect 9217 13821 9229 13824
rect 9263 13821 9275 13855
rect 9508 13852 9536 13883
rect 10410 13880 10416 13892
rect 10468 13880 10474 13932
rect 9582 13852 9588 13864
rect 9495 13824 9588 13852
rect 9217 13815 9275 13821
rect 9582 13812 9588 13824
rect 9640 13852 9646 13864
rect 9858 13852 9864 13864
rect 9640 13824 9864 13852
rect 9640 13812 9646 13824
rect 9858 13812 9864 13824
rect 9916 13812 9922 13864
rect 10321 13855 10379 13861
rect 10321 13821 10333 13855
rect 10367 13852 10379 13855
rect 11164 13852 11192 14028
rect 11992 13988 12020 14028
rect 12342 14016 12348 14068
rect 12400 14056 12406 14068
rect 12621 14059 12679 14065
rect 12621 14056 12633 14059
rect 12400 14028 12633 14056
rect 12400 14016 12406 14028
rect 12621 14025 12633 14028
rect 12667 14025 12679 14059
rect 12621 14019 12679 14025
rect 12434 13988 12440 14000
rect 11992 13960 12440 13988
rect 12434 13948 12440 13960
rect 12492 13988 12498 14000
rect 15930 13988 15936 14000
rect 12492 13960 15936 13988
rect 12492 13948 12498 13960
rect 15930 13948 15936 13960
rect 15988 13948 15994 14000
rect 11517 13923 11575 13929
rect 11517 13889 11529 13923
rect 11563 13920 11575 13923
rect 12342 13920 12348 13932
rect 11563 13892 12348 13920
rect 11563 13889 11575 13892
rect 11517 13883 11575 13889
rect 12342 13880 12348 13892
rect 12400 13880 12406 13932
rect 10367 13824 11192 13852
rect 10367 13821 10379 13824
rect 10321 13815 10379 13821
rect 11330 13812 11336 13864
rect 11388 13852 11394 13864
rect 12437 13855 12495 13861
rect 11388 13824 11433 13852
rect 11388 13812 11394 13824
rect 12437 13821 12449 13855
rect 12483 13852 12495 13855
rect 12710 13852 12716 13864
rect 12483 13824 12716 13852
rect 12483 13821 12495 13824
rect 12437 13815 12495 13821
rect 12710 13812 12716 13824
rect 12768 13812 12774 13864
rect 7190 13784 7196 13796
rect 6135 13756 6960 13784
rect 7151 13756 7196 13784
rect 6135 13753 6147 13756
rect 6089 13747 6147 13753
rect 7190 13744 7196 13756
rect 7248 13744 7254 13796
rect 8205 13787 8263 13793
rect 8205 13753 8217 13787
rect 8251 13784 8263 13787
rect 8570 13784 8576 13796
rect 8251 13756 8576 13784
rect 8251 13753 8263 13756
rect 8205 13747 8263 13753
rect 8570 13744 8576 13756
rect 8628 13744 8634 13796
rect 10229 13787 10287 13793
rect 10229 13753 10241 13787
rect 10275 13784 10287 13787
rect 10778 13784 10784 13796
rect 10275 13756 10784 13784
rect 10275 13753 10287 13756
rect 10229 13747 10287 13753
rect 10778 13744 10784 13756
rect 10836 13744 10842 13796
rect 11256 13756 11560 13784
rect 2682 13676 2688 13728
rect 2740 13716 2746 13728
rect 3697 13719 3755 13725
rect 3697 13716 3709 13719
rect 2740 13688 3709 13716
rect 2740 13676 2746 13688
rect 3697 13685 3709 13688
rect 3743 13685 3755 13719
rect 3697 13679 3755 13685
rect 3878 13676 3884 13728
rect 3936 13716 3942 13728
rect 4157 13719 4215 13725
rect 4157 13716 4169 13719
rect 3936 13688 4169 13716
rect 3936 13676 3942 13688
rect 4157 13685 4169 13688
rect 4203 13685 4215 13719
rect 4706 13716 4712 13728
rect 4667 13688 4712 13716
rect 4157 13679 4215 13685
rect 4706 13676 4712 13688
rect 4764 13676 4770 13728
rect 4798 13676 4804 13728
rect 4856 13716 4862 13728
rect 5077 13719 5135 13725
rect 5077 13716 5089 13719
rect 4856 13688 5089 13716
rect 4856 13676 4862 13688
rect 5077 13685 5089 13688
rect 5123 13685 5135 13719
rect 5077 13679 5135 13685
rect 5534 13676 5540 13728
rect 5592 13716 5598 13728
rect 7282 13716 7288 13728
rect 5592 13688 7288 13716
rect 5592 13676 5598 13688
rect 7282 13676 7288 13688
rect 7340 13676 7346 13728
rect 7926 13676 7932 13728
rect 7984 13716 7990 13728
rect 8938 13716 8944 13728
rect 7984 13688 8944 13716
rect 7984 13676 7990 13688
rect 8938 13676 8944 13688
rect 8996 13676 9002 13728
rect 9306 13676 9312 13728
rect 9364 13716 9370 13728
rect 11256 13725 11284 13756
rect 11241 13719 11299 13725
rect 9364 13688 9409 13716
rect 9364 13676 9370 13688
rect 11241 13685 11253 13719
rect 11287 13685 11299 13719
rect 11532 13716 11560 13756
rect 11606 13716 11612 13728
rect 11532 13688 11612 13716
rect 11241 13679 11299 13685
rect 11606 13676 11612 13688
rect 11664 13676 11670 13728
rect 11885 13719 11943 13725
rect 11885 13685 11897 13719
rect 11931 13716 11943 13719
rect 12434 13716 12440 13728
rect 11931 13688 12440 13716
rect 11931 13685 11943 13688
rect 11885 13679 11943 13685
rect 12434 13676 12440 13688
rect 12492 13676 12498 13728
rect 1104 13626 15824 13648
rect 1104 13574 5912 13626
rect 5964 13574 5976 13626
rect 6028 13574 6040 13626
rect 6092 13574 6104 13626
rect 6156 13574 10843 13626
rect 10895 13574 10907 13626
rect 10959 13574 10971 13626
rect 11023 13574 11035 13626
rect 11087 13574 15824 13626
rect 1104 13552 15824 13574
rect 3421 13515 3479 13521
rect 3421 13481 3433 13515
rect 3467 13512 3479 13515
rect 4338 13512 4344 13524
rect 3467 13484 4344 13512
rect 3467 13481 3479 13484
rect 3421 13475 3479 13481
rect 4338 13472 4344 13484
rect 4396 13472 4402 13524
rect 4617 13515 4675 13521
rect 4617 13481 4629 13515
rect 4663 13512 4675 13515
rect 4890 13512 4896 13524
rect 4663 13484 4896 13512
rect 4663 13481 4675 13484
rect 4617 13475 4675 13481
rect 4890 13472 4896 13484
rect 4948 13472 4954 13524
rect 5261 13515 5319 13521
rect 5261 13481 5273 13515
rect 5307 13512 5319 13515
rect 5350 13512 5356 13524
rect 5307 13484 5356 13512
rect 5307 13481 5319 13484
rect 5261 13475 5319 13481
rect 5350 13472 5356 13484
rect 5408 13472 5414 13524
rect 5629 13515 5687 13521
rect 5629 13481 5641 13515
rect 5675 13512 5687 13515
rect 7466 13512 7472 13524
rect 5675 13484 7472 13512
rect 5675 13481 5687 13484
rect 5629 13475 5687 13481
rect 7466 13472 7472 13484
rect 7524 13472 7530 13524
rect 8757 13515 8815 13521
rect 8757 13481 8769 13515
rect 8803 13512 8815 13515
rect 9950 13512 9956 13524
rect 8803 13484 9956 13512
rect 8803 13481 8815 13484
rect 8757 13475 8815 13481
rect 9950 13472 9956 13484
rect 10008 13472 10014 13524
rect 10137 13515 10195 13521
rect 10137 13481 10149 13515
rect 10183 13512 10195 13515
rect 11057 13515 11115 13521
rect 10183 13484 11008 13512
rect 10183 13481 10195 13484
rect 10137 13475 10195 13481
rect 4706 13444 4712 13456
rect 2240 13416 4712 13444
rect 2240 13385 2268 13416
rect 4706 13404 4712 13416
rect 4764 13404 4770 13456
rect 6914 13444 6920 13456
rect 6288 13416 6920 13444
rect 1489 13379 1547 13385
rect 1489 13345 1501 13379
rect 1535 13376 1547 13379
rect 2225 13379 2283 13385
rect 1535 13348 2176 13376
rect 1535 13345 1547 13348
rect 1489 13339 1547 13345
rect 1670 13308 1676 13320
rect 1631 13280 1676 13308
rect 1670 13268 1676 13280
rect 1728 13268 1734 13320
rect 2148 13308 2176 13348
rect 2225 13345 2237 13379
rect 2271 13345 2283 13379
rect 2225 13339 2283 13345
rect 2501 13379 2559 13385
rect 2501 13345 2513 13379
rect 2547 13376 2559 13379
rect 2866 13376 2872 13388
rect 2547 13348 2872 13376
rect 2547 13345 2559 13348
rect 2501 13339 2559 13345
rect 2866 13336 2872 13348
rect 2924 13336 2930 13388
rect 3050 13336 3056 13388
rect 3108 13376 3114 13388
rect 3329 13379 3387 13385
rect 3329 13376 3341 13379
rect 3108 13348 3341 13376
rect 3108 13336 3114 13348
rect 3329 13345 3341 13348
rect 3375 13345 3387 13379
rect 3329 13339 3387 13345
rect 5534 13336 5540 13388
rect 5592 13376 5598 13388
rect 6288 13385 6316 13416
rect 6914 13404 6920 13416
rect 6972 13404 6978 13456
rect 7926 13404 7932 13456
rect 7984 13444 7990 13456
rect 8202 13444 8208 13456
rect 7984 13416 8208 13444
rect 7984 13404 7990 13416
rect 8202 13404 8208 13416
rect 8260 13444 8266 13456
rect 8297 13447 8355 13453
rect 8297 13444 8309 13447
rect 8260 13416 8309 13444
rect 8260 13404 8266 13416
rect 8297 13413 8309 13416
rect 8343 13413 8355 13447
rect 8297 13407 8355 13413
rect 8570 13404 8576 13456
rect 8628 13444 8634 13456
rect 10042 13444 10048 13456
rect 8628 13416 9904 13444
rect 9955 13416 10048 13444
rect 8628 13404 8634 13416
rect 6273 13379 6331 13385
rect 5592 13348 5856 13376
rect 5592 13336 5598 13348
rect 2958 13308 2964 13320
rect 2148 13280 2964 13308
rect 2958 13268 2964 13280
rect 3016 13268 3022 13320
rect 3605 13311 3663 13317
rect 3605 13277 3617 13311
rect 3651 13308 3663 13311
rect 3970 13308 3976 13320
rect 3651 13280 3976 13308
rect 3651 13277 3663 13280
rect 3605 13271 3663 13277
rect 3970 13268 3976 13280
rect 4028 13268 4034 13320
rect 4706 13308 4712 13320
rect 4667 13280 4712 13308
rect 4706 13268 4712 13280
rect 4764 13268 4770 13320
rect 4893 13311 4951 13317
rect 4893 13277 4905 13311
rect 4939 13277 4951 13311
rect 4893 13271 4951 13277
rect 4908 13240 4936 13271
rect 5074 13268 5080 13320
rect 5132 13308 5138 13320
rect 5828 13317 5856 13348
rect 6273 13345 6285 13379
rect 6319 13345 6331 13379
rect 6273 13339 6331 13345
rect 6540 13379 6598 13385
rect 6540 13345 6552 13379
rect 6586 13376 6598 13379
rect 7650 13376 7656 13388
rect 6586 13348 7656 13376
rect 6586 13345 6598 13348
rect 6540 13339 6598 13345
rect 7650 13336 7656 13348
rect 7708 13336 7714 13388
rect 7834 13336 7840 13388
rect 7892 13376 7898 13388
rect 8389 13379 8447 13385
rect 8389 13376 8401 13379
rect 7892 13348 8401 13376
rect 7892 13336 7898 13348
rect 8389 13345 8401 13348
rect 8435 13376 8447 13379
rect 8662 13376 8668 13388
rect 8435 13348 8668 13376
rect 8435 13345 8447 13348
rect 8389 13339 8447 13345
rect 8662 13336 8668 13348
rect 8720 13336 8726 13388
rect 8941 13379 8999 13385
rect 8941 13345 8953 13379
rect 8987 13376 8999 13379
rect 9122 13376 9128 13388
rect 8987 13348 9128 13376
rect 8987 13345 8999 13348
rect 8941 13339 8999 13345
rect 9122 13336 9128 13348
rect 9180 13336 9186 13388
rect 9876 13376 9904 13416
rect 10042 13404 10048 13416
rect 10100 13444 10106 13456
rect 10870 13444 10876 13456
rect 10100 13416 10876 13444
rect 10100 13404 10106 13416
rect 10870 13404 10876 13416
rect 10928 13404 10934 13456
rect 10980 13444 11008 13484
rect 11057 13481 11069 13515
rect 11103 13512 11115 13515
rect 11330 13512 11336 13524
rect 11103 13484 11336 13512
rect 11103 13481 11115 13484
rect 11057 13475 11115 13481
rect 11330 13472 11336 13484
rect 11388 13472 11394 13524
rect 11698 13512 11704 13524
rect 11659 13484 11704 13512
rect 11698 13472 11704 13484
rect 11756 13472 11762 13524
rect 12158 13512 12164 13524
rect 12119 13484 12164 13512
rect 12158 13472 12164 13484
rect 12216 13472 12222 13524
rect 12894 13444 12900 13456
rect 10980 13416 12900 13444
rect 12894 13404 12900 13416
rect 12952 13404 12958 13456
rect 13998 13444 14004 13456
rect 13959 13416 14004 13444
rect 13998 13404 14004 13416
rect 14056 13404 14062 13456
rect 12069 13379 12127 13385
rect 9876 13348 12020 13376
rect 5721 13311 5779 13317
rect 5721 13308 5733 13311
rect 5132 13280 5733 13308
rect 5132 13268 5138 13280
rect 5721 13277 5733 13280
rect 5767 13277 5779 13311
rect 5721 13271 5779 13277
rect 5813 13311 5871 13317
rect 5813 13277 5825 13311
rect 5859 13277 5871 13311
rect 5813 13271 5871 13277
rect 8573 13311 8631 13317
rect 8573 13277 8585 13311
rect 8619 13308 8631 13311
rect 9214 13308 9220 13320
rect 8619 13280 9220 13308
rect 8619 13277 8631 13280
rect 8573 13271 8631 13277
rect 9214 13268 9220 13280
rect 9272 13268 9278 13320
rect 10042 13308 10048 13320
rect 9692 13280 10048 13308
rect 5534 13240 5540 13252
rect 4908 13212 5540 13240
rect 5534 13200 5540 13212
rect 5592 13200 5598 13252
rect 7929 13243 7987 13249
rect 7929 13209 7941 13243
rect 7975 13240 7987 13243
rect 8757 13243 8815 13249
rect 8757 13240 8769 13243
rect 7975 13212 8769 13240
rect 7975 13209 7987 13212
rect 7929 13203 7987 13209
rect 8757 13209 8769 13212
rect 8803 13209 8815 13243
rect 8757 13203 8815 13209
rect 8938 13200 8944 13252
rect 8996 13240 9002 13252
rect 9692 13249 9720 13280
rect 10042 13268 10048 13280
rect 10100 13268 10106 13320
rect 10321 13311 10379 13317
rect 10321 13277 10333 13311
rect 10367 13277 10379 13311
rect 10321 13271 10379 13277
rect 9125 13243 9183 13249
rect 9125 13240 9137 13243
rect 8996 13212 9137 13240
rect 8996 13200 9002 13212
rect 9125 13209 9137 13212
rect 9171 13209 9183 13243
rect 9125 13203 9183 13209
rect 9677 13243 9735 13249
rect 9677 13209 9689 13243
rect 9723 13209 9735 13243
rect 9677 13203 9735 13209
rect 9858 13200 9864 13252
rect 9916 13240 9922 13252
rect 10336 13240 10364 13271
rect 10410 13268 10416 13320
rect 10468 13308 10474 13320
rect 11149 13311 11207 13317
rect 11149 13308 11161 13311
rect 10468 13280 11161 13308
rect 10468 13268 10474 13280
rect 11149 13277 11161 13280
rect 11195 13277 11207 13311
rect 11330 13308 11336 13320
rect 11291 13280 11336 13308
rect 11149 13271 11207 13277
rect 11330 13268 11336 13280
rect 11388 13268 11394 13320
rect 10962 13240 10968 13252
rect 9916 13212 10968 13240
rect 9916 13200 9922 13212
rect 10962 13200 10968 13212
rect 11020 13200 11026 13252
rect 11054 13200 11060 13252
rect 11112 13240 11118 13252
rect 11422 13240 11428 13252
rect 11112 13212 11428 13240
rect 11112 13200 11118 13212
rect 11422 13200 11428 13212
rect 11480 13200 11486 13252
rect 11992 13240 12020 13348
rect 12069 13345 12081 13379
rect 12115 13376 12127 13379
rect 13078 13376 13084 13388
rect 12115 13348 12480 13376
rect 13039 13348 13084 13376
rect 12115 13345 12127 13348
rect 12069 13339 12127 13345
rect 12158 13268 12164 13320
rect 12216 13308 12222 13320
rect 12253 13311 12311 13317
rect 12253 13308 12265 13311
rect 12216 13280 12265 13308
rect 12216 13268 12222 13280
rect 12253 13277 12265 13280
rect 12299 13277 12311 13311
rect 12452 13308 12480 13348
rect 13078 13336 13084 13348
rect 13136 13336 13142 13388
rect 13725 13379 13783 13385
rect 13725 13376 13737 13379
rect 13556 13348 13737 13376
rect 13170 13308 13176 13320
rect 12452 13280 12664 13308
rect 13131 13280 13176 13308
rect 12253 13271 12311 13277
rect 12342 13240 12348 13252
rect 11992 13212 12348 13240
rect 12342 13200 12348 13212
rect 12400 13200 12406 13252
rect 2961 13175 3019 13181
rect 2961 13141 2973 13175
rect 3007 13172 3019 13175
rect 3142 13172 3148 13184
rect 3007 13144 3148 13172
rect 3007 13141 3019 13144
rect 2961 13135 3019 13141
rect 3142 13132 3148 13144
rect 3200 13132 3206 13184
rect 4154 13132 4160 13184
rect 4212 13172 4218 13184
rect 4249 13175 4307 13181
rect 4249 13172 4261 13175
rect 4212 13144 4261 13172
rect 4212 13132 4218 13144
rect 4249 13141 4261 13144
rect 4295 13141 4307 13175
rect 4249 13135 4307 13141
rect 4430 13132 4436 13184
rect 4488 13172 4494 13184
rect 5166 13172 5172 13184
rect 4488 13144 5172 13172
rect 4488 13132 4494 13144
rect 5166 13132 5172 13144
rect 5224 13132 5230 13184
rect 6546 13132 6552 13184
rect 6604 13172 6610 13184
rect 7653 13175 7711 13181
rect 7653 13172 7665 13175
rect 6604 13144 7665 13172
rect 6604 13132 6610 13144
rect 7653 13141 7665 13144
rect 7699 13141 7711 13175
rect 7653 13135 7711 13141
rect 8202 13132 8208 13184
rect 8260 13172 8266 13184
rect 10689 13175 10747 13181
rect 10689 13172 10701 13175
rect 8260 13144 10701 13172
rect 8260 13132 8266 13144
rect 10689 13141 10701 13144
rect 10735 13141 10747 13175
rect 10689 13135 10747 13141
rect 10778 13132 10784 13184
rect 10836 13172 10842 13184
rect 11514 13172 11520 13184
rect 10836 13144 11520 13172
rect 10836 13132 10842 13144
rect 11514 13132 11520 13144
rect 11572 13132 11578 13184
rect 12636 13172 12664 13280
rect 13170 13268 13176 13280
rect 13228 13268 13234 13320
rect 13357 13311 13415 13317
rect 13357 13277 13369 13311
rect 13403 13308 13415 13311
rect 13446 13308 13452 13320
rect 13403 13280 13452 13308
rect 13403 13277 13415 13280
rect 13357 13271 13415 13277
rect 13446 13268 13452 13280
rect 13504 13268 13510 13320
rect 12713 13243 12771 13249
rect 12713 13209 12725 13243
rect 12759 13240 12771 13243
rect 13556 13240 13584 13348
rect 13725 13345 13737 13348
rect 13771 13345 13783 13379
rect 13725 13339 13783 13345
rect 12759 13212 13584 13240
rect 12759 13209 12771 13212
rect 12713 13203 12771 13209
rect 13722 13172 13728 13184
rect 12636 13144 13728 13172
rect 13722 13132 13728 13144
rect 13780 13132 13786 13184
rect 1104 13082 15824 13104
rect 1104 13030 3447 13082
rect 3499 13030 3511 13082
rect 3563 13030 3575 13082
rect 3627 13030 3639 13082
rect 3691 13030 8378 13082
rect 8430 13030 8442 13082
rect 8494 13030 8506 13082
rect 8558 13030 8570 13082
rect 8622 13030 13308 13082
rect 13360 13030 13372 13082
rect 13424 13030 13436 13082
rect 13488 13030 13500 13082
rect 13552 13030 15824 13082
rect 1104 13008 15824 13030
rect 5994 12928 6000 12980
rect 6052 12968 6058 12980
rect 6549 12971 6607 12977
rect 6549 12968 6561 12971
rect 6052 12940 6561 12968
rect 6052 12928 6058 12940
rect 6549 12937 6561 12940
rect 6595 12937 6607 12971
rect 6549 12931 6607 12937
rect 6641 12971 6699 12977
rect 6641 12937 6653 12971
rect 6687 12968 6699 12971
rect 6822 12968 6828 12980
rect 6687 12940 6828 12968
rect 6687 12937 6699 12940
rect 6641 12931 6699 12937
rect 6822 12928 6828 12940
rect 6880 12928 6886 12980
rect 7006 12928 7012 12980
rect 7064 12968 7070 12980
rect 8205 12971 8263 12977
rect 8205 12968 8217 12971
rect 7064 12940 8217 12968
rect 7064 12928 7070 12940
rect 8205 12937 8217 12940
rect 8251 12937 8263 12971
rect 9490 12968 9496 12980
rect 9451 12940 9496 12968
rect 8205 12931 8263 12937
rect 9490 12928 9496 12940
rect 9548 12928 9554 12980
rect 10042 12928 10048 12980
rect 10100 12968 10106 12980
rect 10413 12971 10471 12977
rect 10413 12968 10425 12971
rect 10100 12940 10425 12968
rect 10100 12928 10106 12940
rect 10413 12937 10425 12940
rect 10459 12937 10471 12971
rect 10413 12931 10471 12937
rect 11054 12928 11060 12980
rect 11112 12968 11118 12980
rect 11701 12971 11759 12977
rect 11701 12968 11713 12971
rect 11112 12940 11713 12968
rect 11112 12928 11118 12940
rect 11701 12937 11713 12940
rect 11747 12937 11759 12971
rect 11701 12931 11759 12937
rect 12158 12928 12164 12980
rect 12216 12968 12222 12980
rect 12216 12940 12848 12968
rect 12216 12928 12222 12940
rect 8478 12900 8484 12912
rect 4356 12872 6868 12900
rect 8439 12872 8484 12900
rect 2317 12835 2375 12841
rect 2317 12801 2329 12835
rect 2363 12832 2375 12835
rect 2866 12832 2872 12844
rect 2363 12804 2872 12832
rect 2363 12801 2375 12804
rect 2317 12795 2375 12801
rect 2866 12792 2872 12804
rect 2924 12792 2930 12844
rect 3142 12832 3148 12844
rect 3103 12804 3148 12832
rect 3142 12792 3148 12804
rect 3200 12792 3206 12844
rect 3237 12835 3295 12841
rect 3237 12801 3249 12835
rect 3283 12801 3295 12835
rect 4154 12832 4160 12844
rect 4115 12804 4160 12832
rect 3237 12795 3295 12801
rect 2590 12724 2596 12776
rect 2648 12764 2654 12776
rect 3252 12764 3280 12795
rect 4154 12792 4160 12804
rect 4212 12792 4218 12844
rect 4356 12841 4384 12872
rect 4341 12835 4399 12841
rect 4341 12801 4353 12835
rect 4387 12801 4399 12835
rect 4341 12795 4399 12801
rect 4890 12792 4896 12844
rect 4948 12832 4954 12844
rect 5261 12835 5319 12841
rect 5261 12832 5273 12835
rect 4948 12804 5273 12832
rect 4948 12792 4954 12804
rect 5261 12801 5273 12804
rect 5307 12801 5319 12835
rect 6362 12832 6368 12844
rect 6275 12804 6368 12832
rect 5261 12795 5319 12801
rect 6362 12792 6368 12804
rect 6420 12832 6426 12844
rect 6546 12832 6552 12844
rect 6420 12804 6552 12832
rect 6420 12792 6426 12804
rect 6546 12792 6552 12804
rect 6604 12792 6610 12844
rect 6840 12832 6868 12872
rect 8478 12860 8484 12872
rect 8536 12860 8542 12912
rect 10226 12900 10232 12912
rect 9508 12872 10232 12900
rect 9508 12844 9536 12872
rect 10226 12860 10232 12872
rect 10284 12860 10290 12912
rect 10505 12903 10563 12909
rect 10505 12869 10517 12903
rect 10551 12900 10563 12903
rect 12066 12900 12072 12912
rect 10551 12872 12072 12900
rect 10551 12869 10563 12872
rect 10505 12863 10563 12869
rect 12066 12860 12072 12872
rect 12124 12860 12130 12912
rect 12434 12900 12440 12912
rect 12395 12872 12440 12900
rect 12434 12860 12440 12872
rect 12492 12860 12498 12912
rect 12820 12900 12848 12940
rect 13078 12928 13084 12980
rect 13136 12968 13142 12980
rect 13449 12971 13507 12977
rect 13449 12968 13461 12971
rect 13136 12940 13461 12968
rect 13136 12928 13142 12940
rect 13449 12937 13461 12940
rect 13495 12937 13507 12971
rect 13449 12931 13507 12937
rect 13814 12900 13820 12912
rect 12820 12872 13124 12900
rect 6840 12804 6960 12832
rect 2648 12736 3280 12764
rect 2648 12724 2654 12736
rect 3694 12724 3700 12776
rect 3752 12764 3758 12776
rect 4065 12767 4123 12773
rect 4065 12764 4077 12767
rect 3752 12736 4077 12764
rect 3752 12724 3758 12736
rect 4065 12733 4077 12736
rect 4111 12733 4123 12767
rect 4430 12764 4436 12776
rect 4065 12727 4123 12733
rect 4172 12736 4436 12764
rect 3053 12699 3111 12705
rect 3053 12665 3065 12699
rect 3099 12696 3111 12699
rect 4172 12696 4200 12736
rect 4430 12724 4436 12736
rect 4488 12724 4494 12776
rect 5077 12767 5135 12773
rect 5077 12733 5089 12767
rect 5123 12764 5135 12767
rect 5718 12764 5724 12776
rect 5123 12736 5724 12764
rect 5123 12733 5135 12736
rect 5077 12727 5135 12733
rect 5718 12724 5724 12736
rect 5776 12724 5782 12776
rect 6178 12764 6184 12776
rect 6139 12736 6184 12764
rect 6178 12724 6184 12736
rect 6236 12724 6242 12776
rect 6733 12767 6791 12773
rect 6733 12733 6745 12767
rect 6779 12764 6791 12767
rect 6825 12767 6883 12773
rect 6825 12764 6837 12767
rect 6779 12736 6837 12764
rect 6779 12733 6791 12736
rect 6733 12727 6791 12733
rect 6825 12733 6837 12736
rect 6871 12733 6883 12767
rect 6932 12764 6960 12804
rect 8294 12792 8300 12844
rect 8352 12832 8358 12844
rect 8941 12835 8999 12841
rect 8941 12832 8953 12835
rect 8352 12804 8953 12832
rect 8352 12792 8358 12804
rect 8941 12801 8953 12804
rect 8987 12801 8999 12835
rect 8941 12795 8999 12801
rect 9033 12835 9091 12841
rect 9033 12801 9045 12835
rect 9079 12832 9091 12835
rect 9214 12832 9220 12844
rect 9079 12804 9220 12832
rect 9079 12801 9091 12804
rect 9033 12795 9091 12801
rect 7081 12767 7139 12773
rect 7081 12764 7093 12767
rect 6932 12736 7093 12764
rect 6825 12727 6883 12733
rect 7081 12733 7093 12736
rect 7127 12733 7139 12767
rect 7081 12727 7139 12733
rect 3099 12668 4200 12696
rect 3099 12665 3111 12668
rect 3053 12659 3111 12665
rect 4246 12656 4252 12708
rect 4304 12696 4310 12708
rect 4304 12668 5764 12696
rect 4304 12656 4310 12668
rect 1578 12588 1584 12640
rect 1636 12628 1642 12640
rect 1673 12631 1731 12637
rect 1673 12628 1685 12631
rect 1636 12600 1685 12628
rect 1636 12588 1642 12600
rect 1673 12597 1685 12600
rect 1719 12597 1731 12631
rect 2038 12628 2044 12640
rect 1999 12600 2044 12628
rect 1673 12591 1731 12597
rect 2038 12588 2044 12600
rect 2096 12588 2102 12640
rect 2133 12631 2191 12637
rect 2133 12597 2145 12631
rect 2179 12628 2191 12631
rect 2685 12631 2743 12637
rect 2685 12628 2697 12631
rect 2179 12600 2697 12628
rect 2179 12597 2191 12600
rect 2133 12591 2191 12597
rect 2685 12597 2697 12600
rect 2731 12597 2743 12631
rect 3694 12628 3700 12640
rect 3655 12600 3700 12628
rect 2685 12591 2743 12597
rect 3694 12588 3700 12600
rect 3752 12588 3758 12640
rect 4154 12588 4160 12640
rect 4212 12628 4218 12640
rect 4709 12631 4767 12637
rect 4709 12628 4721 12631
rect 4212 12600 4721 12628
rect 4212 12588 4218 12600
rect 4709 12597 4721 12600
rect 4755 12597 4767 12631
rect 4709 12591 4767 12597
rect 5169 12631 5227 12637
rect 5169 12597 5181 12631
rect 5215 12628 5227 12631
rect 5442 12628 5448 12640
rect 5215 12600 5448 12628
rect 5215 12597 5227 12600
rect 5169 12591 5227 12597
rect 5442 12588 5448 12600
rect 5500 12588 5506 12640
rect 5736 12637 5764 12668
rect 5994 12656 6000 12708
rect 6052 12696 6058 12708
rect 6089 12699 6147 12705
rect 6089 12696 6101 12699
rect 6052 12668 6101 12696
rect 6052 12656 6058 12668
rect 6089 12665 6101 12668
rect 6135 12665 6147 12699
rect 6089 12659 6147 12665
rect 5721 12631 5779 12637
rect 5721 12597 5733 12631
rect 5767 12597 5779 12631
rect 5721 12591 5779 12597
rect 6641 12631 6699 12637
rect 6641 12597 6653 12631
rect 6687 12628 6699 12631
rect 6822 12628 6828 12640
rect 6687 12600 6828 12628
rect 6687 12597 6699 12600
rect 6641 12591 6699 12597
rect 6822 12588 6828 12600
rect 6880 12588 6886 12640
rect 7107 12628 7135 12727
rect 8754 12724 8760 12776
rect 8812 12764 8818 12776
rect 9048 12764 9076 12795
rect 9214 12792 9220 12804
rect 9272 12792 9278 12844
rect 9490 12792 9496 12844
rect 9548 12792 9554 12844
rect 10042 12832 10048 12844
rect 10003 12804 10048 12832
rect 10042 12792 10048 12804
rect 10100 12792 10106 12844
rect 10686 12792 10692 12844
rect 10744 12832 10750 12844
rect 10965 12835 11023 12841
rect 10965 12832 10977 12835
rect 10744 12804 10977 12832
rect 10744 12792 10750 12804
rect 10965 12801 10977 12804
rect 11011 12801 11023 12835
rect 10965 12795 11023 12801
rect 11054 12792 11060 12844
rect 11112 12832 11118 12844
rect 11149 12835 11207 12841
rect 11149 12832 11161 12835
rect 11112 12804 11161 12832
rect 11112 12792 11118 12804
rect 11149 12801 11161 12804
rect 11195 12832 11207 12835
rect 11698 12832 11704 12844
rect 11195 12804 11704 12832
rect 11195 12801 11207 12804
rect 11149 12795 11207 12801
rect 11698 12792 11704 12804
rect 11756 12792 11762 12844
rect 12158 12792 12164 12844
rect 12216 12832 12222 12844
rect 13096 12841 13124 12872
rect 13188 12872 13820 12900
rect 13081 12835 13139 12841
rect 12216 12804 13032 12832
rect 12216 12792 12222 12804
rect 8812 12736 9076 12764
rect 9861 12767 9919 12773
rect 8812 12724 8818 12736
rect 9861 12733 9873 12767
rect 9907 12764 9919 12767
rect 10873 12767 10931 12773
rect 9907 12736 9976 12764
rect 9907 12733 9919 12736
rect 9861 12727 9919 12733
rect 8849 12699 8907 12705
rect 8849 12665 8861 12699
rect 8895 12696 8907 12699
rect 8938 12696 8944 12708
rect 8895 12668 8944 12696
rect 8895 12665 8907 12668
rect 8849 12659 8907 12665
rect 8938 12656 8944 12668
rect 8996 12656 9002 12708
rect 9122 12656 9128 12708
rect 9180 12696 9186 12708
rect 9582 12696 9588 12708
rect 9180 12668 9588 12696
rect 9180 12656 9186 12668
rect 9582 12656 9588 12668
rect 9640 12656 9646 12708
rect 9948 12696 9976 12736
rect 10873 12733 10885 12767
rect 10919 12764 10931 12767
rect 11238 12764 11244 12776
rect 10919 12736 11244 12764
rect 10919 12733 10931 12736
rect 10873 12727 10931 12733
rect 11238 12724 11244 12736
rect 11296 12724 11302 12776
rect 11517 12767 11575 12773
rect 11517 12733 11529 12767
rect 11563 12733 11575 12767
rect 11517 12727 11575 12733
rect 10962 12696 10968 12708
rect 9948 12668 10968 12696
rect 10962 12656 10968 12668
rect 11020 12696 11026 12708
rect 11422 12696 11428 12708
rect 11020 12668 11428 12696
rect 11020 12656 11026 12668
rect 11422 12656 11428 12668
rect 11480 12656 11486 12708
rect 11532 12696 11560 12727
rect 11974 12724 11980 12776
rect 12032 12764 12038 12776
rect 12253 12767 12311 12773
rect 12253 12764 12265 12767
rect 12032 12736 12265 12764
rect 12032 12724 12038 12736
rect 12253 12733 12265 12736
rect 12299 12733 12311 12767
rect 12894 12764 12900 12776
rect 12253 12727 12311 12733
rect 12544 12736 12756 12764
rect 12855 12736 12900 12764
rect 12544 12696 12572 12736
rect 11532 12668 12572 12696
rect 12728 12696 12756 12736
rect 12894 12724 12900 12736
rect 12952 12724 12958 12776
rect 13004 12764 13032 12804
rect 13081 12801 13093 12835
rect 13127 12801 13139 12835
rect 13081 12795 13139 12801
rect 13188 12764 13216 12872
rect 13814 12860 13820 12872
rect 13872 12900 13878 12912
rect 14366 12900 14372 12912
rect 13872 12872 14372 12900
rect 13872 12860 13878 12872
rect 14366 12860 14372 12872
rect 14424 12860 14430 12912
rect 13262 12792 13268 12844
rect 13320 12832 13326 12844
rect 14001 12835 14059 12841
rect 14001 12832 14013 12835
rect 13320 12804 14013 12832
rect 13320 12792 13326 12804
rect 14001 12801 14013 12804
rect 14047 12801 14059 12835
rect 14001 12795 14059 12801
rect 13004 12736 13216 12764
rect 13817 12767 13875 12773
rect 13817 12733 13829 12767
rect 13863 12764 13875 12767
rect 14182 12764 14188 12776
rect 13863 12736 14188 12764
rect 13863 12733 13875 12736
rect 13817 12727 13875 12733
rect 14182 12724 14188 12736
rect 14240 12724 14246 12776
rect 15378 12696 15384 12708
rect 12728 12668 15384 12696
rect 15378 12656 15384 12668
rect 15436 12656 15442 12708
rect 9490 12628 9496 12640
rect 7107 12600 9496 12628
rect 9490 12588 9496 12600
rect 9548 12588 9554 12640
rect 9953 12631 10011 12637
rect 9953 12597 9965 12631
rect 9999 12628 10011 12631
rect 10318 12628 10324 12640
rect 9999 12600 10324 12628
rect 9999 12597 10011 12600
rect 9953 12591 10011 12597
rect 10318 12588 10324 12600
rect 10376 12588 10382 12640
rect 10413 12631 10471 12637
rect 10413 12597 10425 12631
rect 10459 12628 10471 12631
rect 11238 12628 11244 12640
rect 10459 12600 11244 12628
rect 10459 12597 10471 12600
rect 10413 12591 10471 12597
rect 11238 12588 11244 12600
rect 11296 12588 11302 12640
rect 12069 12631 12127 12637
rect 12069 12597 12081 12631
rect 12115 12628 12127 12631
rect 12158 12628 12164 12640
rect 12115 12600 12164 12628
rect 12115 12597 12127 12600
rect 12069 12591 12127 12597
rect 12158 12588 12164 12600
rect 12216 12588 12222 12640
rect 12802 12628 12808 12640
rect 12763 12600 12808 12628
rect 12802 12588 12808 12600
rect 12860 12588 12866 12640
rect 13446 12588 13452 12640
rect 13504 12628 13510 12640
rect 13722 12628 13728 12640
rect 13504 12600 13728 12628
rect 13504 12588 13510 12600
rect 13722 12588 13728 12600
rect 13780 12588 13786 12640
rect 13909 12631 13967 12637
rect 13909 12597 13921 12631
rect 13955 12628 13967 12631
rect 14918 12628 14924 12640
rect 13955 12600 14924 12628
rect 13955 12597 13967 12600
rect 13909 12591 13967 12597
rect 14918 12588 14924 12600
rect 14976 12588 14982 12640
rect 1104 12538 15824 12560
rect 1104 12486 5912 12538
rect 5964 12486 5976 12538
rect 6028 12486 6040 12538
rect 6092 12486 6104 12538
rect 6156 12486 10843 12538
rect 10895 12486 10907 12538
rect 10959 12486 10971 12538
rect 11023 12486 11035 12538
rect 11087 12486 15824 12538
rect 1104 12464 15824 12486
rect 1949 12427 2007 12433
rect 1949 12393 1961 12427
rect 1995 12424 2007 12427
rect 2038 12424 2044 12436
rect 1995 12396 2044 12424
rect 1995 12393 2007 12396
rect 1949 12387 2007 12393
rect 2038 12384 2044 12396
rect 2096 12384 2102 12436
rect 2961 12427 3019 12433
rect 2961 12393 2973 12427
rect 3007 12424 3019 12427
rect 3234 12424 3240 12436
rect 3007 12396 3240 12424
rect 3007 12393 3019 12396
rect 2961 12387 3019 12393
rect 3234 12384 3240 12396
rect 3292 12384 3298 12436
rect 3421 12427 3479 12433
rect 3421 12393 3433 12427
rect 3467 12424 3479 12427
rect 3694 12424 3700 12436
rect 3467 12396 3700 12424
rect 3467 12393 3479 12396
rect 3421 12387 3479 12393
rect 3694 12384 3700 12396
rect 3752 12384 3758 12436
rect 4062 12424 4068 12436
rect 4023 12396 4068 12424
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 4522 12424 4528 12436
rect 4483 12396 4528 12424
rect 4522 12384 4528 12396
rect 4580 12384 4586 12436
rect 8478 12384 8484 12436
rect 8536 12424 8542 12436
rect 8536 12396 9352 12424
rect 8536 12384 8542 12396
rect 2498 12356 2504 12368
rect 1872 12328 2504 12356
rect 1872 12297 1900 12328
rect 2498 12316 2504 12328
rect 2556 12316 2562 12368
rect 3142 12316 3148 12368
rect 3200 12356 3206 12368
rect 3970 12356 3976 12368
rect 3200 12328 3976 12356
rect 3200 12316 3206 12328
rect 3970 12316 3976 12328
rect 4028 12316 4034 12368
rect 4430 12356 4436 12368
rect 4391 12328 4436 12356
rect 4430 12316 4436 12328
rect 4488 12316 4494 12368
rect 5344 12359 5402 12365
rect 5344 12356 5356 12359
rect 4816 12328 5356 12356
rect 1857 12291 1915 12297
rect 1857 12257 1869 12291
rect 1903 12257 1915 12291
rect 2314 12288 2320 12300
rect 2275 12260 2320 12288
rect 1857 12251 1915 12257
rect 2314 12248 2320 12260
rect 2372 12248 2378 12300
rect 3329 12291 3387 12297
rect 3329 12257 3341 12291
rect 3375 12288 3387 12291
rect 3789 12291 3847 12297
rect 3789 12288 3801 12291
rect 3375 12260 3801 12288
rect 3375 12257 3387 12260
rect 3329 12251 3387 12257
rect 3789 12257 3801 12260
rect 3835 12257 3847 12291
rect 3789 12251 3847 12257
rect 4816 12232 4844 12328
rect 5344 12325 5356 12328
rect 5390 12356 5402 12359
rect 6362 12356 6368 12368
rect 5390 12328 6368 12356
rect 5390 12325 5402 12328
rect 5344 12319 5402 12325
rect 6362 12316 6368 12328
rect 6420 12316 6426 12368
rect 6546 12316 6552 12368
rect 6604 12356 6610 12368
rect 6978 12359 7036 12365
rect 6978 12356 6990 12359
rect 6604 12328 6990 12356
rect 6604 12316 6610 12328
rect 6978 12325 6990 12328
rect 7024 12356 7036 12359
rect 9324 12356 9352 12396
rect 9398 12384 9404 12436
rect 9456 12424 9462 12436
rect 9677 12427 9735 12433
rect 9677 12424 9689 12427
rect 9456 12396 9689 12424
rect 9456 12384 9462 12396
rect 9677 12393 9689 12396
rect 9723 12393 9735 12427
rect 9677 12387 9735 12393
rect 11422 12384 11428 12436
rect 11480 12424 11486 12436
rect 11974 12424 11980 12436
rect 11480 12396 11980 12424
rect 11480 12384 11486 12396
rect 11974 12384 11980 12396
rect 12032 12384 12038 12436
rect 12066 12384 12072 12436
rect 12124 12424 12130 12436
rect 13170 12424 13176 12436
rect 12124 12396 12169 12424
rect 13131 12396 13176 12424
rect 12124 12384 12130 12396
rect 13170 12384 13176 12396
rect 13228 12384 13234 12436
rect 13446 12384 13452 12436
rect 13504 12424 13510 12436
rect 13725 12427 13783 12433
rect 13725 12424 13737 12427
rect 13504 12396 13737 12424
rect 13504 12384 13510 12396
rect 13725 12393 13737 12396
rect 13771 12393 13783 12427
rect 14182 12424 14188 12436
rect 14095 12396 14188 12424
rect 13725 12387 13783 12393
rect 14182 12384 14188 12396
rect 14240 12424 14246 12436
rect 16758 12424 16764 12436
rect 14240 12396 16764 12424
rect 14240 12384 14246 12396
rect 16758 12384 16764 12396
rect 16816 12384 16822 12436
rect 10045 12359 10103 12365
rect 10045 12356 10057 12359
rect 7024 12328 9260 12356
rect 9324 12328 10057 12356
rect 7024 12325 7036 12328
rect 6978 12319 7036 12325
rect 5074 12288 5080 12300
rect 4987 12260 5080 12288
rect 5074 12248 5080 12260
rect 5132 12288 5138 12300
rect 6733 12291 6791 12297
rect 6733 12288 6745 12291
rect 5132 12260 6745 12288
rect 5132 12248 5138 12260
rect 6733 12257 6745 12260
rect 6779 12288 6791 12291
rect 6822 12288 6828 12300
rect 6779 12260 6828 12288
rect 6779 12257 6791 12260
rect 6733 12251 6791 12257
rect 6822 12248 6828 12260
rect 6880 12248 6886 12300
rect 8754 12288 8760 12300
rect 8715 12260 8760 12288
rect 8754 12248 8760 12260
rect 8812 12248 8818 12300
rect 9232 12288 9260 12328
rect 10045 12325 10057 12328
rect 10091 12325 10103 12359
rect 10045 12319 10103 12325
rect 10612 12328 14228 12356
rect 10612 12300 10640 12328
rect 9232 12260 9536 12288
rect 2406 12220 2412 12232
rect 2367 12192 2412 12220
rect 2406 12180 2412 12192
rect 2464 12180 2470 12232
rect 2590 12220 2596 12232
rect 2551 12192 2596 12220
rect 2590 12180 2596 12192
rect 2648 12180 2654 12232
rect 3605 12223 3663 12229
rect 3605 12189 3617 12223
rect 3651 12220 3663 12223
rect 4430 12220 4436 12232
rect 3651 12192 4436 12220
rect 3651 12189 3663 12192
rect 3605 12183 3663 12189
rect 4430 12180 4436 12192
rect 4488 12180 4494 12232
rect 4706 12220 4712 12232
rect 4667 12192 4712 12220
rect 4706 12180 4712 12192
rect 4764 12180 4770 12232
rect 4798 12180 4804 12232
rect 4856 12180 4862 12232
rect 8202 12180 8208 12232
rect 8260 12180 8266 12232
rect 8662 12180 8668 12232
rect 8720 12220 8726 12232
rect 8849 12223 8907 12229
rect 8849 12220 8861 12223
rect 8720 12192 8861 12220
rect 8720 12180 8726 12192
rect 8849 12189 8861 12192
rect 8895 12189 8907 12223
rect 9030 12220 9036 12232
rect 8991 12192 9036 12220
rect 8849 12183 8907 12189
rect 9030 12180 9036 12192
rect 9088 12180 9094 12232
rect 8220 12152 8248 12180
rect 6012 12124 6592 12152
rect 1486 12044 1492 12096
rect 1544 12084 1550 12096
rect 1673 12087 1731 12093
rect 1673 12084 1685 12087
rect 1544 12056 1685 12084
rect 1544 12044 1550 12056
rect 1673 12053 1685 12056
rect 1719 12053 1731 12087
rect 1673 12047 1731 12053
rect 3789 12087 3847 12093
rect 3789 12053 3801 12087
rect 3835 12084 3847 12087
rect 6012 12084 6040 12124
rect 3835 12056 6040 12084
rect 3835 12053 3847 12056
rect 3789 12047 3847 12053
rect 6362 12044 6368 12096
rect 6420 12084 6426 12096
rect 6457 12087 6515 12093
rect 6457 12084 6469 12087
rect 6420 12056 6469 12084
rect 6420 12044 6426 12056
rect 6457 12053 6469 12056
rect 6503 12053 6515 12087
rect 6564 12084 6592 12124
rect 7944 12124 8248 12152
rect 9508 12152 9536 12260
rect 9950 12248 9956 12300
rect 10008 12288 10014 12300
rect 10137 12291 10195 12297
rect 10137 12288 10149 12291
rect 10008 12260 10149 12288
rect 10008 12248 10014 12260
rect 10137 12257 10149 12260
rect 10183 12257 10195 12291
rect 10137 12251 10195 12257
rect 10594 12248 10600 12300
rect 10652 12248 10658 12300
rect 10686 12248 10692 12300
rect 10744 12288 10750 12300
rect 11057 12291 11115 12297
rect 11057 12288 11069 12291
rect 10744 12260 11069 12288
rect 10744 12248 10750 12260
rect 11057 12257 11069 12260
rect 11103 12257 11115 12291
rect 11057 12251 11115 12257
rect 11238 12248 11244 12300
rect 11296 12288 11302 12300
rect 12161 12291 12219 12297
rect 12161 12288 12173 12291
rect 11296 12260 12173 12288
rect 11296 12248 11302 12260
rect 12161 12257 12173 12260
rect 12207 12257 12219 12291
rect 13081 12291 13139 12297
rect 13081 12288 13093 12291
rect 12161 12251 12219 12257
rect 12268 12260 13093 12288
rect 10321 12223 10379 12229
rect 10321 12189 10333 12223
rect 10367 12220 10379 12223
rect 10502 12220 10508 12232
rect 10367 12192 10508 12220
rect 10367 12189 10379 12192
rect 10321 12183 10379 12189
rect 10502 12180 10508 12192
rect 10560 12180 10566 12232
rect 10870 12220 10876 12232
rect 10612 12192 10876 12220
rect 10612 12152 10640 12192
rect 10870 12180 10876 12192
rect 10928 12180 10934 12232
rect 10962 12180 10968 12232
rect 11020 12220 11026 12232
rect 11149 12223 11207 12229
rect 11149 12220 11161 12223
rect 11020 12192 11161 12220
rect 11020 12180 11026 12192
rect 11149 12189 11161 12192
rect 11195 12189 11207 12223
rect 11330 12220 11336 12232
rect 11291 12192 11336 12220
rect 11149 12183 11207 12189
rect 11330 12180 11336 12192
rect 11388 12180 11394 12232
rect 11609 12223 11667 12229
rect 11609 12189 11621 12223
rect 11655 12220 11667 12223
rect 12268 12220 12296 12260
rect 13081 12257 13093 12260
rect 13127 12257 13139 12291
rect 13081 12251 13139 12257
rect 13170 12248 13176 12300
rect 13228 12288 13234 12300
rect 13906 12288 13912 12300
rect 13228 12260 13912 12288
rect 13228 12248 13234 12260
rect 13906 12248 13912 12260
rect 13964 12248 13970 12300
rect 14093 12291 14151 12297
rect 14093 12257 14105 12291
rect 14139 12257 14151 12291
rect 14093 12251 14151 12257
rect 11655 12192 12296 12220
rect 11655 12189 11667 12192
rect 11609 12183 11667 12189
rect 12342 12180 12348 12232
rect 12400 12220 12406 12232
rect 12400 12192 12445 12220
rect 12400 12180 12406 12192
rect 12894 12180 12900 12232
rect 12952 12220 12958 12232
rect 13265 12223 13323 12229
rect 13265 12220 13277 12223
rect 12952 12192 13277 12220
rect 12952 12180 12958 12192
rect 13265 12189 13277 12192
rect 13311 12220 13323 12223
rect 13722 12220 13728 12232
rect 13311 12192 13728 12220
rect 13311 12189 13323 12192
rect 13265 12183 13323 12189
rect 13722 12180 13728 12192
rect 13780 12180 13786 12232
rect 9508 12124 10640 12152
rect 10689 12155 10747 12161
rect 7944 12084 7972 12124
rect 10689 12121 10701 12155
rect 10735 12152 10747 12155
rect 13078 12152 13084 12164
rect 10735 12124 13084 12152
rect 10735 12121 10747 12124
rect 10689 12115 10747 12121
rect 13078 12112 13084 12124
rect 13136 12112 13142 12164
rect 8110 12084 8116 12096
rect 6564 12056 7972 12084
rect 8071 12056 8116 12084
rect 6457 12047 6515 12053
rect 8110 12044 8116 12056
rect 8168 12044 8174 12096
rect 8202 12044 8208 12096
rect 8260 12084 8266 12096
rect 8389 12087 8447 12093
rect 8389 12084 8401 12087
rect 8260 12056 8401 12084
rect 8260 12044 8266 12056
rect 8389 12053 8401 12056
rect 8435 12053 8447 12087
rect 8389 12047 8447 12053
rect 8846 12044 8852 12096
rect 8904 12084 8910 12096
rect 10962 12084 10968 12096
rect 8904 12056 10968 12084
rect 8904 12044 8910 12056
rect 10962 12044 10968 12056
rect 11020 12044 11026 12096
rect 11054 12044 11060 12096
rect 11112 12084 11118 12096
rect 11609 12087 11667 12093
rect 11609 12084 11621 12087
rect 11112 12056 11621 12084
rect 11112 12044 11118 12056
rect 11609 12053 11621 12056
rect 11655 12053 11667 12087
rect 11609 12047 11667 12053
rect 11701 12087 11759 12093
rect 11701 12053 11713 12087
rect 11747 12084 11759 12087
rect 12526 12084 12532 12096
rect 11747 12056 12532 12084
rect 11747 12053 11759 12056
rect 11701 12047 11759 12053
rect 12526 12044 12532 12056
rect 12584 12044 12590 12096
rect 12710 12084 12716 12096
rect 12671 12056 12716 12084
rect 12710 12044 12716 12056
rect 12768 12044 12774 12096
rect 12894 12044 12900 12096
rect 12952 12084 12958 12096
rect 14108 12084 14136 12251
rect 14200 12220 14228 12328
rect 14277 12223 14335 12229
rect 14277 12220 14289 12223
rect 14200 12192 14289 12220
rect 14277 12189 14289 12192
rect 14323 12189 14335 12223
rect 14277 12183 14335 12189
rect 14737 12223 14795 12229
rect 14737 12189 14749 12223
rect 14783 12189 14795 12223
rect 14737 12183 14795 12189
rect 14752 12096 14780 12183
rect 12952 12056 14136 12084
rect 12952 12044 12958 12056
rect 14734 12044 14740 12096
rect 14792 12044 14798 12096
rect 1104 11994 15824 12016
rect 1104 11942 3447 11994
rect 3499 11942 3511 11994
rect 3563 11942 3575 11994
rect 3627 11942 3639 11994
rect 3691 11942 8378 11994
rect 8430 11942 8442 11994
rect 8494 11942 8506 11994
rect 8558 11942 8570 11994
rect 8622 11942 13308 11994
rect 13360 11942 13372 11994
rect 13424 11942 13436 11994
rect 13488 11942 13500 11994
rect 13552 11942 15824 11994
rect 1104 11920 15824 11942
rect 2041 11883 2099 11889
rect 2041 11849 2053 11883
rect 2087 11880 2099 11883
rect 4522 11880 4528 11892
rect 2087 11852 4528 11880
rect 2087 11849 2099 11852
rect 2041 11843 2099 11849
rect 4522 11840 4528 11852
rect 4580 11840 4586 11892
rect 8202 11880 8208 11892
rect 4632 11852 8208 11880
rect 4430 11812 4436 11824
rect 2700 11784 4436 11812
rect 2700 11753 2728 11784
rect 4430 11772 4436 11784
rect 4488 11772 4494 11824
rect 4632 11812 4660 11852
rect 8202 11840 8208 11852
rect 8260 11840 8266 11892
rect 9490 11840 9496 11892
rect 9548 11880 9554 11892
rect 9861 11883 9919 11889
rect 9861 11880 9873 11883
rect 9548 11852 9873 11880
rect 9548 11840 9554 11852
rect 9861 11849 9873 11852
rect 9907 11849 9919 11883
rect 9861 11843 9919 11849
rect 10502 11840 10508 11892
rect 10560 11880 10566 11892
rect 11517 11883 11575 11889
rect 10560 11852 11100 11880
rect 10560 11840 10566 11852
rect 6457 11815 6515 11821
rect 6457 11812 6469 11815
rect 4540 11784 4660 11812
rect 6196 11784 6469 11812
rect 4540 11753 4568 11784
rect 2685 11747 2743 11753
rect 2685 11713 2697 11747
rect 2731 11713 2743 11747
rect 2685 11707 2743 11713
rect 3697 11747 3755 11753
rect 3697 11713 3709 11747
rect 3743 11744 3755 11747
rect 4525 11747 4583 11753
rect 3743 11716 4476 11744
rect 3743 11713 3755 11716
rect 3697 11707 3755 11713
rect 1949 11679 2007 11685
rect 1949 11645 1961 11679
rect 1995 11676 2007 11679
rect 3878 11676 3884 11688
rect 1995 11648 3884 11676
rect 1995 11645 2007 11648
rect 1949 11639 2007 11645
rect 3878 11636 3884 11648
rect 3936 11636 3942 11688
rect 4062 11636 4068 11688
rect 4120 11636 4126 11688
rect 4448 11676 4476 11716
rect 4525 11713 4537 11747
rect 4571 11713 4583 11747
rect 4525 11707 4583 11713
rect 4709 11747 4767 11753
rect 4709 11713 4721 11747
rect 4755 11744 4767 11747
rect 4798 11744 4804 11756
rect 4755 11716 4804 11744
rect 4755 11713 4767 11716
rect 4709 11707 4767 11713
rect 4798 11704 4804 11716
rect 4856 11704 4862 11756
rect 4890 11676 4896 11688
rect 4448 11648 4896 11676
rect 4890 11636 4896 11648
rect 4948 11636 4954 11688
rect 5074 11676 5080 11688
rect 5035 11648 5080 11676
rect 5074 11636 5080 11648
rect 5132 11636 5138 11688
rect 5276 11648 5580 11676
rect 2406 11608 2412 11620
rect 2367 11580 2412 11608
rect 2406 11568 2412 11580
rect 2464 11568 2470 11620
rect 3418 11608 3424 11620
rect 3379 11580 3424 11608
rect 3418 11568 3424 11580
rect 3476 11568 3482 11620
rect 4080 11608 4108 11636
rect 3528 11580 4108 11608
rect 4433 11611 4491 11617
rect 3528 11552 3556 11580
rect 4433 11577 4445 11611
rect 4479 11608 4491 11611
rect 5276 11608 5304 11648
rect 5350 11617 5356 11620
rect 4479 11580 5304 11608
rect 4479 11577 4491 11580
rect 4433 11571 4491 11577
rect 5344 11571 5356 11617
rect 5408 11608 5414 11620
rect 5552 11608 5580 11648
rect 5626 11636 5632 11688
rect 5684 11676 5690 11688
rect 6196 11676 6224 11784
rect 6457 11781 6469 11784
rect 6503 11781 6515 11815
rect 11072 11812 11100 11852
rect 11517 11849 11529 11883
rect 11563 11880 11575 11883
rect 11563 11852 13584 11880
rect 11563 11849 11575 11852
rect 11517 11843 11575 11849
rect 13556 11824 13584 11852
rect 13814 11840 13820 11892
rect 13872 11880 13878 11892
rect 14461 11883 14519 11889
rect 14461 11880 14473 11883
rect 13872 11852 14473 11880
rect 13872 11840 13878 11852
rect 14461 11849 14473 11852
rect 14507 11849 14519 11883
rect 14461 11843 14519 11849
rect 11974 11812 11980 11824
rect 11072 11784 11980 11812
rect 6457 11775 6515 11781
rect 11974 11772 11980 11784
rect 12032 11772 12038 11824
rect 12434 11772 12440 11824
rect 12492 11812 12498 11824
rect 13354 11812 13360 11824
rect 12492 11784 13360 11812
rect 12492 11772 12498 11784
rect 13354 11772 13360 11784
rect 13412 11772 13418 11824
rect 13538 11772 13544 11824
rect 13596 11772 13602 11824
rect 16298 11812 16304 11824
rect 14292 11784 16304 11812
rect 6822 11744 6828 11756
rect 6783 11716 6828 11744
rect 6822 11704 6828 11716
rect 6880 11704 6886 11756
rect 8297 11747 8355 11753
rect 8297 11713 8309 11747
rect 8343 11744 8355 11747
rect 8343 11716 8616 11744
rect 8343 11713 8355 11716
rect 8297 11707 8355 11713
rect 8481 11679 8539 11685
rect 5684 11648 6224 11676
rect 6288 11648 8432 11676
rect 5684 11636 5690 11648
rect 6288 11608 6316 11648
rect 7070 11611 7128 11617
rect 7070 11608 7082 11611
rect 5408 11580 5444 11608
rect 5552 11580 6316 11608
rect 6380 11580 7082 11608
rect 5350 11568 5356 11571
rect 5408 11568 5414 11580
rect 1670 11500 1676 11552
rect 1728 11540 1734 11552
rect 1765 11543 1823 11549
rect 1765 11540 1777 11543
rect 1728 11512 1777 11540
rect 1728 11500 1734 11512
rect 1765 11509 1777 11512
rect 1811 11509 1823 11543
rect 2498 11540 2504 11552
rect 2459 11512 2504 11540
rect 1765 11503 1823 11509
rect 2498 11500 2504 11512
rect 2556 11500 2562 11552
rect 3050 11540 3056 11552
rect 3011 11512 3056 11540
rect 3050 11500 3056 11512
rect 3108 11500 3114 11552
rect 3510 11540 3516 11552
rect 3471 11512 3516 11540
rect 3510 11500 3516 11512
rect 3568 11500 3574 11552
rect 4062 11540 4068 11552
rect 4023 11512 4068 11540
rect 4062 11500 4068 11512
rect 4120 11500 4126 11552
rect 4706 11500 4712 11552
rect 4764 11540 4770 11552
rect 6380 11540 6408 11580
rect 7070 11577 7082 11580
rect 7116 11608 7128 11611
rect 7374 11608 7380 11620
rect 7116 11580 7380 11608
rect 7116 11577 7128 11580
rect 7070 11571 7128 11577
rect 7374 11568 7380 11580
rect 7432 11568 7438 11620
rect 8297 11611 8355 11617
rect 8297 11608 8309 11611
rect 7484 11580 8309 11608
rect 4764 11512 6408 11540
rect 4764 11500 4770 11512
rect 6638 11500 6644 11552
rect 6696 11540 6702 11552
rect 7484 11540 7512 11580
rect 8297 11577 8309 11580
rect 8343 11577 8355 11611
rect 8297 11571 8355 11577
rect 6696 11512 7512 11540
rect 6696 11500 6702 11512
rect 7558 11500 7564 11552
rect 7616 11540 7622 11552
rect 8205 11543 8263 11549
rect 8205 11540 8217 11543
rect 7616 11512 8217 11540
rect 7616 11500 7622 11512
rect 8205 11509 8217 11512
rect 8251 11509 8263 11543
rect 8404 11540 8432 11648
rect 8481 11645 8493 11679
rect 8527 11645 8539 11679
rect 8588 11676 8616 11716
rect 11330 11704 11336 11756
rect 11388 11744 11394 11756
rect 12250 11744 12256 11756
rect 11388 11716 12256 11744
rect 11388 11704 11394 11716
rect 12250 11704 12256 11716
rect 12308 11704 12314 11756
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 12360 11716 13001 11744
rect 12360 11688 12388 11716
rect 12989 11713 13001 11716
rect 13035 11713 13047 11747
rect 12989 11707 13047 11713
rect 13722 11704 13728 11756
rect 13780 11744 13786 11756
rect 14001 11747 14059 11753
rect 14001 11744 14013 11747
rect 13780 11716 14013 11744
rect 13780 11704 13786 11716
rect 14001 11713 14013 11716
rect 14047 11713 14059 11747
rect 14001 11707 14059 11713
rect 8737 11679 8795 11685
rect 8737 11676 8749 11679
rect 8588 11648 8749 11676
rect 8481 11639 8539 11645
rect 8737 11645 8749 11648
rect 8783 11645 8795 11679
rect 8737 11639 8795 11645
rect 10137 11679 10195 11685
rect 10137 11645 10149 11679
rect 10183 11676 10195 11679
rect 10226 11676 10232 11688
rect 10183 11648 10232 11676
rect 10183 11645 10195 11648
rect 10137 11639 10195 11645
rect 8496 11608 8524 11639
rect 10226 11636 10232 11648
rect 10284 11636 10290 11688
rect 12342 11676 12348 11688
rect 10336 11648 12348 11676
rect 9490 11608 9496 11620
rect 8496 11580 9496 11608
rect 9490 11568 9496 11580
rect 9548 11568 9554 11620
rect 9766 11568 9772 11620
rect 9824 11608 9830 11620
rect 10336 11608 10364 11648
rect 12342 11636 12348 11648
rect 12400 11636 12406 11688
rect 12618 11636 12624 11688
rect 12676 11676 12682 11688
rect 13817 11679 13875 11685
rect 13817 11676 13829 11679
rect 12676 11648 13829 11676
rect 12676 11636 12682 11648
rect 13817 11645 13829 11648
rect 13863 11645 13875 11679
rect 13817 11639 13875 11645
rect 13909 11679 13967 11685
rect 13909 11645 13921 11679
rect 13955 11676 13967 11679
rect 14292 11676 14320 11784
rect 15013 11747 15071 11753
rect 15013 11744 15025 11747
rect 13955 11648 14320 11676
rect 14384 11716 15025 11744
rect 13955 11645 13967 11648
rect 13909 11639 13967 11645
rect 10410 11617 10416 11620
rect 9824 11580 10364 11608
rect 9824 11568 9830 11580
rect 10404 11571 10416 11617
rect 10468 11608 10474 11620
rect 10468 11580 10504 11608
rect 10410 11568 10416 11571
rect 10468 11568 10474 11580
rect 11054 11568 11060 11620
rect 11112 11608 11118 11620
rect 12805 11611 12863 11617
rect 12805 11608 12817 11611
rect 11112 11580 12817 11608
rect 11112 11568 11118 11580
rect 12805 11577 12817 11580
rect 12851 11577 12863 11611
rect 14384 11608 14412 11716
rect 15013 11713 15025 11716
rect 15059 11744 15071 11747
rect 15286 11744 15292 11756
rect 15059 11716 15292 11744
rect 15059 11713 15071 11716
rect 15013 11707 15071 11713
rect 15286 11704 15292 11716
rect 15344 11704 15350 11756
rect 14826 11636 14832 11688
rect 14884 11676 14890 11688
rect 14921 11679 14979 11685
rect 14921 11676 14933 11679
rect 14884 11648 14933 11676
rect 14884 11636 14890 11648
rect 14921 11645 14933 11648
rect 14967 11645 14979 11679
rect 14921 11639 14979 11645
rect 12805 11571 12863 11577
rect 13832 11580 14412 11608
rect 14936 11608 14964 11639
rect 15010 11608 15016 11620
rect 14936 11580 15016 11608
rect 13832 11552 13860 11580
rect 15010 11568 15016 11580
rect 15068 11568 15074 11620
rect 15286 11568 15292 11620
rect 15344 11608 15350 11620
rect 15396 11608 15424 11784
rect 16298 11772 16304 11784
rect 16356 11772 16362 11824
rect 15344 11580 15424 11608
rect 15344 11568 15350 11580
rect 10686 11540 10692 11552
rect 8404 11512 10692 11540
rect 8205 11503 8263 11509
rect 10686 11500 10692 11512
rect 10744 11500 10750 11552
rect 11790 11540 11796 11552
rect 11751 11512 11796 11540
rect 11790 11500 11796 11512
rect 11848 11500 11854 11552
rect 12437 11543 12495 11549
rect 12437 11509 12449 11543
rect 12483 11540 12495 11543
rect 12618 11540 12624 11552
rect 12483 11512 12624 11540
rect 12483 11509 12495 11512
rect 12437 11503 12495 11509
rect 12618 11500 12624 11512
rect 12676 11500 12682 11552
rect 12894 11540 12900 11552
rect 12855 11512 12900 11540
rect 12894 11500 12900 11512
rect 12952 11500 12958 11552
rect 13446 11540 13452 11552
rect 13407 11512 13452 11540
rect 13446 11500 13452 11512
rect 13504 11500 13510 11552
rect 13814 11500 13820 11552
rect 13872 11500 13878 11552
rect 14090 11500 14096 11552
rect 14148 11540 14154 11552
rect 14829 11543 14887 11549
rect 14829 11540 14841 11543
rect 14148 11512 14841 11540
rect 14148 11500 14154 11512
rect 14829 11509 14841 11512
rect 14875 11509 14887 11543
rect 14829 11503 14887 11509
rect 1104 11450 15824 11472
rect 1104 11398 5912 11450
rect 5964 11398 5976 11450
rect 6028 11398 6040 11450
rect 6092 11398 6104 11450
rect 6156 11398 10843 11450
rect 10895 11398 10907 11450
rect 10959 11398 10971 11450
rect 11023 11398 11035 11450
rect 11087 11398 15824 11450
rect 1104 11376 15824 11398
rect 1949 11339 2007 11345
rect 1949 11305 1961 11339
rect 1995 11336 2007 11339
rect 2038 11336 2044 11348
rect 1995 11308 2044 11336
rect 1995 11305 2007 11308
rect 1949 11299 2007 11305
rect 2038 11296 2044 11308
rect 2096 11296 2102 11348
rect 2317 11339 2375 11345
rect 2317 11305 2329 11339
rect 2363 11336 2375 11339
rect 3050 11336 3056 11348
rect 2363 11308 3056 11336
rect 2363 11305 2375 11308
rect 2317 11299 2375 11305
rect 3050 11296 3056 11308
rect 3108 11296 3114 11348
rect 3329 11339 3387 11345
rect 3329 11305 3341 11339
rect 3375 11336 3387 11339
rect 4062 11336 4068 11348
rect 3375 11308 4068 11336
rect 3375 11305 3387 11308
rect 3329 11299 3387 11305
rect 4062 11296 4068 11308
rect 4120 11296 4126 11348
rect 5350 11296 5356 11348
rect 5408 11336 5414 11348
rect 5721 11339 5779 11345
rect 5721 11336 5733 11339
rect 5408 11308 5733 11336
rect 5408 11296 5414 11308
rect 5721 11305 5733 11308
rect 5767 11305 5779 11339
rect 6362 11336 6368 11348
rect 5721 11299 5779 11305
rect 5828 11308 6368 11336
rect 3421 11271 3479 11277
rect 3421 11237 3433 11271
rect 3467 11268 3479 11271
rect 4246 11268 4252 11280
rect 3467 11240 4252 11268
rect 3467 11237 3479 11240
rect 3421 11231 3479 11237
rect 4246 11228 4252 11240
rect 4304 11228 4310 11280
rect 5828 11268 5856 11308
rect 6362 11296 6368 11308
rect 6420 11296 6426 11348
rect 7374 11336 7380 11348
rect 7335 11308 7380 11336
rect 7374 11296 7380 11308
rect 7432 11296 7438 11348
rect 9033 11339 9091 11345
rect 9033 11305 9045 11339
rect 9079 11336 9091 11339
rect 9122 11336 9128 11348
rect 9079 11308 9128 11336
rect 9079 11305 9091 11308
rect 9033 11299 9091 11305
rect 9122 11296 9128 11308
rect 9180 11296 9186 11348
rect 9309 11339 9367 11345
rect 9309 11305 9321 11339
rect 9355 11305 9367 11339
rect 9309 11299 9367 11305
rect 4356 11240 5856 11268
rect 6264 11271 6322 11277
rect 4154 11200 4160 11212
rect 2700 11172 4160 11200
rect 1489 11135 1547 11141
rect 1489 11101 1501 11135
rect 1535 11101 1547 11135
rect 1489 11095 1547 11101
rect 2409 11135 2467 11141
rect 2409 11101 2421 11135
rect 2455 11101 2467 11135
rect 2409 11095 2467 11101
rect 1504 11064 1532 11095
rect 1857 11067 1915 11073
rect 1857 11064 1869 11067
rect 1504 11036 1869 11064
rect 1857 11033 1869 11036
rect 1903 11064 1915 11067
rect 2038 11064 2044 11076
rect 1903 11036 2044 11064
rect 1903 11033 1915 11036
rect 1857 11027 1915 11033
rect 2038 11024 2044 11036
rect 2096 11024 2102 11076
rect 2424 11064 2452 11095
rect 2498 11092 2504 11144
rect 2556 11132 2562 11144
rect 2556 11104 2601 11132
rect 2556 11092 2562 11104
rect 2700 11064 2728 11172
rect 4154 11160 4160 11172
rect 4212 11160 4218 11212
rect 4356 11200 4384 11240
rect 6264 11237 6276 11271
rect 6310 11268 6322 11271
rect 8110 11268 8116 11280
rect 6310 11240 8116 11268
rect 6310 11237 6322 11240
rect 6264 11231 6322 11237
rect 8110 11228 8116 11240
rect 8168 11228 8174 11280
rect 8846 11228 8852 11280
rect 8904 11268 8910 11280
rect 9324 11268 9352 11299
rect 10410 11296 10416 11348
rect 10468 11336 10474 11348
rect 10594 11336 10600 11348
rect 10468 11308 10600 11336
rect 10468 11296 10474 11308
rect 10594 11296 10600 11308
rect 10652 11296 10658 11348
rect 11333 11339 11391 11345
rect 11333 11305 11345 11339
rect 11379 11336 11391 11339
rect 11514 11336 11520 11348
rect 11379 11308 11520 11336
rect 11379 11305 11391 11308
rect 11333 11299 11391 11305
rect 11514 11296 11520 11308
rect 11572 11296 11578 11348
rect 11882 11296 11888 11348
rect 11940 11336 11946 11348
rect 12345 11339 12403 11345
rect 12345 11336 12357 11339
rect 11940 11308 12357 11336
rect 11940 11296 11946 11308
rect 12345 11305 12357 11308
rect 12391 11305 12403 11339
rect 12345 11299 12403 11305
rect 12618 11296 12624 11348
rect 12676 11336 12682 11348
rect 12805 11339 12863 11345
rect 12805 11336 12817 11339
rect 12676 11308 12817 11336
rect 12676 11296 12682 11308
rect 12805 11305 12817 11308
rect 12851 11305 12863 11339
rect 13354 11336 13360 11348
rect 13315 11308 13360 11336
rect 12805 11299 12863 11305
rect 13354 11296 13360 11308
rect 13412 11296 13418 11348
rect 13725 11339 13783 11345
rect 13725 11305 13737 11339
rect 13771 11336 13783 11339
rect 14734 11336 14740 11348
rect 13771 11308 14740 11336
rect 13771 11305 13783 11308
rect 13725 11299 13783 11305
rect 14734 11296 14740 11308
rect 14792 11296 14798 11348
rect 8904 11240 9352 11268
rect 8904 11228 8910 11240
rect 11146 11228 11152 11280
rect 11204 11268 11210 11280
rect 11701 11271 11759 11277
rect 11701 11268 11713 11271
rect 11204 11240 11713 11268
rect 11204 11228 11210 11240
rect 11701 11237 11713 11240
rect 11747 11268 11759 11271
rect 12434 11268 12440 11280
rect 11747 11240 12440 11268
rect 11747 11237 11759 11240
rect 11701 11231 11759 11237
rect 12434 11228 12440 11240
rect 12492 11228 12498 11280
rect 12526 11228 12532 11280
rect 12584 11268 12590 11280
rect 12713 11271 12771 11277
rect 12713 11268 12725 11271
rect 12584 11240 12725 11268
rect 12584 11228 12590 11240
rect 12713 11237 12725 11240
rect 12759 11237 12771 11271
rect 12713 11231 12771 11237
rect 12986 11228 12992 11280
rect 13044 11268 13050 11280
rect 14369 11271 14427 11277
rect 14369 11268 14381 11271
rect 13044 11240 14381 11268
rect 13044 11228 13050 11240
rect 14369 11237 14381 11240
rect 14415 11237 14427 11271
rect 14369 11231 14427 11237
rect 4264 11172 4384 11200
rect 3234 11092 3240 11144
rect 3292 11132 3298 11144
rect 3605 11135 3663 11141
rect 3605 11132 3617 11135
rect 3292 11104 3617 11132
rect 3292 11092 3298 11104
rect 3605 11101 3617 11104
rect 3651 11132 3663 11135
rect 4264 11132 4292 11172
rect 4430 11160 4436 11212
rect 4488 11200 4494 11212
rect 4608 11203 4666 11209
rect 4608 11200 4620 11203
rect 4488 11172 4620 11200
rect 4488 11160 4494 11172
rect 4608 11169 4620 11172
rect 4654 11200 4666 11203
rect 5997 11203 6055 11209
rect 4654 11172 5396 11200
rect 4654 11169 4666 11172
rect 4608 11163 4666 11169
rect 3651 11104 4292 11132
rect 4341 11135 4399 11141
rect 3651 11101 3663 11104
rect 3605 11095 3663 11101
rect 4341 11101 4353 11135
rect 4387 11101 4399 11135
rect 5368 11132 5396 11172
rect 5997 11169 6009 11203
rect 6043 11200 6055 11203
rect 6822 11200 6828 11212
rect 6043 11172 6828 11200
rect 6043 11169 6055 11172
rect 5997 11163 6055 11169
rect 6822 11160 6828 11172
rect 6880 11160 6886 11212
rect 7374 11160 7380 11212
rect 7432 11200 7438 11212
rect 7909 11203 7967 11209
rect 7909 11200 7921 11203
rect 7432 11172 7921 11200
rect 7432 11160 7438 11172
rect 7909 11169 7921 11172
rect 7955 11169 7967 11203
rect 7909 11163 7967 11169
rect 8202 11160 8208 11212
rect 8260 11200 8266 11212
rect 9950 11209 9956 11212
rect 9493 11203 9551 11209
rect 9493 11200 9505 11203
rect 8260 11172 9505 11200
rect 8260 11160 8266 11172
rect 9493 11169 9505 11172
rect 9539 11169 9551 11203
rect 9944 11200 9956 11209
rect 9911 11172 9956 11200
rect 9493 11163 9551 11169
rect 9944 11163 9956 11172
rect 9950 11160 9956 11163
rect 10008 11160 10014 11212
rect 10226 11160 10232 11212
rect 10284 11200 10290 11212
rect 11330 11200 11336 11212
rect 10284 11172 11336 11200
rect 10284 11160 10290 11172
rect 11330 11160 11336 11172
rect 11388 11160 11394 11212
rect 11793 11203 11851 11209
rect 11793 11169 11805 11203
rect 11839 11200 11851 11203
rect 12161 11203 12219 11209
rect 12161 11200 12173 11203
rect 11839 11172 12173 11200
rect 11839 11169 11851 11172
rect 11793 11163 11851 11169
rect 12161 11169 12173 11172
rect 12207 11169 12219 11203
rect 12161 11163 12219 11169
rect 13817 11203 13875 11209
rect 13817 11169 13829 11203
rect 13863 11200 13875 11203
rect 14182 11200 14188 11212
rect 13863 11172 14188 11200
rect 13863 11169 13875 11172
rect 13817 11163 13875 11169
rect 14182 11160 14188 11172
rect 14240 11160 14246 11212
rect 15013 11203 15071 11209
rect 15013 11169 15025 11203
rect 15059 11169 15071 11203
rect 15013 11163 15071 11169
rect 7650 11132 7656 11144
rect 5368 11104 6040 11132
rect 7611 11104 7656 11132
rect 4341 11095 4399 11101
rect 2958 11064 2964 11076
rect 2424 11036 2728 11064
rect 2919 11036 2964 11064
rect 2958 11024 2964 11036
rect 3016 11024 3022 11076
rect 3050 11024 3056 11076
rect 3108 11064 3114 11076
rect 3510 11064 3516 11076
rect 3108 11036 3516 11064
rect 3108 11024 3114 11036
rect 3510 11024 3516 11036
rect 3568 11024 3574 11076
rect 4154 11024 4160 11076
rect 4212 11064 4218 11076
rect 4356 11064 4384 11095
rect 4212 11036 4384 11064
rect 4212 11024 4218 11036
rect 6012 10996 6040 11104
rect 7650 11092 7656 11104
rect 7708 11092 7714 11144
rect 8846 11092 8852 11144
rect 8904 11132 8910 11144
rect 9214 11132 9220 11144
rect 8904 11104 9220 11132
rect 8904 11092 8910 11104
rect 9214 11092 9220 11104
rect 9272 11092 9278 11144
rect 9677 11135 9735 11141
rect 9677 11101 9689 11135
rect 9723 11101 9735 11135
rect 11882 11132 11888 11144
rect 11843 11104 11888 11132
rect 9677 11095 9735 11101
rect 7006 11064 7012 11076
rect 6932 11036 7012 11064
rect 6932 10996 6960 11036
rect 7006 11024 7012 11036
rect 7064 11024 7070 11076
rect 6012 10968 6960 10996
rect 7558 10956 7564 11008
rect 7616 10996 7622 11008
rect 8846 10996 8852 11008
rect 7616 10968 8852 10996
rect 7616 10956 7622 10968
rect 8846 10956 8852 10968
rect 8904 10956 8910 11008
rect 9490 10956 9496 11008
rect 9548 10996 9554 11008
rect 9692 10996 9720 11095
rect 11882 11092 11888 11104
rect 11940 11092 11946 11144
rect 12986 11132 12992 11144
rect 12899 11104 12992 11132
rect 12986 11092 12992 11104
rect 13044 11132 13050 11144
rect 13173 11135 13231 11141
rect 13173 11132 13185 11135
rect 13044 11104 13185 11132
rect 13044 11092 13050 11104
rect 13173 11101 13185 11104
rect 13219 11101 13231 11135
rect 13173 11095 13231 11101
rect 13354 11092 13360 11144
rect 13412 11132 13418 11144
rect 13909 11135 13967 11141
rect 13909 11132 13921 11135
rect 13412 11104 13921 11132
rect 13412 11092 13418 11104
rect 13909 11101 13921 11104
rect 13955 11101 13967 11135
rect 13909 11095 13967 11101
rect 14366 11092 14372 11144
rect 14424 11132 14430 11144
rect 15028 11132 15056 11163
rect 14424 11104 15056 11132
rect 14424 11092 14430 11104
rect 14829 11067 14887 11073
rect 14829 11064 14841 11067
rect 10612 11036 12848 11064
rect 10612 10996 10640 11036
rect 11054 10996 11060 11008
rect 9548 10968 10640 10996
rect 11015 10968 11060 10996
rect 9548 10956 9554 10968
rect 11054 10956 11060 10968
rect 11112 10956 11118 11008
rect 11238 10956 11244 11008
rect 11296 10996 11302 11008
rect 12158 10996 12164 11008
rect 11296 10968 12164 10996
rect 11296 10956 11302 10968
rect 12158 10956 12164 10968
rect 12216 10956 12222 11008
rect 12253 10999 12311 11005
rect 12253 10965 12265 10999
rect 12299 10996 12311 10999
rect 12710 10996 12716 11008
rect 12299 10968 12716 10996
rect 12299 10965 12311 10968
rect 12253 10959 12311 10965
rect 12710 10956 12716 10968
rect 12768 10956 12774 11008
rect 12820 10996 12848 11036
rect 13004 11036 14841 11064
rect 13004 10996 13032 11036
rect 14829 11033 14841 11036
rect 14875 11033 14887 11067
rect 14829 11027 14887 11033
rect 12820 10968 13032 10996
rect 13173 10999 13231 11005
rect 13173 10965 13185 10999
rect 13219 10996 13231 10999
rect 15470 10996 15476 11008
rect 13219 10968 15476 10996
rect 13219 10965 13231 10968
rect 13173 10959 13231 10965
rect 15470 10956 15476 10968
rect 15528 10956 15534 11008
rect 1104 10906 15824 10928
rect 1104 10854 3447 10906
rect 3499 10854 3511 10906
rect 3563 10854 3575 10906
rect 3627 10854 3639 10906
rect 3691 10854 8378 10906
rect 8430 10854 8442 10906
rect 8494 10854 8506 10906
rect 8558 10854 8570 10906
rect 8622 10854 13308 10906
rect 13360 10854 13372 10906
rect 13424 10854 13436 10906
rect 13488 10854 13500 10906
rect 13552 10854 15824 10906
rect 1104 10832 15824 10854
rect 4614 10752 4620 10804
rect 4672 10792 4678 10804
rect 7466 10792 7472 10804
rect 4672 10764 7472 10792
rect 4672 10752 4678 10764
rect 7466 10752 7472 10764
rect 7524 10792 7530 10804
rect 8110 10792 8116 10804
rect 7524 10764 8116 10792
rect 7524 10752 7530 10764
rect 8110 10752 8116 10764
rect 8168 10752 8174 10804
rect 11054 10792 11060 10804
rect 8772 10764 11060 10792
rect 3326 10724 3332 10736
rect 1872 10696 3332 10724
rect 1872 10665 1900 10696
rect 3326 10684 3332 10696
rect 3384 10684 3390 10736
rect 4798 10724 4804 10736
rect 4759 10696 4804 10724
rect 4798 10684 4804 10696
rect 4856 10684 4862 10736
rect 6457 10727 6515 10733
rect 6457 10693 6469 10727
rect 6503 10724 6515 10727
rect 6546 10724 6552 10736
rect 6503 10696 6552 10724
rect 6503 10693 6515 10696
rect 6457 10687 6515 10693
rect 6546 10684 6552 10696
rect 6604 10684 6610 10736
rect 7834 10684 7840 10736
rect 7892 10724 7898 10736
rect 8389 10727 8447 10733
rect 8389 10724 8401 10727
rect 7892 10696 8401 10724
rect 7892 10684 7898 10696
rect 8389 10693 8401 10696
rect 8435 10693 8447 10727
rect 8389 10687 8447 10693
rect 8478 10684 8484 10736
rect 8536 10724 8542 10736
rect 8536 10696 8581 10724
rect 8536 10684 8542 10696
rect 1857 10659 1915 10665
rect 1857 10625 1869 10659
rect 1903 10625 1915 10659
rect 1857 10619 1915 10625
rect 2041 10659 2099 10665
rect 2041 10625 2053 10659
rect 2087 10625 2099 10659
rect 2041 10619 2099 10625
rect 1765 10591 1823 10597
rect 1765 10557 1777 10591
rect 1811 10588 1823 10591
rect 1946 10588 1952 10600
rect 1811 10560 1952 10588
rect 1811 10557 1823 10560
rect 1765 10551 1823 10557
rect 1946 10548 1952 10560
rect 2004 10548 2010 10600
rect 2056 10520 2084 10619
rect 2774 10616 2780 10668
rect 2832 10656 2838 10668
rect 2869 10659 2927 10665
rect 2869 10656 2881 10659
rect 2832 10628 2881 10656
rect 2832 10616 2838 10628
rect 2869 10625 2881 10628
rect 2915 10625 2927 10659
rect 2869 10619 2927 10625
rect 3053 10659 3111 10665
rect 3053 10625 3065 10659
rect 3099 10656 3111 10659
rect 3237 10659 3295 10665
rect 3237 10656 3249 10659
rect 3099 10628 3249 10656
rect 3099 10625 3111 10628
rect 3053 10619 3111 10625
rect 3237 10625 3249 10628
rect 3283 10625 3295 10659
rect 6822 10656 6828 10668
rect 6783 10628 6828 10656
rect 3237 10619 3295 10625
rect 6822 10616 6828 10628
rect 6880 10616 6886 10668
rect 2314 10548 2320 10600
rect 2372 10588 2378 10600
rect 3421 10591 3479 10597
rect 3421 10588 3433 10591
rect 2372 10560 3433 10588
rect 2372 10548 2378 10560
rect 3421 10557 3433 10560
rect 3467 10588 3479 10591
rect 4154 10588 4160 10600
rect 3467 10560 4160 10588
rect 3467 10557 3479 10560
rect 3421 10551 3479 10557
rect 4154 10548 4160 10560
rect 4212 10588 4218 10600
rect 5074 10588 5080 10600
rect 4212 10560 5080 10588
rect 4212 10548 4218 10560
rect 5074 10548 5080 10560
rect 5132 10548 5138 10600
rect 5344 10591 5402 10597
rect 5344 10557 5356 10591
rect 5390 10588 5402 10591
rect 5626 10588 5632 10600
rect 5390 10560 5632 10588
rect 5390 10557 5402 10560
rect 5344 10551 5402 10557
rect 5626 10548 5632 10560
rect 5684 10548 5690 10600
rect 8772 10588 8800 10764
rect 11054 10752 11060 10764
rect 11112 10752 11118 10804
rect 11698 10752 11704 10804
rect 11756 10792 11762 10804
rect 14277 10795 14335 10801
rect 11756 10764 14044 10792
rect 11756 10752 11762 10764
rect 10686 10684 10692 10736
rect 10744 10724 10750 10736
rect 11149 10727 11207 10733
rect 11149 10724 11161 10727
rect 10744 10696 11161 10724
rect 10744 10684 10750 10696
rect 11149 10693 11161 10696
rect 11195 10693 11207 10727
rect 11149 10687 11207 10693
rect 11974 10684 11980 10736
rect 12032 10724 12038 10736
rect 12437 10727 12495 10733
rect 12437 10724 12449 10727
rect 12032 10696 12449 10724
rect 12032 10684 12038 10696
rect 12437 10693 12449 10696
rect 12483 10693 12495 10727
rect 12437 10687 12495 10693
rect 12894 10684 12900 10736
rect 12952 10724 12958 10736
rect 13449 10727 13507 10733
rect 13449 10724 13461 10727
rect 12952 10696 13461 10724
rect 12952 10684 12958 10696
rect 13449 10693 13461 10696
rect 13495 10693 13507 10727
rect 13449 10687 13507 10693
rect 9030 10656 9036 10668
rect 8991 10628 9036 10656
rect 9030 10616 9036 10628
rect 9088 10656 9094 10668
rect 9309 10659 9367 10665
rect 9309 10656 9321 10659
rect 9088 10628 9321 10656
rect 9088 10616 9094 10628
rect 9309 10625 9321 10628
rect 9355 10625 9367 10659
rect 9490 10656 9496 10668
rect 9451 10628 9496 10656
rect 9309 10619 9367 10625
rect 9490 10616 9496 10628
rect 9548 10616 9554 10668
rect 10594 10616 10600 10668
rect 10652 10656 10658 10668
rect 11701 10659 11759 10665
rect 11701 10656 11713 10659
rect 10652 10628 11713 10656
rect 10652 10616 10658 10628
rect 11701 10625 11713 10628
rect 11747 10625 11759 10659
rect 11701 10619 11759 10625
rect 11882 10616 11888 10668
rect 11940 10656 11946 10668
rect 12989 10659 13047 10665
rect 12989 10656 13001 10659
rect 11940 10628 13001 10656
rect 11940 10616 11946 10628
rect 12989 10625 13001 10628
rect 13035 10625 13047 10659
rect 12989 10619 13047 10625
rect 13354 10616 13360 10668
rect 13412 10656 13418 10668
rect 14016 10665 14044 10764
rect 14277 10761 14289 10795
rect 14323 10792 14335 10795
rect 14458 10792 14464 10804
rect 14323 10764 14464 10792
rect 14323 10761 14335 10764
rect 14277 10755 14335 10761
rect 14458 10752 14464 10764
rect 14516 10752 14522 10804
rect 14734 10752 14740 10804
rect 14792 10792 14798 10804
rect 15010 10792 15016 10804
rect 14792 10764 15016 10792
rect 14792 10752 14798 10764
rect 15010 10752 15016 10764
rect 15068 10752 15074 10804
rect 13909 10659 13967 10665
rect 13909 10656 13921 10659
rect 13412 10628 13921 10656
rect 13412 10616 13418 10628
rect 13909 10625 13921 10628
rect 13955 10625 13967 10659
rect 13909 10619 13967 10625
rect 14001 10659 14059 10665
rect 14001 10625 14013 10659
rect 14047 10625 14059 10659
rect 15010 10656 15016 10668
rect 14971 10628 15016 10656
rect 14001 10619 14059 10625
rect 15010 10616 15016 10628
rect 15068 10616 15074 10668
rect 11238 10588 11244 10600
rect 6932 10560 8800 10588
rect 9661 10560 11244 10588
rect 3688 10523 3746 10529
rect 3688 10520 3700 10523
rect 2056 10492 3700 10520
rect 3688 10489 3700 10492
rect 3734 10520 3746 10523
rect 6932 10520 6960 10560
rect 7098 10529 7104 10532
rect 7092 10520 7104 10529
rect 3734 10492 6960 10520
rect 7011 10492 7104 10520
rect 3734 10489 3746 10492
rect 3688 10483 3746 10489
rect 7092 10483 7104 10492
rect 7156 10520 7162 10532
rect 7834 10520 7840 10532
rect 7156 10492 7840 10520
rect 7098 10480 7104 10483
rect 7156 10480 7162 10492
rect 7834 10480 7840 10492
rect 7892 10480 7898 10532
rect 8110 10480 8116 10532
rect 8168 10520 8174 10532
rect 9661 10520 9689 10560
rect 11238 10548 11244 10560
rect 11296 10548 11302 10600
rect 11517 10591 11575 10597
rect 11517 10557 11529 10591
rect 11563 10588 11575 10591
rect 11790 10588 11796 10600
rect 11563 10560 11796 10588
rect 11563 10557 11575 10560
rect 11517 10551 11575 10557
rect 11790 10548 11796 10560
rect 11848 10548 11854 10600
rect 12805 10591 12863 10597
rect 12805 10557 12817 10591
rect 12851 10588 12863 10591
rect 15102 10588 15108 10600
rect 12851 10560 15108 10588
rect 12851 10557 12863 10560
rect 12805 10551 12863 10557
rect 15102 10548 15108 10560
rect 15160 10548 15166 10600
rect 9766 10529 9772 10532
rect 9760 10520 9772 10529
rect 8168 10492 9689 10520
rect 9727 10492 9772 10520
rect 8168 10480 8174 10492
rect 9760 10483 9772 10492
rect 9766 10480 9772 10483
rect 9824 10480 9830 10532
rect 12986 10520 12992 10532
rect 10888 10492 12992 10520
rect 1397 10455 1455 10461
rect 1397 10421 1409 10455
rect 1443 10452 1455 10455
rect 2130 10452 2136 10464
rect 1443 10424 2136 10452
rect 1443 10421 1455 10424
rect 1397 10415 1455 10421
rect 2130 10412 2136 10424
rect 2188 10412 2194 10464
rect 2406 10452 2412 10464
rect 2367 10424 2412 10452
rect 2406 10412 2412 10424
rect 2464 10412 2470 10464
rect 2777 10455 2835 10461
rect 2777 10421 2789 10455
rect 2823 10452 2835 10455
rect 3050 10452 3056 10464
rect 2823 10424 3056 10452
rect 2823 10421 2835 10424
rect 2777 10415 2835 10421
rect 3050 10412 3056 10424
rect 3108 10412 3114 10464
rect 3237 10455 3295 10461
rect 3237 10421 3249 10455
rect 3283 10452 3295 10455
rect 4614 10452 4620 10464
rect 3283 10424 4620 10452
rect 3283 10421 3295 10424
rect 3237 10415 3295 10421
rect 4614 10412 4620 10424
rect 4672 10412 4678 10464
rect 6822 10412 6828 10464
rect 6880 10452 6886 10464
rect 8205 10455 8263 10461
rect 8205 10452 8217 10455
rect 6880 10424 8217 10452
rect 6880 10412 6886 10424
rect 8205 10421 8217 10424
rect 8251 10421 8263 10455
rect 8205 10415 8263 10421
rect 8389 10455 8447 10461
rect 8389 10421 8401 10455
rect 8435 10452 8447 10455
rect 8849 10455 8907 10461
rect 8849 10452 8861 10455
rect 8435 10424 8861 10452
rect 8435 10421 8447 10424
rect 8389 10415 8447 10421
rect 8849 10421 8861 10424
rect 8895 10421 8907 10455
rect 8849 10415 8907 10421
rect 8938 10412 8944 10464
rect 8996 10452 9002 10464
rect 9309 10455 9367 10461
rect 8996 10424 9041 10452
rect 8996 10412 9002 10424
rect 9309 10421 9321 10455
rect 9355 10452 9367 10455
rect 10594 10452 10600 10464
rect 9355 10424 10600 10452
rect 9355 10421 9367 10424
rect 9309 10415 9367 10421
rect 10594 10412 10600 10424
rect 10652 10412 10658 10464
rect 10888 10461 10916 10492
rect 12986 10480 12992 10492
rect 13044 10480 13050 10532
rect 13814 10520 13820 10532
rect 13775 10492 13820 10520
rect 13814 10480 13820 10492
rect 13872 10480 13878 10532
rect 14366 10480 14372 10532
rect 14424 10520 14430 10532
rect 14642 10520 14648 10532
rect 14424 10492 14648 10520
rect 14424 10480 14430 10492
rect 14642 10480 14648 10492
rect 14700 10520 14706 10532
rect 14921 10523 14979 10529
rect 14921 10520 14933 10523
rect 14700 10492 14933 10520
rect 14700 10480 14706 10492
rect 14921 10489 14933 10492
rect 14967 10489 14979 10523
rect 14921 10483 14979 10489
rect 10873 10455 10931 10461
rect 10873 10421 10885 10455
rect 10919 10421 10931 10455
rect 10873 10415 10931 10421
rect 11609 10455 11667 10461
rect 11609 10421 11621 10455
rect 11655 10452 11667 10455
rect 11698 10452 11704 10464
rect 11655 10424 11704 10452
rect 11655 10421 11667 10424
rect 11609 10415 11667 10421
rect 11698 10412 11704 10424
rect 11756 10412 11762 10464
rect 12618 10412 12624 10464
rect 12676 10452 12682 10464
rect 12802 10452 12808 10464
rect 12676 10424 12808 10452
rect 12676 10412 12682 10424
rect 12802 10412 12808 10424
rect 12860 10412 12866 10464
rect 12897 10455 12955 10461
rect 12897 10421 12909 10455
rect 12943 10452 12955 10455
rect 13078 10452 13084 10464
rect 12943 10424 13084 10452
rect 12943 10421 12955 10424
rect 12897 10415 12955 10421
rect 13078 10412 13084 10424
rect 13136 10452 13142 10464
rect 14277 10455 14335 10461
rect 14277 10452 14289 10455
rect 13136 10424 14289 10452
rect 13136 10412 13142 10424
rect 14277 10421 14289 10424
rect 14323 10421 14335 10455
rect 14458 10452 14464 10464
rect 14419 10424 14464 10452
rect 14277 10415 14335 10421
rect 14458 10412 14464 10424
rect 14516 10412 14522 10464
rect 14829 10455 14887 10461
rect 14829 10421 14841 10455
rect 14875 10452 14887 10455
rect 15378 10452 15384 10464
rect 14875 10424 15384 10452
rect 14875 10421 14887 10424
rect 14829 10415 14887 10421
rect 15378 10412 15384 10424
rect 15436 10452 15442 10464
rect 15930 10452 15936 10464
rect 15436 10424 15936 10452
rect 15436 10412 15442 10424
rect 15930 10412 15936 10424
rect 15988 10412 15994 10464
rect 1104 10362 15824 10384
rect 1104 10310 5912 10362
rect 5964 10310 5976 10362
rect 6028 10310 6040 10362
rect 6092 10310 6104 10362
rect 6156 10310 10843 10362
rect 10895 10310 10907 10362
rect 10959 10310 10971 10362
rect 11023 10310 11035 10362
rect 11087 10310 15824 10362
rect 1104 10288 15824 10310
rect 5534 10248 5540 10260
rect 5447 10220 5540 10248
rect 5534 10208 5540 10220
rect 5592 10248 5598 10260
rect 6638 10248 6644 10260
rect 5592 10220 6644 10248
rect 5592 10208 5598 10220
rect 6638 10208 6644 10220
rect 6696 10208 6702 10260
rect 7469 10251 7527 10257
rect 7469 10217 7481 10251
rect 7515 10248 7527 10251
rect 9309 10251 9367 10257
rect 7515 10220 9260 10248
rect 7515 10217 7527 10220
rect 7469 10211 7527 10217
rect 1854 10180 1860 10192
rect 1815 10152 1860 10180
rect 1854 10140 1860 10152
rect 1912 10140 1918 10192
rect 2584 10183 2642 10189
rect 2584 10149 2596 10183
rect 2630 10180 2642 10183
rect 3234 10180 3240 10192
rect 2630 10152 3240 10180
rect 2630 10149 2642 10152
rect 2584 10143 2642 10149
rect 3234 10140 3240 10152
rect 3292 10140 3298 10192
rect 4424 10183 4482 10189
rect 4424 10149 4436 10183
rect 4470 10180 4482 10183
rect 6270 10180 6276 10192
rect 4470 10152 6276 10180
rect 4470 10149 4482 10152
rect 4424 10143 4482 10149
rect 6270 10140 6276 10152
rect 6328 10180 6334 10192
rect 6822 10180 6828 10192
rect 6328 10152 6828 10180
rect 6328 10140 6334 10152
rect 6822 10140 6828 10152
rect 6880 10140 6886 10192
rect 8196 10183 8254 10189
rect 8196 10149 8208 10183
rect 8242 10180 8254 10183
rect 9122 10180 9128 10192
rect 8242 10152 9128 10180
rect 8242 10149 8254 10152
rect 8196 10143 8254 10149
rect 9122 10140 9128 10152
rect 9180 10140 9186 10192
rect 9232 10180 9260 10220
rect 9309 10217 9321 10251
rect 9355 10248 9367 10251
rect 9766 10248 9772 10260
rect 9355 10220 9772 10248
rect 9355 10217 9367 10220
rect 9309 10211 9367 10217
rect 9766 10208 9772 10220
rect 9824 10208 9830 10260
rect 9950 10208 9956 10260
rect 10008 10248 10014 10260
rect 12713 10251 12771 10257
rect 12713 10248 12725 10251
rect 10008 10220 12725 10248
rect 10008 10208 10014 10220
rect 12713 10217 12725 10220
rect 12759 10217 12771 10251
rect 12713 10211 12771 10217
rect 12986 10208 12992 10260
rect 13044 10248 13050 10260
rect 13449 10251 13507 10257
rect 13449 10248 13461 10251
rect 13044 10220 13461 10248
rect 13044 10208 13050 10220
rect 13449 10217 13461 10220
rect 13495 10217 13507 10251
rect 13449 10211 13507 10217
rect 13630 10208 13636 10260
rect 13688 10248 13694 10260
rect 14001 10251 14059 10257
rect 14001 10248 14013 10251
rect 13688 10220 14013 10248
rect 13688 10208 13694 10220
rect 14001 10217 14013 10220
rect 14047 10217 14059 10251
rect 14001 10211 14059 10217
rect 10410 10180 10416 10192
rect 9232 10152 10416 10180
rect 10410 10140 10416 10152
rect 10468 10140 10474 10192
rect 11238 10180 11244 10192
rect 10520 10152 11244 10180
rect 1578 10112 1584 10124
rect 1539 10084 1584 10112
rect 1578 10072 1584 10084
rect 1636 10072 1642 10124
rect 4154 10112 4160 10124
rect 4115 10084 4160 10112
rect 4154 10072 4160 10084
rect 4212 10072 4218 10124
rect 6069 10115 6127 10121
rect 6069 10112 6081 10115
rect 4264 10084 6081 10112
rect 1486 10004 1492 10056
rect 1544 10044 1550 10056
rect 2314 10044 2320 10056
rect 1544 10016 2320 10044
rect 1544 10004 1550 10016
rect 2314 10004 2320 10016
rect 2372 10004 2378 10056
rect 3970 10004 3976 10056
rect 4028 10044 4034 10056
rect 4264 10044 4292 10084
rect 6069 10081 6081 10084
rect 6115 10081 6127 10115
rect 6069 10075 6127 10081
rect 7650 10072 7656 10124
rect 7708 10112 7714 10124
rect 7929 10115 7987 10121
rect 7929 10112 7941 10115
rect 7708 10084 7941 10112
rect 7708 10072 7714 10084
rect 7929 10081 7941 10084
rect 7975 10112 7987 10115
rect 9490 10112 9496 10124
rect 7975 10084 9496 10112
rect 7975 10081 7987 10084
rect 7929 10075 7987 10081
rect 9490 10072 9496 10084
rect 9548 10112 9554 10124
rect 9677 10115 9735 10121
rect 9677 10112 9689 10115
rect 9548 10084 9689 10112
rect 9548 10072 9554 10084
rect 9677 10081 9689 10084
rect 9723 10081 9735 10115
rect 9944 10115 10002 10121
rect 9944 10112 9956 10115
rect 9677 10075 9735 10081
rect 9784 10084 9956 10112
rect 4028 10016 4292 10044
rect 4028 10004 4034 10016
rect 5166 10004 5172 10056
rect 5224 10044 5230 10056
rect 5813 10047 5871 10053
rect 5813 10044 5825 10047
rect 5224 10016 5825 10044
rect 5224 10004 5230 10016
rect 5813 10013 5825 10016
rect 5859 10013 5871 10047
rect 5813 10007 5871 10013
rect 9214 10004 9220 10056
rect 9272 10044 9278 10056
rect 9784 10044 9812 10084
rect 9944 10081 9956 10084
rect 9990 10112 10002 10115
rect 10520 10112 10548 10152
rect 11238 10140 11244 10152
rect 11296 10140 11302 10192
rect 12158 10140 12164 10192
rect 12216 10180 12222 10192
rect 12216 10152 14596 10180
rect 12216 10140 12222 10152
rect 9990 10084 10548 10112
rect 9990 10081 10002 10084
rect 9944 10075 10002 10081
rect 11054 10072 11060 10124
rect 11112 10112 11118 10124
rect 11589 10115 11647 10121
rect 11589 10112 11601 10115
rect 11112 10084 11601 10112
rect 11112 10072 11118 10084
rect 11589 10081 11601 10084
rect 11635 10112 11647 10115
rect 11882 10112 11888 10124
rect 11635 10084 11888 10112
rect 11635 10081 11647 10084
rect 11589 10075 11647 10081
rect 11882 10072 11888 10084
rect 11940 10072 11946 10124
rect 12342 10072 12348 10124
rect 12400 10112 12406 10124
rect 13357 10115 13415 10121
rect 13357 10112 13369 10115
rect 12400 10084 13369 10112
rect 12400 10072 12406 10084
rect 13357 10081 13369 10084
rect 13403 10081 13415 10115
rect 13357 10075 13415 10081
rect 13998 10072 14004 10124
rect 14056 10112 14062 10124
rect 14369 10115 14427 10121
rect 14369 10112 14381 10115
rect 14056 10084 14381 10112
rect 14056 10072 14062 10084
rect 11330 10044 11336 10056
rect 9272 10016 9812 10044
rect 11291 10016 11336 10044
rect 9272 10004 9278 10016
rect 11330 10004 11336 10016
rect 11388 10004 11394 10056
rect 13541 10047 13599 10053
rect 13541 10013 13553 10047
rect 13587 10013 13599 10047
rect 13541 10007 13599 10013
rect 10686 9936 10692 9988
rect 10744 9976 10750 9988
rect 13556 9976 13584 10007
rect 10744 9948 11192 9976
rect 10744 9936 10750 9948
rect 3697 9911 3755 9917
rect 3697 9877 3709 9911
rect 3743 9908 3755 9911
rect 3786 9908 3792 9920
rect 3743 9880 3792 9908
rect 3743 9877 3755 9880
rect 3697 9871 3755 9877
rect 3786 9868 3792 9880
rect 3844 9908 3850 9920
rect 6546 9908 6552 9920
rect 3844 9880 6552 9908
rect 3844 9868 3850 9880
rect 6546 9868 6552 9880
rect 6604 9868 6610 9920
rect 7193 9911 7251 9917
rect 7193 9877 7205 9911
rect 7239 9908 7251 9911
rect 7742 9908 7748 9920
rect 7239 9880 7748 9908
rect 7239 9877 7251 9880
rect 7193 9871 7251 9877
rect 7742 9868 7748 9880
rect 7800 9868 7806 9920
rect 7834 9868 7840 9920
rect 7892 9908 7898 9920
rect 11057 9911 11115 9917
rect 11057 9908 11069 9911
rect 7892 9880 11069 9908
rect 7892 9868 7898 9880
rect 11057 9877 11069 9880
rect 11103 9877 11115 9911
rect 11164 9908 11192 9948
rect 12268 9948 13584 9976
rect 12268 9908 12296 9948
rect 11164 9880 12296 9908
rect 11057 9871 11115 9877
rect 12710 9868 12716 9920
rect 12768 9908 12774 9920
rect 12989 9911 13047 9917
rect 12989 9908 13001 9911
rect 12768 9880 13001 9908
rect 12768 9868 12774 9880
rect 12989 9877 13001 9880
rect 13035 9877 13047 9911
rect 14108 9908 14136 10084
rect 14369 10081 14381 10084
rect 14415 10081 14427 10115
rect 14369 10075 14427 10081
rect 14182 10004 14188 10056
rect 14240 10044 14246 10056
rect 14568 10053 14596 10152
rect 14461 10047 14519 10053
rect 14461 10044 14473 10047
rect 14240 10016 14473 10044
rect 14240 10004 14246 10016
rect 14461 10013 14473 10016
rect 14507 10013 14519 10047
rect 14461 10007 14519 10013
rect 14553 10047 14611 10053
rect 14553 10013 14565 10047
rect 14599 10013 14611 10047
rect 14553 10007 14611 10013
rect 14458 9908 14464 9920
rect 14108 9880 14464 9908
rect 12989 9871 13047 9877
rect 14458 9868 14464 9880
rect 14516 9868 14522 9920
rect 1104 9818 15824 9840
rect 1104 9766 3447 9818
rect 3499 9766 3511 9818
rect 3563 9766 3575 9818
rect 3627 9766 3639 9818
rect 3691 9766 8378 9818
rect 8430 9766 8442 9818
rect 8494 9766 8506 9818
rect 8558 9766 8570 9818
rect 8622 9766 13308 9818
rect 13360 9766 13372 9818
rect 13424 9766 13436 9818
rect 13488 9766 13500 9818
rect 13552 9766 15824 9818
rect 1104 9744 15824 9766
rect 4798 9664 4804 9716
rect 4856 9704 4862 9716
rect 8110 9704 8116 9716
rect 4856 9676 8116 9704
rect 4856 9664 4862 9676
rect 8110 9664 8116 9676
rect 8168 9664 8174 9716
rect 9030 9704 9036 9716
rect 8312 9676 9036 9704
rect 7009 9639 7067 9645
rect 7009 9605 7021 9639
rect 7055 9636 7067 9639
rect 7190 9636 7196 9648
rect 7055 9608 7196 9636
rect 7055 9605 7067 9608
rect 7009 9599 7067 9605
rect 7190 9596 7196 9608
rect 7248 9596 7254 9648
rect 7374 9596 7380 9648
rect 7432 9636 7438 9648
rect 8202 9636 8208 9648
rect 7432 9608 8208 9636
rect 7432 9596 7438 9608
rect 8202 9596 8208 9608
rect 8260 9596 8266 9648
rect 1486 9528 1492 9580
rect 1544 9568 1550 9580
rect 1765 9571 1823 9577
rect 1765 9568 1777 9571
rect 1544 9540 1777 9568
rect 1544 9528 1550 9540
rect 1765 9537 1777 9540
rect 1811 9537 1823 9571
rect 5074 9568 5080 9580
rect 5035 9540 5080 9568
rect 1765 9531 1823 9537
rect 1780 9500 1808 9531
rect 5074 9528 5080 9540
rect 5132 9528 5138 9580
rect 6454 9528 6460 9580
rect 6512 9568 6518 9580
rect 6512 9540 7052 9568
rect 6512 9528 6518 9540
rect 2314 9500 2320 9512
rect 1780 9472 2320 9500
rect 2314 9460 2320 9472
rect 2372 9500 2378 9512
rect 3421 9503 3479 9509
rect 3421 9500 3433 9503
rect 2372 9472 3433 9500
rect 2372 9460 2378 9472
rect 3421 9469 3433 9472
rect 3467 9469 3479 9503
rect 7024 9500 7052 9540
rect 7098 9528 7104 9580
rect 7156 9568 7162 9580
rect 7653 9571 7711 9577
rect 7653 9568 7665 9571
rect 7156 9540 7665 9568
rect 7156 9528 7162 9540
rect 7653 9537 7665 9540
rect 7699 9568 7711 9571
rect 8312 9568 8340 9676
rect 9030 9664 9036 9676
rect 9088 9664 9094 9716
rect 9968 9676 10916 9704
rect 9490 9596 9496 9648
rect 9548 9636 9554 9648
rect 9769 9639 9827 9645
rect 9769 9636 9781 9639
rect 9548 9608 9781 9636
rect 9548 9596 9554 9608
rect 9769 9605 9781 9608
rect 9815 9605 9827 9639
rect 9769 9599 9827 9605
rect 9861 9639 9919 9645
rect 9861 9605 9873 9639
rect 9907 9636 9919 9639
rect 9968 9636 9996 9676
rect 9907 9608 9996 9636
rect 10888 9636 10916 9676
rect 10962 9664 10968 9716
rect 11020 9704 11026 9716
rect 11885 9707 11943 9713
rect 11020 9676 11560 9704
rect 11020 9664 11026 9676
rect 11422 9636 11428 9648
rect 10888 9608 11428 9636
rect 9907 9605 9919 9608
rect 9861 9599 9919 9605
rect 11422 9596 11428 9608
rect 11480 9596 11486 9648
rect 11532 9636 11560 9676
rect 11885 9673 11897 9707
rect 11931 9704 11943 9707
rect 15010 9704 15016 9716
rect 11931 9676 15016 9704
rect 11931 9673 11943 9676
rect 11885 9667 11943 9673
rect 15010 9664 15016 9676
rect 15068 9664 15074 9716
rect 11698 9636 11704 9648
rect 11532 9608 11704 9636
rect 11698 9596 11704 9608
rect 11756 9596 11762 9648
rect 14093 9639 14151 9645
rect 14093 9605 14105 9639
rect 14139 9636 14151 9639
rect 14274 9636 14280 9648
rect 14139 9608 14280 9636
rect 14139 9605 14151 9608
rect 14093 9599 14151 9605
rect 14274 9596 14280 9608
rect 14332 9596 14338 9648
rect 11330 9568 11336 9580
rect 7699 9540 8340 9568
rect 11164 9540 11336 9568
rect 7699 9537 7711 9540
rect 7653 9531 7711 9537
rect 7377 9503 7435 9509
rect 7377 9500 7389 9503
rect 7024 9472 7389 9500
rect 3421 9463 3479 9469
rect 7377 9469 7389 9472
rect 7423 9500 7435 9503
rect 7926 9500 7932 9512
rect 7423 9472 7932 9500
rect 7423 9469 7435 9472
rect 7377 9463 7435 9469
rect 7926 9460 7932 9472
rect 7984 9460 7990 9512
rect 8202 9500 8208 9512
rect 8163 9472 8208 9500
rect 8202 9460 8208 9472
rect 8260 9460 8266 9512
rect 8294 9460 8300 9512
rect 8352 9500 8358 9512
rect 9953 9503 10011 9509
rect 8352 9472 9689 9500
rect 8352 9460 8358 9472
rect 2032 9435 2090 9441
rect 2032 9401 2044 9435
rect 2078 9432 2090 9435
rect 3050 9432 3056 9444
rect 2078 9404 3056 9432
rect 2078 9401 2090 9404
rect 2032 9395 2090 9401
rect 3050 9392 3056 9404
rect 3108 9392 3114 9444
rect 3688 9435 3746 9441
rect 3688 9401 3700 9435
rect 3734 9432 3746 9435
rect 3786 9432 3792 9444
rect 3734 9404 3792 9432
rect 3734 9401 3746 9404
rect 3688 9395 3746 9401
rect 3786 9392 3792 9404
rect 3844 9392 3850 9444
rect 5344 9435 5402 9441
rect 5344 9401 5356 9435
rect 5390 9432 5402 9435
rect 5718 9432 5724 9444
rect 5390 9404 5724 9432
rect 5390 9401 5402 9404
rect 5344 9395 5402 9401
rect 5718 9392 5724 9404
rect 5776 9392 5782 9444
rect 8386 9432 8392 9444
rect 6380 9404 8392 9432
rect 2590 9324 2596 9376
rect 2648 9364 2654 9376
rect 3145 9367 3203 9373
rect 3145 9364 3157 9367
rect 2648 9336 3157 9364
rect 2648 9324 2654 9336
rect 3145 9333 3157 9336
rect 3191 9333 3203 9367
rect 3145 9327 3203 9333
rect 4801 9367 4859 9373
rect 4801 9333 4813 9367
rect 4847 9364 4859 9367
rect 6380 9364 6408 9404
rect 8386 9392 8392 9404
rect 8444 9392 8450 9444
rect 8564 9435 8622 9441
rect 8564 9401 8576 9435
rect 8610 9432 8622 9435
rect 8846 9432 8852 9444
rect 8610 9404 8852 9432
rect 8610 9401 8622 9404
rect 8564 9395 8622 9401
rect 8846 9392 8852 9404
rect 8904 9392 8910 9444
rect 9490 9432 9496 9444
rect 9232 9404 9496 9432
rect 4847 9336 6408 9364
rect 6457 9367 6515 9373
rect 4847 9333 4859 9336
rect 4801 9327 4859 9333
rect 6457 9333 6469 9367
rect 6503 9364 6515 9367
rect 6546 9364 6552 9376
rect 6503 9336 6552 9364
rect 6503 9333 6515 9336
rect 6457 9327 6515 9333
rect 6546 9324 6552 9336
rect 6604 9324 6610 9376
rect 7466 9364 7472 9376
rect 7427 9336 7472 9364
rect 7466 9324 7472 9336
rect 7524 9324 7530 9376
rect 8021 9367 8079 9373
rect 8021 9333 8033 9367
rect 8067 9364 8079 9367
rect 9232 9364 9260 9404
rect 9490 9392 9496 9404
rect 9548 9392 9554 9444
rect 9661 9432 9689 9472
rect 9953 9469 9965 9503
rect 9999 9500 10011 9503
rect 11164 9500 11192 9540
rect 11330 9528 11336 9540
rect 11388 9568 11394 9580
rect 12437 9571 12495 9577
rect 12437 9568 12449 9571
rect 11388 9540 12449 9568
rect 11388 9528 11394 9540
rect 12437 9537 12449 9540
rect 12483 9537 12495 9571
rect 12437 9531 12495 9537
rect 13446 9528 13452 9580
rect 13504 9568 13510 9580
rect 14645 9571 14703 9577
rect 14645 9568 14657 9571
rect 13504 9540 14657 9568
rect 13504 9528 13510 9540
rect 14645 9537 14657 9540
rect 14691 9537 14703 9571
rect 15102 9568 15108 9580
rect 15063 9540 15108 9568
rect 14645 9531 14703 9537
rect 15102 9528 15108 9540
rect 15160 9528 15166 9580
rect 9999 9472 11192 9500
rect 9999 9469 10011 9472
rect 9953 9463 10011 9469
rect 11238 9460 11244 9512
rect 11296 9500 11302 9512
rect 11885 9503 11943 9509
rect 11885 9500 11897 9503
rect 11296 9472 11897 9500
rect 11296 9460 11302 9472
rect 11885 9469 11897 9472
rect 11931 9469 11943 9503
rect 11885 9463 11943 9469
rect 11974 9460 11980 9512
rect 12032 9500 12038 9512
rect 12253 9503 12311 9509
rect 12253 9500 12265 9503
rect 12032 9472 12265 9500
rect 12032 9460 12038 9472
rect 12253 9469 12265 9472
rect 12299 9469 12311 9503
rect 12253 9463 12311 9469
rect 12986 9460 12992 9512
rect 13044 9500 13050 9512
rect 13170 9500 13176 9512
rect 13044 9472 13176 9500
rect 13044 9460 13050 9472
rect 13170 9460 13176 9472
rect 13228 9460 13234 9512
rect 10226 9441 10232 9444
rect 10220 9432 10232 9441
rect 9661 9404 9812 9432
rect 10187 9404 10232 9432
rect 8067 9336 9260 9364
rect 8067 9333 8079 9336
rect 8021 9327 8079 9333
rect 9306 9324 9312 9376
rect 9364 9364 9370 9376
rect 9677 9367 9735 9373
rect 9677 9364 9689 9367
rect 9364 9336 9689 9364
rect 9364 9324 9370 9336
rect 9677 9333 9689 9336
rect 9723 9333 9735 9367
rect 9784 9364 9812 9404
rect 10220 9395 10232 9404
rect 10226 9392 10232 9395
rect 10284 9392 10290 9444
rect 11609 9435 11667 9441
rect 10336 9404 11468 9432
rect 10336 9364 10364 9404
rect 9784 9336 10364 9364
rect 9677 9327 9735 9333
rect 11238 9324 11244 9376
rect 11296 9364 11302 9376
rect 11333 9367 11391 9373
rect 11333 9364 11345 9367
rect 11296 9336 11345 9364
rect 11296 9324 11302 9336
rect 11333 9333 11345 9336
rect 11379 9333 11391 9367
rect 11440 9364 11468 9404
rect 11609 9401 11621 9435
rect 11655 9432 11667 9435
rect 12158 9432 12164 9444
rect 11655 9404 12164 9432
rect 11655 9401 11667 9404
rect 11609 9395 11667 9401
rect 12158 9392 12164 9404
rect 12216 9392 12222 9444
rect 12434 9392 12440 9444
rect 12492 9432 12498 9444
rect 12682 9435 12740 9441
rect 12682 9432 12694 9435
rect 12492 9404 12694 9432
rect 12492 9392 12498 9404
rect 12682 9401 12694 9404
rect 12728 9401 12740 9435
rect 12682 9395 12740 9401
rect 12802 9392 12808 9444
rect 12860 9432 12866 9444
rect 14461 9435 14519 9441
rect 14461 9432 14473 9435
rect 12860 9404 14473 9432
rect 12860 9392 12866 9404
rect 14461 9401 14473 9404
rect 14507 9401 14519 9435
rect 14461 9395 14519 9401
rect 12069 9367 12127 9373
rect 12069 9364 12081 9367
rect 11440 9336 12081 9364
rect 11333 9327 11391 9333
rect 12069 9333 12081 9336
rect 12115 9333 12127 9367
rect 12069 9327 12127 9333
rect 13262 9324 13268 9376
rect 13320 9364 13326 9376
rect 13817 9367 13875 9373
rect 13817 9364 13829 9367
rect 13320 9336 13829 9364
rect 13320 9324 13326 9336
rect 13817 9333 13829 9336
rect 13863 9333 13875 9367
rect 13817 9327 13875 9333
rect 13906 9324 13912 9376
rect 13964 9364 13970 9376
rect 14553 9367 14611 9373
rect 14553 9364 14565 9367
rect 13964 9336 14565 9364
rect 13964 9324 13970 9336
rect 14553 9333 14565 9336
rect 14599 9333 14611 9367
rect 14553 9327 14611 9333
rect 1104 9274 15824 9296
rect 1104 9222 5912 9274
rect 5964 9222 5976 9274
rect 6028 9222 6040 9274
rect 6092 9222 6104 9274
rect 6156 9222 10843 9274
rect 10895 9222 10907 9274
rect 10959 9222 10971 9274
rect 11023 9222 11035 9274
rect 11087 9222 15824 9274
rect 1104 9200 15824 9222
rect 2866 9120 2872 9172
rect 2924 9160 2930 9172
rect 3697 9163 3755 9169
rect 3697 9160 3709 9163
rect 2924 9132 3709 9160
rect 2924 9120 2930 9132
rect 3697 9129 3709 9132
rect 3743 9160 3755 9163
rect 3970 9160 3976 9172
rect 3743 9132 3976 9160
rect 3743 9129 3755 9132
rect 3697 9123 3755 9129
rect 3970 9120 3976 9132
rect 4028 9120 4034 9172
rect 4062 9120 4068 9172
rect 4120 9160 4126 9172
rect 4246 9160 4252 9172
rect 4120 9132 4252 9160
rect 4120 9120 4126 9132
rect 4246 9120 4252 9132
rect 4304 9120 4310 9172
rect 5629 9163 5687 9169
rect 5629 9129 5641 9163
rect 5675 9160 5687 9163
rect 7282 9160 7288 9172
rect 5675 9132 7288 9160
rect 5675 9129 5687 9132
rect 5629 9123 5687 9129
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 7558 9120 7564 9172
rect 7616 9160 7622 9172
rect 8202 9160 8208 9172
rect 7616 9132 8208 9160
rect 7616 9120 7622 9132
rect 8202 9120 8208 9132
rect 8260 9160 8266 9172
rect 8665 9163 8723 9169
rect 8665 9160 8677 9163
rect 8260 9132 8677 9160
rect 8260 9120 8266 9132
rect 8665 9129 8677 9132
rect 8711 9129 8723 9163
rect 11057 9163 11115 9169
rect 8665 9123 8723 9129
rect 9784 9132 10263 9160
rect 1854 9092 1860 9104
rect 1815 9064 1860 9092
rect 1854 9052 1860 9064
rect 1912 9052 1918 9104
rect 2590 9101 2596 9104
rect 2584 9092 2596 9101
rect 2551 9064 2596 9092
rect 2584 9055 2596 9064
rect 2590 9052 2596 9055
rect 2648 9052 2654 9104
rect 2682 9052 2688 9104
rect 2740 9052 2746 9104
rect 4516 9095 4574 9101
rect 4516 9061 4528 9095
rect 4562 9092 4574 9095
rect 6546 9092 6552 9104
rect 4562 9064 6552 9092
rect 4562 9061 4574 9064
rect 4516 9055 4574 9061
rect 6546 9052 6552 9064
rect 6604 9052 6610 9104
rect 7377 9095 7435 9101
rect 7377 9061 7389 9095
rect 7423 9092 7435 9095
rect 9784 9092 9812 9132
rect 9950 9101 9956 9104
rect 7423 9064 9812 9092
rect 9933 9095 9956 9101
rect 7423 9061 7435 9064
rect 7377 9055 7435 9061
rect 9933 9061 9945 9095
rect 10008 9092 10014 9104
rect 10134 9092 10140 9104
rect 10008 9064 10140 9092
rect 9933 9055 9956 9061
rect 9950 9052 9956 9055
rect 10008 9052 10014 9064
rect 10134 9052 10140 9064
rect 10192 9052 10198 9104
rect 10235 9092 10263 9132
rect 11057 9129 11069 9163
rect 11103 9160 11115 9163
rect 11238 9160 11244 9172
rect 11103 9132 11244 9160
rect 11103 9129 11115 9132
rect 11057 9123 11115 9129
rect 11238 9120 11244 9132
rect 11296 9120 11302 9172
rect 11330 9120 11336 9172
rect 11388 9160 11394 9172
rect 11388 9132 12020 9160
rect 11388 9120 11394 9132
rect 11790 9092 11796 9104
rect 10235 9064 11796 9092
rect 11790 9052 11796 9064
rect 11848 9052 11854 9104
rect 1581 9027 1639 9033
rect 1581 8993 1593 9027
rect 1627 9024 1639 9027
rect 2700 9024 2728 9052
rect 1627 8996 2728 9024
rect 1627 8993 1639 8996
rect 1581 8987 1639 8993
rect 4154 8984 4160 9036
rect 4212 9024 4218 9036
rect 4249 9027 4307 9033
rect 4249 9024 4261 9027
rect 4212 8996 4261 9024
rect 4212 8984 4218 8996
rect 4249 8993 4261 8996
rect 4295 8993 4307 9027
rect 4249 8987 4307 8993
rect 5074 8984 5080 9036
rect 5132 9024 5138 9036
rect 5721 9027 5779 9033
rect 5721 9024 5733 9027
rect 5132 8996 5733 9024
rect 5132 8984 5138 8996
rect 5721 8993 5733 8996
rect 5767 8993 5779 9027
rect 5721 8987 5779 8993
rect 5988 9027 6046 9033
rect 5988 8993 6000 9027
rect 6034 9024 6046 9027
rect 6034 8996 7604 9024
rect 6034 8993 6046 8996
rect 5988 8987 6046 8993
rect 2314 8956 2320 8968
rect 2275 8928 2320 8956
rect 2314 8916 2320 8928
rect 2372 8916 2378 8968
rect 7576 8956 7604 8996
rect 7650 8984 7656 9036
rect 7708 9024 7714 9036
rect 7708 8996 8984 9024
rect 7708 8984 7714 8996
rect 7834 8956 7840 8968
rect 7576 8928 7840 8956
rect 7834 8916 7840 8928
rect 7892 8916 7898 8968
rect 8956 8956 8984 8996
rect 9214 8984 9220 9036
rect 9272 9024 9278 9036
rect 9677 9027 9735 9033
rect 9677 9024 9689 9027
rect 9272 8996 9689 9024
rect 9272 8984 9278 8996
rect 9677 8993 9689 8996
rect 9723 8993 9735 9027
rect 11054 9024 11060 9036
rect 9677 8987 9735 8993
rect 9775 8996 11060 9024
rect 9775 8956 9803 8996
rect 11054 8984 11060 8996
rect 11112 8984 11118 9036
rect 11330 9024 11336 9036
rect 11291 8996 11336 9024
rect 11330 8984 11336 8996
rect 11388 8984 11394 9036
rect 11600 9027 11658 9033
rect 11600 9024 11612 9027
rect 11440 8996 11612 9024
rect 8956 8928 9803 8956
rect 11146 8916 11152 8968
rect 11204 8956 11210 8968
rect 11440 8956 11468 8996
rect 11600 8993 11612 8996
rect 11646 9024 11658 9027
rect 11882 9024 11888 9036
rect 11646 8996 11888 9024
rect 11646 8993 11658 8996
rect 11600 8987 11658 8993
rect 11882 8984 11888 8996
rect 11940 8984 11946 9036
rect 11992 9024 12020 9132
rect 12158 9120 12164 9172
rect 12216 9160 12222 9172
rect 14369 9163 14427 9169
rect 14369 9160 14381 9163
rect 12216 9132 14381 9160
rect 12216 9120 12222 9132
rect 14369 9129 14381 9132
rect 14415 9129 14427 9163
rect 14369 9123 14427 9129
rect 14550 9120 14556 9172
rect 14608 9160 14614 9172
rect 14645 9163 14703 9169
rect 14645 9160 14657 9163
rect 14608 9132 14657 9160
rect 14608 9120 14614 9132
rect 14645 9129 14657 9132
rect 14691 9129 14703 9163
rect 14645 9123 14703 9129
rect 12710 9052 12716 9104
rect 12768 9092 12774 9104
rect 13722 9092 13728 9104
rect 12768 9064 13728 9092
rect 12768 9052 12774 9064
rect 13722 9052 13728 9064
rect 13780 9052 13786 9104
rect 12989 9027 13047 9033
rect 12989 9024 13001 9027
rect 11992 8996 13001 9024
rect 12989 8993 13001 8996
rect 13035 8993 13047 9027
rect 12989 8987 13047 8993
rect 13256 9027 13314 9033
rect 13256 8993 13268 9027
rect 13302 9024 13314 9027
rect 13302 8996 14044 9024
rect 13302 8993 13314 8996
rect 13256 8987 13314 8993
rect 11204 8928 11468 8956
rect 11204 8916 11210 8928
rect 11330 8888 11336 8900
rect 10980 8860 11336 8888
rect 5350 8780 5356 8832
rect 5408 8820 5414 8832
rect 7101 8823 7159 8829
rect 7101 8820 7113 8823
rect 5408 8792 7113 8820
rect 5408 8780 5414 8792
rect 7101 8789 7113 8792
rect 7147 8789 7159 8823
rect 7101 8783 7159 8789
rect 7926 8780 7932 8832
rect 7984 8820 7990 8832
rect 9122 8820 9128 8832
rect 7984 8792 9128 8820
rect 7984 8780 7990 8792
rect 9122 8780 9128 8792
rect 9180 8780 9186 8832
rect 9306 8780 9312 8832
rect 9364 8820 9370 8832
rect 10980 8820 11008 8860
rect 11330 8848 11336 8860
rect 11388 8848 11394 8900
rect 14016 8888 14044 8996
rect 13924 8860 14044 8888
rect 9364 8792 11008 8820
rect 9364 8780 9370 8792
rect 11054 8780 11060 8832
rect 11112 8820 11118 8832
rect 12434 8820 12440 8832
rect 11112 8792 12440 8820
rect 11112 8780 11118 8792
rect 12434 8780 12440 8792
rect 12492 8780 12498 8832
rect 12710 8820 12716 8832
rect 12671 8792 12716 8820
rect 12710 8780 12716 8792
rect 12768 8780 12774 8832
rect 13722 8780 13728 8832
rect 13780 8820 13786 8832
rect 13924 8820 13952 8860
rect 14090 8848 14096 8900
rect 14148 8888 14154 8900
rect 14274 8888 14280 8900
rect 14148 8860 14280 8888
rect 14148 8848 14154 8860
rect 14274 8848 14280 8860
rect 14332 8848 14338 8900
rect 13780 8792 13952 8820
rect 13780 8780 13786 8792
rect 13998 8780 14004 8832
rect 14056 8820 14062 8832
rect 14734 8820 14740 8832
rect 14056 8792 14740 8820
rect 14056 8780 14062 8792
rect 14734 8780 14740 8792
rect 14792 8780 14798 8832
rect 1104 8730 15824 8752
rect 1104 8678 3447 8730
rect 3499 8678 3511 8730
rect 3563 8678 3575 8730
rect 3627 8678 3639 8730
rect 3691 8678 8378 8730
rect 8430 8678 8442 8730
rect 8494 8678 8506 8730
rect 8558 8678 8570 8730
rect 8622 8678 13308 8730
rect 13360 8678 13372 8730
rect 13424 8678 13436 8730
rect 13488 8678 13500 8730
rect 13552 8678 15824 8730
rect 1104 8656 15824 8678
rect 4801 8619 4859 8625
rect 3344 8588 4384 8616
rect 1670 8440 1676 8492
rect 1728 8480 1734 8492
rect 1765 8483 1823 8489
rect 1765 8480 1777 8483
rect 1728 8452 1777 8480
rect 1728 8440 1734 8452
rect 1765 8449 1777 8452
rect 1811 8449 1823 8483
rect 1765 8443 1823 8449
rect 1780 8344 1808 8443
rect 2032 8415 2090 8421
rect 2032 8381 2044 8415
rect 2078 8412 2090 8415
rect 3344 8412 3372 8588
rect 4356 8548 4384 8588
rect 4801 8585 4813 8619
rect 4847 8616 4859 8619
rect 6914 8616 6920 8628
rect 4847 8588 6920 8616
rect 4847 8585 4859 8588
rect 4801 8579 4859 8585
rect 6914 8576 6920 8588
rect 6972 8576 6978 8628
rect 7009 8619 7067 8625
rect 7009 8585 7021 8619
rect 7055 8616 7067 8619
rect 7098 8616 7104 8628
rect 7055 8588 7104 8616
rect 7055 8585 7067 8588
rect 7009 8579 7067 8585
rect 7098 8576 7104 8588
rect 7156 8576 7162 8628
rect 7374 8616 7380 8628
rect 7335 8588 7380 8616
rect 7374 8576 7380 8588
rect 7432 8576 7438 8628
rect 8202 8616 8208 8628
rect 7944 8588 8208 8616
rect 5074 8548 5080 8560
rect 4356 8520 5080 8548
rect 5074 8508 5080 8520
rect 5132 8508 5138 8560
rect 6457 8551 6515 8557
rect 6457 8517 6469 8551
rect 6503 8548 6515 8551
rect 6503 8520 7788 8548
rect 6503 8517 6515 8520
rect 6457 8511 6515 8517
rect 7466 8480 7472 8492
rect 7116 8452 7472 8480
rect 2078 8384 3372 8412
rect 3421 8415 3479 8421
rect 2078 8381 2090 8384
rect 2032 8375 2090 8381
rect 3421 8381 3433 8415
rect 3467 8381 3479 8415
rect 3421 8375 3479 8381
rect 2314 8344 2320 8356
rect 1780 8316 2320 8344
rect 2314 8304 2320 8316
rect 2372 8344 2378 8356
rect 3326 8344 3332 8356
rect 2372 8316 3332 8344
rect 2372 8304 2378 8316
rect 3326 8304 3332 8316
rect 3384 8344 3390 8356
rect 3436 8344 3464 8375
rect 4614 8372 4620 8424
rect 4672 8412 4678 8424
rect 5077 8415 5135 8421
rect 5077 8412 5089 8415
rect 4672 8384 5089 8412
rect 4672 8372 4678 8384
rect 5077 8381 5089 8384
rect 5123 8381 5135 8415
rect 6850 8415 6908 8421
rect 5077 8375 5135 8381
rect 5276 8384 6592 8412
rect 3384 8316 3464 8344
rect 3688 8347 3746 8353
rect 3384 8304 3390 8316
rect 3688 8313 3700 8347
rect 3734 8344 3746 8347
rect 5276 8344 5304 8384
rect 3734 8316 5304 8344
rect 5333 8347 5391 8353
rect 3734 8313 3746 8316
rect 3688 8307 3746 8313
rect 5333 8313 5345 8347
rect 5379 8313 5391 8347
rect 6564 8344 6592 8384
rect 6850 8381 6862 8415
rect 6896 8412 6908 8415
rect 7116 8412 7144 8452
rect 7466 8440 7472 8452
rect 7524 8440 7530 8492
rect 7558 8412 7564 8424
rect 6896 8384 7144 8412
rect 7519 8384 7564 8412
rect 6896 8381 6908 8384
rect 6850 8375 6908 8381
rect 7558 8372 7564 8384
rect 7616 8372 7622 8424
rect 7760 8412 7788 8520
rect 7944 8492 7972 8588
rect 8202 8576 8208 8588
rect 8260 8576 8266 8628
rect 8662 8576 8668 8628
rect 8720 8616 8726 8628
rect 8846 8616 8852 8628
rect 8720 8588 8852 8616
rect 8720 8576 8726 8588
rect 8846 8576 8852 8588
rect 8904 8576 8910 8628
rect 9122 8576 9128 8628
rect 9180 8616 9186 8628
rect 10873 8619 10931 8625
rect 10873 8616 10885 8619
rect 9180 8588 10885 8616
rect 9180 8576 9186 8588
rect 10873 8585 10885 8588
rect 10919 8585 10931 8619
rect 10873 8579 10931 8585
rect 10962 8576 10968 8628
rect 11020 8616 11026 8628
rect 11020 8588 12480 8616
rect 11020 8576 11026 8588
rect 9309 8551 9367 8557
rect 9309 8548 9321 8551
rect 8956 8520 9321 8548
rect 7926 8480 7932 8492
rect 7839 8452 7932 8480
rect 7926 8440 7932 8452
rect 7984 8440 7990 8492
rect 8018 8412 8024 8424
rect 7760 8384 8024 8412
rect 8018 8372 8024 8384
rect 8076 8372 8082 8424
rect 8202 8421 8208 8424
rect 8196 8375 8208 8421
rect 8260 8412 8266 8424
rect 8260 8384 8296 8412
rect 8202 8372 8208 8375
rect 8260 8372 8266 8384
rect 8570 8372 8576 8424
rect 8628 8412 8634 8424
rect 8956 8412 8984 8520
rect 9309 8517 9321 8520
rect 9355 8517 9367 8551
rect 9309 8511 9367 8517
rect 10686 8508 10692 8560
rect 10744 8548 10750 8560
rect 11514 8548 11520 8560
rect 10744 8520 11520 8548
rect 10744 8508 10750 8520
rect 11514 8508 11520 8520
rect 11572 8508 11578 8560
rect 11790 8508 11796 8560
rect 11848 8548 11854 8560
rect 12342 8548 12348 8560
rect 11848 8520 12348 8548
rect 11848 8508 11854 8520
rect 12342 8508 12348 8520
rect 12400 8508 12406 8560
rect 9214 8440 9220 8492
rect 9272 8480 9278 8492
rect 11422 8480 11428 8492
rect 9272 8452 9444 8480
rect 9272 8440 9278 8452
rect 9416 8421 9444 8452
rect 10520 8452 11428 8480
rect 8628 8384 8984 8412
rect 9401 8415 9459 8421
rect 8628 8372 8634 8384
rect 9401 8381 9413 8415
rect 9447 8412 9459 8415
rect 10134 8412 10140 8424
rect 9447 8384 10140 8412
rect 9447 8381 9459 8384
rect 9401 8375 9459 8381
rect 10134 8372 10140 8384
rect 10192 8372 10198 8424
rect 7742 8344 7748 8356
rect 6564 8316 7748 8344
rect 5333 8307 5391 8313
rect 3145 8279 3203 8285
rect 3145 8245 3157 8279
rect 3191 8276 3203 8279
rect 3878 8276 3884 8288
rect 3191 8248 3884 8276
rect 3191 8245 3203 8248
rect 3145 8239 3203 8245
rect 3878 8236 3884 8248
rect 3936 8236 3942 8288
rect 4798 8236 4804 8288
rect 4856 8276 4862 8288
rect 5348 8276 5376 8307
rect 7742 8304 7748 8316
rect 7800 8304 7806 8356
rect 9214 8344 9220 8356
rect 7944 8316 9220 8344
rect 4856 8248 5376 8276
rect 4856 8236 4862 8248
rect 5442 8236 5448 8288
rect 5500 8276 5506 8288
rect 7006 8276 7012 8288
rect 5500 8248 7012 8276
rect 5500 8236 5506 8248
rect 7006 8236 7012 8248
rect 7064 8236 7070 8288
rect 7282 8236 7288 8288
rect 7340 8276 7346 8288
rect 7944 8276 7972 8316
rect 9214 8304 9220 8316
rect 9272 8344 9278 8356
rect 9646 8347 9704 8353
rect 9646 8344 9658 8347
rect 9272 8316 9658 8344
rect 9272 8304 9278 8316
rect 9646 8313 9658 8316
rect 9692 8313 9704 8347
rect 9646 8307 9704 8313
rect 7340 8248 7972 8276
rect 7340 8236 7346 8248
rect 8018 8236 8024 8288
rect 8076 8276 8082 8288
rect 9950 8276 9956 8288
rect 8076 8248 9956 8276
rect 8076 8236 8082 8248
rect 9950 8236 9956 8248
rect 10008 8276 10014 8288
rect 10520 8276 10548 8452
rect 11422 8440 11428 8452
rect 11480 8440 11486 8492
rect 12452 8480 12480 8588
rect 12618 8576 12624 8628
rect 12676 8616 12682 8628
rect 13814 8616 13820 8628
rect 12676 8588 13492 8616
rect 13775 8588 13820 8616
rect 12676 8576 12682 8588
rect 13464 8560 13492 8588
rect 13814 8576 13820 8588
rect 13872 8576 13878 8628
rect 13924 8588 14504 8616
rect 13446 8508 13452 8560
rect 13504 8508 13510 8560
rect 13924 8548 13952 8588
rect 14090 8548 14096 8560
rect 13556 8520 13952 8548
rect 14051 8520 14096 8548
rect 12452 8452 12572 8480
rect 10594 8372 10600 8424
rect 10652 8372 10658 8424
rect 10778 8372 10784 8424
rect 10836 8412 10842 8424
rect 11241 8415 11299 8421
rect 11241 8412 11253 8415
rect 10836 8384 11253 8412
rect 10836 8372 10842 8384
rect 11241 8381 11253 8384
rect 11287 8381 11299 8415
rect 11241 8375 11299 8381
rect 11514 8372 11520 8424
rect 11572 8412 11578 8424
rect 11885 8415 11943 8421
rect 11885 8412 11897 8415
rect 11572 8384 11897 8412
rect 11572 8372 11578 8384
rect 11885 8381 11897 8384
rect 11931 8381 11943 8415
rect 12434 8412 12440 8424
rect 12395 8384 12440 8412
rect 11885 8375 11943 8381
rect 12434 8372 12440 8384
rect 12492 8372 12498 8424
rect 12544 8412 12572 8452
rect 12693 8415 12751 8421
rect 12693 8412 12705 8415
rect 12544 8384 12705 8412
rect 12693 8381 12705 8384
rect 12739 8412 12751 8415
rect 13556 8412 13584 8520
rect 14090 8508 14096 8520
rect 14148 8508 14154 8560
rect 13630 8440 13636 8492
rect 13688 8480 13694 8492
rect 14476 8480 14504 8588
rect 14645 8483 14703 8489
rect 14645 8480 14657 8483
rect 13688 8452 14412 8480
rect 14476 8452 14657 8480
rect 13688 8440 13694 8452
rect 12739 8384 13584 8412
rect 12739 8381 12751 8384
rect 12693 8375 12751 8381
rect 10008 8248 10548 8276
rect 10612 8276 10640 8372
rect 11333 8347 11391 8353
rect 11333 8313 11345 8347
rect 11379 8344 11391 8347
rect 13998 8344 14004 8356
rect 11379 8316 14004 8344
rect 11379 8313 11391 8316
rect 11333 8307 11391 8313
rect 13998 8304 14004 8316
rect 14056 8304 14062 8356
rect 10781 8279 10839 8285
rect 10781 8276 10793 8279
rect 10612 8248 10793 8276
rect 10008 8236 10014 8248
rect 10781 8245 10793 8248
rect 10827 8245 10839 8279
rect 10781 8239 10839 8245
rect 13078 8236 13084 8288
rect 13136 8276 13142 8288
rect 13722 8276 13728 8288
rect 13136 8248 13728 8276
rect 13136 8236 13142 8248
rect 13722 8236 13728 8248
rect 13780 8236 13786 8288
rect 14384 8276 14412 8452
rect 14645 8449 14657 8452
rect 14691 8449 14703 8483
rect 14645 8443 14703 8449
rect 14550 8344 14556 8356
rect 14511 8316 14556 8344
rect 14550 8304 14556 8316
rect 14608 8304 14614 8356
rect 14461 8279 14519 8285
rect 14461 8276 14473 8279
rect 14384 8248 14473 8276
rect 14461 8245 14473 8248
rect 14507 8245 14519 8279
rect 15102 8276 15108 8288
rect 15063 8248 15108 8276
rect 14461 8239 14519 8245
rect 15102 8236 15108 8248
rect 15160 8236 15166 8288
rect 1104 8186 15824 8208
rect 1104 8134 5912 8186
rect 5964 8134 5976 8186
rect 6028 8134 6040 8186
rect 6092 8134 6104 8186
rect 6156 8134 10843 8186
rect 10895 8134 10907 8186
rect 10959 8134 10971 8186
rect 11023 8134 11035 8186
rect 11087 8134 15824 8186
rect 1104 8112 15824 8134
rect 3694 8072 3700 8084
rect 3655 8044 3700 8072
rect 3694 8032 3700 8044
rect 3752 8032 3758 8084
rect 4890 8072 4896 8084
rect 3988 8044 4896 8072
rect 1581 7939 1639 7945
rect 1581 7905 1593 7939
rect 1627 7936 1639 7939
rect 2130 7936 2136 7948
rect 1627 7908 2136 7936
rect 1627 7905 1639 7908
rect 1581 7899 1639 7905
rect 2130 7896 2136 7908
rect 2188 7896 2194 7948
rect 2314 7896 2320 7948
rect 2372 7936 2378 7948
rect 2584 7939 2642 7945
rect 2372 7908 2417 7936
rect 2372 7896 2378 7908
rect 2584 7905 2596 7939
rect 2630 7936 2642 7939
rect 3988 7936 4016 8044
rect 4890 8032 4896 8044
rect 4948 8032 4954 8084
rect 5997 8075 6055 8081
rect 5997 8041 6009 8075
rect 6043 8072 6055 8075
rect 6914 8072 6920 8084
rect 6043 8044 6920 8072
rect 6043 8041 6055 8044
rect 5997 8035 6055 8041
rect 6914 8032 6920 8044
rect 6972 8032 6978 8084
rect 8202 8032 8208 8084
rect 8260 8072 8266 8084
rect 8938 8072 8944 8084
rect 8260 8044 8944 8072
rect 8260 8032 8266 8044
rect 8938 8032 8944 8044
rect 8996 8032 9002 8084
rect 10502 8072 10508 8084
rect 9140 8044 10508 8072
rect 4154 7964 4160 8016
rect 4212 8004 4218 8016
rect 4341 8007 4399 8013
rect 4341 8004 4353 8007
rect 4212 7976 4353 8004
rect 4212 7964 4218 7976
rect 4341 7973 4353 7976
rect 4387 7973 4399 8007
rect 5534 8004 5540 8016
rect 4341 7967 4399 7973
rect 4816 7976 5540 8004
rect 2630 7908 4016 7936
rect 4065 7939 4123 7945
rect 2630 7905 2642 7908
rect 2584 7899 2642 7905
rect 4065 7905 4077 7939
rect 4111 7936 4123 7939
rect 4816 7936 4844 7976
rect 5534 7964 5540 7976
rect 5592 7964 5598 8016
rect 7926 8004 7932 8016
rect 6104 7976 7236 8004
rect 4111 7908 4844 7936
rect 4884 7939 4942 7945
rect 4111 7905 4123 7908
rect 4065 7899 4123 7905
rect 4884 7905 4896 7939
rect 4930 7936 4942 7939
rect 5166 7936 5172 7948
rect 4930 7908 5172 7936
rect 4930 7905 4942 7908
rect 4884 7899 4942 7905
rect 5166 7896 5172 7908
rect 5224 7896 5230 7948
rect 6104 7945 6132 7976
rect 7208 7948 7236 7976
rect 7576 7976 7932 8004
rect 6089 7939 6147 7945
rect 6089 7905 6101 7939
rect 6135 7905 6147 7939
rect 6089 7899 6147 7905
rect 6356 7939 6414 7945
rect 6356 7905 6368 7939
rect 6402 7936 6414 7939
rect 6638 7936 6644 7948
rect 6402 7908 6644 7936
rect 6402 7905 6414 7908
rect 6356 7899 6414 7905
rect 6638 7896 6644 7908
rect 6696 7896 6702 7948
rect 7190 7896 7196 7948
rect 7248 7936 7254 7948
rect 7576 7945 7604 7976
rect 7926 7964 7932 7976
rect 7984 7964 7990 8016
rect 8570 8004 8576 8016
rect 8036 7976 8576 8004
rect 7561 7939 7619 7945
rect 7561 7936 7573 7939
rect 7248 7908 7573 7936
rect 7248 7896 7254 7908
rect 7561 7905 7573 7908
rect 7607 7905 7619 7939
rect 7561 7899 7619 7905
rect 7650 7896 7656 7948
rect 7708 7936 7714 7948
rect 7817 7939 7875 7945
rect 7817 7936 7829 7939
rect 7708 7908 7829 7936
rect 7708 7896 7714 7908
rect 7817 7905 7829 7908
rect 7863 7936 7875 7939
rect 8036 7936 8064 7976
rect 8570 7964 8576 7976
rect 8628 7964 8634 8016
rect 7863 7908 8064 7936
rect 7863 7905 7875 7908
rect 7817 7899 7875 7905
rect 8110 7896 8116 7948
rect 8168 7936 8174 7948
rect 9033 7939 9091 7945
rect 9033 7936 9045 7939
rect 8168 7908 9045 7936
rect 8168 7896 8174 7908
rect 9033 7905 9045 7908
rect 9079 7905 9091 7939
rect 9033 7899 9091 7905
rect 1762 7868 1768 7880
rect 1723 7840 1768 7868
rect 1762 7828 1768 7840
rect 1820 7828 1826 7880
rect 3326 7828 3332 7880
rect 3384 7868 3390 7880
rect 4614 7868 4620 7880
rect 3384 7840 4620 7868
rect 3384 7828 3390 7840
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 7282 7828 7288 7880
rect 7340 7868 7346 7880
rect 7668 7868 7696 7896
rect 7340 7840 7696 7868
rect 7340 7828 7346 7840
rect 8570 7828 8576 7880
rect 8628 7868 8634 7880
rect 9140 7868 9168 8044
rect 10502 8032 10508 8044
rect 10560 8032 10566 8084
rect 12526 8032 12532 8084
rect 12584 8072 12590 8084
rect 14369 8075 14427 8081
rect 14369 8072 14381 8075
rect 12584 8044 14381 8072
rect 12584 8032 12590 8044
rect 14369 8041 14381 8044
rect 14415 8041 14427 8075
rect 14369 8035 14427 8041
rect 10134 8004 10140 8016
rect 9692 7976 10140 8004
rect 9692 7945 9720 7976
rect 10134 7964 10140 7976
rect 10192 8004 10198 8016
rect 11600 8007 11658 8013
rect 10192 7976 11376 8004
rect 10192 7964 10198 7976
rect 9950 7945 9956 7948
rect 9677 7939 9735 7945
rect 9677 7905 9689 7939
rect 9723 7905 9735 7939
rect 9944 7936 9956 7945
rect 9911 7908 9956 7936
rect 9677 7899 9735 7905
rect 9944 7899 9956 7908
rect 9950 7896 9956 7899
rect 10008 7896 10014 7948
rect 11348 7945 11376 7976
rect 11600 7973 11612 8007
rect 11646 8004 11658 8007
rect 11698 8004 11704 8016
rect 11646 7976 11704 8004
rect 11646 7973 11658 7976
rect 11600 7967 11658 7973
rect 11698 7964 11704 7976
rect 11756 7964 11762 8016
rect 12618 7964 12624 8016
rect 12676 8004 12682 8016
rect 13449 8007 13507 8013
rect 13449 8004 13461 8007
rect 12676 7976 13461 8004
rect 12676 7964 12682 7976
rect 13449 7973 13461 7976
rect 13495 8004 13507 8007
rect 14642 8004 14648 8016
rect 13495 7976 14648 8004
rect 13495 7973 13507 7976
rect 13449 7967 13507 7973
rect 14642 7964 14648 7976
rect 14700 7964 14706 8016
rect 11333 7939 11391 7945
rect 11333 7905 11345 7939
rect 11379 7936 11391 7939
rect 12434 7936 12440 7948
rect 11379 7908 12440 7936
rect 11379 7905 11391 7908
rect 11333 7899 11391 7905
rect 12434 7896 12440 7908
rect 12492 7936 12498 7948
rect 13170 7936 13176 7948
rect 12492 7908 13176 7936
rect 12492 7896 12498 7908
rect 13170 7896 13176 7908
rect 13228 7896 13234 7948
rect 13357 7939 13415 7945
rect 13357 7905 13369 7939
rect 13403 7936 13415 7939
rect 14461 7939 14519 7945
rect 14461 7936 14473 7939
rect 13403 7908 13768 7936
rect 13403 7905 13415 7908
rect 13357 7899 13415 7905
rect 8628 7840 9168 7868
rect 9217 7871 9275 7877
rect 8628 7828 8634 7840
rect 9217 7837 9229 7871
rect 9263 7837 9275 7871
rect 9217 7831 9275 7837
rect 9232 7800 9260 7831
rect 12342 7828 12348 7880
rect 12400 7868 12406 7880
rect 13541 7871 13599 7877
rect 13541 7868 13553 7871
rect 12400 7840 13553 7868
rect 12400 7828 12406 7840
rect 13541 7837 13553 7840
rect 13587 7837 13599 7871
rect 13541 7831 13599 7837
rect 13740 7800 13768 7908
rect 14108 7908 14473 7936
rect 13814 7800 13820 7812
rect 7015 7772 7604 7800
rect 1302 7692 1308 7744
rect 1360 7732 1366 7744
rect 7015 7732 7043 7772
rect 7466 7732 7472 7744
rect 1360 7704 7043 7732
rect 7427 7704 7472 7732
rect 1360 7692 1366 7704
rect 7466 7692 7472 7704
rect 7524 7692 7530 7744
rect 7576 7732 7604 7772
rect 8496 7772 9260 7800
rect 12268 7772 13124 7800
rect 13740 7772 13820 7800
rect 8496 7732 8524 7772
rect 8938 7732 8944 7744
rect 7576 7704 8524 7732
rect 8899 7704 8944 7732
rect 8938 7692 8944 7704
rect 8996 7692 9002 7744
rect 9214 7692 9220 7744
rect 9272 7732 9278 7744
rect 11057 7735 11115 7741
rect 11057 7732 11069 7735
rect 9272 7704 11069 7732
rect 9272 7692 9278 7704
rect 11057 7701 11069 7704
rect 11103 7701 11115 7735
rect 11057 7695 11115 7701
rect 11146 7692 11152 7744
rect 11204 7732 11210 7744
rect 12268 7732 12296 7772
rect 12710 7732 12716 7744
rect 11204 7704 12296 7732
rect 12671 7704 12716 7732
rect 11204 7692 11210 7704
rect 12710 7692 12716 7704
rect 12768 7692 12774 7744
rect 12802 7692 12808 7744
rect 12860 7732 12866 7744
rect 12989 7735 13047 7741
rect 12989 7732 13001 7735
rect 12860 7704 13001 7732
rect 12860 7692 12866 7704
rect 12989 7701 13001 7704
rect 13035 7701 13047 7735
rect 13096 7732 13124 7772
rect 13814 7760 13820 7772
rect 13872 7760 13878 7812
rect 13998 7800 14004 7812
rect 13959 7772 14004 7800
rect 13998 7760 14004 7772
rect 14056 7760 14062 7812
rect 14108 7732 14136 7908
rect 14461 7905 14473 7908
rect 14507 7905 14519 7939
rect 14461 7899 14519 7905
rect 14274 7828 14280 7880
rect 14332 7868 14338 7880
rect 14553 7871 14611 7877
rect 14553 7868 14565 7871
rect 14332 7840 14565 7868
rect 14332 7828 14338 7840
rect 14553 7837 14565 7840
rect 14599 7837 14611 7871
rect 14553 7831 14611 7837
rect 13096 7704 14136 7732
rect 12989 7695 13047 7701
rect 1104 7642 15824 7664
rect 1104 7590 3447 7642
rect 3499 7590 3511 7642
rect 3563 7590 3575 7642
rect 3627 7590 3639 7642
rect 3691 7590 8378 7642
rect 8430 7590 8442 7642
rect 8494 7590 8506 7642
rect 8558 7590 8570 7642
rect 8622 7590 13308 7642
rect 13360 7590 13372 7642
rect 13424 7590 13436 7642
rect 13488 7590 13500 7642
rect 13552 7590 15824 7642
rect 1104 7568 15824 7590
rect 3237 7531 3295 7537
rect 3237 7497 3249 7531
rect 3283 7528 3295 7531
rect 5810 7528 5816 7540
rect 3283 7500 5816 7528
rect 3283 7497 3295 7500
rect 3237 7491 3295 7497
rect 5810 7488 5816 7500
rect 5868 7528 5874 7540
rect 8205 7531 8263 7537
rect 8205 7528 8217 7531
rect 5868 7500 8217 7528
rect 5868 7488 5874 7500
rect 8205 7497 8217 7500
rect 8251 7497 8263 7531
rect 9214 7528 9220 7540
rect 8205 7491 8263 7497
rect 8496 7500 9220 7528
rect 4798 7460 4804 7472
rect 4759 7432 4804 7460
rect 4798 7420 4804 7432
rect 4856 7420 4862 7472
rect 8018 7420 8024 7472
rect 8076 7460 8082 7472
rect 8496 7460 8524 7500
rect 9214 7488 9220 7500
rect 9272 7488 9278 7540
rect 9861 7531 9919 7537
rect 9861 7497 9873 7531
rect 9907 7528 9919 7531
rect 12161 7531 12219 7537
rect 12161 7528 12173 7531
rect 9907 7500 12173 7528
rect 9907 7497 9919 7500
rect 9861 7491 9919 7497
rect 12161 7497 12173 7500
rect 12207 7497 12219 7531
rect 13265 7531 13323 7537
rect 13265 7528 13277 7531
rect 12161 7491 12219 7497
rect 12360 7500 13277 7528
rect 8076 7432 8524 7460
rect 8076 7420 8082 7432
rect 2041 7395 2099 7401
rect 2041 7361 2053 7395
rect 2087 7392 2099 7395
rect 3053 7395 3111 7401
rect 2087 7364 3004 7392
rect 2087 7361 2099 7364
rect 2041 7355 2099 7361
rect 1765 7327 1823 7333
rect 1765 7293 1777 7327
rect 1811 7324 1823 7327
rect 2222 7324 2228 7336
rect 1811 7296 2228 7324
rect 1811 7293 1823 7296
rect 1765 7287 1823 7293
rect 2222 7284 2228 7296
rect 2280 7324 2286 7336
rect 2774 7324 2780 7336
rect 2280 7296 2780 7324
rect 2280 7284 2286 7296
rect 2774 7284 2780 7296
rect 2832 7284 2838 7336
rect 2869 7259 2927 7265
rect 2869 7256 2881 7259
rect 1412 7228 2881 7256
rect 1412 7197 1440 7228
rect 2869 7225 2881 7228
rect 2915 7225 2927 7259
rect 2976 7256 3004 7364
rect 3053 7361 3065 7395
rect 3099 7392 3111 7395
rect 3237 7395 3295 7401
rect 3237 7392 3249 7395
rect 3099 7364 3249 7392
rect 3099 7361 3111 7364
rect 3053 7355 3111 7361
rect 3237 7361 3249 7364
rect 3283 7361 3295 7395
rect 3237 7355 3295 7361
rect 4614 7352 4620 7404
rect 4672 7392 4678 7404
rect 5077 7395 5135 7401
rect 5077 7392 5089 7395
rect 4672 7364 5089 7392
rect 4672 7352 4678 7364
rect 5077 7361 5089 7364
rect 5123 7361 5135 7395
rect 5077 7355 5135 7361
rect 6086 7352 6092 7404
rect 6144 7392 6150 7404
rect 6144 7364 6951 7392
rect 6144 7352 6150 7364
rect 3326 7284 3332 7336
rect 3384 7324 3390 7336
rect 3421 7327 3479 7333
rect 3421 7324 3433 7327
rect 3384 7296 3433 7324
rect 3384 7284 3390 7296
rect 3421 7293 3433 7296
rect 3467 7293 3479 7327
rect 3421 7287 3479 7293
rect 3685 7284 3691 7336
rect 3743 7324 3749 7336
rect 6822 7324 6828 7336
rect 3743 7296 3788 7324
rect 6783 7296 6828 7324
rect 3743 7284 3749 7296
rect 6822 7284 6828 7296
rect 6880 7284 6886 7336
rect 6923 7324 6951 7364
rect 7926 7352 7932 7404
rect 7984 7392 7990 7404
rect 8481 7395 8539 7401
rect 8481 7392 8493 7395
rect 7984 7364 8493 7392
rect 7984 7352 7990 7364
rect 8481 7361 8493 7364
rect 8527 7361 8539 7395
rect 8481 7355 8539 7361
rect 9876 7324 9904 7491
rect 11330 7420 11336 7472
rect 11388 7460 11394 7472
rect 11977 7463 12035 7469
rect 11977 7460 11989 7463
rect 11388 7432 11989 7460
rect 11388 7420 11394 7432
rect 11977 7429 11989 7432
rect 12023 7429 12035 7463
rect 11977 7423 12035 7429
rect 12066 7420 12072 7472
rect 12124 7460 12130 7472
rect 12360 7460 12388 7500
rect 13265 7497 13277 7500
rect 13311 7497 13323 7531
rect 13265 7491 13323 7497
rect 13998 7488 14004 7540
rect 14056 7528 14062 7540
rect 14369 7531 14427 7537
rect 14369 7528 14381 7531
rect 14056 7500 14381 7528
rect 14056 7488 14062 7500
rect 14369 7497 14381 7500
rect 14415 7497 14427 7531
rect 14369 7491 14427 7497
rect 12124 7432 12388 7460
rect 12437 7463 12495 7469
rect 12124 7420 12130 7432
rect 12437 7429 12449 7463
rect 12483 7460 12495 7463
rect 12526 7460 12532 7472
rect 12483 7432 12532 7460
rect 12483 7429 12495 7432
rect 12437 7423 12495 7429
rect 12526 7420 12532 7432
rect 12584 7420 12590 7472
rect 14090 7460 14096 7472
rect 13924 7432 14096 7460
rect 10134 7392 10140 7404
rect 10095 7364 10140 7392
rect 10134 7352 10140 7364
rect 10192 7352 10198 7404
rect 11422 7352 11428 7404
rect 11480 7392 11486 7404
rect 12342 7392 12348 7404
rect 11480 7364 12348 7392
rect 11480 7352 11486 7364
rect 12342 7352 12348 7364
rect 12400 7392 12406 7404
rect 12989 7395 13047 7401
rect 12989 7392 13001 7395
rect 12400 7364 13001 7392
rect 12400 7352 12406 7364
rect 12989 7361 13001 7364
rect 13035 7361 13047 7395
rect 12989 7355 13047 7361
rect 13078 7352 13084 7404
rect 13136 7392 13142 7404
rect 13924 7401 13952 7432
rect 14090 7420 14096 7432
rect 14148 7460 14154 7472
rect 14458 7460 14464 7472
rect 14148 7432 14464 7460
rect 14148 7420 14154 7432
rect 14458 7420 14464 7432
rect 14516 7420 14522 7472
rect 13909 7395 13967 7401
rect 13136 7364 13860 7392
rect 13136 7352 13142 7364
rect 6923 7296 9904 7324
rect 10404 7327 10462 7333
rect 10404 7293 10416 7327
rect 10450 7324 10462 7327
rect 10962 7324 10968 7336
rect 10450 7296 10968 7324
rect 10450 7293 10462 7296
rect 10404 7287 10462 7293
rect 10962 7284 10968 7296
rect 11020 7284 11026 7336
rect 11793 7327 11851 7333
rect 11793 7324 11805 7327
rect 11256 7296 11805 7324
rect 4706 7256 4712 7268
rect 2976 7228 4712 7256
rect 2869 7219 2927 7225
rect 4706 7216 4712 7228
rect 4764 7216 4770 7268
rect 5344 7259 5402 7265
rect 5344 7256 5356 7259
rect 5092 7228 5356 7256
rect 5092 7200 5120 7228
rect 5344 7225 5356 7228
rect 5390 7256 5402 7259
rect 6086 7256 6092 7268
rect 5390 7228 6092 7256
rect 5390 7225 5402 7228
rect 5344 7219 5402 7225
rect 6086 7216 6092 7228
rect 6144 7216 6150 7268
rect 6362 7216 6368 7268
rect 6420 7256 6426 7268
rect 7070 7259 7128 7265
rect 7070 7256 7082 7259
rect 6420 7228 7082 7256
rect 6420 7216 6426 7228
rect 7070 7225 7082 7228
rect 7116 7256 7128 7259
rect 7466 7256 7472 7268
rect 7116 7228 7472 7256
rect 7116 7225 7128 7228
rect 7070 7219 7128 7225
rect 7466 7216 7472 7228
rect 7524 7216 7530 7268
rect 7558 7216 7564 7268
rect 7616 7256 7622 7268
rect 8570 7256 8576 7268
rect 7616 7228 8576 7256
rect 7616 7216 7622 7228
rect 8570 7216 8576 7228
rect 8628 7216 8634 7268
rect 8748 7259 8806 7265
rect 8748 7225 8760 7259
rect 8794 7256 8806 7259
rect 8938 7256 8944 7268
rect 8794 7228 8944 7256
rect 8794 7225 8806 7228
rect 8748 7219 8806 7225
rect 8938 7216 8944 7228
rect 8996 7216 9002 7268
rect 11146 7256 11152 7268
rect 9048 7228 11152 7256
rect 1397 7191 1455 7197
rect 1397 7157 1409 7191
rect 1443 7157 1455 7191
rect 1854 7188 1860 7200
rect 1815 7160 1860 7188
rect 1397 7151 1455 7157
rect 1854 7148 1860 7160
rect 1912 7148 1918 7200
rect 2406 7188 2412 7200
rect 2367 7160 2412 7188
rect 2406 7148 2412 7160
rect 2464 7148 2470 7200
rect 2777 7191 2835 7197
rect 2777 7157 2789 7191
rect 2823 7188 2835 7191
rect 4614 7188 4620 7200
rect 2823 7160 4620 7188
rect 2823 7157 2835 7160
rect 2777 7151 2835 7157
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 5074 7148 5080 7200
rect 5132 7148 5138 7200
rect 5718 7148 5724 7200
rect 5776 7188 5782 7200
rect 6457 7191 6515 7197
rect 6457 7188 6469 7191
rect 5776 7160 6469 7188
rect 5776 7148 5782 7160
rect 6457 7157 6469 7160
rect 6503 7188 6515 7191
rect 7282 7188 7288 7200
rect 6503 7160 7288 7188
rect 6503 7157 6515 7160
rect 6457 7151 6515 7157
rect 7282 7148 7288 7160
rect 7340 7148 7346 7200
rect 8662 7148 8668 7200
rect 8720 7188 8726 7200
rect 9048 7188 9076 7228
rect 11146 7216 11152 7228
rect 11204 7216 11210 7268
rect 8720 7160 9076 7188
rect 8720 7148 8726 7160
rect 10318 7148 10324 7200
rect 10376 7188 10382 7200
rect 11256 7188 11284 7296
rect 11793 7293 11805 7296
rect 11839 7293 11851 7327
rect 12618 7324 12624 7336
rect 11793 7287 11851 7293
rect 11900 7296 12624 7324
rect 11422 7216 11428 7268
rect 11480 7256 11486 7268
rect 11900 7256 11928 7296
rect 12618 7284 12624 7296
rect 12676 7284 12682 7336
rect 13265 7327 13323 7333
rect 13265 7293 13277 7327
rect 13311 7324 13323 7327
rect 13832 7324 13860 7364
rect 13909 7361 13921 7395
rect 13955 7361 13967 7395
rect 13909 7355 13967 7361
rect 14001 7395 14059 7401
rect 14001 7361 14013 7395
rect 14047 7392 14059 7395
rect 14274 7392 14280 7404
rect 14047 7364 14280 7392
rect 14047 7361 14059 7364
rect 14001 7355 14059 7361
rect 14016 7324 14044 7355
rect 14274 7352 14280 7364
rect 14332 7352 14338 7404
rect 15010 7392 15016 7404
rect 14971 7364 15016 7392
rect 15010 7352 15016 7364
rect 15068 7352 15074 7404
rect 14550 7324 14556 7336
rect 13311 7296 13768 7324
rect 13832 7296 14044 7324
rect 14200 7296 14556 7324
rect 13311 7293 13323 7296
rect 13265 7287 13323 7293
rect 11480 7228 11928 7256
rect 12161 7259 12219 7265
rect 11480 7216 11486 7228
rect 12161 7225 12173 7259
rect 12207 7225 12219 7259
rect 12161 7219 12219 7225
rect 10376 7160 11284 7188
rect 10376 7148 10382 7160
rect 11330 7148 11336 7200
rect 11388 7188 11394 7200
rect 11517 7191 11575 7197
rect 11517 7188 11529 7191
rect 11388 7160 11529 7188
rect 11388 7148 11394 7160
rect 11517 7157 11529 7160
rect 11563 7157 11575 7191
rect 12176 7188 12204 7219
rect 12342 7216 12348 7268
rect 12400 7256 12406 7268
rect 12805 7259 12863 7265
rect 12805 7256 12817 7259
rect 12400 7228 12817 7256
rect 12400 7216 12406 7228
rect 12805 7225 12817 7228
rect 12851 7256 12863 7259
rect 13354 7256 13360 7268
rect 12851 7228 13360 7256
rect 12851 7225 12863 7228
rect 12805 7219 12863 7225
rect 13354 7216 13360 7228
rect 13412 7216 13418 7268
rect 13740 7256 13768 7296
rect 14090 7256 14096 7268
rect 13740 7228 14096 7256
rect 14090 7216 14096 7228
rect 14148 7216 14154 7268
rect 12618 7188 12624 7200
rect 12176 7160 12624 7188
rect 11517 7151 11575 7157
rect 12618 7148 12624 7160
rect 12676 7148 12682 7200
rect 12894 7188 12900 7200
rect 12855 7160 12900 7188
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 13446 7188 13452 7200
rect 13407 7160 13452 7188
rect 13446 7148 13452 7160
rect 13504 7148 13510 7200
rect 13817 7191 13875 7197
rect 13817 7157 13829 7191
rect 13863 7188 13875 7191
rect 14200 7188 14228 7296
rect 14550 7284 14556 7296
rect 14608 7324 14614 7336
rect 15102 7324 15108 7336
rect 14608 7296 15108 7324
rect 14608 7284 14614 7296
rect 15102 7284 15108 7296
rect 15160 7284 15166 7336
rect 14274 7216 14280 7268
rect 14332 7256 14338 7268
rect 14921 7259 14979 7265
rect 14921 7256 14933 7259
rect 14332 7228 14933 7256
rect 14332 7216 14338 7228
rect 14921 7225 14933 7228
rect 14967 7225 14979 7259
rect 14921 7219 14979 7225
rect 13863 7160 14228 7188
rect 14369 7191 14427 7197
rect 13863 7157 13875 7160
rect 13817 7151 13875 7157
rect 14369 7157 14381 7191
rect 14415 7188 14427 7191
rect 14461 7191 14519 7197
rect 14461 7188 14473 7191
rect 14415 7160 14473 7188
rect 14415 7157 14427 7160
rect 14369 7151 14427 7157
rect 14461 7157 14473 7160
rect 14507 7157 14519 7191
rect 14826 7188 14832 7200
rect 14787 7160 14832 7188
rect 14461 7151 14519 7157
rect 14826 7148 14832 7160
rect 14884 7148 14890 7200
rect 1104 7098 15824 7120
rect 1104 7046 5912 7098
rect 5964 7046 5976 7098
rect 6028 7046 6040 7098
rect 6092 7046 6104 7098
rect 6156 7046 10843 7098
rect 10895 7046 10907 7098
rect 10959 7046 10971 7098
rect 11023 7046 11035 7098
rect 11087 7046 15824 7098
rect 1104 7024 15824 7046
rect 2406 6944 2412 6996
rect 2464 6984 2470 6996
rect 4985 6987 5043 6993
rect 4985 6984 4997 6987
rect 2464 6956 4997 6984
rect 2464 6944 2470 6956
rect 4985 6953 4997 6956
rect 5031 6953 5043 6987
rect 4985 6947 5043 6953
rect 5353 6987 5411 6993
rect 5353 6953 5365 6987
rect 5399 6984 5411 6987
rect 8846 6984 8852 6996
rect 5399 6956 8852 6984
rect 5399 6953 5411 6956
rect 5353 6947 5411 6953
rect 8846 6944 8852 6956
rect 8904 6944 8910 6996
rect 9030 6984 9036 6996
rect 8991 6956 9036 6984
rect 9030 6944 9036 6956
rect 9088 6944 9094 6996
rect 9493 6987 9551 6993
rect 9493 6953 9505 6987
rect 9539 6984 9551 6987
rect 10134 6984 10140 6996
rect 9539 6956 10140 6984
rect 9539 6953 9551 6956
rect 9493 6947 9551 6953
rect 10134 6944 10140 6956
rect 10192 6944 10198 6996
rect 11330 6944 11336 6996
rect 11388 6984 11394 6996
rect 11701 6987 11759 6993
rect 11388 6956 11433 6984
rect 11388 6944 11394 6956
rect 11701 6953 11713 6987
rect 11747 6984 11759 6987
rect 11882 6984 11888 6996
rect 11747 6956 11888 6984
rect 11747 6953 11759 6956
rect 11701 6947 11759 6953
rect 11882 6944 11888 6956
rect 11940 6984 11946 6996
rect 12342 6984 12348 6996
rect 11940 6956 12348 6984
rect 11940 6944 11946 6956
rect 12342 6944 12348 6956
rect 12400 6944 12406 6996
rect 12894 6944 12900 6996
rect 12952 6984 12958 6996
rect 13725 6987 13783 6993
rect 13725 6984 13737 6987
rect 12952 6956 13737 6984
rect 12952 6944 12958 6956
rect 13725 6953 13737 6956
rect 13771 6953 13783 6987
rect 13725 6947 13783 6953
rect 13817 6987 13875 6993
rect 13817 6953 13829 6987
rect 13863 6984 13875 6987
rect 14090 6984 14096 6996
rect 13863 6956 14096 6984
rect 13863 6953 13875 6956
rect 13817 6947 13875 6953
rect 14090 6944 14096 6956
rect 14148 6944 14154 6996
rect 14921 6987 14979 6993
rect 14921 6953 14933 6987
rect 14967 6953 14979 6987
rect 14921 6947 14979 6953
rect 2498 6876 2504 6928
rect 2556 6925 2562 6928
rect 2556 6919 2620 6925
rect 2556 6885 2574 6919
rect 2608 6885 2620 6919
rect 2556 6879 2620 6885
rect 4893 6919 4951 6925
rect 4893 6885 4905 6919
rect 4939 6916 4951 6919
rect 5626 6916 5632 6928
rect 4939 6888 5632 6916
rect 4939 6885 4951 6888
rect 4893 6879 4951 6885
rect 2556 6876 2562 6879
rect 5626 6876 5632 6888
rect 5684 6876 5690 6928
rect 6822 6916 6828 6928
rect 5736 6888 6828 6916
rect 1581 6851 1639 6857
rect 1581 6817 1593 6851
rect 1627 6848 1639 6851
rect 1946 6848 1952 6860
rect 1627 6820 1952 6848
rect 1627 6817 1639 6820
rect 1581 6811 1639 6817
rect 1946 6808 1952 6820
rect 2004 6808 2010 6860
rect 2314 6848 2320 6860
rect 2275 6820 2320 6848
rect 2314 6808 2320 6820
rect 2372 6808 2378 6860
rect 4798 6808 4804 6860
rect 4856 6848 4862 6860
rect 5353 6851 5411 6857
rect 5353 6848 5365 6851
rect 4856 6820 5365 6848
rect 4856 6808 4862 6820
rect 5353 6817 5365 6820
rect 5399 6817 5411 6851
rect 5353 6811 5411 6817
rect 5537 6851 5595 6857
rect 5537 6817 5549 6851
rect 5583 6848 5595 6851
rect 5736 6848 5764 6888
rect 6822 6876 6828 6888
rect 6880 6876 6886 6928
rect 7006 6876 7012 6928
rect 7064 6916 7070 6928
rect 7064 6888 8524 6916
rect 7064 6876 7070 6888
rect 5810 6857 5816 6860
rect 5583 6820 5764 6848
rect 5583 6817 5595 6820
rect 5537 6811 5595 6817
rect 5804 6811 5816 6857
rect 5868 6848 5874 6860
rect 7190 6848 7196 6860
rect 5868 6820 5904 6848
rect 7151 6820 7196 6848
rect 5810 6808 5816 6811
rect 5868 6808 5874 6820
rect 7190 6808 7196 6820
rect 7248 6808 7254 6860
rect 7282 6808 7288 6860
rect 7340 6848 7346 6860
rect 7449 6851 7507 6857
rect 7449 6848 7461 6851
rect 7340 6820 7461 6848
rect 7340 6808 7346 6820
rect 7449 6817 7461 6820
rect 7495 6817 7507 6851
rect 7449 6811 7507 6817
rect 7742 6808 7748 6860
rect 7800 6848 7806 6860
rect 8496 6848 8524 6888
rect 9306 6876 9312 6928
rect 9364 6916 9370 6928
rect 11790 6916 11796 6928
rect 9364 6888 10088 6916
rect 9364 6876 9370 6888
rect 8938 6848 8944 6860
rect 7800 6820 8239 6848
rect 8496 6820 8944 6848
rect 7800 6808 7806 6820
rect 1762 6780 1768 6792
rect 1723 6752 1768 6780
rect 1762 6740 1768 6752
rect 1820 6740 1826 6792
rect 4062 6780 4068 6792
rect 4023 6752 4068 6780
rect 4062 6740 4068 6752
rect 4120 6740 4126 6792
rect 5166 6780 5172 6792
rect 5079 6752 5172 6780
rect 5166 6740 5172 6752
rect 5224 6780 5230 6792
rect 8211 6780 8239 6820
rect 8938 6808 8944 6820
rect 8996 6848 9002 6860
rect 9950 6857 9956 6860
rect 9125 6851 9183 6857
rect 9125 6848 9137 6851
rect 8996 6820 9137 6848
rect 8996 6808 9002 6820
rect 9125 6817 9137 6820
rect 9171 6817 9183 6851
rect 9125 6811 9183 6817
rect 9493 6851 9551 6857
rect 9493 6817 9505 6851
rect 9539 6848 9551 6851
rect 9677 6851 9735 6857
rect 9677 6848 9689 6851
rect 9539 6820 9689 6848
rect 9539 6817 9551 6820
rect 9493 6811 9551 6817
rect 9677 6817 9689 6820
rect 9723 6817 9735 6851
rect 9944 6848 9956 6857
rect 9911 6820 9956 6848
rect 9677 6811 9735 6817
rect 9944 6811 9956 6820
rect 9950 6808 9956 6811
rect 10008 6808 10014 6860
rect 10060 6848 10088 6888
rect 10419 6888 11796 6916
rect 10419 6848 10447 6888
rect 11790 6876 11796 6888
rect 11848 6876 11854 6928
rect 12158 6876 12164 6928
rect 12216 6916 12222 6928
rect 12713 6919 12771 6925
rect 12713 6916 12725 6919
rect 12216 6888 12725 6916
rect 12216 6876 12222 6888
rect 12713 6885 12725 6888
rect 12759 6916 12771 6919
rect 13906 6916 13912 6928
rect 12759 6888 13912 6916
rect 12759 6885 12771 6888
rect 12713 6879 12771 6885
rect 13906 6876 13912 6888
rect 13964 6876 13970 6928
rect 14936 6916 14964 6947
rect 14016 6888 14964 6916
rect 10060 6820 10447 6848
rect 10778 6808 10784 6860
rect 10836 6848 10842 6860
rect 10836 6820 11928 6848
rect 10836 6808 10842 6820
rect 9217 6783 9275 6789
rect 9217 6780 9229 6783
rect 5224 6752 5488 6780
rect 8211 6752 9229 6780
rect 5224 6740 5230 6752
rect 3697 6647 3755 6653
rect 3697 6613 3709 6647
rect 3743 6644 3755 6647
rect 3878 6644 3884 6656
rect 3743 6616 3884 6644
rect 3743 6613 3755 6616
rect 3697 6607 3755 6613
rect 3878 6604 3884 6616
rect 3936 6604 3942 6656
rect 3970 6604 3976 6656
rect 4028 6644 4034 6656
rect 4525 6647 4583 6653
rect 4525 6644 4537 6647
rect 4028 6616 4537 6644
rect 4028 6604 4034 6616
rect 4525 6613 4537 6616
rect 4571 6613 4583 6647
rect 5460 6644 5488 6752
rect 9217 6749 9229 6752
rect 9263 6749 9275 6783
rect 9217 6743 9275 6749
rect 10686 6740 10692 6792
rect 10744 6780 10750 6792
rect 11422 6780 11428 6792
rect 10744 6752 11428 6780
rect 10744 6740 10750 6752
rect 11422 6740 11428 6752
rect 11480 6740 11486 6792
rect 11900 6789 11928 6820
rect 12342 6808 12348 6860
rect 12400 6848 12406 6860
rect 12805 6851 12863 6857
rect 12805 6848 12817 6851
rect 12400 6820 12817 6848
rect 12400 6808 12406 6820
rect 12805 6817 12817 6820
rect 12851 6848 12863 6851
rect 13078 6848 13084 6860
rect 12851 6820 13084 6848
rect 12851 6817 12863 6820
rect 12805 6811 12863 6817
rect 13078 6808 13084 6820
rect 13136 6808 13142 6860
rect 13170 6808 13176 6860
rect 13228 6848 13234 6860
rect 14016 6848 14044 6888
rect 13228 6820 14044 6848
rect 13228 6808 13234 6820
rect 14182 6808 14188 6860
rect 14240 6848 14246 6860
rect 14369 6851 14427 6857
rect 14369 6848 14381 6851
rect 14240 6820 14381 6848
rect 14240 6808 14246 6820
rect 14369 6817 14381 6820
rect 14415 6848 14427 6851
rect 14458 6848 14464 6860
rect 14415 6820 14464 6848
rect 14415 6817 14427 6820
rect 14369 6811 14427 6817
rect 14458 6808 14464 6820
rect 14516 6808 14522 6860
rect 15105 6851 15163 6857
rect 15105 6817 15117 6851
rect 15151 6848 15163 6851
rect 15194 6848 15200 6860
rect 15151 6820 15200 6848
rect 15151 6817 15163 6820
rect 15105 6811 15163 6817
rect 15194 6808 15200 6820
rect 15252 6808 15258 6860
rect 11885 6783 11943 6789
rect 11885 6749 11897 6783
rect 11931 6749 11943 6783
rect 11885 6743 11943 6749
rect 11974 6740 11980 6792
rect 12032 6780 12038 6792
rect 12710 6780 12716 6792
rect 12032 6752 12716 6780
rect 12032 6740 12038 6752
rect 12710 6740 12716 6752
rect 12768 6740 12774 6792
rect 12894 6780 12900 6792
rect 12855 6752 12900 6780
rect 12894 6740 12900 6752
rect 12952 6740 12958 6792
rect 13909 6783 13967 6789
rect 13909 6780 13921 6783
rect 13004 6752 13921 6780
rect 6638 6672 6644 6724
rect 6696 6712 6702 6724
rect 6696 6684 7144 6712
rect 6696 6672 6702 6684
rect 6917 6647 6975 6653
rect 6917 6644 6929 6647
rect 5460 6616 6929 6644
rect 4525 6607 4583 6613
rect 6917 6613 6929 6616
rect 6963 6613 6975 6647
rect 7116 6644 7144 6684
rect 8202 6672 8208 6724
rect 8260 6712 8266 6724
rect 8665 6715 8723 6721
rect 8665 6712 8677 6715
rect 8260 6684 8677 6712
rect 8260 6672 8266 6684
rect 8665 6681 8677 6684
rect 8711 6681 8723 6715
rect 12345 6715 12403 6721
rect 12345 6712 12357 6715
rect 8665 6675 8723 6681
rect 10980 6684 12357 6712
rect 8573 6647 8631 6653
rect 8573 6644 8585 6647
rect 7116 6616 8585 6644
rect 6917 6607 6975 6613
rect 8573 6613 8585 6616
rect 8619 6613 8631 6647
rect 8573 6607 8631 6613
rect 9858 6604 9864 6656
rect 9916 6644 9922 6656
rect 10980 6644 11008 6684
rect 12345 6681 12357 6684
rect 12391 6681 12403 6715
rect 13004 6712 13032 6752
rect 13909 6749 13921 6752
rect 13955 6780 13967 6783
rect 15010 6780 15016 6792
rect 13955 6752 15016 6780
rect 13955 6749 13967 6752
rect 13909 6743 13967 6749
rect 15010 6740 15016 6752
rect 15068 6740 15074 6792
rect 12345 6675 12403 6681
rect 12452 6684 13032 6712
rect 9916 6616 11008 6644
rect 11057 6647 11115 6653
rect 9916 6604 9922 6616
rect 11057 6613 11069 6647
rect 11103 6644 11115 6647
rect 11698 6644 11704 6656
rect 11103 6616 11704 6644
rect 11103 6613 11115 6616
rect 11057 6607 11115 6613
rect 11698 6604 11704 6616
rect 11756 6604 11762 6656
rect 11882 6604 11888 6656
rect 11940 6644 11946 6656
rect 12452 6644 12480 6684
rect 13170 6672 13176 6724
rect 13228 6712 13234 6724
rect 13357 6715 13415 6721
rect 13357 6712 13369 6715
rect 13228 6684 13369 6712
rect 13228 6672 13234 6684
rect 13357 6681 13369 6684
rect 13403 6681 13415 6715
rect 13357 6675 13415 6681
rect 13446 6672 13452 6724
rect 13504 6672 13510 6724
rect 11940 6616 12480 6644
rect 11940 6604 11946 6616
rect 12710 6604 12716 6656
rect 12768 6644 12774 6656
rect 13464 6644 13492 6672
rect 12768 6616 13492 6644
rect 12768 6604 12774 6616
rect 14182 6604 14188 6656
rect 14240 6644 14246 6656
rect 14553 6647 14611 6653
rect 14553 6644 14565 6647
rect 14240 6616 14565 6644
rect 14240 6604 14246 6616
rect 14553 6613 14565 6616
rect 14599 6613 14611 6647
rect 14553 6607 14611 6613
rect 1104 6554 15824 6576
rect 1104 6502 3447 6554
rect 3499 6502 3511 6554
rect 3563 6502 3575 6554
rect 3627 6502 3639 6554
rect 3691 6502 8378 6554
rect 8430 6502 8442 6554
rect 8494 6502 8506 6554
rect 8558 6502 8570 6554
rect 8622 6502 13308 6554
rect 13360 6502 13372 6554
rect 13424 6502 13436 6554
rect 13488 6502 13500 6554
rect 13552 6502 15824 6554
rect 1104 6480 15824 6502
rect 2409 6443 2467 6449
rect 2409 6409 2421 6443
rect 2455 6440 2467 6443
rect 4154 6440 4160 6452
rect 2455 6412 4160 6440
rect 2455 6409 2467 6412
rect 2409 6403 2467 6409
rect 4154 6400 4160 6412
rect 4212 6400 4218 6452
rect 5350 6440 5356 6452
rect 5092 6412 5356 6440
rect 4522 6332 4528 6384
rect 4580 6372 4586 6384
rect 4801 6375 4859 6381
rect 4801 6372 4813 6375
rect 4580 6344 4813 6372
rect 4580 6332 4586 6344
rect 4801 6341 4813 6344
rect 4847 6372 4859 6375
rect 4985 6375 5043 6381
rect 4985 6372 4997 6375
rect 4847 6344 4997 6372
rect 4847 6341 4859 6344
rect 4801 6335 4859 6341
rect 4985 6341 4997 6344
rect 5031 6341 5043 6375
rect 4985 6335 5043 6341
rect 2041 6307 2099 6313
rect 2041 6273 2053 6307
rect 2087 6304 2099 6307
rect 2682 6304 2688 6316
rect 2087 6276 2688 6304
rect 2087 6273 2099 6276
rect 2041 6267 2099 6273
rect 2682 6264 2688 6276
rect 2740 6264 2746 6316
rect 2961 6307 3019 6313
rect 2961 6273 2973 6307
rect 3007 6304 3019 6307
rect 3007 6276 3280 6304
rect 3007 6273 3019 6276
rect 2961 6267 3019 6273
rect 2869 6239 2927 6245
rect 2869 6205 2881 6239
rect 2915 6236 2927 6239
rect 3050 6236 3056 6248
rect 2915 6208 3056 6236
rect 2915 6205 2927 6208
rect 2869 6199 2927 6205
rect 3050 6196 3056 6208
rect 3108 6196 3114 6248
rect 3252 6236 3280 6276
rect 3326 6264 3332 6316
rect 3384 6304 3390 6316
rect 3421 6307 3479 6313
rect 3421 6304 3433 6307
rect 3384 6276 3433 6304
rect 3384 6264 3390 6276
rect 3421 6273 3433 6276
rect 3467 6273 3479 6307
rect 5092 6304 5120 6412
rect 5350 6400 5356 6412
rect 5408 6400 5414 6452
rect 5442 6400 5448 6452
rect 5500 6440 5506 6452
rect 9858 6440 9864 6452
rect 5500 6412 9864 6440
rect 5500 6400 5506 6412
rect 9858 6400 9864 6412
rect 9916 6400 9922 6452
rect 9953 6443 10011 6449
rect 9953 6409 9965 6443
rect 9999 6440 10011 6443
rect 10042 6440 10048 6452
rect 9999 6412 10048 6440
rect 9999 6409 10011 6412
rect 9953 6403 10011 6409
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 10137 6443 10195 6449
rect 10137 6409 10149 6443
rect 10183 6440 10195 6443
rect 11330 6440 11336 6452
rect 10183 6412 11336 6440
rect 10183 6409 10195 6412
rect 10137 6403 10195 6409
rect 11330 6400 11336 6412
rect 11388 6400 11394 6452
rect 12710 6440 12716 6452
rect 11440 6412 12716 6440
rect 11238 6332 11244 6384
rect 11296 6372 11302 6384
rect 11440 6372 11468 6412
rect 12710 6400 12716 6412
rect 12768 6400 12774 6452
rect 13449 6443 13507 6449
rect 13449 6409 13461 6443
rect 13495 6440 13507 6443
rect 13630 6440 13636 6452
rect 13495 6412 13636 6440
rect 13495 6409 13507 6412
rect 13449 6403 13507 6409
rect 13630 6400 13636 6412
rect 13688 6400 13694 6452
rect 14461 6443 14519 6449
rect 14461 6409 14473 6443
rect 14507 6440 14519 6443
rect 14918 6440 14924 6452
rect 14507 6412 14924 6440
rect 14507 6409 14519 6412
rect 14461 6403 14519 6409
rect 14918 6400 14924 6412
rect 14976 6400 14982 6452
rect 11296 6344 11468 6372
rect 11609 6375 11667 6381
rect 11296 6332 11302 6344
rect 11609 6341 11621 6375
rect 11655 6372 11667 6375
rect 12161 6375 12219 6381
rect 12161 6372 12173 6375
rect 11655 6344 12173 6372
rect 11655 6341 11667 6344
rect 11609 6335 11667 6341
rect 12161 6341 12173 6344
rect 12207 6341 12219 6375
rect 12161 6335 12219 6341
rect 12342 6332 12348 6384
rect 12400 6372 12406 6384
rect 12894 6372 12900 6384
rect 12400 6344 12900 6372
rect 12400 6332 12406 6344
rect 12894 6332 12900 6344
rect 12952 6332 12958 6384
rect 13265 6375 13323 6381
rect 13265 6341 13277 6375
rect 13311 6372 13323 6375
rect 13311 6344 14044 6372
rect 13311 6341 13323 6344
rect 13265 6335 13323 6341
rect 6270 6304 6276 6316
rect 5092 6276 5212 6304
rect 3421 6267 3479 6273
rect 4430 6236 4436 6248
rect 3252 6208 4436 6236
rect 4430 6196 4436 6208
rect 4488 6196 4494 6248
rect 4706 6196 4712 6248
rect 4764 6236 4770 6248
rect 5077 6239 5135 6245
rect 5077 6236 5089 6239
rect 4764 6208 5089 6236
rect 4764 6196 4770 6208
rect 5077 6205 5089 6208
rect 5123 6205 5135 6239
rect 5184 6236 5212 6276
rect 6104 6276 6276 6304
rect 5333 6239 5391 6245
rect 5333 6236 5345 6239
rect 5184 6208 5345 6236
rect 5077 6199 5135 6205
rect 5333 6205 5345 6208
rect 5379 6205 5391 6239
rect 5333 6199 5391 6205
rect 5718 6196 5724 6248
rect 5776 6236 5782 6248
rect 6104 6236 6132 6276
rect 6270 6264 6276 6276
rect 6328 6264 6334 6316
rect 6822 6264 6828 6316
rect 6880 6304 6886 6316
rect 6917 6307 6975 6313
rect 6917 6304 6929 6307
rect 6880 6276 6929 6304
rect 6880 6264 6886 6276
rect 6917 6273 6929 6276
rect 6963 6273 6975 6307
rect 6917 6267 6975 6273
rect 7926 6264 7932 6316
rect 7984 6304 7990 6316
rect 8294 6304 8300 6316
rect 7984 6276 8300 6304
rect 7984 6264 7990 6276
rect 8294 6264 8300 6276
rect 8352 6304 8358 6316
rect 8573 6307 8631 6313
rect 8573 6304 8585 6307
rect 8352 6276 8585 6304
rect 8352 6264 8358 6276
rect 8573 6273 8585 6276
rect 8619 6273 8631 6307
rect 8573 6267 8631 6273
rect 10134 6264 10140 6316
rect 10192 6304 10198 6316
rect 10229 6307 10287 6313
rect 10229 6304 10241 6307
rect 10192 6276 10241 6304
rect 10192 6264 10198 6276
rect 10229 6273 10241 6276
rect 10275 6273 10287 6307
rect 10229 6267 10287 6273
rect 11698 6264 11704 6316
rect 11756 6304 11762 6316
rect 12989 6307 13047 6313
rect 12989 6304 13001 6307
rect 11756 6276 13001 6304
rect 11756 6264 11762 6276
rect 12989 6273 13001 6276
rect 13035 6273 13047 6307
rect 12989 6267 13047 6273
rect 13078 6264 13084 6316
rect 13136 6304 13142 6316
rect 14016 6313 14044 6344
rect 14734 6332 14740 6384
rect 14792 6372 14798 6384
rect 14792 6344 14872 6372
rect 14792 6332 14798 6344
rect 13909 6307 13967 6313
rect 13909 6304 13921 6307
rect 13136 6276 13921 6304
rect 13136 6264 13142 6276
rect 13909 6273 13921 6276
rect 13955 6273 13967 6307
rect 13909 6267 13967 6273
rect 14001 6307 14059 6313
rect 14001 6273 14013 6307
rect 14047 6273 14059 6307
rect 14001 6267 14059 6273
rect 10485 6239 10543 6245
rect 10485 6236 10497 6239
rect 5776 6208 6132 6236
rect 6196 6208 10497 6236
rect 5776 6196 5782 6208
rect 1765 6171 1823 6177
rect 1765 6137 1777 6171
rect 1811 6168 1823 6171
rect 1811 6140 2268 6168
rect 1811 6137 1823 6140
rect 1765 6131 1823 6137
rect 1394 6100 1400 6112
rect 1355 6072 1400 6100
rect 1394 6060 1400 6072
rect 1452 6060 1458 6112
rect 1670 6060 1676 6112
rect 1728 6100 1734 6112
rect 1857 6103 1915 6109
rect 1857 6100 1869 6103
rect 1728 6072 1869 6100
rect 1728 6060 1734 6072
rect 1857 6069 1869 6072
rect 1903 6069 1915 6103
rect 2240 6100 2268 6140
rect 2774 6128 2780 6180
rect 2832 6168 2838 6180
rect 2832 6140 2877 6168
rect 2832 6128 2838 6140
rect 3234 6128 3240 6180
rect 3292 6168 3298 6180
rect 3694 6177 3700 6180
rect 3666 6171 3700 6177
rect 3666 6168 3678 6171
rect 3292 6140 3678 6168
rect 3292 6128 3298 6140
rect 3666 6137 3678 6140
rect 3666 6131 3700 6137
rect 3694 6128 3700 6131
rect 3752 6128 3758 6180
rect 3786 6128 3792 6180
rect 3844 6168 3850 6180
rect 4985 6171 5043 6177
rect 3844 6140 4927 6168
rect 3844 6128 3850 6140
rect 3050 6100 3056 6112
rect 2240 6072 3056 6100
rect 1857 6063 1915 6069
rect 3050 6060 3056 6072
rect 3108 6060 3114 6112
rect 4899 6100 4927 6140
rect 4985 6137 4997 6171
rect 5031 6168 5043 6171
rect 6196 6168 6224 6208
rect 10485 6205 10497 6208
rect 10531 6205 10543 6239
rect 11793 6239 11851 6245
rect 10485 6199 10543 6205
rect 10796 6208 11744 6236
rect 5031 6140 6224 6168
rect 5031 6137 5043 6140
rect 4985 6131 5043 6137
rect 6270 6128 6276 6180
rect 6328 6168 6334 6180
rect 7184 6171 7242 6177
rect 7184 6168 7196 6171
rect 6328 6140 7196 6168
rect 6328 6128 6334 6140
rect 7184 6137 7196 6140
rect 7230 6168 7242 6171
rect 7282 6168 7288 6180
rect 7230 6140 7288 6168
rect 7230 6137 7242 6140
rect 7184 6131 7242 6137
rect 7282 6128 7288 6140
rect 7340 6128 7346 6180
rect 8840 6171 8898 6177
rect 8840 6137 8852 6171
rect 8886 6168 8898 6171
rect 9030 6168 9036 6180
rect 8886 6140 9036 6168
rect 8886 6137 8898 6140
rect 8840 6131 8898 6137
rect 9030 6128 9036 6140
rect 9088 6128 9094 6180
rect 10796 6168 10824 6208
rect 9876 6140 10824 6168
rect 9876 6112 9904 6140
rect 11330 6128 11336 6180
rect 11388 6168 11394 6180
rect 11514 6168 11520 6180
rect 11388 6140 11520 6168
rect 11388 6128 11394 6140
rect 11514 6128 11520 6140
rect 11572 6128 11578 6180
rect 11716 6168 11744 6208
rect 11793 6205 11805 6239
rect 11839 6236 11851 6239
rect 11882 6236 11888 6248
rect 11839 6208 11888 6236
rect 11839 6205 11851 6208
rect 11793 6199 11851 6205
rect 11882 6196 11888 6208
rect 11940 6196 11946 6248
rect 12066 6196 12072 6248
rect 12124 6236 12130 6248
rect 12161 6239 12219 6245
rect 12161 6236 12173 6239
rect 12124 6208 12173 6236
rect 12124 6196 12130 6208
rect 12161 6205 12173 6208
rect 12207 6205 12219 6239
rect 12161 6199 12219 6205
rect 12434 6196 12440 6248
rect 12492 6236 12498 6248
rect 12710 6236 12716 6248
rect 12492 6208 12716 6236
rect 12492 6196 12498 6208
rect 12710 6196 12716 6208
rect 12768 6196 12774 6248
rect 12897 6239 12955 6245
rect 12897 6205 12909 6239
rect 12943 6236 12955 6239
rect 13170 6236 13176 6248
rect 12943 6208 13176 6236
rect 12943 6205 12955 6208
rect 12897 6199 12955 6205
rect 13170 6196 13176 6208
rect 13228 6196 13234 6248
rect 13262 6196 13268 6248
rect 13320 6236 13326 6248
rect 13320 6208 13365 6236
rect 13320 6196 13326 6208
rect 13814 6196 13820 6248
rect 13872 6236 13878 6248
rect 14734 6236 14740 6248
rect 13872 6208 14740 6236
rect 13872 6196 13878 6208
rect 14734 6196 14740 6208
rect 14792 6196 14798 6248
rect 13906 6168 13912 6180
rect 11716 6140 13912 6168
rect 13906 6128 13912 6140
rect 13964 6128 13970 6180
rect 14844 6177 14872 6344
rect 15010 6304 15016 6316
rect 14971 6276 15016 6304
rect 15010 6264 15016 6276
rect 15068 6264 15074 6316
rect 14829 6171 14887 6177
rect 14829 6137 14841 6171
rect 14875 6168 14887 6171
rect 15470 6168 15476 6180
rect 14875 6140 15476 6168
rect 14875 6137 14887 6140
rect 14829 6131 14887 6137
rect 15470 6128 15476 6140
rect 15528 6128 15534 6180
rect 6457 6103 6515 6109
rect 6457 6100 6469 6103
rect 4899 6072 6469 6100
rect 6457 6069 6469 6072
rect 6503 6069 6515 6103
rect 6457 6063 6515 6069
rect 8297 6103 8355 6109
rect 8297 6069 8309 6103
rect 8343 6100 8355 6103
rect 9858 6100 9864 6112
rect 8343 6072 9864 6100
rect 8343 6069 8355 6072
rect 8297 6063 8355 6069
rect 9858 6060 9864 6072
rect 9916 6060 9922 6112
rect 9950 6060 9956 6112
rect 10008 6100 10014 6112
rect 10137 6103 10195 6109
rect 10137 6100 10149 6103
rect 10008 6072 10149 6100
rect 10008 6060 10014 6072
rect 10137 6069 10149 6072
rect 10183 6069 10195 6103
rect 10137 6063 10195 6069
rect 10226 6060 10232 6112
rect 10284 6100 10290 6112
rect 11701 6103 11759 6109
rect 11701 6100 11713 6103
rect 10284 6072 11713 6100
rect 10284 6060 10290 6072
rect 11701 6069 11713 6072
rect 11747 6069 11759 6103
rect 11882 6100 11888 6112
rect 11843 6072 11888 6100
rect 11701 6063 11759 6069
rect 11882 6060 11888 6072
rect 11940 6060 11946 6112
rect 12434 6100 12440 6112
rect 12395 6072 12440 6100
rect 12434 6060 12440 6072
rect 12492 6060 12498 6112
rect 12805 6103 12863 6109
rect 12805 6069 12817 6103
rect 12851 6100 12863 6103
rect 13446 6100 13452 6112
rect 12851 6072 13452 6100
rect 12851 6069 12863 6072
rect 12805 6063 12863 6069
rect 13446 6060 13452 6072
rect 13504 6060 13510 6112
rect 13814 6100 13820 6112
rect 13775 6072 13820 6100
rect 13814 6060 13820 6072
rect 13872 6060 13878 6112
rect 14642 6060 14648 6112
rect 14700 6100 14706 6112
rect 14921 6103 14979 6109
rect 14921 6100 14933 6103
rect 14700 6072 14933 6100
rect 14700 6060 14706 6072
rect 14921 6069 14933 6072
rect 14967 6069 14979 6103
rect 14921 6063 14979 6069
rect 1104 6010 15824 6032
rect 1104 5958 5912 6010
rect 5964 5958 5976 6010
rect 6028 5958 6040 6010
rect 6092 5958 6104 6010
rect 6156 5958 10843 6010
rect 10895 5958 10907 6010
rect 10959 5958 10971 6010
rect 11023 5958 11035 6010
rect 11087 5958 15824 6010
rect 1104 5936 15824 5958
rect 1394 5856 1400 5908
rect 1452 5896 1458 5908
rect 2409 5899 2467 5905
rect 2409 5896 2421 5899
rect 1452 5868 2421 5896
rect 1452 5856 1458 5868
rect 2409 5865 2421 5868
rect 2455 5865 2467 5899
rect 2409 5859 2467 5865
rect 3789 5899 3847 5905
rect 3789 5865 3801 5899
rect 3835 5896 3847 5899
rect 8110 5896 8116 5908
rect 3835 5868 8116 5896
rect 3835 5865 3847 5868
rect 3789 5859 3847 5865
rect 8110 5856 8116 5868
rect 8168 5856 8174 5908
rect 8570 5856 8576 5908
rect 8628 5896 8634 5908
rect 8665 5899 8723 5905
rect 8665 5896 8677 5899
rect 8628 5868 8677 5896
rect 8628 5856 8634 5868
rect 8665 5865 8677 5868
rect 8711 5865 8723 5899
rect 8665 5859 8723 5865
rect 8938 5856 8944 5908
rect 8996 5896 9002 5908
rect 9125 5899 9183 5905
rect 9125 5896 9137 5899
rect 8996 5868 9137 5896
rect 8996 5856 9002 5868
rect 9125 5865 9137 5868
rect 9171 5865 9183 5899
rect 9125 5859 9183 5865
rect 9306 5856 9312 5908
rect 9364 5896 9370 5908
rect 9364 5868 10180 5896
rect 9364 5856 9370 5868
rect 4617 5831 4675 5837
rect 2608 5800 4568 5828
rect 1394 5760 1400 5772
rect 1355 5732 1400 5760
rect 1394 5720 1400 5732
rect 1452 5720 1458 5772
rect 1762 5720 1768 5772
rect 1820 5760 1826 5772
rect 2317 5763 2375 5769
rect 2317 5760 2329 5763
rect 1820 5732 2329 5760
rect 1820 5720 1826 5732
rect 2317 5729 2329 5732
rect 2363 5729 2375 5763
rect 2317 5723 2375 5729
rect 2608 5701 2636 5800
rect 3326 5760 3332 5772
rect 3287 5732 3332 5760
rect 3326 5720 3332 5732
rect 3384 5720 3390 5772
rect 3421 5763 3479 5769
rect 3421 5729 3433 5763
rect 3467 5760 3479 5763
rect 3786 5760 3792 5772
rect 3467 5732 3792 5760
rect 3467 5729 3479 5732
rect 3421 5723 3479 5729
rect 3786 5720 3792 5732
rect 3844 5720 3850 5772
rect 4062 5760 4068 5772
rect 4023 5732 4068 5760
rect 4062 5720 4068 5732
rect 4120 5720 4126 5772
rect 4540 5760 4568 5800
rect 4617 5797 4629 5831
rect 4663 5828 4675 5831
rect 10045 5831 10103 5837
rect 10045 5828 10057 5831
rect 4663 5800 10057 5828
rect 4663 5797 4675 5800
rect 4617 5791 4675 5797
rect 10045 5797 10057 5800
rect 10091 5797 10103 5831
rect 10152 5828 10180 5868
rect 10226 5856 10232 5908
rect 10284 5896 10290 5908
rect 10594 5896 10600 5908
rect 10284 5868 10600 5896
rect 10284 5856 10290 5868
rect 10594 5856 10600 5868
rect 10652 5856 10658 5908
rect 11149 5899 11207 5905
rect 11149 5865 11161 5899
rect 11195 5896 11207 5899
rect 11238 5896 11244 5908
rect 11195 5868 11244 5896
rect 11195 5865 11207 5868
rect 11149 5859 11207 5865
rect 11238 5856 11244 5868
rect 11296 5856 11302 5908
rect 11609 5899 11667 5905
rect 11609 5865 11621 5899
rect 11655 5896 11667 5899
rect 11701 5899 11759 5905
rect 11701 5896 11713 5899
rect 11655 5868 11713 5896
rect 11655 5865 11667 5868
rect 11609 5859 11667 5865
rect 11701 5865 11713 5868
rect 11747 5865 11759 5899
rect 11701 5859 11759 5865
rect 11790 5856 11796 5908
rect 11848 5896 11854 5908
rect 12434 5896 12440 5908
rect 11848 5868 12440 5896
rect 11848 5856 11854 5868
rect 12434 5856 12440 5868
rect 12492 5856 12498 5908
rect 12529 5899 12587 5905
rect 12529 5865 12541 5899
rect 12575 5896 12587 5899
rect 13081 5899 13139 5905
rect 13081 5896 13093 5899
rect 12575 5868 13093 5896
rect 12575 5865 12587 5868
rect 12529 5859 12587 5865
rect 13081 5865 13093 5868
rect 13127 5896 13139 5899
rect 13722 5896 13728 5908
rect 13127 5868 13728 5896
rect 13127 5865 13139 5868
rect 13081 5859 13139 5865
rect 13722 5856 13728 5868
rect 13780 5856 13786 5908
rect 14090 5896 14096 5908
rect 14051 5868 14096 5896
rect 14090 5856 14096 5868
rect 14148 5856 14154 5908
rect 14734 5896 14740 5908
rect 14695 5868 14740 5896
rect 14734 5856 14740 5868
rect 14792 5856 14798 5908
rect 10686 5828 10692 5840
rect 10152 5800 10692 5828
rect 10045 5791 10103 5797
rect 10686 5788 10692 5800
rect 10744 5788 10750 5840
rect 10962 5828 10968 5840
rect 10888 5800 10968 5828
rect 5241 5763 5299 5769
rect 5241 5760 5253 5763
rect 4540 5732 5253 5760
rect 5241 5729 5253 5732
rect 5287 5760 5299 5763
rect 6454 5760 6460 5772
rect 5287 5732 6460 5760
rect 5287 5729 5299 5732
rect 5241 5723 5299 5729
rect 6454 5720 6460 5732
rect 6512 5720 6518 5772
rect 6914 5769 6920 5772
rect 6908 5760 6920 5769
rect 6875 5732 6920 5760
rect 6908 5723 6920 5732
rect 6914 5720 6920 5723
rect 6972 5720 6978 5772
rect 8110 5720 8116 5772
rect 8168 5760 8174 5772
rect 8846 5760 8852 5772
rect 8168 5732 8852 5760
rect 8168 5720 8174 5732
rect 8846 5720 8852 5732
rect 8904 5720 8910 5772
rect 9490 5760 9496 5772
rect 9451 5732 9496 5760
rect 9490 5720 9496 5732
rect 9548 5720 9554 5772
rect 10137 5763 10195 5769
rect 10137 5729 10149 5763
rect 10183 5760 10195 5763
rect 10888 5760 10916 5800
rect 10962 5788 10968 5800
rect 11020 5788 11026 5840
rect 11057 5831 11115 5837
rect 11057 5797 11069 5831
rect 11103 5828 11115 5831
rect 11514 5828 11520 5840
rect 11103 5800 11520 5828
rect 11103 5797 11115 5800
rect 11057 5791 11115 5797
rect 11514 5788 11520 5800
rect 11572 5788 11578 5840
rect 11974 5828 11980 5840
rect 11900 5800 11980 5828
rect 11900 5760 11928 5800
rect 11974 5788 11980 5800
rect 12032 5788 12038 5840
rect 12069 5831 12127 5837
rect 12069 5797 12081 5831
rect 12115 5828 12127 5831
rect 12115 5800 12756 5828
rect 12115 5797 12127 5800
rect 12069 5791 12127 5797
rect 12728 5760 12756 5800
rect 12802 5788 12808 5840
rect 12860 5828 12866 5840
rect 12860 5800 14320 5828
rect 12860 5788 12866 5800
rect 13998 5760 14004 5772
rect 10183 5732 10916 5760
rect 10980 5732 11928 5760
rect 11992 5732 12296 5760
rect 12728 5732 14004 5760
rect 10183 5729 10195 5732
rect 10137 5723 10195 5729
rect 2593 5695 2651 5701
rect 2593 5661 2605 5695
rect 2639 5661 2651 5695
rect 3602 5692 3608 5704
rect 3563 5664 3608 5692
rect 2593 5655 2651 5661
rect 3602 5652 3608 5664
rect 3660 5652 3666 5704
rect 3694 5652 3700 5704
rect 3752 5692 3758 5704
rect 4249 5695 4307 5701
rect 4249 5692 4261 5695
rect 3752 5664 4261 5692
rect 3752 5652 3758 5664
rect 4249 5661 4261 5664
rect 4295 5661 4307 5695
rect 4249 5655 4307 5661
rect 4706 5652 4712 5704
rect 4764 5692 4770 5704
rect 4985 5695 5043 5701
rect 4985 5692 4997 5695
rect 4764 5664 4997 5692
rect 4764 5652 4770 5664
rect 4985 5661 4997 5664
rect 5031 5661 5043 5695
rect 4985 5655 5043 5661
rect 6641 5695 6699 5701
rect 6641 5661 6653 5695
rect 6687 5661 6699 5695
rect 6641 5655 6699 5661
rect 8757 5695 8815 5701
rect 8757 5661 8769 5695
rect 8803 5661 8815 5695
rect 8757 5655 8815 5661
rect 8941 5695 8999 5701
rect 8941 5661 8953 5695
rect 8987 5692 8999 5695
rect 9214 5692 9220 5704
rect 8987 5664 9220 5692
rect 8987 5661 8999 5664
rect 8941 5655 8999 5661
rect 1946 5624 1952 5636
rect 1907 5596 1952 5624
rect 1946 5584 1952 5596
rect 2004 5584 2010 5636
rect 2682 5584 2688 5636
rect 2740 5624 2746 5636
rect 4338 5624 4344 5636
rect 2740 5596 4344 5624
rect 2740 5584 2746 5596
rect 4338 5584 4344 5596
rect 4396 5584 4402 5636
rect 1581 5559 1639 5565
rect 1581 5525 1593 5559
rect 1627 5556 1639 5559
rect 2406 5556 2412 5568
rect 1627 5528 2412 5556
rect 1627 5525 1639 5528
rect 1581 5519 1639 5525
rect 2406 5516 2412 5528
rect 2464 5516 2470 5568
rect 2961 5559 3019 5565
rect 2961 5525 2973 5559
rect 3007 5556 3019 5559
rect 3789 5559 3847 5565
rect 3789 5556 3801 5559
rect 3007 5528 3801 5556
rect 3007 5525 3019 5528
rect 2961 5519 3019 5525
rect 3789 5525 3801 5528
rect 3835 5525 3847 5559
rect 3789 5519 3847 5525
rect 4154 5516 4160 5568
rect 4212 5556 4218 5568
rect 5718 5556 5724 5568
rect 4212 5528 5724 5556
rect 4212 5516 4218 5528
rect 5718 5516 5724 5528
rect 5776 5516 5782 5568
rect 6362 5556 6368 5568
rect 6323 5528 6368 5556
rect 6362 5516 6368 5528
rect 6420 5516 6426 5568
rect 6656 5556 6684 5655
rect 8297 5627 8355 5633
rect 8297 5624 8309 5627
rect 7576 5596 8309 5624
rect 7576 5568 7604 5596
rect 8297 5593 8309 5596
rect 8343 5593 8355 5627
rect 8297 5587 8355 5593
rect 8772 5624 8800 5655
rect 9214 5652 9220 5664
rect 9272 5652 9278 5704
rect 9306 5652 9312 5704
rect 9364 5692 9370 5704
rect 10321 5695 10379 5701
rect 10321 5692 10333 5695
rect 9364 5664 10333 5692
rect 9364 5652 9370 5664
rect 10321 5661 10333 5664
rect 10367 5661 10379 5695
rect 10778 5692 10784 5704
rect 10321 5655 10379 5661
rect 10419 5664 10784 5692
rect 9125 5627 9183 5633
rect 9125 5624 9137 5627
rect 8772 5596 9137 5624
rect 8772 5568 8800 5596
rect 9125 5593 9137 5596
rect 9171 5593 9183 5627
rect 9125 5587 9183 5593
rect 9324 5596 10180 5624
rect 6822 5556 6828 5568
rect 6656 5528 6828 5556
rect 6822 5516 6828 5528
rect 6880 5516 6886 5568
rect 7558 5516 7564 5568
rect 7616 5516 7622 5568
rect 7834 5516 7840 5568
rect 7892 5556 7898 5568
rect 8021 5559 8079 5565
rect 8021 5556 8033 5559
rect 7892 5528 8033 5556
rect 7892 5516 7898 5528
rect 8021 5525 8033 5528
rect 8067 5525 8079 5559
rect 8021 5519 8079 5525
rect 8754 5516 8760 5568
rect 8812 5516 8818 5568
rect 9324 5565 9352 5596
rect 9309 5559 9367 5565
rect 9309 5525 9321 5559
rect 9355 5525 9367 5559
rect 9309 5519 9367 5525
rect 9674 5516 9680 5568
rect 9732 5556 9738 5568
rect 10152 5556 10180 5596
rect 10226 5584 10232 5636
rect 10284 5624 10290 5636
rect 10419 5624 10447 5664
rect 10778 5652 10784 5664
rect 10836 5652 10842 5704
rect 10980 5624 11008 5732
rect 11992 5704 12020 5732
rect 11054 5652 11060 5704
rect 11112 5692 11118 5704
rect 11333 5695 11391 5701
rect 11112 5664 11284 5692
rect 11112 5652 11118 5664
rect 10284 5596 10447 5624
rect 10520 5596 11008 5624
rect 11256 5624 11284 5664
rect 11333 5661 11345 5695
rect 11379 5692 11391 5695
rect 11422 5692 11428 5704
rect 11379 5664 11428 5692
rect 11379 5661 11391 5664
rect 11333 5655 11391 5661
rect 11422 5652 11428 5664
rect 11480 5652 11486 5704
rect 11514 5652 11520 5704
rect 11572 5692 11578 5704
rect 11572 5664 11744 5692
rect 11572 5652 11578 5664
rect 11716 5624 11744 5664
rect 11974 5652 11980 5704
rect 12032 5652 12038 5704
rect 12268 5701 12296 5732
rect 13998 5720 14004 5732
rect 14056 5720 14062 5772
rect 12161 5695 12219 5701
rect 12161 5661 12173 5695
rect 12207 5661 12219 5695
rect 12161 5655 12219 5661
rect 12253 5695 12311 5701
rect 12253 5661 12265 5695
rect 12299 5661 12311 5695
rect 12253 5655 12311 5661
rect 12176 5624 12204 5655
rect 12894 5652 12900 5704
rect 12952 5692 12958 5704
rect 13173 5695 13231 5701
rect 13173 5692 13185 5695
rect 12952 5664 13185 5692
rect 12952 5652 12958 5664
rect 13173 5661 13185 5664
rect 13219 5661 13231 5695
rect 13173 5655 13231 5661
rect 13262 5652 13268 5704
rect 13320 5692 13326 5704
rect 13320 5664 13365 5692
rect 13320 5652 13326 5664
rect 13446 5652 13452 5704
rect 13504 5692 13510 5704
rect 14090 5692 14096 5704
rect 13504 5664 14096 5692
rect 13504 5652 13510 5664
rect 14090 5652 14096 5664
rect 14148 5652 14154 5704
rect 14292 5701 14320 5800
rect 14185 5695 14243 5701
rect 14185 5661 14197 5695
rect 14231 5661 14243 5695
rect 14185 5655 14243 5661
rect 14277 5695 14335 5701
rect 14277 5661 14289 5695
rect 14323 5661 14335 5695
rect 14277 5655 14335 5661
rect 11256 5596 11652 5624
rect 11716 5596 12204 5624
rect 10284 5584 10290 5596
rect 10520 5556 10548 5596
rect 10686 5556 10692 5568
rect 9732 5528 9777 5556
rect 10152 5528 10548 5556
rect 10647 5528 10692 5556
rect 9732 5516 9738 5528
rect 10686 5516 10692 5528
rect 10744 5516 10750 5568
rect 10778 5516 10784 5568
rect 10836 5556 10842 5568
rect 11517 5559 11575 5565
rect 11517 5556 11529 5559
rect 10836 5528 11529 5556
rect 10836 5516 10842 5528
rect 11517 5525 11529 5528
rect 11563 5525 11575 5559
rect 11624 5556 11652 5596
rect 12434 5584 12440 5636
rect 12492 5624 12498 5636
rect 14200 5624 14228 5655
rect 12492 5596 14228 5624
rect 12492 5584 12498 5596
rect 12529 5559 12587 5565
rect 12529 5556 12541 5559
rect 11624 5528 12541 5556
rect 11517 5519 11575 5525
rect 12529 5525 12541 5528
rect 12575 5525 12587 5559
rect 12710 5556 12716 5568
rect 12671 5528 12716 5556
rect 12529 5519 12587 5525
rect 12710 5516 12716 5528
rect 12768 5516 12774 5568
rect 13725 5559 13783 5565
rect 13725 5525 13737 5559
rect 13771 5556 13783 5559
rect 13998 5556 14004 5568
rect 13771 5528 14004 5556
rect 13771 5525 13783 5528
rect 13725 5519 13783 5525
rect 13998 5516 14004 5528
rect 14056 5516 14062 5568
rect 1104 5466 15824 5488
rect 1104 5414 3447 5466
rect 3499 5414 3511 5466
rect 3563 5414 3575 5466
rect 3627 5414 3639 5466
rect 3691 5414 8378 5466
rect 8430 5414 8442 5466
rect 8494 5414 8506 5466
rect 8558 5414 8570 5466
rect 8622 5414 13308 5466
rect 13360 5414 13372 5466
rect 13424 5414 13436 5466
rect 13488 5414 13500 5466
rect 13552 5414 15824 5466
rect 1104 5392 15824 5414
rect 2130 5312 2136 5364
rect 2188 5352 2194 5364
rect 3053 5355 3111 5361
rect 3053 5352 3065 5355
rect 2188 5324 3065 5352
rect 2188 5312 2194 5324
rect 3053 5321 3065 5324
rect 3099 5321 3111 5355
rect 3053 5315 3111 5321
rect 3326 5312 3332 5364
rect 3384 5352 3390 5364
rect 4065 5355 4123 5361
rect 4065 5352 4077 5355
rect 3384 5324 4077 5352
rect 3384 5312 3390 5324
rect 4065 5321 4077 5324
rect 4111 5321 4123 5355
rect 4065 5315 4123 5321
rect 4154 5312 4160 5364
rect 4212 5352 4218 5364
rect 10137 5355 10195 5361
rect 10137 5352 10149 5355
rect 4212 5324 4660 5352
rect 4212 5312 4218 5324
rect 1673 5287 1731 5293
rect 1673 5253 1685 5287
rect 1719 5284 1731 5287
rect 2590 5284 2596 5296
rect 1719 5256 2596 5284
rect 1719 5253 1731 5256
rect 1673 5247 1731 5253
rect 2590 5244 2596 5256
rect 2648 5244 2654 5296
rect 3878 5284 3884 5296
rect 3712 5256 3884 5284
rect 2501 5219 2559 5225
rect 2501 5185 2513 5219
rect 2547 5216 2559 5219
rect 2866 5216 2872 5228
rect 2547 5188 2872 5216
rect 2547 5185 2559 5188
rect 2501 5179 2559 5185
rect 2866 5176 2872 5188
rect 2924 5176 2930 5228
rect 2961 5219 3019 5225
rect 2961 5185 2973 5219
rect 3007 5216 3019 5219
rect 3510 5216 3516 5228
rect 3007 5188 3516 5216
rect 3007 5185 3019 5188
rect 2961 5179 3019 5185
rect 3510 5176 3516 5188
rect 3568 5176 3574 5228
rect 3712 5225 3740 5256
rect 3878 5244 3884 5256
rect 3936 5244 3942 5296
rect 4430 5284 4436 5296
rect 4264 5256 4436 5284
rect 3697 5219 3755 5225
rect 3697 5185 3709 5219
rect 3743 5185 3755 5219
rect 3697 5179 3755 5185
rect 1489 5151 1547 5157
rect 1489 5117 1501 5151
rect 1535 5148 1547 5151
rect 1535 5120 3556 5148
rect 1535 5117 1547 5120
rect 1489 5111 1547 5117
rect 2225 5083 2283 5089
rect 2225 5049 2237 5083
rect 2271 5080 2283 5083
rect 2774 5080 2780 5092
rect 2271 5052 2780 5080
rect 2271 5049 2283 5052
rect 2225 5043 2283 5049
rect 2774 5040 2780 5052
rect 2832 5040 2838 5092
rect 3528 5080 3556 5120
rect 4264 5080 4292 5256
rect 4430 5244 4436 5256
rect 4488 5244 4494 5296
rect 4632 5225 4660 5324
rect 5000 5324 10149 5352
rect 4617 5219 4675 5225
rect 4617 5185 4629 5219
rect 4663 5185 4675 5219
rect 4617 5179 4675 5185
rect 4433 5151 4491 5157
rect 4433 5117 4445 5151
rect 4479 5148 4491 5151
rect 5000 5148 5028 5324
rect 10137 5321 10149 5324
rect 10183 5321 10195 5355
rect 10137 5315 10195 5321
rect 10235 5324 11376 5352
rect 6454 5284 6460 5296
rect 6415 5256 6460 5284
rect 6454 5244 6460 5256
rect 6512 5244 6518 5296
rect 7834 5244 7840 5296
rect 7892 5284 7898 5296
rect 8297 5287 8355 5293
rect 8297 5284 8309 5287
rect 7892 5256 8309 5284
rect 7892 5244 7898 5256
rect 8297 5253 8309 5256
rect 8343 5253 8355 5287
rect 8297 5247 8355 5253
rect 9861 5287 9919 5293
rect 9861 5253 9873 5287
rect 9907 5253 9919 5287
rect 9861 5247 9919 5253
rect 9953 5287 10011 5293
rect 9953 5253 9965 5287
rect 9999 5284 10011 5287
rect 10235 5284 10263 5324
rect 10502 5284 10508 5296
rect 9999 5256 10263 5284
rect 9999 5253 10011 5256
rect 9953 5247 10011 5253
rect 6822 5216 6828 5228
rect 6288 5188 6828 5216
rect 4479 5120 5028 5148
rect 5077 5151 5135 5157
rect 4479 5117 4491 5120
rect 4433 5111 4491 5117
rect 5077 5117 5089 5151
rect 5123 5148 5135 5151
rect 5902 5148 5908 5160
rect 5123 5120 5908 5148
rect 5123 5117 5135 5120
rect 5077 5111 5135 5117
rect 5902 5108 5908 5120
rect 5960 5148 5966 5160
rect 6288 5148 6316 5188
rect 6822 5176 6828 5188
rect 6880 5176 6886 5228
rect 8386 5176 8392 5228
rect 8444 5216 8450 5228
rect 8481 5219 8539 5225
rect 8481 5216 8493 5219
rect 8444 5188 8493 5216
rect 8444 5176 8450 5188
rect 8481 5185 8493 5188
rect 8527 5185 8539 5219
rect 8481 5179 8539 5185
rect 5960 5120 6316 5148
rect 5960 5108 5966 5120
rect 6362 5108 6368 5160
rect 6420 5148 6426 5160
rect 6420 5120 7236 5148
rect 6420 5108 6426 5120
rect 3528 5052 4292 5080
rect 4338 5040 4344 5092
rect 4396 5080 4402 5092
rect 5258 5080 5264 5092
rect 4396 5052 5264 5080
rect 4396 5040 4402 5052
rect 5258 5040 5264 5052
rect 5316 5089 5322 5092
rect 5316 5083 5380 5089
rect 5316 5049 5334 5083
rect 5368 5049 5380 5083
rect 5316 5043 5380 5049
rect 5316 5040 5322 5043
rect 7006 5040 7012 5092
rect 7064 5089 7070 5092
rect 7064 5083 7128 5089
rect 7064 5049 7082 5083
rect 7116 5049 7128 5083
rect 7208 5080 7236 5120
rect 7926 5108 7932 5160
rect 7984 5148 7990 5160
rect 9876 5148 9904 5247
rect 10500 5244 10508 5284
rect 10560 5244 10566 5296
rect 10500 5157 10528 5244
rect 10796 5225 10824 5324
rect 10870 5244 10876 5296
rect 10928 5284 10934 5296
rect 11348 5284 11376 5324
rect 12250 5312 12256 5364
rect 12308 5352 12314 5364
rect 14458 5352 14464 5364
rect 12308 5324 14464 5352
rect 12308 5312 12314 5324
rect 14458 5312 14464 5324
rect 14516 5312 14522 5364
rect 12342 5284 12348 5296
rect 10928 5256 11284 5284
rect 11348 5256 12348 5284
rect 10928 5244 10934 5256
rect 10597 5219 10655 5225
rect 10597 5185 10609 5219
rect 10643 5185 10655 5219
rect 10597 5179 10655 5185
rect 10781 5219 10839 5225
rect 10781 5185 10793 5219
rect 10827 5185 10839 5219
rect 10781 5179 10839 5185
rect 10500 5151 10563 5157
rect 7984 5120 10456 5148
rect 10500 5120 10517 5151
rect 7984 5108 7990 5120
rect 8726 5083 8784 5089
rect 8726 5080 8738 5083
rect 7208 5052 8738 5080
rect 7064 5043 7128 5049
rect 8726 5049 8738 5052
rect 8772 5049 8784 5083
rect 8726 5043 8784 5049
rect 7064 5040 7070 5043
rect 8846 5040 8852 5092
rect 8904 5080 8910 5092
rect 9122 5080 9128 5092
rect 8904 5052 9128 5080
rect 8904 5040 8910 5052
rect 9122 5040 9128 5052
rect 9180 5040 9186 5092
rect 9214 5040 9220 5092
rect 9272 5080 9278 5092
rect 9398 5080 9404 5092
rect 9272 5052 9404 5080
rect 9272 5040 9278 5052
rect 9398 5040 9404 5052
rect 9456 5040 9462 5092
rect 9490 5040 9496 5092
rect 9548 5080 9554 5092
rect 10226 5080 10232 5092
rect 9548 5052 10232 5080
rect 9548 5040 9554 5052
rect 10226 5040 10232 5052
rect 10284 5040 10290 5092
rect 10428 5024 10456 5120
rect 10505 5117 10517 5120
rect 10551 5117 10563 5151
rect 10612 5148 10640 5179
rect 10962 5176 10968 5228
rect 11020 5216 11026 5228
rect 11256 5216 11284 5256
rect 12342 5244 12348 5256
rect 12400 5244 12406 5296
rect 12894 5244 12900 5296
rect 12952 5284 12958 5296
rect 12952 5256 13216 5284
rect 12952 5244 12958 5256
rect 11698 5216 11704 5228
rect 11020 5188 11192 5216
rect 11256 5188 11704 5216
rect 11020 5176 11026 5188
rect 11164 5148 11192 5188
rect 11698 5176 11704 5188
rect 11756 5216 11762 5228
rect 11882 5216 11888 5228
rect 11756 5188 11888 5216
rect 11756 5176 11762 5188
rect 11882 5176 11888 5188
rect 11940 5176 11946 5228
rect 12526 5176 12532 5228
rect 12584 5216 12590 5228
rect 13081 5219 13139 5225
rect 13081 5216 13093 5219
rect 12584 5188 13093 5216
rect 12584 5176 12590 5188
rect 13081 5185 13093 5188
rect 13127 5185 13139 5219
rect 13188 5216 13216 5256
rect 13722 5244 13728 5296
rect 13780 5284 13786 5296
rect 16758 5284 16764 5296
rect 13780 5256 16764 5284
rect 13780 5244 13786 5256
rect 16758 5244 16764 5256
rect 16816 5244 16822 5296
rect 13814 5216 13820 5228
rect 13188 5188 13820 5216
rect 13081 5179 13139 5185
rect 13814 5176 13820 5188
rect 13872 5176 13878 5228
rect 13906 5176 13912 5228
rect 13964 5216 13970 5228
rect 14001 5219 14059 5225
rect 14001 5216 14013 5219
rect 13964 5188 14013 5216
rect 13964 5176 13970 5188
rect 14001 5185 14013 5188
rect 14047 5185 14059 5219
rect 14001 5179 14059 5185
rect 14918 5176 14924 5228
rect 14976 5216 14982 5228
rect 15013 5219 15071 5225
rect 15013 5216 15025 5219
rect 14976 5188 15025 5216
rect 14976 5176 14982 5188
rect 15013 5185 15025 5188
rect 15059 5185 15071 5219
rect 15013 5179 15071 5185
rect 11517 5151 11575 5157
rect 11517 5148 11529 5151
rect 10612 5120 10916 5148
rect 11164 5120 11529 5148
rect 10505 5111 10563 5117
rect 10594 5040 10600 5092
rect 10652 5080 10658 5092
rect 10778 5080 10784 5092
rect 10652 5052 10784 5080
rect 10652 5040 10658 5052
rect 10778 5040 10784 5052
rect 10836 5040 10842 5092
rect 10888 5080 10916 5120
rect 11517 5117 11529 5120
rect 11563 5117 11575 5151
rect 11517 5111 11575 5117
rect 11609 5151 11667 5157
rect 11609 5117 11621 5151
rect 11655 5148 11667 5151
rect 12618 5148 12624 5160
rect 11655 5120 12624 5148
rect 11655 5117 11667 5120
rect 11609 5111 11667 5117
rect 12618 5108 12624 5120
rect 12676 5108 12682 5160
rect 11238 5080 11244 5092
rect 10888 5052 11244 5080
rect 11238 5040 11244 5052
rect 11296 5040 11302 5092
rect 12805 5083 12863 5089
rect 12805 5080 12817 5083
rect 11440 5052 12817 5080
rect 1854 5012 1860 5024
rect 1815 4984 1860 5012
rect 1854 4972 1860 4984
rect 1912 4972 1918 5024
rect 2317 5015 2375 5021
rect 2317 4981 2329 5015
rect 2363 5012 2375 5015
rect 2958 5012 2964 5024
rect 2363 4984 2964 5012
rect 2363 4981 2375 4984
rect 2317 4975 2375 4981
rect 2958 4972 2964 4984
rect 3016 5012 3022 5024
rect 3326 5012 3332 5024
rect 3016 4984 3332 5012
rect 3016 4972 3022 4984
rect 3326 4972 3332 4984
rect 3384 4972 3390 5024
rect 3421 5015 3479 5021
rect 3421 4981 3433 5015
rect 3467 5012 3479 5015
rect 4430 5012 4436 5024
rect 3467 4984 4436 5012
rect 3467 4981 3479 4984
rect 3421 4975 3479 4981
rect 4430 4972 4436 4984
rect 4488 4972 4494 5024
rect 4525 5015 4583 5021
rect 4525 4981 4537 5015
rect 4571 5012 4583 5015
rect 6270 5012 6276 5024
rect 4571 4984 6276 5012
rect 4571 4981 4583 4984
rect 4525 4975 4583 4981
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 8018 4972 8024 5024
rect 8076 5012 8082 5024
rect 8205 5015 8263 5021
rect 8205 5012 8217 5015
rect 8076 4984 8217 5012
rect 8076 4972 8082 4984
rect 8205 4981 8217 4984
rect 8251 4981 8263 5015
rect 8205 4975 8263 4981
rect 8297 5015 8355 5021
rect 8297 4981 8309 5015
rect 8343 5012 8355 5015
rect 9582 5012 9588 5024
rect 8343 4984 9588 5012
rect 8343 4981 8355 4984
rect 8297 4975 8355 4981
rect 9582 4972 9588 4984
rect 9640 5012 9646 5024
rect 9953 5015 10011 5021
rect 9953 5012 9965 5015
rect 9640 4984 9965 5012
rect 9640 4972 9646 4984
rect 9953 4981 9965 4984
rect 9999 4981 10011 5015
rect 9953 4975 10011 4981
rect 10410 4972 10416 5024
rect 10468 4972 10474 5024
rect 11149 5015 11207 5021
rect 11149 4981 11161 5015
rect 11195 5012 11207 5015
rect 11440 5012 11468 5052
rect 12805 5049 12817 5052
rect 12851 5049 12863 5083
rect 12805 5043 12863 5049
rect 13078 5040 13084 5092
rect 13136 5080 13142 5092
rect 13998 5080 14004 5092
rect 13136 5052 14004 5080
rect 13136 5040 13142 5052
rect 13998 5040 14004 5052
rect 14056 5040 14062 5092
rect 14829 5083 14887 5089
rect 14829 5049 14841 5083
rect 14875 5080 14887 5083
rect 15010 5080 15016 5092
rect 14875 5052 15016 5080
rect 14875 5049 14887 5052
rect 14829 5043 14887 5049
rect 15010 5040 15016 5052
rect 15068 5080 15074 5092
rect 16298 5080 16304 5092
rect 15068 5052 16304 5080
rect 15068 5040 15074 5052
rect 16298 5040 16304 5052
rect 16356 5040 16362 5092
rect 11195 4984 11468 5012
rect 11195 4981 11207 4984
rect 11149 4975 11207 4981
rect 11790 4972 11796 5024
rect 11848 5012 11854 5024
rect 12437 5015 12495 5021
rect 12437 5012 12449 5015
rect 11848 4984 12449 5012
rect 11848 4972 11854 4984
rect 12437 4981 12449 4984
rect 12483 4981 12495 5015
rect 12437 4975 12495 4981
rect 12526 4972 12532 5024
rect 12584 5012 12590 5024
rect 12897 5015 12955 5021
rect 12897 5012 12909 5015
rect 12584 4984 12909 5012
rect 12584 4972 12590 4984
rect 12897 4981 12909 4984
rect 12943 4981 12955 5015
rect 12897 4975 12955 4981
rect 13262 4972 13268 5024
rect 13320 5012 13326 5024
rect 13449 5015 13507 5021
rect 13449 5012 13461 5015
rect 13320 4984 13461 5012
rect 13320 4972 13326 4984
rect 13449 4981 13461 4984
rect 13495 4981 13507 5015
rect 13814 5012 13820 5024
rect 13775 4984 13820 5012
rect 13449 4975 13507 4981
rect 13814 4972 13820 4984
rect 13872 4972 13878 5024
rect 13906 4972 13912 5024
rect 13964 5012 13970 5024
rect 14458 5012 14464 5024
rect 13964 4984 14009 5012
rect 14419 4984 14464 5012
rect 13964 4972 13970 4984
rect 14458 4972 14464 4984
rect 14516 4972 14522 5024
rect 14642 4972 14648 5024
rect 14700 5012 14706 5024
rect 14921 5015 14979 5021
rect 14921 5012 14933 5015
rect 14700 4984 14933 5012
rect 14700 4972 14706 4984
rect 14921 4981 14933 4984
rect 14967 4981 14979 5015
rect 14921 4975 14979 4981
rect 1104 4922 15824 4944
rect 1104 4870 5912 4922
rect 5964 4870 5976 4922
rect 6028 4870 6040 4922
rect 6092 4870 6104 4922
rect 6156 4870 10843 4922
rect 10895 4870 10907 4922
rect 10959 4870 10971 4922
rect 11023 4870 11035 4922
rect 11087 4870 15824 4922
rect 1104 4848 15824 4870
rect 2314 4768 2320 4820
rect 2372 4808 2378 4820
rect 2682 4808 2688 4820
rect 2372 4780 2688 4808
rect 2372 4768 2378 4780
rect 2682 4768 2688 4780
rect 2740 4768 2746 4820
rect 3329 4811 3387 4817
rect 3329 4777 3341 4811
rect 3375 4808 3387 4811
rect 4154 4808 4160 4820
rect 3375 4780 4160 4808
rect 3375 4777 3387 4780
rect 3329 4771 3387 4777
rect 4154 4768 4160 4780
rect 4212 4768 4218 4820
rect 4709 4811 4767 4817
rect 4709 4777 4721 4811
rect 4755 4777 4767 4811
rect 4709 4771 4767 4777
rect 5077 4811 5135 4817
rect 5077 4777 5089 4811
rect 5123 4808 5135 4811
rect 5442 4808 5448 4820
rect 5123 4780 5448 4808
rect 5123 4777 5135 4780
rect 5077 4771 5135 4777
rect 2409 4743 2467 4749
rect 2409 4709 2421 4743
rect 2455 4740 2467 4743
rect 3878 4740 3884 4752
rect 2455 4712 3884 4740
rect 2455 4709 2467 4712
rect 2409 4703 2467 4709
rect 3878 4700 3884 4712
rect 3936 4700 3942 4752
rect 4724 4740 4752 4771
rect 5442 4768 5448 4780
rect 5500 4768 5506 4820
rect 5626 4768 5632 4820
rect 5684 4808 5690 4820
rect 5721 4811 5779 4817
rect 5721 4808 5733 4811
rect 5684 4780 5733 4808
rect 5684 4768 5690 4780
rect 5721 4777 5733 4780
rect 5767 4777 5779 4811
rect 5721 4771 5779 4777
rect 6089 4811 6147 4817
rect 6089 4777 6101 4811
rect 6135 4808 6147 4811
rect 9674 4808 9680 4820
rect 6135 4780 9680 4808
rect 6135 4777 6147 4780
rect 6089 4771 6147 4777
rect 9674 4768 9680 4780
rect 9732 4768 9738 4820
rect 9858 4768 9864 4820
rect 9916 4808 9922 4820
rect 10045 4811 10103 4817
rect 10045 4808 10057 4811
rect 9916 4780 10057 4808
rect 9916 4768 9922 4780
rect 10045 4777 10057 4780
rect 10091 4777 10103 4811
rect 10045 4771 10103 4777
rect 10137 4811 10195 4817
rect 10137 4777 10149 4811
rect 10183 4808 10195 4811
rect 10318 4808 10324 4820
rect 10183 4780 10324 4808
rect 10183 4777 10195 4780
rect 10137 4771 10195 4777
rect 10318 4768 10324 4780
rect 10376 4768 10382 4820
rect 10502 4768 10508 4820
rect 10560 4808 10566 4820
rect 10689 4811 10747 4817
rect 10689 4808 10701 4811
rect 10560 4780 10701 4808
rect 10560 4768 10566 4780
rect 10689 4777 10701 4780
rect 10735 4777 10747 4811
rect 11330 4808 11336 4820
rect 10689 4771 10747 4777
rect 11072 4780 11336 4808
rect 4080 4712 4752 4740
rect 1394 4672 1400 4684
rect 1355 4644 1400 4672
rect 1394 4632 1400 4644
rect 1452 4632 1458 4684
rect 2314 4672 2320 4684
rect 2275 4644 2320 4672
rect 2314 4632 2320 4644
rect 2372 4632 2378 4684
rect 2866 4632 2872 4684
rect 2924 4672 2930 4684
rect 2924 4644 3556 4672
rect 2924 4632 2930 4644
rect 2593 4607 2651 4613
rect 2593 4573 2605 4607
rect 2639 4604 2651 4607
rect 3142 4604 3148 4616
rect 2639 4576 3148 4604
rect 2639 4573 2651 4576
rect 2593 4567 2651 4573
rect 3142 4564 3148 4576
rect 3200 4564 3206 4616
rect 3528 4613 3556 4644
rect 3694 4632 3700 4684
rect 3752 4672 3758 4684
rect 4080 4672 4108 4712
rect 5902 4700 5908 4752
rect 5960 4740 5966 4752
rect 6362 4740 6368 4752
rect 5960 4712 6368 4740
rect 5960 4700 5966 4712
rect 6362 4700 6368 4712
rect 6420 4700 6426 4752
rect 7098 4700 7104 4752
rect 7156 4740 7162 4752
rect 8570 4740 8576 4752
rect 7156 4712 8576 4740
rect 7156 4700 7162 4712
rect 8570 4700 8576 4712
rect 8628 4700 8634 4752
rect 8757 4743 8815 4749
rect 8757 4709 8769 4743
rect 8803 4740 8815 4743
rect 9122 4740 9128 4752
rect 8803 4712 9128 4740
rect 8803 4709 8815 4712
rect 8757 4703 8815 4709
rect 9122 4700 9128 4712
rect 9180 4700 9186 4752
rect 10410 4700 10416 4752
rect 10468 4740 10474 4752
rect 10962 4740 10968 4752
rect 10468 4712 10968 4740
rect 10468 4700 10474 4712
rect 10962 4700 10968 4712
rect 11020 4700 11026 4752
rect 11072 4749 11100 4780
rect 11330 4768 11336 4780
rect 11388 4768 11394 4820
rect 11698 4808 11704 4820
rect 11659 4780 11704 4808
rect 11698 4768 11704 4780
rect 11756 4768 11762 4820
rect 12526 4808 12532 4820
rect 11808 4780 12532 4808
rect 11057 4743 11115 4749
rect 11057 4709 11069 4743
rect 11103 4709 11115 4743
rect 11057 4703 11115 4709
rect 11149 4743 11207 4749
rect 11149 4709 11161 4743
rect 11195 4709 11207 4743
rect 11149 4703 11207 4709
rect 3752 4644 4108 4672
rect 4157 4675 4215 4681
rect 3752 4632 3758 4644
rect 4157 4641 4169 4675
rect 4203 4672 4215 4675
rect 4982 4672 4988 4684
rect 4203 4644 4988 4672
rect 4203 4641 4215 4644
rect 4157 4635 4215 4641
rect 4982 4632 4988 4644
rect 5040 4632 5046 4684
rect 5169 4675 5227 4681
rect 5169 4641 5181 4675
rect 5215 4672 5227 4675
rect 6733 4675 6791 4681
rect 5215 4644 5764 4672
rect 5215 4641 5227 4644
rect 5169 4635 5227 4641
rect 5736 4616 5764 4644
rect 6196 4644 6592 4672
rect 3421 4607 3479 4613
rect 3421 4573 3433 4607
rect 3467 4573 3479 4607
rect 3421 4567 3479 4573
rect 3513 4607 3571 4613
rect 3513 4573 3525 4607
rect 3559 4573 3571 4607
rect 3513 4567 3571 4573
rect 1581 4539 1639 4545
rect 1581 4505 1593 4539
rect 1627 4536 1639 4539
rect 2958 4536 2964 4548
rect 1627 4508 2735 4536
rect 2919 4508 2964 4536
rect 1627 4505 1639 4508
rect 1581 4499 1639 4505
rect 1946 4468 1952 4480
rect 1907 4440 1952 4468
rect 1946 4428 1952 4440
rect 2004 4428 2010 4480
rect 2707 4468 2735 4508
rect 2958 4496 2964 4508
rect 3016 4496 3022 4548
rect 3436 4536 3464 4567
rect 3602 4564 3608 4616
rect 3660 4604 3666 4616
rect 5350 4604 5356 4616
rect 3660 4576 5212 4604
rect 5311 4576 5356 4604
rect 3660 4564 3666 4576
rect 4706 4536 4712 4548
rect 3436 4508 4712 4536
rect 4706 4496 4712 4508
rect 4764 4496 4770 4548
rect 5184 4536 5212 4576
rect 5350 4564 5356 4576
rect 5408 4564 5414 4616
rect 5718 4564 5724 4616
rect 5776 4564 5782 4616
rect 5810 4564 5816 4616
rect 5868 4604 5874 4616
rect 6196 4613 6224 4644
rect 6181 4607 6239 4613
rect 5868 4576 6132 4604
rect 5868 4564 5874 4576
rect 5442 4536 5448 4548
rect 5184 4508 5448 4536
rect 5442 4496 5448 4508
rect 5500 4496 5506 4548
rect 3142 4468 3148 4480
rect 2707 4440 3148 4468
rect 3142 4428 3148 4440
rect 3200 4428 3206 4480
rect 3786 4428 3792 4480
rect 3844 4468 3850 4480
rect 4341 4471 4399 4477
rect 4341 4468 4353 4471
rect 3844 4440 4353 4468
rect 3844 4428 3850 4440
rect 4341 4437 4353 4440
rect 4387 4437 4399 4471
rect 4341 4431 4399 4437
rect 5258 4428 5264 4480
rect 5316 4468 5322 4480
rect 5994 4468 6000 4480
rect 5316 4440 6000 4468
rect 5316 4428 5322 4440
rect 5994 4428 6000 4440
rect 6052 4428 6058 4480
rect 6104 4468 6132 4576
rect 6181 4573 6193 4607
rect 6227 4573 6239 4607
rect 6181 4567 6239 4573
rect 6273 4607 6331 4613
rect 6273 4573 6285 4607
rect 6319 4573 6331 4607
rect 6273 4567 6331 4573
rect 6288 4468 6316 4567
rect 6104 4440 6316 4468
rect 6564 4468 6592 4644
rect 6733 4641 6745 4675
rect 6779 4672 6791 4675
rect 6822 4672 6828 4684
rect 6779 4644 6828 4672
rect 6779 4641 6791 4644
rect 6733 4635 6791 4641
rect 6822 4632 6828 4644
rect 6880 4632 6886 4684
rect 7000 4675 7058 4681
rect 7000 4641 7012 4675
rect 7046 4672 7058 4675
rect 7926 4672 7932 4684
rect 7046 4644 7932 4672
rect 7046 4641 7058 4644
rect 7000 4635 7058 4641
rect 7926 4632 7932 4644
rect 7984 4632 7990 4684
rect 9950 4672 9956 4684
rect 8036 4644 9956 4672
rect 8036 4536 8064 4644
rect 9950 4632 9956 4644
rect 10008 4632 10014 4684
rect 10870 4672 10876 4684
rect 10336 4644 10876 4672
rect 8110 4564 8116 4616
rect 8168 4604 8174 4616
rect 8297 4607 8355 4613
rect 8297 4604 8309 4607
rect 8168 4576 8309 4604
rect 8168 4564 8174 4576
rect 8297 4573 8309 4576
rect 8343 4573 8355 4607
rect 8297 4567 8355 4573
rect 8849 4607 8907 4613
rect 8849 4573 8861 4607
rect 8895 4573 8907 4607
rect 8849 4567 8907 4573
rect 9033 4607 9091 4613
rect 9033 4573 9045 4607
rect 9079 4604 9091 4607
rect 9306 4604 9312 4616
rect 9079 4576 9312 4604
rect 9079 4573 9091 4576
rect 9033 4567 9091 4573
rect 7944 4508 8064 4536
rect 7944 4468 7972 4508
rect 8570 4496 8576 4548
rect 8628 4496 8634 4548
rect 8855 4536 8883 4567
rect 9306 4564 9312 4576
rect 9364 4564 9370 4616
rect 9766 4564 9772 4616
rect 9824 4604 9830 4616
rect 10229 4607 10287 4613
rect 10229 4604 10241 4607
rect 9824 4576 10241 4604
rect 9824 4564 9830 4576
rect 10229 4573 10241 4576
rect 10275 4573 10287 4607
rect 10229 4567 10287 4573
rect 9214 4536 9220 4548
rect 8855 4508 9220 4536
rect 9214 4496 9220 4508
rect 9272 4496 9278 4548
rect 9677 4539 9735 4545
rect 9677 4505 9689 4539
rect 9723 4536 9735 4539
rect 10336 4536 10364 4644
rect 10870 4632 10876 4644
rect 10928 4632 10934 4684
rect 11164 4672 11192 4703
rect 11238 4700 11244 4752
rect 11296 4740 11302 4752
rect 11808 4740 11836 4780
rect 12526 4768 12532 4780
rect 12584 4768 12590 4820
rect 12618 4768 12624 4820
rect 12676 4808 12682 4820
rect 14185 4811 14243 4817
rect 14185 4808 14197 4811
rect 12676 4780 14197 4808
rect 12676 4768 12682 4780
rect 14185 4777 14197 4780
rect 14231 4808 14243 4811
rect 15286 4808 15292 4820
rect 14231 4780 15292 4808
rect 14231 4777 14243 4780
rect 14185 4771 14243 4777
rect 15286 4768 15292 4780
rect 15344 4768 15350 4820
rect 12250 4740 12256 4752
rect 11296 4712 11836 4740
rect 11900 4712 12256 4740
rect 11296 4700 11302 4712
rect 11900 4672 11928 4712
rect 12250 4700 12256 4712
rect 12308 4700 12314 4752
rect 13170 4740 13176 4752
rect 12360 4712 13176 4740
rect 11164 4644 11928 4672
rect 11974 4632 11980 4684
rect 12032 4672 12038 4684
rect 12069 4675 12127 4681
rect 12069 4672 12081 4675
rect 12032 4644 12081 4672
rect 12032 4632 12038 4644
rect 12069 4641 12081 4644
rect 12115 4641 12127 4675
rect 12069 4635 12127 4641
rect 10594 4564 10600 4616
rect 10652 4604 10658 4616
rect 11330 4604 11336 4616
rect 10652 4576 11192 4604
rect 11291 4576 11336 4604
rect 10652 4564 10658 4576
rect 9723 4508 10364 4536
rect 11164 4536 11192 4576
rect 11330 4564 11336 4576
rect 11388 4564 11394 4616
rect 12161 4607 12219 4613
rect 12161 4604 12173 4607
rect 11440 4576 12173 4604
rect 11440 4536 11468 4576
rect 12161 4573 12173 4576
rect 12207 4573 12219 4607
rect 12161 4567 12219 4573
rect 12253 4607 12311 4613
rect 12253 4573 12265 4607
rect 12299 4573 12311 4607
rect 12253 4567 12311 4573
rect 11164 4508 11468 4536
rect 9723 4505 9735 4508
rect 9677 4499 9735 4505
rect 11606 4496 11612 4548
rect 11664 4536 11670 4548
rect 12268 4536 12296 4567
rect 11664 4508 12296 4536
rect 11664 4496 11670 4508
rect 8110 4468 8116 4480
rect 6564 4440 7972 4468
rect 8071 4440 8116 4468
rect 8110 4428 8116 4440
rect 8168 4428 8174 4480
rect 8297 4471 8355 4477
rect 8297 4437 8309 4471
rect 8343 4468 8355 4471
rect 8389 4471 8447 4477
rect 8389 4468 8401 4471
rect 8343 4440 8401 4468
rect 8343 4437 8355 4440
rect 8297 4431 8355 4437
rect 8389 4437 8401 4440
rect 8435 4437 8447 4471
rect 8588 4468 8616 4496
rect 10962 4468 10968 4480
rect 8588 4440 10968 4468
rect 8389 4431 8447 4437
rect 10962 4428 10968 4440
rect 11020 4428 11026 4480
rect 11054 4428 11060 4480
rect 11112 4468 11118 4480
rect 11330 4468 11336 4480
rect 11112 4440 11336 4468
rect 11112 4428 11118 4440
rect 11330 4428 11336 4440
rect 11388 4468 11394 4480
rect 12360 4468 12388 4712
rect 13170 4700 13176 4712
rect 13228 4700 13234 4752
rect 12894 4672 12900 4684
rect 12855 4644 12900 4672
rect 12894 4632 12900 4644
rect 12952 4632 12958 4684
rect 13538 4672 13544 4684
rect 13499 4644 13544 4672
rect 13538 4632 13544 4644
rect 13596 4672 13602 4684
rect 14093 4675 14151 4681
rect 14093 4672 14105 4675
rect 13596 4644 14105 4672
rect 13596 4632 13602 4644
rect 14093 4641 14105 4644
rect 14139 4641 14151 4675
rect 14093 4635 14151 4641
rect 12986 4604 12992 4616
rect 12947 4576 12992 4604
rect 12986 4564 12992 4576
rect 13044 4564 13050 4616
rect 13081 4607 13139 4613
rect 13081 4573 13093 4607
rect 13127 4573 13139 4607
rect 13081 4567 13139 4573
rect 12894 4496 12900 4548
rect 12952 4536 12958 4548
rect 13096 4536 13124 4567
rect 13722 4564 13728 4616
rect 13780 4604 13786 4616
rect 14277 4607 14335 4613
rect 14277 4604 14289 4607
rect 13780 4576 14289 4604
rect 13780 4564 13786 4576
rect 14277 4573 14289 4576
rect 14323 4604 14335 4607
rect 14918 4604 14924 4616
rect 14323 4576 14924 4604
rect 14323 4573 14335 4576
rect 14277 4567 14335 4573
rect 14918 4564 14924 4576
rect 14976 4564 14982 4616
rect 12952 4508 13124 4536
rect 12952 4496 12958 4508
rect 12526 4468 12532 4480
rect 11388 4440 12388 4468
rect 12487 4440 12532 4468
rect 11388 4428 11394 4440
rect 12526 4428 12532 4440
rect 12584 4428 12590 4480
rect 12618 4428 12624 4480
rect 12676 4468 12682 4480
rect 13725 4471 13783 4477
rect 13725 4468 13737 4471
rect 12676 4440 13737 4468
rect 12676 4428 12682 4440
rect 13725 4437 13737 4440
rect 13771 4437 13783 4471
rect 13725 4431 13783 4437
rect 1104 4378 15824 4400
rect 1104 4326 3447 4378
rect 3499 4326 3511 4378
rect 3563 4326 3575 4378
rect 3627 4326 3639 4378
rect 3691 4326 8378 4378
rect 8430 4326 8442 4378
rect 8494 4326 8506 4378
rect 8558 4326 8570 4378
rect 8622 4326 13308 4378
rect 13360 4326 13372 4378
rect 13424 4326 13436 4378
rect 13488 4326 13500 4378
rect 13552 4326 15824 4378
rect 1104 4304 15824 4326
rect 2222 4224 2228 4276
rect 2280 4264 2286 4276
rect 2280 4236 4108 4264
rect 2280 4224 2286 4236
rect 4080 4205 4108 4236
rect 4706 4224 4712 4276
rect 4764 4264 4770 4276
rect 5350 4264 5356 4276
rect 4764 4236 5356 4264
rect 4764 4224 4770 4236
rect 4065 4199 4123 4205
rect 4065 4165 4077 4199
rect 4111 4196 4123 4199
rect 4338 4196 4344 4208
rect 4111 4168 4344 4196
rect 4111 4165 4123 4168
rect 4065 4159 4123 4165
rect 4338 4156 4344 4168
rect 4396 4156 4402 4208
rect 2317 4131 2375 4137
rect 2317 4097 2329 4131
rect 2363 4128 2375 4131
rect 2363 4100 2820 4128
rect 2363 4097 2375 4100
rect 2317 4091 2375 4097
rect 2041 4063 2099 4069
rect 2041 4029 2053 4063
rect 2087 4060 2099 4063
rect 2130 4060 2136 4072
rect 2087 4032 2136 4060
rect 2087 4029 2099 4032
rect 2041 4023 2099 4029
rect 2130 4020 2136 4032
rect 2188 4020 2194 4072
rect 2682 4060 2688 4072
rect 2643 4032 2688 4060
rect 2682 4020 2688 4032
rect 2740 4020 2746 4072
rect 2792 4060 2820 4100
rect 4154 4088 4160 4140
rect 4212 4128 4218 4140
rect 4890 4128 4896 4140
rect 4212 4100 4896 4128
rect 4212 4088 4218 4100
rect 4890 4088 4896 4100
rect 4948 4088 4954 4140
rect 5184 4137 5212 4236
rect 5350 4224 5356 4236
rect 5408 4224 5414 4276
rect 5442 4224 5448 4276
rect 5500 4264 5506 4276
rect 5537 4267 5595 4273
rect 5537 4264 5549 4267
rect 5500 4236 5549 4264
rect 5500 4224 5506 4236
rect 5537 4233 5549 4236
rect 5583 4233 5595 4267
rect 5718 4264 5724 4276
rect 5679 4236 5724 4264
rect 5537 4227 5595 4233
rect 5718 4224 5724 4236
rect 5776 4224 5782 4276
rect 6362 4224 6368 4276
rect 6420 4264 6426 4276
rect 8481 4267 8539 4273
rect 8481 4264 8493 4267
rect 6420 4236 8493 4264
rect 6420 4224 6426 4236
rect 8481 4233 8493 4236
rect 8527 4233 8539 4267
rect 8481 4227 8539 4233
rect 8938 4224 8944 4276
rect 8996 4264 9002 4276
rect 9309 4267 9367 4273
rect 9309 4264 9321 4267
rect 8996 4236 9321 4264
rect 8996 4224 9002 4236
rect 9309 4233 9321 4236
rect 9355 4233 9367 4267
rect 9490 4264 9496 4276
rect 9451 4236 9496 4264
rect 9309 4227 9367 4233
rect 9490 4224 9496 4236
rect 9548 4224 9554 4276
rect 9766 4224 9772 4276
rect 9824 4264 9830 4276
rect 9824 4236 10916 4264
rect 9824 4224 9830 4236
rect 5902 4196 5908 4208
rect 5368 4168 5908 4196
rect 5368 4137 5396 4168
rect 5902 4156 5908 4168
rect 5960 4156 5966 4208
rect 6730 4196 6736 4208
rect 6472 4168 6736 4196
rect 5169 4131 5227 4137
rect 5169 4097 5181 4131
rect 5215 4097 5227 4131
rect 5169 4091 5227 4097
rect 5353 4131 5411 4137
rect 5353 4097 5365 4131
rect 5399 4097 5411 4131
rect 5353 4091 5411 4097
rect 5537 4131 5595 4137
rect 5537 4097 5549 4131
rect 5583 4128 5595 4131
rect 5810 4128 5816 4140
rect 5583 4100 5816 4128
rect 5583 4097 5595 4100
rect 5537 4091 5595 4097
rect 5810 4088 5816 4100
rect 5868 4088 5874 4140
rect 6362 4128 6368 4140
rect 6323 4100 6368 4128
rect 6362 4088 6368 4100
rect 6420 4088 6426 4140
rect 4617 4063 4675 4069
rect 2792 4032 3648 4060
rect 2148 3992 2176 4020
rect 3620 4004 3648 4032
rect 4617 4029 4629 4063
rect 4663 4060 4675 4063
rect 6181 4063 6239 4069
rect 4663 4032 6132 4060
rect 4663 4029 4675 4032
rect 4617 4023 4675 4029
rect 2148 3964 2735 3992
rect 1670 3924 1676 3936
rect 1631 3896 1676 3924
rect 1670 3884 1676 3896
rect 1728 3884 1734 3936
rect 2130 3884 2136 3936
rect 2188 3924 2194 3936
rect 2707 3924 2735 3964
rect 2774 3952 2780 4004
rect 2832 3992 2838 4004
rect 2930 3995 2988 4001
rect 2930 3992 2942 3995
rect 2832 3964 2942 3992
rect 2832 3952 2838 3964
rect 2930 3961 2942 3964
rect 2976 3961 2988 3995
rect 2930 3955 2988 3961
rect 3602 3952 3608 4004
rect 3660 3952 3666 4004
rect 5718 3992 5724 4004
rect 4724 3964 5724 3992
rect 4154 3924 4160 3936
rect 2188 3896 2233 3924
rect 2707 3896 4160 3924
rect 2188 3884 2194 3896
rect 4154 3884 4160 3896
rect 4212 3884 4218 3936
rect 4246 3884 4252 3936
rect 4304 3924 4310 3936
rect 4724 3933 4752 3964
rect 5718 3952 5724 3964
rect 5776 3952 5782 4004
rect 6104 3992 6132 4032
rect 6181 4029 6193 4063
rect 6227 4060 6239 4063
rect 6472 4060 6500 4168
rect 6730 4156 6736 4168
rect 6788 4156 6794 4208
rect 8110 4156 8116 4208
rect 8168 4196 8174 4208
rect 10318 4196 10324 4208
rect 8168 4168 10180 4196
rect 8168 4156 8174 4168
rect 10152 4140 10180 4168
rect 10235 4168 10324 4196
rect 6822 4128 6828 4140
rect 6783 4100 6828 4128
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 8754 4088 8760 4140
rect 8812 4128 8818 4140
rect 8938 4128 8944 4140
rect 8812 4100 8944 4128
rect 8812 4088 8818 4100
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 9125 4131 9183 4137
rect 9125 4097 9137 4131
rect 9171 4128 9183 4131
rect 9582 4128 9588 4140
rect 9171 4100 9588 4128
rect 9171 4097 9183 4100
rect 9125 4091 9183 4097
rect 9582 4088 9588 4100
rect 9640 4088 9646 4140
rect 10134 4128 10140 4140
rect 10095 4100 10140 4128
rect 10134 4088 10140 4100
rect 10192 4088 10198 4140
rect 7374 4060 7380 4072
rect 6227 4032 6500 4060
rect 6932 4032 7380 4060
rect 6227 4029 6239 4032
rect 6181 4023 6239 4029
rect 6932 3992 6960 4032
rect 7374 4020 7380 4032
rect 7432 4020 7438 4072
rect 7650 4020 7656 4072
rect 7708 4060 7714 4072
rect 9766 4060 9772 4072
rect 7708 4032 9772 4060
rect 7708 4020 7714 4032
rect 9766 4020 9772 4032
rect 9824 4020 9830 4072
rect 9861 4063 9919 4069
rect 9861 4029 9873 4063
rect 9907 4060 9919 4063
rect 10235 4060 10263 4168
rect 10318 4156 10324 4168
rect 10376 4156 10382 4208
rect 10502 4196 10508 4208
rect 10463 4168 10508 4196
rect 10502 4156 10508 4168
rect 10560 4156 10566 4208
rect 10888 4196 10916 4236
rect 10962 4224 10968 4276
rect 11020 4264 11026 4276
rect 12066 4264 12072 4276
rect 11020 4236 12072 4264
rect 11020 4224 11026 4236
rect 12066 4224 12072 4236
rect 12124 4224 12130 4276
rect 12360 4236 13860 4264
rect 11054 4196 11060 4208
rect 10888 4168 11060 4196
rect 11054 4156 11060 4168
rect 11112 4156 11118 4208
rect 11330 4196 11336 4208
rect 11164 4168 11336 4196
rect 11164 4137 11192 4168
rect 11330 4156 11336 4168
rect 11388 4196 11394 4208
rect 11606 4196 11612 4208
rect 11388 4168 11612 4196
rect 11388 4156 11394 4168
rect 11606 4156 11612 4168
rect 11664 4156 11670 4208
rect 10413 4131 10471 4137
rect 10413 4097 10425 4131
rect 10459 4128 10471 4131
rect 11149 4131 11207 4137
rect 10459 4100 11008 4128
rect 10459 4097 10471 4100
rect 10413 4091 10471 4097
rect 9907 4032 10263 4060
rect 9907 4029 9919 4032
rect 9861 4023 9919 4029
rect 10318 4020 10324 4072
rect 10376 4060 10382 4072
rect 10594 4060 10600 4072
rect 10376 4032 10600 4060
rect 10376 4020 10382 4032
rect 10594 4020 10600 4032
rect 10652 4020 10658 4072
rect 10778 4020 10784 4072
rect 10836 4060 10842 4072
rect 10873 4063 10931 4069
rect 10873 4060 10885 4063
rect 10836 4032 10885 4060
rect 10836 4020 10842 4032
rect 10873 4029 10885 4032
rect 10919 4029 10931 4063
rect 10980 4060 11008 4100
rect 11149 4097 11161 4131
rect 11195 4097 11207 4131
rect 11149 4091 11207 4097
rect 11422 4088 11428 4140
rect 11480 4088 11486 4140
rect 12360 4128 12388 4236
rect 12802 4156 12808 4208
rect 12860 4196 12866 4208
rect 13832 4196 13860 4236
rect 13906 4224 13912 4276
rect 13964 4264 13970 4276
rect 14461 4267 14519 4273
rect 14461 4264 14473 4267
rect 13964 4236 14473 4264
rect 13964 4224 13970 4236
rect 14461 4233 14473 4236
rect 14507 4233 14519 4267
rect 14461 4227 14519 4233
rect 15194 4196 15200 4208
rect 12860 4168 13032 4196
rect 13832 4168 15200 4196
rect 12860 4156 12866 4168
rect 11624 4100 12388 4128
rect 11440 4060 11468 4088
rect 10980 4032 11468 4060
rect 11523 4063 11581 4069
rect 10873 4023 10931 4029
rect 11523 4029 11535 4063
rect 11569 4060 11581 4063
rect 11624 4060 11652 4100
rect 12434 4088 12440 4140
rect 12492 4128 12498 4140
rect 13004 4137 13032 4168
rect 12989 4131 13047 4137
rect 12492 4100 12848 4128
rect 12492 4088 12498 4100
rect 12710 4060 12716 4072
rect 11569 4032 11652 4060
rect 11716 4032 12716 4060
rect 11569 4029 11581 4032
rect 11523 4023 11581 4029
rect 7098 4001 7104 4004
rect 7092 3992 7104 4001
rect 6104 3964 6960 3992
rect 7059 3964 7104 3992
rect 7092 3955 7104 3964
rect 7098 3952 7104 3955
rect 7156 3952 7162 4004
rect 7466 3952 7472 4004
rect 7524 3992 7530 4004
rect 8849 3995 8907 4001
rect 7524 3964 8340 3992
rect 7524 3952 7530 3964
rect 4433 3927 4491 3933
rect 4433 3924 4445 3927
rect 4304 3896 4445 3924
rect 4304 3884 4310 3896
rect 4433 3893 4445 3896
rect 4479 3893 4491 3927
rect 4433 3887 4491 3893
rect 4709 3927 4767 3933
rect 4709 3893 4721 3927
rect 4755 3893 4767 3927
rect 4709 3887 4767 3893
rect 4890 3884 4896 3936
rect 4948 3924 4954 3936
rect 5077 3927 5135 3933
rect 5077 3924 5089 3927
rect 4948 3896 5089 3924
rect 4948 3884 4954 3896
rect 5077 3893 5089 3896
rect 5123 3924 5135 3927
rect 5537 3927 5595 3933
rect 5537 3924 5549 3927
rect 5123 3896 5549 3924
rect 5123 3893 5135 3896
rect 5077 3887 5135 3893
rect 5537 3893 5549 3896
rect 5583 3893 5595 3927
rect 5537 3887 5595 3893
rect 5629 3927 5687 3933
rect 5629 3893 5641 3927
rect 5675 3924 5687 3927
rect 6089 3927 6147 3933
rect 6089 3924 6101 3927
rect 5675 3896 6101 3924
rect 5675 3893 5687 3896
rect 5629 3887 5687 3893
rect 6089 3893 6101 3896
rect 6135 3893 6147 3927
rect 6089 3887 6147 3893
rect 6270 3884 6276 3936
rect 6328 3924 6334 3936
rect 8110 3924 8116 3936
rect 6328 3896 8116 3924
rect 6328 3884 6334 3896
rect 8110 3884 8116 3896
rect 8168 3924 8174 3936
rect 8205 3927 8263 3933
rect 8205 3924 8217 3927
rect 8168 3896 8217 3924
rect 8168 3884 8174 3896
rect 8205 3893 8217 3896
rect 8251 3893 8263 3927
rect 8312 3924 8340 3964
rect 8849 3961 8861 3995
rect 8895 3992 8907 3995
rect 9309 3995 9367 4001
rect 9309 3992 9321 3995
rect 8895 3964 9321 3992
rect 8895 3961 8907 3964
rect 8849 3955 8907 3961
rect 9309 3961 9321 3964
rect 9355 3992 9367 3995
rect 9490 3992 9496 4004
rect 9355 3964 9496 3992
rect 9355 3961 9367 3964
rect 9309 3955 9367 3961
rect 9490 3952 9496 3964
rect 9548 3952 9554 4004
rect 9953 3995 10011 4001
rect 9953 3961 9965 3995
rect 9999 3992 10011 3995
rect 11716 3992 11744 4032
rect 12710 4020 12716 4032
rect 12768 4020 12774 4072
rect 12820 4060 12848 4100
rect 12989 4097 13001 4131
rect 13035 4097 13047 4131
rect 12989 4091 13047 4097
rect 13538 4088 13544 4140
rect 13596 4128 13602 4140
rect 14001 4131 14059 4137
rect 14001 4128 14013 4131
rect 13596 4100 14013 4128
rect 13596 4088 13602 4100
rect 14001 4097 14013 4100
rect 14047 4097 14059 4131
rect 14001 4091 14059 4097
rect 13354 4060 13360 4072
rect 12820 4032 13360 4060
rect 13354 4020 13360 4032
rect 13412 4020 13418 4072
rect 13906 4060 13912 4072
rect 13867 4032 13912 4060
rect 13906 4020 13912 4032
rect 13964 4020 13970 4072
rect 9999 3964 11744 3992
rect 9999 3961 10011 3964
rect 9953 3955 10011 3961
rect 11790 3952 11796 4004
rect 11848 3992 11854 4004
rect 14844 4001 14872 4168
rect 15194 4156 15200 4168
rect 15252 4156 15258 4208
rect 14918 4088 14924 4140
rect 14976 4128 14982 4140
rect 15013 4131 15071 4137
rect 15013 4128 15025 4131
rect 14976 4100 15025 4128
rect 14976 4088 14982 4100
rect 15013 4097 15025 4100
rect 15059 4097 15071 4131
rect 15013 4091 15071 4097
rect 12805 3995 12863 4001
rect 12805 3992 12817 3995
rect 11848 3964 12817 3992
rect 11848 3952 11854 3964
rect 12805 3961 12817 3964
rect 12851 3961 12863 3995
rect 12805 3955 12863 3961
rect 14829 3995 14887 4001
rect 14829 3961 14841 3995
rect 14875 3961 14887 3995
rect 14829 3955 14887 3961
rect 8941 3927 8999 3933
rect 8941 3924 8953 3927
rect 8312 3896 8953 3924
rect 8205 3887 8263 3893
rect 8941 3893 8953 3896
rect 8987 3893 8999 3927
rect 8941 3887 8999 3893
rect 9122 3884 9128 3936
rect 9180 3924 9186 3936
rect 9766 3924 9772 3936
rect 9180 3896 9772 3924
rect 9180 3884 9186 3896
rect 9766 3884 9772 3896
rect 9824 3884 9830 3936
rect 9858 3884 9864 3936
rect 9916 3924 9922 3936
rect 10413 3927 10471 3933
rect 10413 3924 10425 3927
rect 9916 3896 10425 3924
rect 9916 3884 9922 3896
rect 10413 3893 10425 3896
rect 10459 3893 10471 3927
rect 10413 3887 10471 3893
rect 10594 3884 10600 3936
rect 10652 3924 10658 3936
rect 10965 3927 11023 3933
rect 10965 3924 10977 3927
rect 10652 3896 10977 3924
rect 10652 3884 10658 3896
rect 10965 3893 10977 3896
rect 11011 3893 11023 3927
rect 10965 3887 11023 3893
rect 11422 3884 11428 3936
rect 11480 3924 11486 3936
rect 11701 3927 11759 3933
rect 11701 3924 11713 3927
rect 11480 3896 11713 3924
rect 11480 3884 11486 3896
rect 11701 3893 11713 3896
rect 11747 3893 11759 3927
rect 11701 3887 11759 3893
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 12492 3896 12537 3924
rect 12492 3884 12498 3896
rect 12710 3884 12716 3936
rect 12768 3924 12774 3936
rect 12897 3927 12955 3933
rect 12897 3924 12909 3927
rect 12768 3896 12909 3924
rect 12768 3884 12774 3896
rect 12897 3893 12909 3896
rect 12943 3893 12955 3927
rect 12897 3887 12955 3893
rect 12986 3884 12992 3936
rect 13044 3924 13050 3936
rect 13449 3927 13507 3933
rect 13449 3924 13461 3927
rect 13044 3896 13461 3924
rect 13044 3884 13050 3896
rect 13449 3893 13461 3896
rect 13495 3893 13507 3927
rect 13449 3887 13507 3893
rect 13722 3884 13728 3936
rect 13780 3924 13786 3936
rect 13817 3927 13875 3933
rect 13817 3924 13829 3927
rect 13780 3896 13829 3924
rect 13780 3884 13786 3896
rect 13817 3893 13829 3896
rect 13863 3893 13875 3927
rect 13817 3887 13875 3893
rect 14550 3884 14556 3936
rect 14608 3924 14614 3936
rect 14921 3927 14979 3933
rect 14921 3924 14933 3927
rect 14608 3896 14933 3924
rect 14608 3884 14614 3896
rect 14921 3893 14933 3896
rect 14967 3924 14979 3927
rect 15102 3924 15108 3936
rect 14967 3896 15108 3924
rect 14967 3893 14979 3896
rect 14921 3887 14979 3893
rect 15102 3884 15108 3896
rect 15160 3884 15166 3936
rect 1104 3834 15824 3856
rect 1104 3782 5912 3834
rect 5964 3782 5976 3834
rect 6028 3782 6040 3834
rect 6092 3782 6104 3834
rect 6156 3782 10843 3834
rect 10895 3782 10907 3834
rect 10959 3782 10971 3834
rect 11023 3782 11035 3834
rect 11087 3782 15824 3834
rect 1104 3760 15824 3782
rect 1949 3723 2007 3729
rect 1949 3689 1961 3723
rect 1995 3689 2007 3723
rect 1949 3683 2007 3689
rect 2961 3723 3019 3729
rect 2961 3689 2973 3723
rect 3007 3720 3019 3723
rect 3050 3720 3056 3732
rect 3007 3692 3056 3720
rect 3007 3689 3019 3692
rect 2961 3683 3019 3689
rect 1964 3652 1992 3683
rect 3050 3680 3056 3692
rect 3108 3680 3114 3732
rect 3418 3720 3424 3732
rect 3379 3692 3424 3720
rect 3418 3680 3424 3692
rect 3476 3680 3482 3732
rect 4798 3720 4804 3732
rect 4759 3692 4804 3720
rect 4798 3680 4804 3692
rect 4856 3680 4862 3732
rect 5442 3680 5448 3732
rect 5500 3720 5506 3732
rect 6270 3720 6276 3732
rect 5500 3692 6276 3720
rect 5500 3680 5506 3692
rect 6270 3680 6276 3692
rect 6328 3680 6334 3732
rect 6457 3723 6515 3729
rect 6457 3689 6469 3723
rect 6503 3720 6515 3723
rect 6822 3720 6828 3732
rect 6503 3692 6828 3720
rect 6503 3689 6515 3692
rect 6457 3683 6515 3689
rect 6822 3680 6828 3692
rect 6880 3680 6886 3732
rect 7101 3723 7159 3729
rect 7101 3720 7113 3723
rect 7011 3692 7113 3720
rect 7101 3689 7113 3692
rect 7147 3720 7159 3723
rect 7282 3720 7288 3732
rect 7147 3692 7288 3720
rect 7147 3689 7159 3692
rect 7101 3683 7159 3689
rect 1964 3624 3096 3652
rect 1394 3584 1400 3596
rect 1355 3556 1400 3584
rect 1394 3544 1400 3556
rect 1452 3544 1458 3596
rect 2317 3587 2375 3593
rect 2317 3553 2329 3587
rect 2363 3584 2375 3587
rect 2866 3584 2872 3596
rect 2363 3556 2872 3584
rect 2363 3553 2375 3556
rect 2317 3547 2375 3553
rect 2866 3544 2872 3556
rect 2924 3544 2930 3596
rect 2409 3519 2467 3525
rect 2409 3485 2421 3519
rect 2455 3485 2467 3519
rect 2409 3479 2467 3485
rect 2593 3519 2651 3525
rect 2593 3485 2605 3519
rect 2639 3516 2651 3519
rect 2958 3516 2964 3528
rect 2639 3488 2964 3516
rect 2639 3485 2651 3488
rect 2593 3479 2651 3485
rect 2424 3448 2452 3479
rect 2958 3476 2964 3488
rect 3016 3476 3022 3528
rect 3068 3516 3096 3624
rect 4614 3612 4620 3664
rect 4672 3652 4678 3664
rect 4709 3655 4767 3661
rect 4709 3652 4721 3655
rect 4672 3624 4721 3652
rect 4672 3612 4678 3624
rect 4709 3621 4721 3624
rect 4755 3621 4767 3655
rect 4709 3615 4767 3621
rect 5626 3612 5632 3664
rect 5684 3652 5690 3664
rect 5721 3655 5779 3661
rect 5721 3652 5733 3655
rect 5684 3624 5733 3652
rect 5684 3612 5690 3624
rect 5721 3621 5733 3624
rect 5767 3621 5779 3655
rect 5721 3615 5779 3621
rect 5810 3612 5816 3664
rect 5868 3652 5874 3664
rect 7116 3652 7144 3683
rect 7282 3680 7288 3692
rect 7340 3680 7346 3732
rect 7742 3720 7748 3732
rect 7703 3692 7748 3720
rect 7742 3680 7748 3692
rect 7800 3680 7806 3732
rect 7834 3680 7840 3732
rect 7892 3720 7898 3732
rect 7892 3692 9260 3720
rect 7892 3680 7898 3692
rect 5868 3624 7144 3652
rect 7193 3655 7251 3661
rect 5868 3612 5874 3624
rect 7193 3621 7205 3655
rect 7239 3652 7251 3655
rect 8938 3652 8944 3664
rect 7239 3624 8944 3652
rect 7239 3621 7251 3624
rect 7193 3615 7251 3621
rect 3326 3584 3332 3596
rect 3287 3556 3332 3584
rect 3326 3544 3332 3556
rect 3384 3544 3390 3596
rect 4062 3584 4068 3596
rect 3436 3556 4068 3584
rect 3436 3516 3464 3556
rect 4062 3544 4068 3556
rect 4120 3544 4126 3596
rect 4246 3544 4252 3596
rect 4304 3584 4310 3596
rect 6641 3587 6699 3593
rect 6641 3584 6653 3587
rect 4304 3556 6653 3584
rect 4304 3544 4310 3556
rect 6641 3553 6653 3556
rect 6687 3553 6699 3587
rect 7208 3584 7236 3615
rect 8938 3612 8944 3624
rect 8996 3652 9002 3664
rect 9122 3652 9128 3664
rect 8996 3624 9128 3652
rect 8996 3612 9002 3624
rect 9122 3612 9128 3624
rect 9180 3612 9186 3664
rect 9232 3652 9260 3692
rect 9674 3680 9680 3732
rect 9732 3720 9738 3732
rect 9732 3692 9777 3720
rect 9732 3680 9738 3692
rect 9950 3680 9956 3732
rect 10008 3720 10014 3732
rect 10318 3720 10324 3732
rect 10008 3692 10324 3720
rect 10008 3680 10014 3692
rect 10318 3680 10324 3692
rect 10376 3680 10382 3732
rect 10410 3680 10416 3732
rect 10468 3720 10474 3732
rect 11057 3723 11115 3729
rect 11057 3720 11069 3723
rect 10468 3692 11069 3720
rect 10468 3680 10474 3692
rect 11057 3689 11069 3692
rect 11103 3689 11115 3723
rect 11057 3683 11115 3689
rect 11146 3680 11152 3732
rect 11204 3720 11210 3732
rect 11606 3720 11612 3732
rect 11204 3692 11612 3720
rect 11204 3680 11210 3692
rect 11606 3680 11612 3692
rect 11664 3680 11670 3732
rect 11701 3723 11759 3729
rect 11701 3689 11713 3723
rect 11747 3720 11759 3723
rect 11790 3720 11796 3732
rect 11747 3692 11796 3720
rect 11747 3689 11759 3692
rect 11701 3683 11759 3689
rect 11790 3680 11796 3692
rect 11848 3680 11854 3732
rect 12161 3723 12219 3729
rect 12161 3689 12173 3723
rect 12207 3720 12219 3723
rect 12250 3720 12256 3732
rect 12207 3692 12256 3720
rect 12207 3689 12219 3692
rect 12161 3683 12219 3689
rect 12250 3680 12256 3692
rect 12308 3680 12314 3732
rect 12526 3680 12532 3732
rect 12584 3720 12590 3732
rect 12710 3720 12716 3732
rect 12584 3692 12716 3720
rect 12584 3680 12590 3692
rect 12710 3680 12716 3692
rect 12768 3680 12774 3732
rect 12894 3680 12900 3732
rect 12952 3720 12958 3732
rect 13170 3720 13176 3732
rect 12952 3692 13176 3720
rect 12952 3680 12958 3692
rect 13170 3680 13176 3692
rect 13228 3680 13234 3732
rect 13354 3680 13360 3732
rect 13412 3720 13418 3732
rect 13725 3723 13783 3729
rect 13725 3720 13737 3723
rect 13412 3692 13737 3720
rect 13412 3680 13418 3692
rect 13725 3689 13737 3692
rect 13771 3689 13783 3723
rect 13725 3683 13783 3689
rect 14093 3723 14151 3729
rect 14093 3689 14105 3723
rect 14139 3720 14151 3723
rect 14550 3720 14556 3732
rect 14139 3692 14556 3720
rect 14139 3689 14151 3692
rect 14093 3683 14151 3689
rect 14550 3680 14556 3692
rect 14608 3720 14614 3732
rect 14826 3720 14832 3732
rect 14608 3692 14832 3720
rect 14608 3680 14614 3692
rect 14826 3680 14832 3692
rect 14884 3680 14890 3732
rect 9858 3652 9864 3664
rect 9232 3624 9864 3652
rect 9858 3612 9864 3624
rect 9916 3612 9922 3664
rect 10045 3655 10103 3661
rect 10045 3621 10057 3655
rect 10091 3652 10103 3655
rect 13906 3652 13912 3664
rect 10091 3624 13912 3652
rect 10091 3621 10103 3624
rect 10045 3615 10103 3621
rect 6641 3547 6699 3553
rect 6748 3556 7236 3584
rect 3602 3516 3608 3528
rect 3068 3488 3464 3516
rect 3563 3488 3608 3516
rect 3602 3476 3608 3488
rect 3660 3476 3666 3528
rect 4982 3516 4988 3528
rect 4943 3488 4988 3516
rect 4982 3476 4988 3488
rect 5040 3476 5046 3528
rect 5350 3476 5356 3528
rect 5408 3516 5414 3528
rect 5810 3516 5816 3528
rect 5408 3488 5672 3516
rect 5771 3488 5816 3516
rect 5408 3476 5414 3488
rect 3234 3448 3240 3460
rect 2424 3420 3240 3448
rect 3234 3408 3240 3420
rect 3292 3408 3298 3460
rect 4154 3408 4160 3460
rect 4212 3448 4218 3460
rect 5644 3448 5672 3488
rect 5810 3476 5816 3488
rect 5868 3476 5874 3528
rect 5997 3519 6055 3525
rect 5997 3485 6009 3519
rect 6043 3516 6055 3519
rect 6546 3516 6552 3528
rect 6043 3488 6552 3516
rect 6043 3485 6055 3488
rect 5997 3479 6055 3485
rect 6546 3476 6552 3488
rect 6604 3476 6610 3528
rect 6748 3516 6776 3556
rect 7650 3544 7656 3596
rect 7708 3584 7714 3596
rect 8113 3587 8171 3593
rect 8113 3584 8125 3587
rect 7708 3556 8125 3584
rect 7708 3544 7714 3556
rect 8113 3553 8125 3556
rect 8159 3584 8171 3587
rect 8757 3587 8815 3593
rect 8159 3556 8708 3584
rect 8159 3553 8171 3556
rect 8113 3547 8171 3553
rect 7285 3519 7343 3525
rect 7285 3516 7297 3519
rect 6656 3488 6776 3516
rect 7208 3488 7297 3516
rect 6656 3448 6684 3488
rect 4212 3420 5580 3448
rect 5644 3420 6684 3448
rect 4212 3408 4218 3420
rect 198 3340 204 3392
rect 256 3380 262 3392
rect 1581 3383 1639 3389
rect 1581 3380 1593 3383
rect 256 3352 1593 3380
rect 256 3340 262 3352
rect 1581 3349 1593 3352
rect 1627 3349 1639 3383
rect 1581 3343 1639 3349
rect 2498 3340 2504 3392
rect 2556 3380 2562 3392
rect 4246 3380 4252 3392
rect 2556 3352 4252 3380
rect 2556 3340 2562 3352
rect 4246 3340 4252 3352
rect 4304 3340 4310 3392
rect 4341 3383 4399 3389
rect 4341 3349 4353 3383
rect 4387 3380 4399 3383
rect 4982 3380 4988 3392
rect 4387 3352 4988 3380
rect 4387 3349 4399 3352
rect 4341 3343 4399 3349
rect 4982 3340 4988 3352
rect 5040 3340 5046 3392
rect 5350 3380 5356 3392
rect 5311 3352 5356 3380
rect 5350 3340 5356 3352
rect 5408 3340 5414 3392
rect 5552 3380 5580 3420
rect 6730 3408 6736 3460
rect 6788 3448 6794 3460
rect 6788 3420 6833 3448
rect 6788 3408 6794 3420
rect 6914 3408 6920 3460
rect 6972 3448 6978 3460
rect 7208 3448 7236 3488
rect 7285 3485 7297 3488
rect 7331 3485 7343 3519
rect 8205 3519 8263 3525
rect 8205 3516 8217 3519
rect 7285 3479 7343 3485
rect 7392 3488 8217 3516
rect 6972 3420 7236 3448
rect 6972 3408 6978 3420
rect 7392 3380 7420 3488
rect 8205 3485 8217 3488
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 8294 3476 8300 3528
rect 8352 3516 8358 3528
rect 8680 3516 8708 3556
rect 8757 3553 8769 3587
rect 8803 3584 8815 3587
rect 10060 3584 10088 3615
rect 13906 3612 13912 3624
rect 13964 3612 13970 3664
rect 14185 3655 14243 3661
rect 14185 3621 14197 3655
rect 14231 3652 14243 3655
rect 14274 3652 14280 3664
rect 14231 3624 14280 3652
rect 14231 3621 14243 3624
rect 14185 3615 14243 3621
rect 14274 3612 14280 3624
rect 14332 3612 14338 3664
rect 14918 3612 14924 3664
rect 14976 3612 14982 3664
rect 11330 3584 11336 3596
rect 8803 3556 10088 3584
rect 10336 3556 11336 3584
rect 8803 3553 8815 3556
rect 8757 3547 8815 3553
rect 9214 3516 9220 3528
rect 8352 3488 8397 3516
rect 8680 3488 9220 3516
rect 8352 3476 8358 3488
rect 9214 3476 9220 3488
rect 9272 3476 9278 3528
rect 9306 3476 9312 3528
rect 9364 3516 9370 3528
rect 10336 3525 10364 3556
rect 11330 3544 11336 3556
rect 11388 3544 11394 3596
rect 11882 3544 11888 3596
rect 11940 3584 11946 3596
rect 12069 3587 12127 3593
rect 12069 3584 12081 3587
rect 11940 3556 12081 3584
rect 11940 3544 11946 3556
rect 12069 3553 12081 3556
rect 12115 3553 12127 3587
rect 13081 3587 13139 3593
rect 13081 3584 13093 3587
rect 12069 3547 12127 3553
rect 12544 3556 13093 3584
rect 10137 3519 10195 3525
rect 9364 3488 9812 3516
rect 9364 3476 9370 3488
rect 7650 3408 7656 3460
rect 7708 3448 7714 3460
rect 8941 3451 8999 3457
rect 8941 3448 8953 3451
rect 7708 3420 8953 3448
rect 7708 3408 7714 3420
rect 8941 3417 8953 3420
rect 8987 3417 8999 3451
rect 9582 3448 9588 3460
rect 8941 3411 8999 3417
rect 9232 3420 9588 3448
rect 7466 3380 7472 3392
rect 5552 3352 7472 3380
rect 7466 3340 7472 3352
rect 7524 3340 7530 3392
rect 7834 3340 7840 3392
rect 7892 3380 7898 3392
rect 9232 3380 9260 3420
rect 9582 3408 9588 3420
rect 9640 3408 9646 3460
rect 9784 3448 9812 3488
rect 10137 3485 10149 3519
rect 10183 3485 10195 3519
rect 10137 3479 10195 3485
rect 10321 3519 10379 3525
rect 10321 3485 10333 3519
rect 10367 3485 10379 3519
rect 10321 3479 10379 3485
rect 10152 3448 10180 3479
rect 10778 3476 10784 3528
rect 10836 3516 10842 3528
rect 11241 3519 11299 3525
rect 11241 3516 11253 3519
rect 10836 3488 11253 3516
rect 10836 3476 10842 3488
rect 11241 3485 11253 3488
rect 11287 3485 11299 3519
rect 11609 3519 11667 3525
rect 11609 3516 11621 3519
rect 11241 3479 11299 3485
rect 11440 3488 11621 3516
rect 10410 3448 10416 3460
rect 9784 3420 10416 3448
rect 10410 3408 10416 3420
rect 10468 3408 10474 3460
rect 10689 3451 10747 3457
rect 10689 3417 10701 3451
rect 10735 3448 10747 3451
rect 11440 3448 11468 3488
rect 11609 3485 11621 3488
rect 11655 3485 11667 3519
rect 11609 3479 11667 3485
rect 11790 3476 11796 3528
rect 11848 3516 11854 3528
rect 12253 3519 12311 3525
rect 12253 3516 12265 3519
rect 11848 3488 12265 3516
rect 11848 3476 11854 3488
rect 12253 3485 12265 3488
rect 12299 3485 12311 3519
rect 12253 3479 12311 3485
rect 12342 3476 12348 3528
rect 12400 3516 12406 3528
rect 12544 3516 12572 3556
rect 13081 3553 13093 3556
rect 13127 3553 13139 3587
rect 13081 3547 13139 3553
rect 13170 3544 13176 3596
rect 13228 3584 13234 3596
rect 14936 3584 14964 3612
rect 13228 3556 13273 3584
rect 14292 3556 14964 3584
rect 13228 3544 13234 3556
rect 12400 3488 12572 3516
rect 12621 3519 12679 3525
rect 12400 3476 12406 3488
rect 12621 3485 12633 3519
rect 12667 3516 12679 3519
rect 13357 3519 13415 3525
rect 12667 3488 12848 3516
rect 12667 3485 12679 3488
rect 12621 3479 12679 3485
rect 12529 3451 12587 3457
rect 12529 3448 12541 3451
rect 10735 3420 11468 3448
rect 11532 3420 12541 3448
rect 10735 3417 10747 3420
rect 10689 3411 10747 3417
rect 7892 3352 9260 3380
rect 7892 3340 7898 3352
rect 9306 3340 9312 3392
rect 9364 3380 9370 3392
rect 11532 3380 11560 3420
rect 12529 3417 12541 3420
rect 12575 3417 12587 3451
rect 12710 3448 12716 3460
rect 12671 3420 12716 3448
rect 12529 3411 12587 3417
rect 12710 3408 12716 3420
rect 12768 3408 12774 3460
rect 12820 3448 12848 3488
rect 13357 3485 13369 3519
rect 13403 3516 13415 3519
rect 13538 3516 13544 3528
rect 13403 3488 13544 3516
rect 13403 3485 13415 3488
rect 13357 3479 13415 3485
rect 13538 3476 13544 3488
rect 13596 3516 13602 3528
rect 13906 3516 13912 3528
rect 13596 3488 13912 3516
rect 13596 3476 13602 3488
rect 13906 3476 13912 3488
rect 13964 3476 13970 3528
rect 13998 3476 14004 3528
rect 14056 3516 14062 3528
rect 14292 3525 14320 3556
rect 14277 3519 14335 3525
rect 14277 3516 14289 3519
rect 14056 3488 14289 3516
rect 14056 3476 14062 3488
rect 14277 3485 14289 3488
rect 14323 3485 14335 3519
rect 14277 3479 14335 3485
rect 13262 3448 13268 3460
rect 12820 3420 13268 3448
rect 13262 3408 13268 3420
rect 13320 3408 13326 3460
rect 9364 3352 11560 3380
rect 11609 3383 11667 3389
rect 9364 3340 9370 3352
rect 11609 3349 11621 3383
rect 11655 3380 11667 3383
rect 12802 3380 12808 3392
rect 11655 3352 12808 3380
rect 11655 3349 11667 3352
rect 11609 3343 11667 3349
rect 12802 3340 12808 3352
rect 12860 3340 12866 3392
rect 1104 3290 15824 3312
rect 1104 3238 3447 3290
rect 3499 3238 3511 3290
rect 3563 3238 3575 3290
rect 3627 3238 3639 3290
rect 3691 3238 8378 3290
rect 8430 3238 8442 3290
rect 8494 3238 8506 3290
rect 8558 3238 8570 3290
rect 8622 3238 13308 3290
rect 13360 3238 13372 3290
rect 13424 3238 13436 3290
rect 13488 3238 13500 3290
rect 13552 3238 15824 3290
rect 1104 3216 15824 3238
rect 1578 3136 1584 3188
rect 1636 3176 1642 3188
rect 1673 3179 1731 3185
rect 1673 3176 1685 3179
rect 1636 3148 1685 3176
rect 1636 3136 1642 3148
rect 1673 3145 1685 3148
rect 1719 3145 1731 3179
rect 1673 3139 1731 3145
rect 2130 3136 2136 3188
rect 2188 3176 2194 3188
rect 2685 3179 2743 3185
rect 2685 3176 2697 3179
rect 2188 3148 2697 3176
rect 2188 3136 2194 3148
rect 2685 3145 2697 3148
rect 2731 3145 2743 3179
rect 2685 3139 2743 3145
rect 3234 3136 3240 3188
rect 3292 3176 3298 3188
rect 3697 3179 3755 3185
rect 3697 3176 3709 3179
rect 3292 3148 3709 3176
rect 3292 3136 3298 3148
rect 3697 3145 3709 3148
rect 3743 3145 3755 3179
rect 3697 3139 3755 3145
rect 3878 3136 3884 3188
rect 3936 3176 3942 3188
rect 4709 3179 4767 3185
rect 4709 3176 4721 3179
rect 3936 3148 4721 3176
rect 3936 3136 3942 3148
rect 4709 3145 4721 3148
rect 4755 3145 4767 3179
rect 4709 3139 4767 3145
rect 5074 3136 5080 3188
rect 5132 3176 5138 3188
rect 5442 3176 5448 3188
rect 5132 3148 5448 3176
rect 5132 3136 5138 3148
rect 5442 3136 5448 3148
rect 5500 3136 5506 3188
rect 5534 3136 5540 3188
rect 5592 3176 5598 3188
rect 5721 3179 5779 3185
rect 5721 3176 5733 3179
rect 5592 3148 5733 3176
rect 5592 3136 5598 3148
rect 5721 3145 5733 3148
rect 5767 3145 5779 3179
rect 5721 3139 5779 3145
rect 5810 3136 5816 3188
rect 5868 3176 5874 3188
rect 6825 3179 6883 3185
rect 6825 3176 6837 3179
rect 5868 3148 6837 3176
rect 5868 3136 5874 3148
rect 6825 3145 6837 3148
rect 6871 3145 6883 3179
rect 6825 3139 6883 3145
rect 7006 3136 7012 3188
rect 7064 3176 7070 3188
rect 7834 3176 7840 3188
rect 7064 3148 7840 3176
rect 7064 3136 7070 3148
rect 7834 3136 7840 3148
rect 7892 3136 7898 3188
rect 10686 3176 10692 3188
rect 8128 3148 10692 3176
rect 1854 3068 1860 3120
rect 1912 3108 1918 3120
rect 2406 3108 2412 3120
rect 1912 3080 2412 3108
rect 1912 3068 1918 3080
rect 2406 3068 2412 3080
rect 2464 3068 2470 3120
rect 3344 3080 4384 3108
rect 2222 3040 2228 3052
rect 2183 3012 2228 3040
rect 2222 3000 2228 3012
rect 2280 3000 2286 3052
rect 3344 3049 3372 3080
rect 3329 3043 3387 3049
rect 3329 3009 3341 3043
rect 3375 3009 3387 3043
rect 4246 3040 4252 3052
rect 4207 3012 4252 3040
rect 3329 3003 3387 3009
rect 4246 3000 4252 3012
rect 4304 3000 4310 3052
rect 4356 3040 4384 3080
rect 4982 3068 4988 3120
rect 5040 3108 5046 3120
rect 5040 3080 6224 3108
rect 5040 3068 5046 3080
rect 4522 3040 4528 3052
rect 4356 3012 4528 3040
rect 4522 3000 4528 3012
rect 4580 3000 4586 3052
rect 5166 3040 5172 3052
rect 5127 3012 5172 3040
rect 5166 3000 5172 3012
rect 5224 3000 5230 3052
rect 5353 3043 5411 3049
rect 5353 3009 5365 3043
rect 5399 3040 5411 3043
rect 5442 3040 5448 3052
rect 5399 3012 5448 3040
rect 5399 3009 5411 3012
rect 5353 3003 5411 3009
rect 5442 3000 5448 3012
rect 5500 3000 5506 3052
rect 6196 3049 6224 3080
rect 6181 3043 6239 3049
rect 6181 3009 6193 3043
rect 6227 3009 6239 3043
rect 6181 3003 6239 3009
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3040 6423 3043
rect 6454 3040 6460 3052
rect 6411 3012 6460 3040
rect 6411 3009 6423 3012
rect 6365 3003 6423 3009
rect 6454 3000 6460 3012
rect 6512 3000 6518 3052
rect 7469 3043 7527 3049
rect 7469 3009 7481 3043
rect 7515 3040 7527 3043
rect 7558 3040 7564 3052
rect 7515 3012 7564 3040
rect 7515 3009 7527 3012
rect 7469 3003 7527 3009
rect 7558 3000 7564 3012
rect 7616 3000 7622 3052
rect 2133 2975 2191 2981
rect 2133 2941 2145 2975
rect 2179 2972 2191 2975
rect 3145 2975 3203 2981
rect 3145 2972 3157 2975
rect 2179 2944 3157 2972
rect 2179 2941 2191 2944
rect 2133 2935 2191 2941
rect 3145 2941 3157 2944
rect 3191 2972 3203 2975
rect 6270 2972 6276 2984
rect 3191 2944 6276 2972
rect 3191 2941 3203 2944
rect 3145 2935 3203 2941
rect 6270 2932 6276 2944
rect 6328 2932 6334 2984
rect 7193 2975 7251 2981
rect 7193 2941 7205 2975
rect 7239 2972 7251 2975
rect 8128 2972 8156 3148
rect 10686 3136 10692 3148
rect 10744 3136 10750 3188
rect 10873 3179 10931 3185
rect 10873 3145 10885 3179
rect 10919 3176 10931 3179
rect 10919 3148 12112 3176
rect 10919 3145 10931 3148
rect 10873 3139 10931 3145
rect 8757 3111 8815 3117
rect 8757 3108 8769 3111
rect 8404 3080 8769 3108
rect 8404 3040 8432 3080
rect 8757 3077 8769 3080
rect 8803 3077 8815 3111
rect 9861 3111 9919 3117
rect 8757 3071 8815 3077
rect 9508 3080 9689 3108
rect 7239 2944 8156 2972
rect 8220 3012 8432 3040
rect 8481 3043 8539 3049
rect 7239 2941 7251 2944
rect 7193 2935 7251 2941
rect 2958 2864 2964 2916
rect 3016 2904 3022 2916
rect 4157 2907 4215 2913
rect 4157 2904 4169 2907
rect 3016 2876 4169 2904
rect 3016 2864 3022 2876
rect 4157 2873 4169 2876
rect 4203 2873 4215 2907
rect 4157 2867 4215 2873
rect 5077 2907 5135 2913
rect 5077 2873 5089 2907
rect 5123 2904 5135 2907
rect 5626 2904 5632 2916
rect 5123 2876 5632 2904
rect 5123 2873 5135 2876
rect 5077 2867 5135 2873
rect 5626 2864 5632 2876
rect 5684 2864 5690 2916
rect 6089 2907 6147 2913
rect 6089 2873 6101 2907
rect 6135 2904 6147 2907
rect 7098 2904 7104 2916
rect 6135 2876 7104 2904
rect 6135 2873 6147 2876
rect 6089 2867 6147 2873
rect 7098 2864 7104 2876
rect 7156 2864 7162 2916
rect 7285 2907 7343 2913
rect 7285 2873 7297 2907
rect 7331 2904 7343 2907
rect 8220 2904 8248 3012
rect 8481 3009 8493 3043
rect 8527 3040 8539 3043
rect 8527 3012 9260 3040
rect 8527 3009 8539 3012
rect 8481 3003 8539 3009
rect 8297 2975 8355 2981
rect 8297 2941 8309 2975
rect 8343 2972 8355 2975
rect 8386 2972 8392 2984
rect 8343 2944 8392 2972
rect 8343 2941 8355 2944
rect 8297 2935 8355 2941
rect 8386 2932 8392 2944
rect 8444 2972 8450 2984
rect 8662 2972 8668 2984
rect 8444 2944 8668 2972
rect 8444 2932 8450 2944
rect 8662 2932 8668 2944
rect 8720 2932 8726 2984
rect 8757 2975 8815 2981
rect 8757 2941 8769 2975
rect 8803 2972 8815 2975
rect 8846 2972 8852 2984
rect 8803 2944 8852 2972
rect 8803 2941 8815 2944
rect 8757 2935 8815 2941
rect 8846 2932 8852 2944
rect 8904 2932 8910 2984
rect 9232 2972 9260 3012
rect 9306 3000 9312 3052
rect 9364 3040 9370 3052
rect 9508 3049 9536 3080
rect 9661 3052 9689 3080
rect 9861 3077 9873 3111
rect 9907 3077 9919 3111
rect 9861 3071 9919 3077
rect 9493 3043 9551 3049
rect 9364 3012 9409 3040
rect 9364 3000 9370 3012
rect 9493 3009 9505 3043
rect 9539 3009 9551 3043
rect 9661 3012 9680 3052
rect 9493 3003 9551 3009
rect 9674 3000 9680 3012
rect 9732 3000 9738 3052
rect 9876 3040 9904 3071
rect 10410 3068 10416 3120
rect 10468 3108 10474 3120
rect 12084 3108 12112 3148
rect 12250 3136 12256 3188
rect 12308 3176 12314 3188
rect 12437 3179 12495 3185
rect 12437 3176 12449 3179
rect 12308 3148 12449 3176
rect 12308 3136 12314 3148
rect 12437 3145 12449 3148
rect 12483 3145 12495 3179
rect 13630 3176 13636 3188
rect 13591 3148 13636 3176
rect 12437 3139 12495 3145
rect 13630 3136 13636 3148
rect 13688 3136 13694 3188
rect 12526 3108 12532 3120
rect 10468 3080 12020 3108
rect 12084 3080 12532 3108
rect 10468 3068 10474 3080
rect 9950 3040 9956 3052
rect 9876 3012 9956 3040
rect 9950 3000 9956 3012
rect 10008 3000 10014 3052
rect 10318 3040 10324 3052
rect 10279 3012 10324 3040
rect 10318 3000 10324 3012
rect 10376 3000 10382 3052
rect 10505 3043 10563 3049
rect 10505 3009 10517 3043
rect 10551 3040 10563 3043
rect 10686 3040 10692 3052
rect 10551 3012 10692 3040
rect 10551 3009 10563 3012
rect 10505 3003 10563 3009
rect 10686 3000 10692 3012
rect 10744 3000 10750 3052
rect 11238 3000 11244 3052
rect 11296 3040 11302 3052
rect 11425 3043 11483 3049
rect 11425 3040 11437 3043
rect 11296 3012 11437 3040
rect 11296 3000 11302 3012
rect 11425 3009 11437 3012
rect 11471 3040 11483 3043
rect 11790 3040 11796 3052
rect 11471 3012 11796 3040
rect 11471 3009 11483 3012
rect 11425 3003 11483 3009
rect 11790 3000 11796 3012
rect 11848 3000 11854 3052
rect 10042 2972 10048 2984
rect 9232 2944 10048 2972
rect 10042 2932 10048 2944
rect 10100 2932 10106 2984
rect 10229 2975 10287 2981
rect 10229 2941 10241 2975
rect 10275 2972 10287 2975
rect 11992 2972 12020 3080
rect 12526 3068 12532 3080
rect 12584 3068 12590 3120
rect 12802 3068 12808 3120
rect 12860 3108 12866 3120
rect 12860 3080 12940 3108
rect 12860 3068 12866 3080
rect 12158 3000 12164 3052
rect 12216 3040 12222 3052
rect 12618 3040 12624 3052
rect 12216 3012 12624 3040
rect 12216 3000 12222 3012
rect 12618 3000 12624 3012
rect 12676 3000 12682 3052
rect 12912 3049 12940 3080
rect 13262 3068 13268 3120
rect 13320 3108 13326 3120
rect 14185 3111 14243 3117
rect 14185 3108 14197 3111
rect 13320 3080 14197 3108
rect 13320 3068 13326 3080
rect 14185 3077 14197 3080
rect 14231 3077 14243 3111
rect 14185 3071 14243 3077
rect 12897 3043 12955 3049
rect 12897 3009 12909 3043
rect 12943 3009 12955 3043
rect 12897 3003 12955 3009
rect 13081 3043 13139 3049
rect 13081 3009 13093 3043
rect 13127 3040 13139 3043
rect 13127 3012 13676 3040
rect 13127 3009 13139 3012
rect 13081 3003 13139 3009
rect 12526 2972 12532 2984
rect 10275 2944 11836 2972
rect 11992 2944 12532 2972
rect 10275 2941 10287 2944
rect 10229 2935 10287 2941
rect 7331 2876 8248 2904
rect 7331 2873 7343 2876
rect 7285 2867 7343 2873
rect 9950 2864 9956 2916
rect 10008 2904 10014 2916
rect 10594 2904 10600 2916
rect 10008 2876 10600 2904
rect 10008 2864 10014 2876
rect 10594 2864 10600 2876
rect 10652 2864 10658 2916
rect 10778 2864 10784 2916
rect 10836 2864 10842 2916
rect 11333 2907 11391 2913
rect 11333 2873 11345 2907
rect 11379 2904 11391 2907
rect 11698 2904 11704 2916
rect 11379 2876 11704 2904
rect 11379 2873 11391 2876
rect 11333 2867 11391 2873
rect 11698 2864 11704 2876
rect 11756 2864 11762 2916
rect 11808 2904 11836 2944
rect 12526 2932 12532 2944
rect 12584 2972 12590 2984
rect 12805 2975 12863 2981
rect 12805 2972 12817 2975
rect 12584 2944 12817 2972
rect 12584 2932 12590 2944
rect 12805 2941 12817 2944
rect 12851 2941 12863 2975
rect 13096 2972 13124 3003
rect 13262 2972 13268 2984
rect 13096 2944 13268 2972
rect 12805 2935 12863 2941
rect 13262 2932 13268 2944
rect 13320 2932 13326 2984
rect 13446 2972 13452 2984
rect 13407 2944 13452 2972
rect 13446 2932 13452 2944
rect 13504 2932 13510 2984
rect 13648 2972 13676 3012
rect 13722 3000 13728 3052
rect 13780 3040 13786 3052
rect 13780 3012 14596 3040
rect 13780 3000 13786 3012
rect 13906 2972 13912 2984
rect 13648 2944 13912 2972
rect 13906 2932 13912 2944
rect 13964 2932 13970 2984
rect 14001 2975 14059 2981
rect 14001 2941 14013 2975
rect 14047 2972 14059 2975
rect 14366 2972 14372 2984
rect 14047 2944 14372 2972
rect 14047 2941 14059 2944
rect 14001 2935 14059 2941
rect 14366 2932 14372 2944
rect 14424 2932 14430 2984
rect 14568 2981 14596 3012
rect 14553 2975 14611 2981
rect 14553 2941 14565 2975
rect 14599 2941 14611 2975
rect 14553 2935 14611 2941
rect 11808 2876 12572 2904
rect 1394 2796 1400 2848
rect 1452 2836 1458 2848
rect 2041 2839 2099 2845
rect 2041 2836 2053 2839
rect 1452 2808 2053 2836
rect 1452 2796 1458 2808
rect 2041 2805 2053 2808
rect 2087 2836 2099 2839
rect 3053 2839 3111 2845
rect 3053 2836 3065 2839
rect 2087 2808 3065 2836
rect 2087 2805 2099 2808
rect 2041 2799 2099 2805
rect 3053 2805 3065 2808
rect 3099 2836 3111 2839
rect 3878 2836 3884 2848
rect 3099 2808 3884 2836
rect 3099 2805 3111 2808
rect 3053 2799 3111 2805
rect 3878 2796 3884 2808
rect 3936 2796 3942 2848
rect 4062 2836 4068 2848
rect 4023 2808 4068 2836
rect 4062 2796 4068 2808
rect 4120 2796 4126 2848
rect 5718 2796 5724 2848
rect 5776 2836 5782 2848
rect 6914 2836 6920 2848
rect 5776 2808 6920 2836
rect 5776 2796 5782 2808
rect 6914 2796 6920 2808
rect 6972 2796 6978 2848
rect 7742 2796 7748 2848
rect 7800 2836 7806 2848
rect 7837 2839 7895 2845
rect 7837 2836 7849 2839
rect 7800 2808 7849 2836
rect 7800 2796 7806 2808
rect 7837 2805 7849 2808
rect 7883 2805 7895 2839
rect 8202 2836 8208 2848
rect 8163 2808 8208 2836
rect 7837 2799 7895 2805
rect 8202 2796 8208 2808
rect 8260 2796 8266 2848
rect 8294 2796 8300 2848
rect 8352 2836 8358 2848
rect 8849 2839 8907 2845
rect 8849 2836 8861 2839
rect 8352 2808 8861 2836
rect 8352 2796 8358 2808
rect 8849 2805 8861 2808
rect 8895 2805 8907 2839
rect 8849 2799 8907 2805
rect 9217 2839 9275 2845
rect 9217 2805 9229 2839
rect 9263 2836 9275 2839
rect 9306 2836 9312 2848
rect 9263 2808 9312 2836
rect 9263 2805 9275 2808
rect 9217 2799 9275 2805
rect 9306 2796 9312 2808
rect 9364 2796 9370 2848
rect 9398 2796 9404 2848
rect 9456 2836 9462 2848
rect 10796 2836 10824 2864
rect 9456 2808 10824 2836
rect 11241 2839 11299 2845
rect 9456 2796 9462 2808
rect 11241 2805 11253 2839
rect 11287 2836 11299 2839
rect 11514 2836 11520 2848
rect 11287 2808 11520 2836
rect 11287 2805 11299 2808
rect 11241 2799 11299 2805
rect 11514 2796 11520 2808
rect 11572 2796 11578 2848
rect 11885 2839 11943 2845
rect 11885 2805 11897 2839
rect 11931 2836 11943 2839
rect 12342 2836 12348 2848
rect 11931 2808 12348 2836
rect 11931 2805 11943 2808
rect 11885 2799 11943 2805
rect 12342 2796 12348 2808
rect 12400 2796 12406 2848
rect 12544 2836 12572 2876
rect 12618 2864 12624 2916
rect 12676 2904 12682 2916
rect 13464 2904 13492 2932
rect 12676 2876 13492 2904
rect 12676 2864 12682 2876
rect 12894 2836 12900 2848
rect 12544 2808 12900 2836
rect 12894 2796 12900 2808
rect 12952 2796 12958 2848
rect 14734 2836 14740 2848
rect 14695 2808 14740 2836
rect 14734 2796 14740 2808
rect 14792 2796 14798 2848
rect 1104 2746 15824 2768
rect 1104 2694 5912 2746
rect 5964 2694 5976 2746
rect 6028 2694 6040 2746
rect 6092 2694 6104 2746
rect 6156 2694 10843 2746
rect 10895 2694 10907 2746
rect 10959 2694 10971 2746
rect 11023 2694 11035 2746
rect 11087 2694 15824 2746
rect 1104 2672 15824 2694
rect 2958 2632 2964 2644
rect 2919 2604 2964 2632
rect 2958 2592 2964 2604
rect 3016 2592 3022 2644
rect 3421 2635 3479 2641
rect 3421 2601 3433 2635
rect 3467 2632 3479 2635
rect 4062 2632 4068 2644
rect 3467 2604 4068 2632
rect 3467 2601 3479 2604
rect 3421 2595 3479 2601
rect 4062 2592 4068 2604
rect 4120 2592 4126 2644
rect 4801 2635 4859 2641
rect 4801 2601 4813 2635
rect 4847 2601 4859 2635
rect 5166 2632 5172 2644
rect 5127 2604 5172 2632
rect 4801 2595 4859 2601
rect 2869 2567 2927 2573
rect 2869 2564 2881 2567
rect 2240 2536 2881 2564
rect 1489 2499 1547 2505
rect 1489 2465 1501 2499
rect 1535 2496 1547 2499
rect 1946 2496 1952 2508
rect 1535 2468 1952 2496
rect 1535 2465 1547 2468
rect 1489 2459 1547 2465
rect 1946 2456 1952 2468
rect 2004 2456 2010 2508
rect 2240 2505 2268 2536
rect 2869 2533 2881 2536
rect 2915 2533 2927 2567
rect 2869 2527 2927 2533
rect 3329 2567 3387 2573
rect 3329 2533 3341 2567
rect 3375 2564 3387 2567
rect 4816 2564 4844 2595
rect 5166 2592 5172 2604
rect 5224 2592 5230 2644
rect 5261 2635 5319 2641
rect 5261 2601 5273 2635
rect 5307 2632 5319 2635
rect 5442 2632 5448 2644
rect 5307 2604 5448 2632
rect 5307 2601 5319 2604
rect 5261 2595 5319 2601
rect 5442 2592 5448 2604
rect 5500 2632 5506 2644
rect 5629 2635 5687 2641
rect 5629 2632 5641 2635
rect 5500 2604 5641 2632
rect 5500 2592 5506 2604
rect 5629 2601 5641 2604
rect 5675 2601 5687 2635
rect 5629 2595 5687 2601
rect 5813 2635 5871 2641
rect 5813 2601 5825 2635
rect 5859 2601 5871 2635
rect 6270 2632 6276 2644
rect 6183 2604 6276 2632
rect 5813 2595 5871 2601
rect 3375 2536 4844 2564
rect 3375 2533 3387 2536
rect 3329 2527 3387 2533
rect 4890 2524 4896 2576
rect 4948 2564 4954 2576
rect 5828 2564 5856 2595
rect 6270 2592 6276 2604
rect 6328 2632 6334 2644
rect 8386 2632 8392 2644
rect 6328 2604 8392 2632
rect 6328 2592 6334 2604
rect 8386 2592 8392 2604
rect 8444 2592 8450 2644
rect 8481 2635 8539 2641
rect 8481 2601 8493 2635
rect 8527 2632 8539 2635
rect 10502 2632 10508 2644
rect 8527 2604 10508 2632
rect 8527 2601 8539 2604
rect 8481 2595 8539 2601
rect 10502 2592 10508 2604
rect 10560 2592 10566 2644
rect 11149 2635 11207 2641
rect 11149 2601 11161 2635
rect 11195 2632 11207 2635
rect 12710 2632 12716 2644
rect 11195 2604 12716 2632
rect 11195 2601 11207 2604
rect 11149 2595 11207 2601
rect 12710 2592 12716 2604
rect 12768 2592 12774 2644
rect 12805 2635 12863 2641
rect 12805 2601 12817 2635
rect 12851 2632 12863 2635
rect 12894 2632 12900 2644
rect 12851 2604 12900 2632
rect 12851 2601 12863 2604
rect 12805 2595 12863 2601
rect 12894 2592 12900 2604
rect 12952 2592 12958 2644
rect 13170 2592 13176 2644
rect 13228 2632 13234 2644
rect 13633 2635 13691 2641
rect 13633 2632 13645 2635
rect 13228 2604 13645 2632
rect 13228 2592 13234 2604
rect 13633 2601 13645 2604
rect 13679 2601 13691 2635
rect 13633 2595 13691 2601
rect 4948 2536 5856 2564
rect 4948 2524 4954 2536
rect 5902 2524 5908 2576
rect 5960 2564 5966 2576
rect 7561 2567 7619 2573
rect 7561 2564 7573 2567
rect 5960 2536 7573 2564
rect 5960 2524 5966 2536
rect 7561 2533 7573 2536
rect 7607 2533 7619 2567
rect 7561 2527 7619 2533
rect 8573 2567 8631 2573
rect 8573 2533 8585 2567
rect 8619 2564 8631 2567
rect 9493 2567 9551 2573
rect 9493 2564 9505 2567
rect 8619 2536 9505 2564
rect 8619 2533 8631 2536
rect 8573 2527 8631 2533
rect 9493 2533 9505 2536
rect 9539 2533 9551 2567
rect 9493 2527 9551 2533
rect 9585 2567 9643 2573
rect 9585 2533 9597 2567
rect 9631 2564 9643 2567
rect 10686 2564 10692 2576
rect 9631 2536 10692 2564
rect 9631 2533 9643 2536
rect 9585 2527 9643 2533
rect 10686 2524 10692 2536
rect 10744 2524 10750 2576
rect 11241 2567 11299 2573
rect 11241 2533 11253 2567
rect 11287 2564 11299 2567
rect 12986 2564 12992 2576
rect 11287 2536 12992 2564
rect 11287 2533 11299 2536
rect 11241 2527 11299 2533
rect 12986 2524 12992 2536
rect 13044 2524 13050 2576
rect 14918 2564 14924 2576
rect 13096 2536 14924 2564
rect 2225 2499 2283 2505
rect 2225 2465 2237 2499
rect 2271 2465 2283 2499
rect 2225 2459 2283 2465
rect 3970 2456 3976 2508
rect 4028 2496 4034 2508
rect 4065 2499 4123 2505
rect 4065 2496 4077 2499
rect 4028 2468 4077 2496
rect 4028 2456 4034 2468
rect 4065 2465 4077 2468
rect 4111 2465 4123 2499
rect 6178 2496 6184 2508
rect 6139 2468 6184 2496
rect 4065 2459 4123 2465
rect 6178 2456 6184 2468
rect 6236 2456 6242 2508
rect 7469 2499 7527 2505
rect 7469 2496 7481 2499
rect 6288 2468 7481 2496
rect 1670 2428 1676 2440
rect 1631 2400 1676 2428
rect 1670 2388 1676 2400
rect 1728 2388 1734 2440
rect 2406 2428 2412 2440
rect 2367 2400 2412 2428
rect 2406 2388 2412 2400
rect 2464 2388 2470 2440
rect 3510 2428 3516 2440
rect 3471 2400 3516 2428
rect 3510 2388 3516 2400
rect 3568 2388 3574 2440
rect 3602 2388 3608 2440
rect 3660 2428 3666 2440
rect 4249 2431 4307 2437
rect 4249 2428 4261 2431
rect 3660 2400 4261 2428
rect 3660 2388 3666 2400
rect 4249 2397 4261 2400
rect 4295 2397 4307 2431
rect 5442 2428 5448 2440
rect 5403 2400 5448 2428
rect 4249 2391 4307 2397
rect 5442 2388 5448 2400
rect 5500 2388 5506 2440
rect 5629 2431 5687 2437
rect 5629 2397 5641 2431
rect 5675 2428 5687 2431
rect 6288 2428 6316 2468
rect 7469 2465 7481 2468
rect 7515 2496 7527 2499
rect 7834 2496 7840 2508
rect 7515 2468 7840 2496
rect 7515 2465 7527 2468
rect 7469 2459 7527 2465
rect 7834 2456 7840 2468
rect 7892 2456 7898 2508
rect 8018 2456 8024 2508
rect 8076 2496 8082 2508
rect 8076 2468 9076 2496
rect 8076 2456 8082 2468
rect 5675 2400 6316 2428
rect 6457 2431 6515 2437
rect 5675 2397 5687 2400
rect 5629 2391 5687 2397
rect 6457 2397 6469 2431
rect 6503 2428 6515 2431
rect 6638 2428 6644 2440
rect 6503 2400 6644 2428
rect 6503 2397 6515 2400
rect 6457 2391 6515 2397
rect 6638 2388 6644 2400
rect 6696 2388 6702 2440
rect 7745 2431 7803 2437
rect 7745 2397 7757 2431
rect 7791 2428 7803 2431
rect 7926 2428 7932 2440
rect 7791 2400 7932 2428
rect 7791 2397 7803 2400
rect 7745 2391 7803 2397
rect 7926 2388 7932 2400
rect 7984 2388 7990 2440
rect 8757 2431 8815 2437
rect 8757 2397 8769 2431
rect 8803 2428 8815 2431
rect 8938 2428 8944 2440
rect 8803 2400 8944 2428
rect 8803 2397 8815 2400
rect 8757 2391 8815 2397
rect 8938 2388 8944 2400
rect 8996 2388 9002 2440
rect 9048 2428 9076 2468
rect 9122 2456 9128 2508
rect 9180 2496 9186 2508
rect 10134 2496 10140 2508
rect 9180 2468 9225 2496
rect 9462 2468 9812 2496
rect 10095 2468 10140 2496
rect 9180 2456 9186 2468
rect 9462 2428 9490 2468
rect 9048 2400 9490 2428
rect 1026 2320 1032 2372
rect 1084 2360 1090 2372
rect 9309 2363 9367 2369
rect 9309 2360 9321 2363
rect 1084 2332 9321 2360
rect 1084 2320 1090 2332
rect 9309 2329 9321 2332
rect 9355 2329 9367 2363
rect 9784 2360 9812 2468
rect 10134 2456 10140 2468
rect 10192 2456 10198 2508
rect 10229 2499 10287 2505
rect 10229 2465 10241 2499
rect 10275 2496 10287 2499
rect 11790 2496 11796 2508
rect 10275 2468 11652 2496
rect 11751 2468 11796 2496
rect 10275 2465 10287 2468
rect 10229 2459 10287 2465
rect 10410 2428 10416 2440
rect 10371 2400 10416 2428
rect 10410 2388 10416 2400
rect 10468 2428 10474 2440
rect 11146 2428 11152 2440
rect 10468 2400 11152 2428
rect 10468 2388 10474 2400
rect 11146 2388 11152 2400
rect 11204 2388 11210 2440
rect 11333 2431 11391 2437
rect 11333 2428 11345 2431
rect 11256 2400 11345 2428
rect 11256 2360 11284 2400
rect 11333 2397 11345 2400
rect 11379 2397 11391 2431
rect 11624 2428 11652 2468
rect 11790 2456 11796 2468
rect 11848 2456 11854 2508
rect 12621 2499 12679 2505
rect 12621 2465 12633 2499
rect 12667 2496 12679 2499
rect 13096 2496 13124 2536
rect 14918 2524 14924 2536
rect 14976 2524 14982 2576
rect 12667 2468 13124 2496
rect 12667 2465 12679 2468
rect 12621 2459 12679 2465
rect 13170 2456 13176 2508
rect 13228 2496 13234 2508
rect 13633 2499 13691 2505
rect 13228 2468 13273 2496
rect 13228 2456 13234 2468
rect 13633 2465 13645 2499
rect 13679 2496 13691 2499
rect 13725 2499 13783 2505
rect 13725 2496 13737 2499
rect 13679 2468 13737 2496
rect 13679 2465 13691 2468
rect 13633 2459 13691 2465
rect 13725 2465 13737 2468
rect 13771 2465 13783 2499
rect 13725 2459 13783 2465
rect 14277 2499 14335 2505
rect 14277 2465 14289 2499
rect 14323 2465 14335 2499
rect 14277 2459 14335 2465
rect 14829 2499 14887 2505
rect 14829 2465 14841 2499
rect 14875 2496 14887 2499
rect 15286 2496 15292 2508
rect 14875 2468 15292 2496
rect 14875 2465 14887 2468
rect 14829 2459 14887 2465
rect 13078 2428 13084 2440
rect 11624 2400 13084 2428
rect 11333 2391 11391 2397
rect 13078 2388 13084 2400
rect 13136 2388 13142 2440
rect 9784 2332 11284 2360
rect 9309 2323 9367 2329
rect 11422 2320 11428 2372
rect 11480 2360 11486 2372
rect 13357 2363 13415 2369
rect 13357 2360 13369 2363
rect 11480 2332 13369 2360
rect 11480 2320 11486 2332
rect 13357 2329 13369 2332
rect 13403 2329 13415 2363
rect 13357 2323 13415 2329
rect 13446 2320 13452 2372
rect 13504 2360 13510 2372
rect 14292 2360 14320 2459
rect 15286 2456 15292 2468
rect 15344 2456 15350 2508
rect 13504 2332 14320 2360
rect 13504 2320 13510 2332
rect 2869 2295 2927 2301
rect 2869 2261 2881 2295
rect 2915 2292 2927 2295
rect 5350 2292 5356 2304
rect 2915 2264 5356 2292
rect 2915 2261 2927 2264
rect 2869 2255 2927 2261
rect 5350 2252 5356 2264
rect 5408 2252 5414 2304
rect 7098 2292 7104 2304
rect 7059 2264 7104 2292
rect 7098 2252 7104 2264
rect 7156 2252 7162 2304
rect 8110 2292 8116 2304
rect 8071 2264 8116 2292
rect 8110 2252 8116 2264
rect 8168 2252 8174 2304
rect 9766 2292 9772 2304
rect 9727 2264 9772 2292
rect 9766 2252 9772 2264
rect 9824 2252 9830 2304
rect 10594 2252 10600 2304
rect 10652 2292 10658 2304
rect 10781 2295 10839 2301
rect 10781 2292 10793 2295
rect 10652 2264 10793 2292
rect 10652 2252 10658 2264
rect 10781 2261 10793 2264
rect 10827 2261 10839 2295
rect 11974 2292 11980 2304
rect 11935 2264 11980 2292
rect 10781 2255 10839 2261
rect 11974 2252 11980 2264
rect 12032 2252 12038 2304
rect 13906 2292 13912 2304
rect 13867 2264 13912 2292
rect 13906 2252 13912 2264
rect 13964 2252 13970 2304
rect 14458 2292 14464 2304
rect 14419 2264 14464 2292
rect 14458 2252 14464 2264
rect 14516 2252 14522 2304
rect 14550 2252 14556 2304
rect 14608 2292 14614 2304
rect 15013 2295 15071 2301
rect 15013 2292 15025 2295
rect 14608 2264 15025 2292
rect 14608 2252 14614 2264
rect 15013 2261 15025 2264
rect 15059 2261 15071 2295
rect 15013 2255 15071 2261
rect 1104 2202 15824 2224
rect 1104 2150 3447 2202
rect 3499 2150 3511 2202
rect 3563 2150 3575 2202
rect 3627 2150 3639 2202
rect 3691 2150 8378 2202
rect 8430 2150 8442 2202
rect 8494 2150 8506 2202
rect 8558 2150 8570 2202
rect 8622 2150 13308 2202
rect 13360 2150 13372 2202
rect 13424 2150 13436 2202
rect 13488 2150 13500 2202
rect 13552 2150 15824 2202
rect 1104 2128 15824 2150
rect 4062 2048 4068 2100
rect 4120 2088 4126 2100
rect 7282 2088 7288 2100
rect 4120 2060 7288 2088
rect 4120 2048 4126 2060
rect 7282 2048 7288 2060
rect 7340 2048 7346 2100
rect 7374 2048 7380 2100
rect 7432 2088 7438 2100
rect 14458 2088 14464 2100
rect 7432 2060 14464 2088
rect 7432 2048 7438 2060
rect 14458 2048 14464 2060
rect 14516 2048 14522 2100
rect 1762 1980 1768 2032
rect 1820 2020 1826 2032
rect 8202 2020 8208 2032
rect 1820 1992 8208 2020
rect 1820 1980 1826 1992
rect 8202 1980 8208 1992
rect 8260 1980 8266 2032
rect 11698 1980 11704 2032
rect 11756 2020 11762 2032
rect 12618 2020 12624 2032
rect 11756 1992 12624 2020
rect 11756 1980 11762 1992
rect 12618 1980 12624 1992
rect 12676 1980 12682 2032
rect 6546 1912 6552 1964
rect 6604 1952 6610 1964
rect 13906 1952 13912 1964
rect 6604 1924 13912 1952
rect 6604 1912 6610 1924
rect 13906 1912 13912 1924
rect 13964 1912 13970 1964
rect 4430 1844 4436 1896
rect 4488 1884 4494 1896
rect 12894 1884 12900 1896
rect 4488 1856 12900 1884
rect 4488 1844 4494 1856
rect 12894 1844 12900 1856
rect 12952 1844 12958 1896
rect 5442 1776 5448 1828
rect 5500 1816 5506 1828
rect 9398 1816 9404 1828
rect 5500 1788 9404 1816
rect 5500 1776 5506 1788
rect 9398 1776 9404 1788
rect 9456 1776 9462 1828
rect 10134 1776 10140 1828
rect 10192 1816 10198 1828
rect 12434 1816 12440 1828
rect 10192 1788 12440 1816
rect 10192 1776 10198 1788
rect 12434 1776 12440 1788
rect 12492 1816 12498 1828
rect 13354 1816 13360 1828
rect 12492 1788 13360 1816
rect 12492 1776 12498 1788
rect 13354 1776 13360 1788
rect 13412 1776 13418 1828
rect 566 1708 572 1760
rect 624 1748 630 1760
rect 11974 1748 11980 1760
rect 624 1720 11980 1748
rect 624 1708 630 1720
rect 11974 1708 11980 1720
rect 12032 1708 12038 1760
rect 3326 1640 3332 1692
rect 3384 1680 3390 1692
rect 8113 1683 8171 1689
rect 8113 1680 8125 1683
rect 3384 1652 8125 1680
rect 3384 1640 3390 1652
rect 8113 1649 8125 1652
rect 8159 1649 8171 1683
rect 8113 1643 8171 1649
rect 8202 1640 8208 1692
rect 8260 1680 8266 1692
rect 14090 1680 14096 1692
rect 8260 1652 14096 1680
rect 8260 1640 8266 1652
rect 14090 1640 14096 1652
rect 14148 1640 14154 1692
rect 6086 1572 6092 1624
rect 6144 1612 6150 1624
rect 11422 1612 11428 1624
rect 6144 1584 11428 1612
rect 6144 1572 6150 1584
rect 11422 1572 11428 1584
rect 11480 1572 11486 1624
rect 5534 1504 5540 1556
rect 5592 1544 5598 1556
rect 9766 1544 9772 1556
rect 5592 1516 9772 1544
rect 5592 1504 5598 1516
rect 9766 1504 9772 1516
rect 9824 1504 9830 1556
rect 2866 1436 2872 1488
rect 2924 1476 2930 1488
rect 10594 1476 10600 1488
rect 2924 1448 10600 1476
rect 2924 1436 2930 1448
rect 10594 1436 10600 1448
rect 10652 1436 10658 1488
rect 3970 1368 3976 1420
rect 4028 1408 4034 1420
rect 7650 1408 7656 1420
rect 4028 1380 7656 1408
rect 4028 1368 4034 1380
rect 7650 1368 7656 1380
rect 7708 1368 7714 1420
rect 7834 1368 7840 1420
rect 7892 1408 7898 1420
rect 14550 1408 14556 1420
rect 7892 1380 14556 1408
rect 7892 1368 7898 1380
rect 14550 1368 14556 1380
rect 14608 1368 14614 1420
rect 7742 1300 7748 1352
rect 7800 1340 7806 1352
rect 13170 1340 13176 1352
rect 7800 1312 13176 1340
rect 7800 1300 7806 1312
rect 13170 1300 13176 1312
rect 13228 1300 13234 1352
rect 7466 1232 7472 1284
rect 7524 1272 7530 1284
rect 14274 1272 14280 1284
rect 7524 1244 14280 1272
rect 7524 1232 7530 1244
rect 9508 1216 9536 1244
rect 14274 1232 14280 1244
rect 14332 1232 14338 1284
rect 9490 1164 9496 1216
rect 9548 1164 9554 1216
rect 10410 1164 10416 1216
rect 10468 1204 10474 1216
rect 15102 1204 15108 1216
rect 10468 1176 15108 1204
rect 10468 1164 10474 1176
rect 15102 1164 15108 1176
rect 15160 1164 15166 1216
rect 9306 1096 9312 1148
rect 9364 1136 9370 1148
rect 12158 1136 12164 1148
rect 9364 1108 12164 1136
rect 9364 1096 9370 1108
rect 12158 1096 12164 1108
rect 12216 1096 12222 1148
rect 8113 935 8171 941
rect 8113 901 8125 935
rect 8159 932 8171 935
rect 12894 932 12900 944
rect 8159 904 12900 932
rect 8159 901 8171 904
rect 8113 895 8171 901
rect 12894 892 12900 904
rect 12952 932 12958 944
rect 13722 932 13728 944
rect 12952 904 13728 932
rect 12952 892 12958 904
rect 13722 892 13728 904
rect 13780 892 13786 944
rect 1854 552 1860 604
rect 1912 592 1918 604
rect 11330 592 11336 604
rect 1912 564 11336 592
rect 1912 552 1918 564
rect 11330 552 11336 564
rect 11388 552 11394 604
<< via1 >>
rect 7472 16124 7524 16176
rect 9128 16124 9180 16176
rect 8116 16056 8168 16108
rect 8668 16056 8720 16108
rect 7012 15988 7064 16040
rect 9404 15988 9456 16040
rect 1032 15920 1084 15972
rect 3332 15920 3384 15972
rect 4252 15920 4304 15972
rect 11796 15920 11848 15972
rect 3148 15852 3200 15904
rect 4068 15852 4120 15904
rect 6644 15852 6696 15904
rect 9864 15852 9916 15904
rect 5912 15750 5964 15802
rect 5976 15750 6028 15802
rect 6040 15750 6092 15802
rect 6104 15750 6156 15802
rect 10843 15750 10895 15802
rect 10907 15750 10959 15802
rect 10971 15750 11023 15802
rect 11035 15750 11087 15802
rect 3608 15648 3660 15700
rect 5264 15648 5316 15700
rect 2044 15580 2096 15632
rect 8208 15648 8260 15700
rect 9404 15648 9456 15700
rect 3792 15512 3844 15564
rect 4252 15555 4304 15564
rect 4252 15521 4261 15555
rect 4261 15521 4295 15555
rect 4295 15521 4304 15555
rect 4252 15512 4304 15521
rect 5816 15512 5868 15564
rect 6184 15555 6236 15564
rect 6184 15521 6193 15555
rect 6193 15521 6227 15555
rect 6227 15521 6236 15555
rect 6184 15512 6236 15521
rect 2780 15444 2832 15496
rect 5632 15444 5684 15496
rect 7472 15555 7524 15564
rect 7472 15521 7481 15555
rect 7481 15521 7515 15555
rect 7515 15521 7524 15555
rect 7472 15512 7524 15521
rect 6644 15444 6696 15496
rect 2688 15376 2740 15428
rect 5448 15376 5500 15428
rect 9036 15512 9088 15564
rect 10048 15512 10100 15564
rect 11152 15512 11204 15564
rect 8668 15487 8720 15496
rect 8668 15453 8677 15487
rect 8677 15453 8711 15487
rect 8711 15453 8720 15487
rect 8668 15444 8720 15453
rect 8760 15444 8812 15496
rect 9956 15444 10008 15496
rect 9312 15376 9364 15428
rect 10416 15376 10468 15428
rect 13912 15376 13964 15428
rect 3056 15308 3108 15360
rect 6644 15308 6696 15360
rect 7104 15351 7156 15360
rect 7104 15317 7113 15351
rect 7113 15317 7147 15351
rect 7147 15317 7156 15351
rect 7104 15308 7156 15317
rect 7196 15308 7248 15360
rect 10324 15308 10376 15360
rect 13820 15308 13872 15360
rect 3447 15206 3499 15258
rect 3511 15206 3563 15258
rect 3575 15206 3627 15258
rect 3639 15206 3691 15258
rect 8378 15206 8430 15258
rect 8442 15206 8494 15258
rect 8506 15206 8558 15258
rect 8570 15206 8622 15258
rect 13308 15206 13360 15258
rect 13372 15206 13424 15258
rect 13436 15206 13488 15258
rect 13500 15206 13552 15258
rect 1400 15104 1452 15156
rect 3056 15104 3108 15156
rect 3148 15104 3200 15156
rect 6552 15104 6604 15156
rect 572 15036 624 15088
rect 3332 15036 3384 15088
rect 1860 14968 1912 15020
rect 5540 15036 5592 15088
rect 2228 14943 2280 14952
rect 2228 14909 2237 14943
rect 2237 14909 2271 14943
rect 2271 14909 2280 14943
rect 2228 14900 2280 14909
rect 2780 14943 2832 14952
rect 2780 14909 2789 14943
rect 2789 14909 2823 14943
rect 2823 14909 2832 14943
rect 2780 14900 2832 14909
rect 3240 14900 3292 14952
rect 3700 14900 3752 14952
rect 3976 14900 4028 14952
rect 6092 14968 6144 15020
rect 6276 15036 6328 15088
rect 6368 15011 6420 15020
rect 6368 14977 6377 15011
rect 6377 14977 6411 15011
rect 6411 14977 6420 15011
rect 6368 14968 6420 14977
rect 6920 15036 6972 15088
rect 12164 15104 12216 15156
rect 4988 14900 5040 14952
rect 5724 14900 5776 14952
rect 6276 14900 6328 14952
rect 6460 14900 6512 14952
rect 4068 14832 4120 14884
rect 7288 14968 7340 15020
rect 8668 14968 8720 15020
rect 7380 14900 7432 14952
rect 7656 14900 7708 14952
rect 7932 14900 7984 14952
rect 8024 14900 8076 14952
rect 14188 15036 14240 15088
rect 14740 15036 14792 15088
rect 10508 14968 10560 15020
rect 4804 14764 4856 14816
rect 5172 14764 5224 14816
rect 5816 14764 5868 14816
rect 6736 14764 6788 14816
rect 8944 14832 8996 14884
rect 10232 14832 10284 14884
rect 10600 14900 10652 14952
rect 10784 14900 10836 14952
rect 12992 14900 13044 14952
rect 7656 14807 7708 14816
rect 7656 14773 7665 14807
rect 7665 14773 7699 14807
rect 7699 14773 7708 14807
rect 7656 14764 7708 14773
rect 8208 14764 8260 14816
rect 8668 14807 8720 14816
rect 8668 14773 8677 14807
rect 8677 14773 8711 14807
rect 8711 14773 8720 14807
rect 8668 14764 8720 14773
rect 9036 14807 9088 14816
rect 9036 14773 9045 14807
rect 9045 14773 9079 14807
rect 9079 14773 9088 14807
rect 9036 14764 9088 14773
rect 11244 14807 11296 14816
rect 11244 14773 11253 14807
rect 11253 14773 11287 14807
rect 11287 14773 11296 14807
rect 11244 14764 11296 14773
rect 11336 14764 11388 14816
rect 11888 14764 11940 14816
rect 5912 14662 5964 14714
rect 5976 14662 6028 14714
rect 6040 14662 6092 14714
rect 6104 14662 6156 14714
rect 10843 14662 10895 14714
rect 10907 14662 10959 14714
rect 10971 14662 11023 14714
rect 11035 14662 11087 14714
rect 204 14560 256 14612
rect 3792 14560 3844 14612
rect 5724 14603 5776 14612
rect 5724 14569 5733 14603
rect 5733 14569 5767 14603
rect 5767 14569 5776 14603
rect 5724 14560 5776 14569
rect 7104 14560 7156 14612
rect 7564 14560 7616 14612
rect 8484 14560 8536 14612
rect 8852 14603 8904 14612
rect 8852 14569 8861 14603
rect 8861 14569 8895 14603
rect 8895 14569 8904 14603
rect 8852 14560 8904 14569
rect 8944 14560 8996 14612
rect 9588 14560 9640 14612
rect 12808 14560 12860 14612
rect 1860 14467 1912 14476
rect 1860 14433 1869 14467
rect 1869 14433 1903 14467
rect 1903 14433 1912 14467
rect 1860 14424 1912 14433
rect 4436 14492 4488 14544
rect 2964 14467 3016 14476
rect 2964 14433 2973 14467
rect 2973 14433 3007 14467
rect 3007 14433 3016 14467
rect 2964 14424 3016 14433
rect 3332 14424 3384 14476
rect 6552 14492 6604 14544
rect 8576 14492 8628 14544
rect 10600 14492 10652 14544
rect 14556 14492 14608 14544
rect 4712 14467 4764 14476
rect 4712 14433 4721 14467
rect 4721 14433 4755 14467
rect 4755 14433 4764 14467
rect 4712 14424 4764 14433
rect 3148 14399 3200 14408
rect 3148 14365 3157 14399
rect 3157 14365 3191 14399
rect 3191 14365 3200 14399
rect 3148 14356 3200 14365
rect 4620 14356 4672 14408
rect 5540 14356 5592 14408
rect 7012 14424 7064 14476
rect 7748 14467 7800 14476
rect 7748 14433 7757 14467
rect 7757 14433 7791 14467
rect 7791 14433 7800 14467
rect 7748 14424 7800 14433
rect 9496 14424 9548 14476
rect 5080 14288 5132 14340
rect 6828 14288 6880 14340
rect 2780 14220 2832 14272
rect 3884 14220 3936 14272
rect 4344 14263 4396 14272
rect 4344 14229 4353 14263
rect 4353 14229 4387 14263
rect 4387 14229 4396 14263
rect 4344 14220 4396 14229
rect 5356 14263 5408 14272
rect 5356 14229 5365 14263
rect 5365 14229 5399 14263
rect 5399 14229 5408 14263
rect 5356 14220 5408 14229
rect 5540 14220 5592 14272
rect 5816 14220 5868 14272
rect 7104 14288 7156 14340
rect 7472 14220 7524 14272
rect 8576 14288 8628 14340
rect 8760 14288 8812 14340
rect 9404 14356 9456 14408
rect 9772 14424 9824 14476
rect 9864 14424 9916 14476
rect 10232 14424 10284 14476
rect 9680 14356 9732 14408
rect 10508 14356 10560 14408
rect 10692 14424 10744 14476
rect 11704 14467 11756 14476
rect 11704 14433 11713 14467
rect 11713 14433 11747 14467
rect 11747 14433 11756 14467
rect 11704 14424 11756 14433
rect 13820 14424 13872 14476
rect 14464 14356 14516 14408
rect 15476 14356 15528 14408
rect 9772 14288 9824 14340
rect 10416 14288 10468 14340
rect 9404 14220 9456 14272
rect 9588 14220 9640 14272
rect 12256 14263 12308 14272
rect 12256 14229 12265 14263
rect 12265 14229 12299 14263
rect 12299 14229 12308 14263
rect 12256 14220 12308 14229
rect 14188 14220 14240 14272
rect 3447 14118 3499 14170
rect 3511 14118 3563 14170
rect 3575 14118 3627 14170
rect 3639 14118 3691 14170
rect 8378 14118 8430 14170
rect 8442 14118 8494 14170
rect 8506 14118 8558 14170
rect 8570 14118 8622 14170
rect 13308 14118 13360 14170
rect 13372 14118 13424 14170
rect 13436 14118 13488 14170
rect 13500 14118 13552 14170
rect 2964 14016 3016 14068
rect 6828 14059 6880 14068
rect 6828 14025 6837 14059
rect 6837 14025 6871 14059
rect 6871 14025 6880 14059
rect 6828 14016 6880 14025
rect 7012 14016 7064 14068
rect 8208 14016 8260 14068
rect 2780 13948 2832 14000
rect 2228 13880 2280 13932
rect 2136 13855 2188 13864
rect 2136 13821 2145 13855
rect 2145 13821 2179 13855
rect 2179 13821 2188 13855
rect 2136 13812 2188 13821
rect 2780 13812 2832 13864
rect 4068 13948 4120 14000
rect 5356 13948 5408 14000
rect 3056 13923 3108 13932
rect 3056 13889 3065 13923
rect 3065 13889 3099 13923
rect 3099 13889 3108 13923
rect 3056 13880 3108 13889
rect 3792 13880 3844 13932
rect 4528 13880 4580 13932
rect 5080 13880 5132 13932
rect 5264 13923 5316 13932
rect 5264 13889 5273 13923
rect 5273 13889 5307 13923
rect 5307 13889 5316 13923
rect 5264 13880 5316 13889
rect 6276 13923 6328 13932
rect 6276 13889 6285 13923
rect 6285 13889 6319 13923
rect 6319 13889 6328 13923
rect 6276 13880 6328 13889
rect 8668 13948 8720 14000
rect 9588 13948 9640 14000
rect 9772 13948 9824 14000
rect 3240 13744 3292 13796
rect 5356 13812 5408 13864
rect 5724 13744 5776 13796
rect 7656 13812 7708 13864
rect 8116 13812 8168 13864
rect 8944 13880 8996 13932
rect 9404 13880 9456 13932
rect 10416 13923 10468 13932
rect 9128 13812 9180 13864
rect 10416 13889 10425 13923
rect 10425 13889 10459 13923
rect 10459 13889 10468 13923
rect 10416 13880 10468 13889
rect 9588 13812 9640 13864
rect 9864 13812 9916 13864
rect 12348 14016 12400 14068
rect 12440 13948 12492 14000
rect 15936 13948 15988 14000
rect 12348 13880 12400 13932
rect 11336 13855 11388 13864
rect 11336 13821 11345 13855
rect 11345 13821 11379 13855
rect 11379 13821 11388 13855
rect 11336 13812 11388 13821
rect 12716 13812 12768 13864
rect 7196 13787 7248 13796
rect 7196 13753 7205 13787
rect 7205 13753 7239 13787
rect 7239 13753 7248 13787
rect 7196 13744 7248 13753
rect 8576 13744 8628 13796
rect 10784 13744 10836 13796
rect 2688 13676 2740 13728
rect 3884 13676 3936 13728
rect 4712 13719 4764 13728
rect 4712 13685 4721 13719
rect 4721 13685 4755 13719
rect 4755 13685 4764 13719
rect 4712 13676 4764 13685
rect 4804 13676 4856 13728
rect 5540 13676 5592 13728
rect 7288 13676 7340 13728
rect 7932 13676 7984 13728
rect 8944 13676 8996 13728
rect 9312 13719 9364 13728
rect 9312 13685 9321 13719
rect 9321 13685 9355 13719
rect 9355 13685 9364 13719
rect 9312 13676 9364 13685
rect 11612 13676 11664 13728
rect 12440 13676 12492 13728
rect 5912 13574 5964 13626
rect 5976 13574 6028 13626
rect 6040 13574 6092 13626
rect 6104 13574 6156 13626
rect 10843 13574 10895 13626
rect 10907 13574 10959 13626
rect 10971 13574 11023 13626
rect 11035 13574 11087 13626
rect 4344 13472 4396 13524
rect 4896 13472 4948 13524
rect 5356 13472 5408 13524
rect 7472 13472 7524 13524
rect 9956 13472 10008 13524
rect 4712 13404 4764 13456
rect 1676 13311 1728 13320
rect 1676 13277 1685 13311
rect 1685 13277 1719 13311
rect 1719 13277 1728 13311
rect 1676 13268 1728 13277
rect 2872 13336 2924 13388
rect 3056 13336 3108 13388
rect 5540 13336 5592 13388
rect 6920 13404 6972 13456
rect 7932 13404 7984 13456
rect 8208 13404 8260 13456
rect 8576 13404 8628 13456
rect 10048 13447 10100 13456
rect 2964 13268 3016 13320
rect 3976 13268 4028 13320
rect 4712 13311 4764 13320
rect 4712 13277 4721 13311
rect 4721 13277 4755 13311
rect 4755 13277 4764 13311
rect 4712 13268 4764 13277
rect 5080 13268 5132 13320
rect 7656 13336 7708 13388
rect 7840 13336 7892 13388
rect 8668 13336 8720 13388
rect 9128 13336 9180 13388
rect 10048 13413 10057 13447
rect 10057 13413 10091 13447
rect 10091 13413 10100 13447
rect 10048 13404 10100 13413
rect 10876 13404 10928 13456
rect 11336 13472 11388 13524
rect 11704 13515 11756 13524
rect 11704 13481 11713 13515
rect 11713 13481 11747 13515
rect 11747 13481 11756 13515
rect 11704 13472 11756 13481
rect 12164 13515 12216 13524
rect 12164 13481 12173 13515
rect 12173 13481 12207 13515
rect 12207 13481 12216 13515
rect 12164 13472 12216 13481
rect 12900 13404 12952 13456
rect 14004 13447 14056 13456
rect 14004 13413 14013 13447
rect 14013 13413 14047 13447
rect 14047 13413 14056 13447
rect 14004 13404 14056 13413
rect 9220 13268 9272 13320
rect 5540 13200 5592 13252
rect 8944 13200 8996 13252
rect 10048 13268 10100 13320
rect 9864 13200 9916 13252
rect 10416 13268 10468 13320
rect 11336 13311 11388 13320
rect 11336 13277 11345 13311
rect 11345 13277 11379 13311
rect 11379 13277 11388 13311
rect 11336 13268 11388 13277
rect 10968 13200 11020 13252
rect 11060 13200 11112 13252
rect 11428 13200 11480 13252
rect 13084 13379 13136 13388
rect 12164 13268 12216 13320
rect 13084 13345 13093 13379
rect 13093 13345 13127 13379
rect 13127 13345 13136 13379
rect 13084 13336 13136 13345
rect 13176 13311 13228 13320
rect 12348 13200 12400 13252
rect 3148 13132 3200 13184
rect 4160 13132 4212 13184
rect 4436 13132 4488 13184
rect 5172 13132 5224 13184
rect 6552 13132 6604 13184
rect 8208 13132 8260 13184
rect 10784 13132 10836 13184
rect 11520 13132 11572 13184
rect 13176 13277 13185 13311
rect 13185 13277 13219 13311
rect 13219 13277 13228 13311
rect 13176 13268 13228 13277
rect 13452 13268 13504 13320
rect 13728 13132 13780 13184
rect 3447 13030 3499 13082
rect 3511 13030 3563 13082
rect 3575 13030 3627 13082
rect 3639 13030 3691 13082
rect 8378 13030 8430 13082
rect 8442 13030 8494 13082
rect 8506 13030 8558 13082
rect 8570 13030 8622 13082
rect 13308 13030 13360 13082
rect 13372 13030 13424 13082
rect 13436 13030 13488 13082
rect 13500 13030 13552 13082
rect 6000 12928 6052 12980
rect 6828 12928 6880 12980
rect 7012 12928 7064 12980
rect 9496 12971 9548 12980
rect 9496 12937 9505 12971
rect 9505 12937 9539 12971
rect 9539 12937 9548 12971
rect 9496 12928 9548 12937
rect 10048 12928 10100 12980
rect 11060 12928 11112 12980
rect 12164 12928 12216 12980
rect 8484 12903 8536 12912
rect 2872 12792 2924 12844
rect 3148 12835 3200 12844
rect 3148 12801 3157 12835
rect 3157 12801 3191 12835
rect 3191 12801 3200 12835
rect 3148 12792 3200 12801
rect 4160 12835 4212 12844
rect 2596 12724 2648 12776
rect 4160 12801 4169 12835
rect 4169 12801 4203 12835
rect 4203 12801 4212 12835
rect 4160 12792 4212 12801
rect 4896 12792 4948 12844
rect 6368 12835 6420 12844
rect 6368 12801 6377 12835
rect 6377 12801 6411 12835
rect 6411 12801 6420 12835
rect 6368 12792 6420 12801
rect 6552 12792 6604 12844
rect 8484 12869 8493 12903
rect 8493 12869 8527 12903
rect 8527 12869 8536 12903
rect 8484 12860 8536 12869
rect 10232 12860 10284 12912
rect 12072 12860 12124 12912
rect 12440 12903 12492 12912
rect 12440 12869 12449 12903
rect 12449 12869 12483 12903
rect 12483 12869 12492 12903
rect 12440 12860 12492 12869
rect 13084 12928 13136 12980
rect 3700 12724 3752 12776
rect 4436 12724 4488 12776
rect 5724 12724 5776 12776
rect 6184 12767 6236 12776
rect 6184 12733 6193 12767
rect 6193 12733 6227 12767
rect 6227 12733 6236 12767
rect 6184 12724 6236 12733
rect 8300 12792 8352 12844
rect 4252 12656 4304 12708
rect 1584 12588 1636 12640
rect 2044 12631 2096 12640
rect 2044 12597 2053 12631
rect 2053 12597 2087 12631
rect 2087 12597 2096 12631
rect 2044 12588 2096 12597
rect 3700 12631 3752 12640
rect 3700 12597 3709 12631
rect 3709 12597 3743 12631
rect 3743 12597 3752 12631
rect 3700 12588 3752 12597
rect 4160 12588 4212 12640
rect 5448 12588 5500 12640
rect 6000 12656 6052 12708
rect 6828 12588 6880 12640
rect 8760 12724 8812 12776
rect 9220 12792 9272 12844
rect 9496 12792 9548 12844
rect 10048 12835 10100 12844
rect 10048 12801 10057 12835
rect 10057 12801 10091 12835
rect 10091 12801 10100 12835
rect 10048 12792 10100 12801
rect 10692 12792 10744 12844
rect 11060 12792 11112 12844
rect 11704 12792 11756 12844
rect 12164 12792 12216 12844
rect 8944 12656 8996 12708
rect 9128 12656 9180 12708
rect 9588 12656 9640 12708
rect 11244 12724 11296 12776
rect 10968 12656 11020 12708
rect 11428 12656 11480 12708
rect 11980 12724 12032 12776
rect 12900 12767 12952 12776
rect 12900 12733 12909 12767
rect 12909 12733 12943 12767
rect 12943 12733 12952 12767
rect 12900 12724 12952 12733
rect 13820 12860 13872 12912
rect 14372 12860 14424 12912
rect 13268 12792 13320 12844
rect 14188 12724 14240 12776
rect 15384 12656 15436 12708
rect 9496 12588 9548 12640
rect 10324 12588 10376 12640
rect 11244 12588 11296 12640
rect 12164 12588 12216 12640
rect 12808 12631 12860 12640
rect 12808 12597 12817 12631
rect 12817 12597 12851 12631
rect 12851 12597 12860 12631
rect 12808 12588 12860 12597
rect 13452 12588 13504 12640
rect 13728 12588 13780 12640
rect 14924 12588 14976 12640
rect 5912 12486 5964 12538
rect 5976 12486 6028 12538
rect 6040 12486 6092 12538
rect 6104 12486 6156 12538
rect 10843 12486 10895 12538
rect 10907 12486 10959 12538
rect 10971 12486 11023 12538
rect 11035 12486 11087 12538
rect 2044 12384 2096 12436
rect 3240 12384 3292 12436
rect 3700 12384 3752 12436
rect 4068 12427 4120 12436
rect 4068 12393 4077 12427
rect 4077 12393 4111 12427
rect 4111 12393 4120 12427
rect 4068 12384 4120 12393
rect 4528 12427 4580 12436
rect 4528 12393 4537 12427
rect 4537 12393 4571 12427
rect 4571 12393 4580 12427
rect 4528 12384 4580 12393
rect 8484 12384 8536 12436
rect 2504 12316 2556 12368
rect 3148 12316 3200 12368
rect 3976 12316 4028 12368
rect 4436 12359 4488 12368
rect 4436 12325 4445 12359
rect 4445 12325 4479 12359
rect 4479 12325 4488 12359
rect 4436 12316 4488 12325
rect 2320 12291 2372 12300
rect 2320 12257 2329 12291
rect 2329 12257 2363 12291
rect 2363 12257 2372 12291
rect 2320 12248 2372 12257
rect 6368 12316 6420 12368
rect 6552 12316 6604 12368
rect 9404 12384 9456 12436
rect 11428 12384 11480 12436
rect 11980 12384 12032 12436
rect 12072 12427 12124 12436
rect 12072 12393 12081 12427
rect 12081 12393 12115 12427
rect 12115 12393 12124 12427
rect 13176 12427 13228 12436
rect 12072 12384 12124 12393
rect 13176 12393 13185 12427
rect 13185 12393 13219 12427
rect 13219 12393 13228 12427
rect 13176 12384 13228 12393
rect 13452 12384 13504 12436
rect 14188 12427 14240 12436
rect 14188 12393 14197 12427
rect 14197 12393 14231 12427
rect 14231 12393 14240 12427
rect 14188 12384 14240 12393
rect 16764 12384 16816 12436
rect 5080 12291 5132 12300
rect 5080 12257 5089 12291
rect 5089 12257 5123 12291
rect 5123 12257 5132 12291
rect 5080 12248 5132 12257
rect 6828 12248 6880 12300
rect 8760 12291 8812 12300
rect 8760 12257 8769 12291
rect 8769 12257 8803 12291
rect 8803 12257 8812 12291
rect 8760 12248 8812 12257
rect 2412 12223 2464 12232
rect 2412 12189 2421 12223
rect 2421 12189 2455 12223
rect 2455 12189 2464 12223
rect 2412 12180 2464 12189
rect 2596 12223 2648 12232
rect 2596 12189 2605 12223
rect 2605 12189 2639 12223
rect 2639 12189 2648 12223
rect 2596 12180 2648 12189
rect 4436 12180 4488 12232
rect 4712 12223 4764 12232
rect 4712 12189 4721 12223
rect 4721 12189 4755 12223
rect 4755 12189 4764 12223
rect 4712 12180 4764 12189
rect 4804 12180 4856 12232
rect 8208 12180 8260 12232
rect 8668 12180 8720 12232
rect 9036 12223 9088 12232
rect 9036 12189 9045 12223
rect 9045 12189 9079 12223
rect 9079 12189 9088 12223
rect 9036 12180 9088 12189
rect 1492 12044 1544 12096
rect 6368 12044 6420 12096
rect 9956 12248 10008 12300
rect 10600 12248 10652 12300
rect 10692 12248 10744 12300
rect 11244 12248 11296 12300
rect 10508 12180 10560 12232
rect 10876 12180 10928 12232
rect 10968 12180 11020 12232
rect 11336 12223 11388 12232
rect 11336 12189 11345 12223
rect 11345 12189 11379 12223
rect 11379 12189 11388 12223
rect 11336 12180 11388 12189
rect 13176 12248 13228 12300
rect 13912 12248 13964 12300
rect 12348 12223 12400 12232
rect 12348 12189 12357 12223
rect 12357 12189 12391 12223
rect 12391 12189 12400 12223
rect 12348 12180 12400 12189
rect 12900 12180 12952 12232
rect 13728 12180 13780 12232
rect 13084 12112 13136 12164
rect 8116 12087 8168 12096
rect 8116 12053 8125 12087
rect 8125 12053 8159 12087
rect 8159 12053 8168 12087
rect 8116 12044 8168 12053
rect 8208 12044 8260 12096
rect 8852 12044 8904 12096
rect 10968 12044 11020 12096
rect 11060 12044 11112 12096
rect 12532 12044 12584 12096
rect 12716 12087 12768 12096
rect 12716 12053 12725 12087
rect 12725 12053 12759 12087
rect 12759 12053 12768 12087
rect 12716 12044 12768 12053
rect 12900 12044 12952 12096
rect 14740 12044 14792 12096
rect 3447 11942 3499 11994
rect 3511 11942 3563 11994
rect 3575 11942 3627 11994
rect 3639 11942 3691 11994
rect 8378 11942 8430 11994
rect 8442 11942 8494 11994
rect 8506 11942 8558 11994
rect 8570 11942 8622 11994
rect 13308 11942 13360 11994
rect 13372 11942 13424 11994
rect 13436 11942 13488 11994
rect 13500 11942 13552 11994
rect 4528 11840 4580 11892
rect 4436 11772 4488 11824
rect 8208 11840 8260 11892
rect 9496 11840 9548 11892
rect 10508 11840 10560 11892
rect 3884 11636 3936 11688
rect 4068 11636 4120 11688
rect 4804 11704 4856 11756
rect 4896 11636 4948 11688
rect 5080 11679 5132 11688
rect 5080 11645 5089 11679
rect 5089 11645 5123 11679
rect 5123 11645 5132 11679
rect 5080 11636 5132 11645
rect 2412 11611 2464 11620
rect 2412 11577 2421 11611
rect 2421 11577 2455 11611
rect 2455 11577 2464 11611
rect 2412 11568 2464 11577
rect 3424 11611 3476 11620
rect 3424 11577 3433 11611
rect 3433 11577 3467 11611
rect 3467 11577 3476 11611
rect 3424 11568 3476 11577
rect 5356 11611 5408 11620
rect 5356 11577 5390 11611
rect 5390 11577 5408 11611
rect 5632 11636 5684 11688
rect 13820 11840 13872 11892
rect 11980 11772 12032 11824
rect 12440 11772 12492 11824
rect 13360 11772 13412 11824
rect 13544 11772 13596 11824
rect 6828 11747 6880 11756
rect 6828 11713 6837 11747
rect 6837 11713 6871 11747
rect 6871 11713 6880 11747
rect 6828 11704 6880 11713
rect 5356 11568 5408 11577
rect 1676 11500 1728 11552
rect 2504 11543 2556 11552
rect 2504 11509 2513 11543
rect 2513 11509 2547 11543
rect 2547 11509 2556 11543
rect 2504 11500 2556 11509
rect 3056 11543 3108 11552
rect 3056 11509 3065 11543
rect 3065 11509 3099 11543
rect 3099 11509 3108 11543
rect 3056 11500 3108 11509
rect 3516 11543 3568 11552
rect 3516 11509 3525 11543
rect 3525 11509 3559 11543
rect 3559 11509 3568 11543
rect 3516 11500 3568 11509
rect 4068 11543 4120 11552
rect 4068 11509 4077 11543
rect 4077 11509 4111 11543
rect 4111 11509 4120 11543
rect 4068 11500 4120 11509
rect 4712 11500 4764 11552
rect 7380 11568 7432 11620
rect 6644 11500 6696 11552
rect 7564 11500 7616 11552
rect 11336 11704 11388 11756
rect 12256 11704 12308 11756
rect 13728 11704 13780 11756
rect 10232 11636 10284 11688
rect 9496 11568 9548 11620
rect 9772 11568 9824 11620
rect 12348 11636 12400 11688
rect 12624 11636 12676 11688
rect 10416 11611 10468 11620
rect 10416 11577 10450 11611
rect 10450 11577 10468 11611
rect 10416 11568 10468 11577
rect 11060 11568 11112 11620
rect 15292 11704 15344 11756
rect 14832 11636 14884 11688
rect 15016 11568 15068 11620
rect 15292 11568 15344 11620
rect 16304 11772 16356 11824
rect 10692 11500 10744 11552
rect 11796 11543 11848 11552
rect 11796 11509 11805 11543
rect 11805 11509 11839 11543
rect 11839 11509 11848 11543
rect 11796 11500 11848 11509
rect 12624 11500 12676 11552
rect 12900 11543 12952 11552
rect 12900 11509 12909 11543
rect 12909 11509 12943 11543
rect 12943 11509 12952 11543
rect 12900 11500 12952 11509
rect 13452 11543 13504 11552
rect 13452 11509 13461 11543
rect 13461 11509 13495 11543
rect 13495 11509 13504 11543
rect 13452 11500 13504 11509
rect 13820 11500 13872 11552
rect 14096 11500 14148 11552
rect 5912 11398 5964 11450
rect 5976 11398 6028 11450
rect 6040 11398 6092 11450
rect 6104 11398 6156 11450
rect 10843 11398 10895 11450
rect 10907 11398 10959 11450
rect 10971 11398 11023 11450
rect 11035 11398 11087 11450
rect 2044 11296 2096 11348
rect 3056 11296 3108 11348
rect 4068 11296 4120 11348
rect 5356 11296 5408 11348
rect 4252 11228 4304 11280
rect 6368 11296 6420 11348
rect 7380 11339 7432 11348
rect 7380 11305 7389 11339
rect 7389 11305 7423 11339
rect 7423 11305 7432 11339
rect 7380 11296 7432 11305
rect 9128 11296 9180 11348
rect 2044 11024 2096 11076
rect 2504 11135 2556 11144
rect 2504 11101 2513 11135
rect 2513 11101 2547 11135
rect 2547 11101 2556 11135
rect 2504 11092 2556 11101
rect 4160 11160 4212 11212
rect 8116 11228 8168 11280
rect 8852 11228 8904 11280
rect 10416 11296 10468 11348
rect 10600 11296 10652 11348
rect 11520 11296 11572 11348
rect 11888 11296 11940 11348
rect 12624 11296 12676 11348
rect 13360 11339 13412 11348
rect 13360 11305 13369 11339
rect 13369 11305 13403 11339
rect 13403 11305 13412 11339
rect 13360 11296 13412 11305
rect 14740 11296 14792 11348
rect 11152 11228 11204 11280
rect 12440 11228 12492 11280
rect 12532 11228 12584 11280
rect 12992 11228 13044 11280
rect 3240 11092 3292 11144
rect 4436 11160 4488 11212
rect 6828 11160 6880 11212
rect 7380 11160 7432 11212
rect 8208 11160 8260 11212
rect 9956 11203 10008 11212
rect 9956 11169 9990 11203
rect 9990 11169 10008 11203
rect 9956 11160 10008 11169
rect 10232 11160 10284 11212
rect 11336 11160 11388 11212
rect 14188 11160 14240 11212
rect 7656 11135 7708 11144
rect 2964 11067 3016 11076
rect 2964 11033 2973 11067
rect 2973 11033 3007 11067
rect 3007 11033 3016 11067
rect 2964 11024 3016 11033
rect 3056 11024 3108 11076
rect 3516 11024 3568 11076
rect 4160 11024 4212 11076
rect 7656 11101 7665 11135
rect 7665 11101 7699 11135
rect 7699 11101 7708 11135
rect 7656 11092 7708 11101
rect 8852 11092 8904 11144
rect 9220 11092 9272 11144
rect 11888 11135 11940 11144
rect 7012 11024 7064 11076
rect 7564 10956 7616 11008
rect 8852 10956 8904 11008
rect 9496 10956 9548 11008
rect 11888 11101 11897 11135
rect 11897 11101 11931 11135
rect 11931 11101 11940 11135
rect 11888 11092 11940 11101
rect 12992 11135 13044 11144
rect 12992 11101 13001 11135
rect 13001 11101 13035 11135
rect 13035 11101 13044 11135
rect 12992 11092 13044 11101
rect 13360 11092 13412 11144
rect 14372 11092 14424 11144
rect 11060 10999 11112 11008
rect 11060 10965 11069 10999
rect 11069 10965 11103 10999
rect 11103 10965 11112 10999
rect 11060 10956 11112 10965
rect 11244 10956 11296 11008
rect 12164 10956 12216 11008
rect 12716 10956 12768 11008
rect 15476 10956 15528 11008
rect 3447 10854 3499 10906
rect 3511 10854 3563 10906
rect 3575 10854 3627 10906
rect 3639 10854 3691 10906
rect 8378 10854 8430 10906
rect 8442 10854 8494 10906
rect 8506 10854 8558 10906
rect 8570 10854 8622 10906
rect 13308 10854 13360 10906
rect 13372 10854 13424 10906
rect 13436 10854 13488 10906
rect 13500 10854 13552 10906
rect 4620 10752 4672 10804
rect 7472 10752 7524 10804
rect 8116 10752 8168 10804
rect 3332 10684 3384 10736
rect 4804 10727 4856 10736
rect 4804 10693 4813 10727
rect 4813 10693 4847 10727
rect 4847 10693 4856 10727
rect 4804 10684 4856 10693
rect 6552 10684 6604 10736
rect 7840 10684 7892 10736
rect 8484 10727 8536 10736
rect 8484 10693 8493 10727
rect 8493 10693 8527 10727
rect 8527 10693 8536 10727
rect 8484 10684 8536 10693
rect 1952 10548 2004 10600
rect 2780 10616 2832 10668
rect 6828 10659 6880 10668
rect 6828 10625 6837 10659
rect 6837 10625 6871 10659
rect 6871 10625 6880 10659
rect 6828 10616 6880 10625
rect 2320 10548 2372 10600
rect 4160 10548 4212 10600
rect 5080 10591 5132 10600
rect 5080 10557 5089 10591
rect 5089 10557 5123 10591
rect 5123 10557 5132 10591
rect 5080 10548 5132 10557
rect 5632 10548 5684 10600
rect 11060 10752 11112 10804
rect 11704 10752 11756 10804
rect 10692 10684 10744 10736
rect 11980 10684 12032 10736
rect 12900 10684 12952 10736
rect 9036 10659 9088 10668
rect 9036 10625 9045 10659
rect 9045 10625 9079 10659
rect 9079 10625 9088 10659
rect 9036 10616 9088 10625
rect 9496 10659 9548 10668
rect 9496 10625 9505 10659
rect 9505 10625 9539 10659
rect 9539 10625 9548 10659
rect 9496 10616 9548 10625
rect 10600 10616 10652 10668
rect 11888 10616 11940 10668
rect 13360 10616 13412 10668
rect 14464 10752 14516 10804
rect 14740 10752 14792 10804
rect 15016 10752 15068 10804
rect 15016 10659 15068 10668
rect 15016 10625 15025 10659
rect 15025 10625 15059 10659
rect 15059 10625 15068 10659
rect 15016 10616 15068 10625
rect 7104 10523 7156 10532
rect 7104 10489 7138 10523
rect 7138 10489 7156 10523
rect 7104 10480 7156 10489
rect 7840 10480 7892 10532
rect 8116 10480 8168 10532
rect 11244 10548 11296 10600
rect 11796 10548 11848 10600
rect 15108 10548 15160 10600
rect 9772 10523 9824 10532
rect 9772 10489 9806 10523
rect 9806 10489 9824 10523
rect 9772 10480 9824 10489
rect 2136 10412 2188 10464
rect 2412 10455 2464 10464
rect 2412 10421 2421 10455
rect 2421 10421 2455 10455
rect 2455 10421 2464 10455
rect 2412 10412 2464 10421
rect 3056 10412 3108 10464
rect 4620 10412 4672 10464
rect 6828 10412 6880 10464
rect 8944 10455 8996 10464
rect 8944 10421 8953 10455
rect 8953 10421 8987 10455
rect 8987 10421 8996 10455
rect 8944 10412 8996 10421
rect 10600 10412 10652 10464
rect 12992 10480 13044 10532
rect 13820 10523 13872 10532
rect 13820 10489 13829 10523
rect 13829 10489 13863 10523
rect 13863 10489 13872 10523
rect 13820 10480 13872 10489
rect 14372 10480 14424 10532
rect 14648 10480 14700 10532
rect 11704 10412 11756 10464
rect 12624 10412 12676 10464
rect 12808 10412 12860 10464
rect 13084 10412 13136 10464
rect 14464 10455 14516 10464
rect 14464 10421 14473 10455
rect 14473 10421 14507 10455
rect 14507 10421 14516 10455
rect 14464 10412 14516 10421
rect 15384 10412 15436 10464
rect 15936 10412 15988 10464
rect 5912 10310 5964 10362
rect 5976 10310 6028 10362
rect 6040 10310 6092 10362
rect 6104 10310 6156 10362
rect 10843 10310 10895 10362
rect 10907 10310 10959 10362
rect 10971 10310 11023 10362
rect 11035 10310 11087 10362
rect 5540 10251 5592 10260
rect 5540 10217 5549 10251
rect 5549 10217 5583 10251
rect 5583 10217 5592 10251
rect 5540 10208 5592 10217
rect 6644 10208 6696 10260
rect 1860 10183 1912 10192
rect 1860 10149 1869 10183
rect 1869 10149 1903 10183
rect 1903 10149 1912 10183
rect 1860 10140 1912 10149
rect 3240 10140 3292 10192
rect 6276 10140 6328 10192
rect 6828 10140 6880 10192
rect 9128 10140 9180 10192
rect 9772 10208 9824 10260
rect 9956 10208 10008 10260
rect 12992 10208 13044 10260
rect 13636 10208 13688 10260
rect 10416 10140 10468 10192
rect 1584 10115 1636 10124
rect 1584 10081 1593 10115
rect 1593 10081 1627 10115
rect 1627 10081 1636 10115
rect 1584 10072 1636 10081
rect 4160 10115 4212 10124
rect 4160 10081 4169 10115
rect 4169 10081 4203 10115
rect 4203 10081 4212 10115
rect 4160 10072 4212 10081
rect 1492 10004 1544 10056
rect 2320 10047 2372 10056
rect 2320 10013 2329 10047
rect 2329 10013 2363 10047
rect 2363 10013 2372 10047
rect 2320 10004 2372 10013
rect 3976 10004 4028 10056
rect 7656 10072 7708 10124
rect 9496 10072 9548 10124
rect 5172 10004 5224 10056
rect 9220 10004 9272 10056
rect 11244 10140 11296 10192
rect 12164 10140 12216 10192
rect 11060 10072 11112 10124
rect 11888 10072 11940 10124
rect 12348 10072 12400 10124
rect 14004 10072 14056 10124
rect 11336 10047 11388 10056
rect 11336 10013 11345 10047
rect 11345 10013 11379 10047
rect 11379 10013 11388 10047
rect 11336 10004 11388 10013
rect 10692 9936 10744 9988
rect 3792 9868 3844 9920
rect 6552 9868 6604 9920
rect 7748 9868 7800 9920
rect 7840 9868 7892 9920
rect 12716 9868 12768 9920
rect 14188 10004 14240 10056
rect 14464 9868 14516 9920
rect 3447 9766 3499 9818
rect 3511 9766 3563 9818
rect 3575 9766 3627 9818
rect 3639 9766 3691 9818
rect 8378 9766 8430 9818
rect 8442 9766 8494 9818
rect 8506 9766 8558 9818
rect 8570 9766 8622 9818
rect 13308 9766 13360 9818
rect 13372 9766 13424 9818
rect 13436 9766 13488 9818
rect 13500 9766 13552 9818
rect 4804 9664 4856 9716
rect 8116 9664 8168 9716
rect 7196 9596 7248 9648
rect 7380 9596 7432 9648
rect 8208 9596 8260 9648
rect 1492 9528 1544 9580
rect 5080 9571 5132 9580
rect 5080 9537 5089 9571
rect 5089 9537 5123 9571
rect 5123 9537 5132 9571
rect 5080 9528 5132 9537
rect 6460 9528 6512 9580
rect 2320 9460 2372 9512
rect 7104 9528 7156 9580
rect 9036 9664 9088 9716
rect 9496 9596 9548 9648
rect 10968 9664 11020 9716
rect 11428 9596 11480 9648
rect 15016 9664 15068 9716
rect 11704 9596 11756 9648
rect 14280 9596 14332 9648
rect 7932 9460 7984 9512
rect 8208 9503 8260 9512
rect 8208 9469 8217 9503
rect 8217 9469 8251 9503
rect 8251 9469 8260 9503
rect 8208 9460 8260 9469
rect 8300 9503 8352 9512
rect 8300 9469 8309 9503
rect 8309 9469 8343 9503
rect 8343 9469 8352 9503
rect 8300 9460 8352 9469
rect 3056 9392 3108 9444
rect 3792 9392 3844 9444
rect 5724 9392 5776 9444
rect 2596 9324 2648 9376
rect 8392 9392 8444 9444
rect 8852 9392 8904 9444
rect 6552 9324 6604 9376
rect 7472 9367 7524 9376
rect 7472 9333 7481 9367
rect 7481 9333 7515 9367
rect 7515 9333 7524 9367
rect 7472 9324 7524 9333
rect 9496 9392 9548 9444
rect 11336 9528 11388 9580
rect 13452 9528 13504 9580
rect 15108 9571 15160 9580
rect 15108 9537 15117 9571
rect 15117 9537 15151 9571
rect 15151 9537 15160 9571
rect 15108 9528 15160 9537
rect 11244 9460 11296 9512
rect 11980 9460 12032 9512
rect 12992 9460 13044 9512
rect 13176 9460 13228 9512
rect 10232 9435 10284 9444
rect 9312 9324 9364 9376
rect 10232 9401 10266 9435
rect 10266 9401 10284 9435
rect 10232 9392 10284 9401
rect 11244 9324 11296 9376
rect 12164 9392 12216 9444
rect 12440 9392 12492 9444
rect 12808 9392 12860 9444
rect 13268 9324 13320 9376
rect 13912 9324 13964 9376
rect 5912 9222 5964 9274
rect 5976 9222 6028 9274
rect 6040 9222 6092 9274
rect 6104 9222 6156 9274
rect 10843 9222 10895 9274
rect 10907 9222 10959 9274
rect 10971 9222 11023 9274
rect 11035 9222 11087 9274
rect 2872 9120 2924 9172
rect 3976 9120 4028 9172
rect 4068 9120 4120 9172
rect 4252 9120 4304 9172
rect 7288 9120 7340 9172
rect 7564 9120 7616 9172
rect 8208 9120 8260 9172
rect 1860 9095 1912 9104
rect 1860 9061 1869 9095
rect 1869 9061 1903 9095
rect 1903 9061 1912 9095
rect 1860 9052 1912 9061
rect 2596 9095 2648 9104
rect 2596 9061 2630 9095
rect 2630 9061 2648 9095
rect 2596 9052 2648 9061
rect 2688 9052 2740 9104
rect 6552 9052 6604 9104
rect 9956 9095 10008 9104
rect 9956 9061 9979 9095
rect 9979 9061 10008 9095
rect 9956 9052 10008 9061
rect 10140 9052 10192 9104
rect 11244 9120 11296 9172
rect 11336 9120 11388 9172
rect 11796 9052 11848 9104
rect 4160 8984 4212 9036
rect 5080 8984 5132 9036
rect 2320 8959 2372 8968
rect 2320 8925 2329 8959
rect 2329 8925 2363 8959
rect 2363 8925 2372 8959
rect 2320 8916 2372 8925
rect 7656 8984 7708 9036
rect 7840 8916 7892 8968
rect 9220 8984 9272 9036
rect 11060 8984 11112 9036
rect 11336 9027 11388 9036
rect 11336 8993 11345 9027
rect 11345 8993 11379 9027
rect 11379 8993 11388 9027
rect 11336 8984 11388 8993
rect 11152 8916 11204 8968
rect 11888 8984 11940 9036
rect 12164 9120 12216 9172
rect 14556 9120 14608 9172
rect 12716 9052 12768 9104
rect 13728 9052 13780 9104
rect 5356 8780 5408 8832
rect 7932 8780 7984 8832
rect 9128 8780 9180 8832
rect 9312 8780 9364 8832
rect 11336 8848 11388 8900
rect 11060 8780 11112 8832
rect 12440 8780 12492 8832
rect 12716 8823 12768 8832
rect 12716 8789 12725 8823
rect 12725 8789 12759 8823
rect 12759 8789 12768 8823
rect 12716 8780 12768 8789
rect 13728 8780 13780 8832
rect 14096 8848 14148 8900
rect 14280 8848 14332 8900
rect 14004 8780 14056 8832
rect 14740 8780 14792 8832
rect 3447 8678 3499 8730
rect 3511 8678 3563 8730
rect 3575 8678 3627 8730
rect 3639 8678 3691 8730
rect 8378 8678 8430 8730
rect 8442 8678 8494 8730
rect 8506 8678 8558 8730
rect 8570 8678 8622 8730
rect 13308 8678 13360 8730
rect 13372 8678 13424 8730
rect 13436 8678 13488 8730
rect 13500 8678 13552 8730
rect 1676 8440 1728 8492
rect 6920 8576 6972 8628
rect 7104 8576 7156 8628
rect 7380 8619 7432 8628
rect 7380 8585 7389 8619
rect 7389 8585 7423 8619
rect 7423 8585 7432 8619
rect 7380 8576 7432 8585
rect 5080 8508 5132 8560
rect 2320 8304 2372 8356
rect 3332 8304 3384 8356
rect 4620 8372 4672 8424
rect 7472 8440 7524 8492
rect 7564 8415 7616 8424
rect 7564 8381 7573 8415
rect 7573 8381 7607 8415
rect 7607 8381 7616 8415
rect 7564 8372 7616 8381
rect 8208 8576 8260 8628
rect 8668 8576 8720 8628
rect 8852 8576 8904 8628
rect 9128 8576 9180 8628
rect 10968 8576 11020 8628
rect 7932 8483 7984 8492
rect 7932 8449 7941 8483
rect 7941 8449 7975 8483
rect 7975 8449 7984 8483
rect 7932 8440 7984 8449
rect 8024 8372 8076 8424
rect 8208 8415 8260 8424
rect 8208 8381 8242 8415
rect 8242 8381 8260 8415
rect 8208 8372 8260 8381
rect 8576 8372 8628 8424
rect 10692 8508 10744 8560
rect 11520 8508 11572 8560
rect 11796 8508 11848 8560
rect 12348 8508 12400 8560
rect 9220 8440 9272 8492
rect 11428 8483 11480 8492
rect 10140 8372 10192 8424
rect 3884 8236 3936 8288
rect 4804 8236 4856 8288
rect 7748 8304 7800 8356
rect 5448 8236 5500 8288
rect 7012 8236 7064 8288
rect 7288 8236 7340 8288
rect 9220 8304 9272 8356
rect 8024 8236 8076 8288
rect 9956 8236 10008 8288
rect 11428 8449 11437 8483
rect 11437 8449 11471 8483
rect 11471 8449 11480 8483
rect 11428 8440 11480 8449
rect 12624 8576 12676 8628
rect 13820 8619 13872 8628
rect 13820 8585 13829 8619
rect 13829 8585 13863 8619
rect 13863 8585 13872 8619
rect 13820 8576 13872 8585
rect 13452 8508 13504 8560
rect 14096 8551 14148 8560
rect 10600 8372 10652 8424
rect 10784 8372 10836 8424
rect 11520 8372 11572 8424
rect 12440 8415 12492 8424
rect 12440 8381 12449 8415
rect 12449 8381 12483 8415
rect 12483 8381 12492 8415
rect 12440 8372 12492 8381
rect 14096 8517 14105 8551
rect 14105 8517 14139 8551
rect 14139 8517 14148 8551
rect 14096 8508 14148 8517
rect 13636 8440 13688 8492
rect 14004 8304 14056 8356
rect 13084 8236 13136 8288
rect 13728 8236 13780 8288
rect 14556 8347 14608 8356
rect 14556 8313 14565 8347
rect 14565 8313 14599 8347
rect 14599 8313 14608 8347
rect 14556 8304 14608 8313
rect 15108 8279 15160 8288
rect 15108 8245 15117 8279
rect 15117 8245 15151 8279
rect 15151 8245 15160 8279
rect 15108 8236 15160 8245
rect 5912 8134 5964 8186
rect 5976 8134 6028 8186
rect 6040 8134 6092 8186
rect 6104 8134 6156 8186
rect 10843 8134 10895 8186
rect 10907 8134 10959 8186
rect 10971 8134 11023 8186
rect 11035 8134 11087 8186
rect 3700 8075 3752 8084
rect 3700 8041 3709 8075
rect 3709 8041 3743 8075
rect 3743 8041 3752 8075
rect 3700 8032 3752 8041
rect 2136 7896 2188 7948
rect 2320 7939 2372 7948
rect 2320 7905 2329 7939
rect 2329 7905 2363 7939
rect 2363 7905 2372 7939
rect 2320 7896 2372 7905
rect 4896 8032 4948 8084
rect 6920 8032 6972 8084
rect 8208 8032 8260 8084
rect 8944 8032 8996 8084
rect 4160 7964 4212 8016
rect 5540 7964 5592 8016
rect 5172 7896 5224 7948
rect 6644 7896 6696 7948
rect 7196 7896 7248 7948
rect 7932 7964 7984 8016
rect 7656 7896 7708 7948
rect 8576 7964 8628 8016
rect 8116 7896 8168 7948
rect 1768 7871 1820 7880
rect 1768 7837 1777 7871
rect 1777 7837 1811 7871
rect 1811 7837 1820 7871
rect 1768 7828 1820 7837
rect 3332 7828 3384 7880
rect 4620 7871 4672 7880
rect 4620 7837 4629 7871
rect 4629 7837 4663 7871
rect 4663 7837 4672 7871
rect 4620 7828 4672 7837
rect 7288 7828 7340 7880
rect 8576 7828 8628 7880
rect 10508 8032 10560 8084
rect 12532 8032 12584 8084
rect 10140 7964 10192 8016
rect 9956 7939 10008 7948
rect 9956 7905 9990 7939
rect 9990 7905 10008 7939
rect 9956 7896 10008 7905
rect 11704 7964 11756 8016
rect 12624 7964 12676 8016
rect 14648 7964 14700 8016
rect 12440 7896 12492 7948
rect 13176 7896 13228 7948
rect 12348 7828 12400 7880
rect 1308 7692 1360 7744
rect 7472 7735 7524 7744
rect 7472 7701 7481 7735
rect 7481 7701 7515 7735
rect 7515 7701 7524 7735
rect 7472 7692 7524 7701
rect 8944 7735 8996 7744
rect 8944 7701 8953 7735
rect 8953 7701 8987 7735
rect 8987 7701 8996 7735
rect 8944 7692 8996 7701
rect 9220 7692 9272 7744
rect 11152 7692 11204 7744
rect 12716 7735 12768 7744
rect 12716 7701 12725 7735
rect 12725 7701 12759 7735
rect 12759 7701 12768 7735
rect 12716 7692 12768 7701
rect 12808 7692 12860 7744
rect 13820 7760 13872 7812
rect 14004 7803 14056 7812
rect 14004 7769 14013 7803
rect 14013 7769 14047 7803
rect 14047 7769 14056 7803
rect 14004 7760 14056 7769
rect 14280 7828 14332 7880
rect 3447 7590 3499 7642
rect 3511 7590 3563 7642
rect 3575 7590 3627 7642
rect 3639 7590 3691 7642
rect 8378 7590 8430 7642
rect 8442 7590 8494 7642
rect 8506 7590 8558 7642
rect 8570 7590 8622 7642
rect 13308 7590 13360 7642
rect 13372 7590 13424 7642
rect 13436 7590 13488 7642
rect 13500 7590 13552 7642
rect 5816 7488 5868 7540
rect 4804 7463 4856 7472
rect 4804 7429 4813 7463
rect 4813 7429 4847 7463
rect 4847 7429 4856 7463
rect 4804 7420 4856 7429
rect 8024 7420 8076 7472
rect 9220 7488 9272 7540
rect 2228 7284 2280 7336
rect 2780 7284 2832 7336
rect 4620 7352 4672 7404
rect 6092 7352 6144 7404
rect 3332 7284 3384 7336
rect 3691 7327 3743 7336
rect 3691 7293 3700 7327
rect 3700 7293 3734 7327
rect 3734 7293 3743 7327
rect 6828 7327 6880 7336
rect 3691 7284 3743 7293
rect 6828 7293 6837 7327
rect 6837 7293 6871 7327
rect 6871 7293 6880 7327
rect 6828 7284 6880 7293
rect 7932 7352 7984 7404
rect 11336 7420 11388 7472
rect 12072 7420 12124 7472
rect 14004 7488 14056 7540
rect 12532 7420 12584 7472
rect 10140 7395 10192 7404
rect 10140 7361 10149 7395
rect 10149 7361 10183 7395
rect 10183 7361 10192 7395
rect 10140 7352 10192 7361
rect 11428 7352 11480 7404
rect 12348 7352 12400 7404
rect 13084 7352 13136 7404
rect 14096 7420 14148 7472
rect 14464 7420 14516 7472
rect 10968 7284 11020 7336
rect 4712 7216 4764 7268
rect 6092 7216 6144 7268
rect 6368 7216 6420 7268
rect 7472 7216 7524 7268
rect 7564 7216 7616 7268
rect 8576 7216 8628 7268
rect 8944 7216 8996 7268
rect 1860 7191 1912 7200
rect 1860 7157 1869 7191
rect 1869 7157 1903 7191
rect 1903 7157 1912 7191
rect 1860 7148 1912 7157
rect 2412 7191 2464 7200
rect 2412 7157 2421 7191
rect 2421 7157 2455 7191
rect 2455 7157 2464 7191
rect 2412 7148 2464 7157
rect 4620 7148 4672 7200
rect 5080 7148 5132 7200
rect 5724 7148 5776 7200
rect 7288 7148 7340 7200
rect 8668 7148 8720 7200
rect 11152 7216 11204 7268
rect 10324 7148 10376 7200
rect 11428 7216 11480 7268
rect 12624 7284 12676 7336
rect 14280 7352 14332 7404
rect 15016 7395 15068 7404
rect 15016 7361 15025 7395
rect 15025 7361 15059 7395
rect 15059 7361 15068 7395
rect 15016 7352 15068 7361
rect 11336 7148 11388 7200
rect 12348 7216 12400 7268
rect 13360 7216 13412 7268
rect 14096 7216 14148 7268
rect 12624 7148 12676 7200
rect 12900 7191 12952 7200
rect 12900 7157 12909 7191
rect 12909 7157 12943 7191
rect 12943 7157 12952 7191
rect 12900 7148 12952 7157
rect 13452 7191 13504 7200
rect 13452 7157 13461 7191
rect 13461 7157 13495 7191
rect 13495 7157 13504 7191
rect 13452 7148 13504 7157
rect 14556 7284 14608 7336
rect 15108 7284 15160 7336
rect 14280 7216 14332 7268
rect 14832 7191 14884 7200
rect 14832 7157 14841 7191
rect 14841 7157 14875 7191
rect 14875 7157 14884 7191
rect 14832 7148 14884 7157
rect 5912 7046 5964 7098
rect 5976 7046 6028 7098
rect 6040 7046 6092 7098
rect 6104 7046 6156 7098
rect 10843 7046 10895 7098
rect 10907 7046 10959 7098
rect 10971 7046 11023 7098
rect 11035 7046 11087 7098
rect 2412 6944 2464 6996
rect 8852 6944 8904 6996
rect 9036 6987 9088 6996
rect 9036 6953 9045 6987
rect 9045 6953 9079 6987
rect 9079 6953 9088 6987
rect 9036 6944 9088 6953
rect 10140 6944 10192 6996
rect 11336 6987 11388 6996
rect 11336 6953 11345 6987
rect 11345 6953 11379 6987
rect 11379 6953 11388 6987
rect 11336 6944 11388 6953
rect 11888 6944 11940 6996
rect 12348 6944 12400 6996
rect 12900 6944 12952 6996
rect 14096 6944 14148 6996
rect 2504 6876 2556 6928
rect 5632 6876 5684 6928
rect 1952 6808 2004 6860
rect 2320 6851 2372 6860
rect 2320 6817 2329 6851
rect 2329 6817 2363 6851
rect 2363 6817 2372 6851
rect 2320 6808 2372 6817
rect 4804 6808 4856 6860
rect 6828 6876 6880 6928
rect 7012 6876 7064 6928
rect 5816 6851 5868 6860
rect 5816 6817 5850 6851
rect 5850 6817 5868 6851
rect 7196 6851 7248 6860
rect 5816 6808 5868 6817
rect 7196 6817 7205 6851
rect 7205 6817 7239 6851
rect 7239 6817 7248 6851
rect 7196 6808 7248 6817
rect 7288 6808 7340 6860
rect 7748 6808 7800 6860
rect 9312 6876 9364 6928
rect 11796 6919 11848 6928
rect 1768 6783 1820 6792
rect 1768 6749 1777 6783
rect 1777 6749 1811 6783
rect 1811 6749 1820 6783
rect 1768 6740 1820 6749
rect 4068 6783 4120 6792
rect 4068 6749 4077 6783
rect 4077 6749 4111 6783
rect 4111 6749 4120 6783
rect 4068 6740 4120 6749
rect 5172 6783 5224 6792
rect 5172 6749 5181 6783
rect 5181 6749 5215 6783
rect 5215 6749 5224 6783
rect 8944 6808 8996 6860
rect 9956 6851 10008 6860
rect 9956 6817 9990 6851
rect 9990 6817 10008 6851
rect 9956 6808 10008 6817
rect 11796 6885 11805 6919
rect 11805 6885 11839 6919
rect 11839 6885 11848 6919
rect 11796 6876 11848 6885
rect 12164 6876 12216 6928
rect 13912 6876 13964 6928
rect 10784 6808 10836 6860
rect 5172 6740 5224 6749
rect 3884 6604 3936 6656
rect 3976 6604 4028 6656
rect 10692 6740 10744 6792
rect 11428 6740 11480 6792
rect 12348 6808 12400 6860
rect 13084 6808 13136 6860
rect 13176 6808 13228 6860
rect 14188 6808 14240 6860
rect 14464 6808 14516 6860
rect 15200 6808 15252 6860
rect 11980 6740 12032 6792
rect 12716 6740 12768 6792
rect 12900 6783 12952 6792
rect 12900 6749 12909 6783
rect 12909 6749 12943 6783
rect 12943 6749 12952 6783
rect 12900 6740 12952 6749
rect 6644 6672 6696 6724
rect 8208 6672 8260 6724
rect 9864 6604 9916 6656
rect 15016 6740 15068 6792
rect 11704 6604 11756 6656
rect 11888 6604 11940 6656
rect 13176 6672 13228 6724
rect 13452 6672 13504 6724
rect 12716 6604 12768 6656
rect 14188 6604 14240 6656
rect 3447 6502 3499 6554
rect 3511 6502 3563 6554
rect 3575 6502 3627 6554
rect 3639 6502 3691 6554
rect 8378 6502 8430 6554
rect 8442 6502 8494 6554
rect 8506 6502 8558 6554
rect 8570 6502 8622 6554
rect 13308 6502 13360 6554
rect 13372 6502 13424 6554
rect 13436 6502 13488 6554
rect 13500 6502 13552 6554
rect 4160 6400 4212 6452
rect 4528 6332 4580 6384
rect 2688 6264 2740 6316
rect 3056 6196 3108 6248
rect 3332 6264 3384 6316
rect 5356 6400 5408 6452
rect 5448 6400 5500 6452
rect 9864 6400 9916 6452
rect 10048 6400 10100 6452
rect 11336 6400 11388 6452
rect 11244 6332 11296 6384
rect 12716 6400 12768 6452
rect 13636 6400 13688 6452
rect 14924 6400 14976 6452
rect 12348 6332 12400 6384
rect 12900 6332 12952 6384
rect 4436 6196 4488 6248
rect 4712 6196 4764 6248
rect 5724 6196 5776 6248
rect 6276 6264 6328 6316
rect 6828 6264 6880 6316
rect 7932 6264 7984 6316
rect 8300 6264 8352 6316
rect 10140 6264 10192 6316
rect 11704 6264 11756 6316
rect 13084 6264 13136 6316
rect 14740 6332 14792 6384
rect 1400 6103 1452 6112
rect 1400 6069 1409 6103
rect 1409 6069 1443 6103
rect 1443 6069 1452 6103
rect 1400 6060 1452 6069
rect 1676 6060 1728 6112
rect 2780 6171 2832 6180
rect 2780 6137 2789 6171
rect 2789 6137 2823 6171
rect 2823 6137 2832 6171
rect 2780 6128 2832 6137
rect 3240 6128 3292 6180
rect 3700 6171 3752 6180
rect 3700 6137 3712 6171
rect 3712 6137 3752 6171
rect 3700 6128 3752 6137
rect 3792 6128 3844 6180
rect 3056 6060 3108 6112
rect 6276 6128 6328 6180
rect 7288 6128 7340 6180
rect 9036 6128 9088 6180
rect 11336 6128 11388 6180
rect 11520 6128 11572 6180
rect 11888 6196 11940 6248
rect 12072 6196 12124 6248
rect 12440 6196 12492 6248
rect 12716 6196 12768 6248
rect 13176 6196 13228 6248
rect 13268 6239 13320 6248
rect 13268 6205 13277 6239
rect 13277 6205 13311 6239
rect 13311 6205 13320 6239
rect 13268 6196 13320 6205
rect 13820 6196 13872 6248
rect 14740 6196 14792 6248
rect 13912 6128 13964 6180
rect 15016 6307 15068 6316
rect 15016 6273 15025 6307
rect 15025 6273 15059 6307
rect 15059 6273 15068 6307
rect 15016 6264 15068 6273
rect 15476 6128 15528 6180
rect 9864 6060 9916 6112
rect 9956 6060 10008 6112
rect 10232 6060 10284 6112
rect 11888 6103 11940 6112
rect 11888 6069 11897 6103
rect 11897 6069 11931 6103
rect 11931 6069 11940 6103
rect 11888 6060 11940 6069
rect 12440 6103 12492 6112
rect 12440 6069 12449 6103
rect 12449 6069 12483 6103
rect 12483 6069 12492 6103
rect 12440 6060 12492 6069
rect 13452 6060 13504 6112
rect 13820 6103 13872 6112
rect 13820 6069 13829 6103
rect 13829 6069 13863 6103
rect 13863 6069 13872 6103
rect 13820 6060 13872 6069
rect 14648 6060 14700 6112
rect 5912 5958 5964 6010
rect 5976 5958 6028 6010
rect 6040 5958 6092 6010
rect 6104 5958 6156 6010
rect 10843 5958 10895 6010
rect 10907 5958 10959 6010
rect 10971 5958 11023 6010
rect 11035 5958 11087 6010
rect 1400 5856 1452 5908
rect 8116 5856 8168 5908
rect 8576 5856 8628 5908
rect 8944 5856 8996 5908
rect 9312 5856 9364 5908
rect 1400 5763 1452 5772
rect 1400 5729 1409 5763
rect 1409 5729 1443 5763
rect 1443 5729 1452 5763
rect 1400 5720 1452 5729
rect 1768 5720 1820 5772
rect 3332 5763 3384 5772
rect 3332 5729 3341 5763
rect 3341 5729 3375 5763
rect 3375 5729 3384 5763
rect 3332 5720 3384 5729
rect 3792 5720 3844 5772
rect 4068 5763 4120 5772
rect 4068 5729 4077 5763
rect 4077 5729 4111 5763
rect 4111 5729 4120 5763
rect 4068 5720 4120 5729
rect 10232 5856 10284 5908
rect 10600 5856 10652 5908
rect 11244 5856 11296 5908
rect 11796 5856 11848 5908
rect 12440 5856 12492 5908
rect 13728 5856 13780 5908
rect 14096 5899 14148 5908
rect 14096 5865 14105 5899
rect 14105 5865 14139 5899
rect 14139 5865 14148 5899
rect 14096 5856 14148 5865
rect 14740 5899 14792 5908
rect 14740 5865 14749 5899
rect 14749 5865 14783 5899
rect 14783 5865 14792 5899
rect 14740 5856 14792 5865
rect 10692 5788 10744 5840
rect 6460 5720 6512 5772
rect 6920 5763 6972 5772
rect 6920 5729 6954 5763
rect 6954 5729 6972 5763
rect 6920 5720 6972 5729
rect 8116 5720 8168 5772
rect 8852 5720 8904 5772
rect 9496 5763 9548 5772
rect 9496 5729 9505 5763
rect 9505 5729 9539 5763
rect 9539 5729 9548 5763
rect 9496 5720 9548 5729
rect 10968 5788 11020 5840
rect 11520 5788 11572 5840
rect 11980 5788 12032 5840
rect 12808 5788 12860 5840
rect 3608 5695 3660 5704
rect 3608 5661 3617 5695
rect 3617 5661 3651 5695
rect 3651 5661 3660 5695
rect 3608 5652 3660 5661
rect 3700 5652 3752 5704
rect 4712 5652 4764 5704
rect 1952 5627 2004 5636
rect 1952 5593 1961 5627
rect 1961 5593 1995 5627
rect 1995 5593 2004 5627
rect 1952 5584 2004 5593
rect 2688 5584 2740 5636
rect 4344 5584 4396 5636
rect 2412 5516 2464 5568
rect 4160 5516 4212 5568
rect 5724 5516 5776 5568
rect 6368 5559 6420 5568
rect 6368 5525 6377 5559
rect 6377 5525 6411 5559
rect 6411 5525 6420 5559
rect 6368 5516 6420 5525
rect 9220 5652 9272 5704
rect 9312 5652 9364 5704
rect 6828 5516 6880 5568
rect 7564 5516 7616 5568
rect 7840 5516 7892 5568
rect 8760 5516 8812 5568
rect 9680 5559 9732 5568
rect 9680 5525 9689 5559
rect 9689 5525 9723 5559
rect 9723 5525 9732 5559
rect 10232 5584 10284 5636
rect 10784 5652 10836 5704
rect 11060 5652 11112 5704
rect 11428 5652 11480 5704
rect 11520 5652 11572 5704
rect 11980 5652 12032 5704
rect 14004 5720 14056 5772
rect 12900 5652 12952 5704
rect 13268 5695 13320 5704
rect 13268 5661 13277 5695
rect 13277 5661 13311 5695
rect 13311 5661 13320 5695
rect 13268 5652 13320 5661
rect 13452 5652 13504 5704
rect 14096 5652 14148 5704
rect 10692 5559 10744 5568
rect 9680 5516 9732 5525
rect 10692 5525 10701 5559
rect 10701 5525 10735 5559
rect 10735 5525 10744 5559
rect 10692 5516 10744 5525
rect 10784 5516 10836 5568
rect 12440 5584 12492 5636
rect 12716 5559 12768 5568
rect 12716 5525 12725 5559
rect 12725 5525 12759 5559
rect 12759 5525 12768 5559
rect 12716 5516 12768 5525
rect 14004 5516 14056 5568
rect 3447 5414 3499 5466
rect 3511 5414 3563 5466
rect 3575 5414 3627 5466
rect 3639 5414 3691 5466
rect 8378 5414 8430 5466
rect 8442 5414 8494 5466
rect 8506 5414 8558 5466
rect 8570 5414 8622 5466
rect 13308 5414 13360 5466
rect 13372 5414 13424 5466
rect 13436 5414 13488 5466
rect 13500 5414 13552 5466
rect 2136 5312 2188 5364
rect 3332 5312 3384 5364
rect 4160 5312 4212 5364
rect 2596 5244 2648 5296
rect 2872 5176 2924 5228
rect 3516 5219 3568 5228
rect 3516 5185 3525 5219
rect 3525 5185 3559 5219
rect 3559 5185 3568 5219
rect 3516 5176 3568 5185
rect 3884 5244 3936 5296
rect 2780 5040 2832 5092
rect 4436 5244 4488 5296
rect 6460 5287 6512 5296
rect 6460 5253 6469 5287
rect 6469 5253 6503 5287
rect 6503 5253 6512 5287
rect 6460 5244 6512 5253
rect 7840 5244 7892 5296
rect 6828 5219 6880 5228
rect 5908 5108 5960 5160
rect 6828 5185 6837 5219
rect 6837 5185 6871 5219
rect 6871 5185 6880 5219
rect 6828 5176 6880 5185
rect 8392 5176 8444 5228
rect 6368 5108 6420 5160
rect 4344 5040 4396 5092
rect 5264 5040 5316 5092
rect 7012 5040 7064 5092
rect 7932 5108 7984 5160
rect 10508 5244 10560 5296
rect 10876 5244 10928 5296
rect 12256 5312 12308 5364
rect 14464 5312 14516 5364
rect 8852 5040 8904 5092
rect 9128 5040 9180 5092
rect 9220 5040 9272 5092
rect 9404 5040 9456 5092
rect 9496 5040 9548 5092
rect 10232 5040 10284 5092
rect 10968 5176 11020 5228
rect 12348 5244 12400 5296
rect 12900 5244 12952 5296
rect 11704 5219 11756 5228
rect 11704 5185 11713 5219
rect 11713 5185 11747 5219
rect 11747 5185 11756 5219
rect 11704 5176 11756 5185
rect 11888 5176 11940 5228
rect 12532 5176 12584 5228
rect 13728 5244 13780 5296
rect 16764 5244 16816 5296
rect 13820 5176 13872 5228
rect 13912 5176 13964 5228
rect 14924 5176 14976 5228
rect 10600 5040 10652 5092
rect 10784 5040 10836 5092
rect 12624 5108 12676 5160
rect 11244 5040 11296 5092
rect 1860 5015 1912 5024
rect 1860 4981 1869 5015
rect 1869 4981 1903 5015
rect 1903 4981 1912 5015
rect 1860 4972 1912 4981
rect 2964 4972 3016 5024
rect 3332 4972 3384 5024
rect 4436 4972 4488 5024
rect 6276 4972 6328 5024
rect 8024 4972 8076 5024
rect 9588 4972 9640 5024
rect 10416 4972 10468 5024
rect 13084 5040 13136 5092
rect 14004 5040 14056 5092
rect 15016 5040 15068 5092
rect 16304 5040 16356 5092
rect 11796 4972 11848 5024
rect 12532 4972 12584 5024
rect 13268 4972 13320 5024
rect 13820 5015 13872 5024
rect 13820 4981 13829 5015
rect 13829 4981 13863 5015
rect 13863 4981 13872 5015
rect 13820 4972 13872 4981
rect 13912 5015 13964 5024
rect 13912 4981 13921 5015
rect 13921 4981 13955 5015
rect 13955 4981 13964 5015
rect 14464 5015 14516 5024
rect 13912 4972 13964 4981
rect 14464 4981 14473 5015
rect 14473 4981 14507 5015
rect 14507 4981 14516 5015
rect 14464 4972 14516 4981
rect 14648 4972 14700 5024
rect 5912 4870 5964 4922
rect 5976 4870 6028 4922
rect 6040 4870 6092 4922
rect 6104 4870 6156 4922
rect 10843 4870 10895 4922
rect 10907 4870 10959 4922
rect 10971 4870 11023 4922
rect 11035 4870 11087 4922
rect 2320 4768 2372 4820
rect 2688 4768 2740 4820
rect 4160 4768 4212 4820
rect 3884 4700 3936 4752
rect 5448 4768 5500 4820
rect 5632 4768 5684 4820
rect 9680 4768 9732 4820
rect 9864 4768 9916 4820
rect 10324 4768 10376 4820
rect 10508 4768 10560 4820
rect 1400 4675 1452 4684
rect 1400 4641 1409 4675
rect 1409 4641 1443 4675
rect 1443 4641 1452 4675
rect 1400 4632 1452 4641
rect 2320 4675 2372 4684
rect 2320 4641 2329 4675
rect 2329 4641 2363 4675
rect 2363 4641 2372 4675
rect 2320 4632 2372 4641
rect 2872 4632 2924 4684
rect 3148 4564 3200 4616
rect 3700 4632 3752 4684
rect 5908 4700 5960 4752
rect 6368 4700 6420 4752
rect 7104 4700 7156 4752
rect 8576 4700 8628 4752
rect 9128 4700 9180 4752
rect 10416 4700 10468 4752
rect 10968 4700 11020 4752
rect 11336 4768 11388 4820
rect 11704 4811 11756 4820
rect 11704 4777 11713 4811
rect 11713 4777 11747 4811
rect 11747 4777 11756 4811
rect 11704 4768 11756 4777
rect 4988 4632 5040 4684
rect 2964 4539 3016 4548
rect 1952 4471 2004 4480
rect 1952 4437 1961 4471
rect 1961 4437 1995 4471
rect 1995 4437 2004 4471
rect 1952 4428 2004 4437
rect 2964 4505 2973 4539
rect 2973 4505 3007 4539
rect 3007 4505 3016 4539
rect 2964 4496 3016 4505
rect 3608 4564 3660 4616
rect 5356 4607 5408 4616
rect 4712 4496 4764 4548
rect 5356 4573 5365 4607
rect 5365 4573 5399 4607
rect 5399 4573 5408 4607
rect 5356 4564 5408 4573
rect 5724 4564 5776 4616
rect 5816 4564 5868 4616
rect 5448 4496 5500 4548
rect 3148 4428 3200 4480
rect 3792 4428 3844 4480
rect 5264 4428 5316 4480
rect 6000 4428 6052 4480
rect 6828 4632 6880 4684
rect 7932 4632 7984 4684
rect 9956 4632 10008 4684
rect 8116 4564 8168 4616
rect 8576 4496 8628 4548
rect 9312 4564 9364 4616
rect 9772 4564 9824 4616
rect 9220 4496 9272 4548
rect 10876 4632 10928 4684
rect 11244 4700 11296 4752
rect 12532 4768 12584 4820
rect 12624 4768 12676 4820
rect 15292 4768 15344 4820
rect 12256 4700 12308 4752
rect 11980 4632 12032 4684
rect 10600 4564 10652 4616
rect 11336 4607 11388 4616
rect 11336 4573 11345 4607
rect 11345 4573 11379 4607
rect 11379 4573 11388 4607
rect 11336 4564 11388 4573
rect 11612 4496 11664 4548
rect 8116 4471 8168 4480
rect 8116 4437 8125 4471
rect 8125 4437 8159 4471
rect 8159 4437 8168 4471
rect 8116 4428 8168 4437
rect 10968 4428 11020 4480
rect 11060 4428 11112 4480
rect 11336 4428 11388 4480
rect 13176 4700 13228 4752
rect 12900 4675 12952 4684
rect 12900 4641 12909 4675
rect 12909 4641 12943 4675
rect 12943 4641 12952 4675
rect 12900 4632 12952 4641
rect 13544 4675 13596 4684
rect 13544 4641 13553 4675
rect 13553 4641 13587 4675
rect 13587 4641 13596 4675
rect 13544 4632 13596 4641
rect 12992 4607 13044 4616
rect 12992 4573 13001 4607
rect 13001 4573 13035 4607
rect 13035 4573 13044 4607
rect 12992 4564 13044 4573
rect 12900 4496 12952 4548
rect 13728 4564 13780 4616
rect 14924 4564 14976 4616
rect 12532 4471 12584 4480
rect 12532 4437 12541 4471
rect 12541 4437 12575 4471
rect 12575 4437 12584 4471
rect 12532 4428 12584 4437
rect 12624 4428 12676 4480
rect 3447 4326 3499 4378
rect 3511 4326 3563 4378
rect 3575 4326 3627 4378
rect 3639 4326 3691 4378
rect 8378 4326 8430 4378
rect 8442 4326 8494 4378
rect 8506 4326 8558 4378
rect 8570 4326 8622 4378
rect 13308 4326 13360 4378
rect 13372 4326 13424 4378
rect 13436 4326 13488 4378
rect 13500 4326 13552 4378
rect 2228 4224 2280 4276
rect 4712 4224 4764 4276
rect 4344 4156 4396 4208
rect 2136 4020 2188 4072
rect 2688 4063 2740 4072
rect 2688 4029 2697 4063
rect 2697 4029 2731 4063
rect 2731 4029 2740 4063
rect 2688 4020 2740 4029
rect 4160 4088 4212 4140
rect 4896 4088 4948 4140
rect 5356 4224 5408 4276
rect 5448 4224 5500 4276
rect 5724 4267 5776 4276
rect 5724 4233 5733 4267
rect 5733 4233 5767 4267
rect 5767 4233 5776 4267
rect 5724 4224 5776 4233
rect 6368 4224 6420 4276
rect 8944 4224 8996 4276
rect 9496 4267 9548 4276
rect 9496 4233 9505 4267
rect 9505 4233 9539 4267
rect 9539 4233 9548 4267
rect 9496 4224 9548 4233
rect 9772 4224 9824 4276
rect 5908 4156 5960 4208
rect 5816 4088 5868 4140
rect 6368 4131 6420 4140
rect 6368 4097 6377 4131
rect 6377 4097 6411 4131
rect 6411 4097 6420 4131
rect 6368 4088 6420 4097
rect 1676 3927 1728 3936
rect 1676 3893 1685 3927
rect 1685 3893 1719 3927
rect 1719 3893 1728 3927
rect 1676 3884 1728 3893
rect 2136 3927 2188 3936
rect 2136 3893 2145 3927
rect 2145 3893 2179 3927
rect 2179 3893 2188 3927
rect 2780 3952 2832 4004
rect 3608 3952 3660 4004
rect 2136 3884 2188 3893
rect 4160 3884 4212 3936
rect 4252 3884 4304 3936
rect 5724 3952 5776 4004
rect 6736 4156 6788 4208
rect 8116 4156 8168 4208
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 6828 4088 6880 4097
rect 8760 4088 8812 4140
rect 8944 4088 8996 4140
rect 9588 4088 9640 4140
rect 10140 4131 10192 4140
rect 10140 4097 10149 4131
rect 10149 4097 10183 4131
rect 10183 4097 10192 4131
rect 10140 4088 10192 4097
rect 7380 4020 7432 4072
rect 7656 4020 7708 4072
rect 9772 4020 9824 4072
rect 10324 4156 10376 4208
rect 10508 4199 10560 4208
rect 10508 4165 10517 4199
rect 10517 4165 10551 4199
rect 10551 4165 10560 4199
rect 10508 4156 10560 4165
rect 10968 4224 11020 4276
rect 12072 4224 12124 4276
rect 11060 4156 11112 4208
rect 11336 4156 11388 4208
rect 11612 4156 11664 4208
rect 10324 4020 10376 4072
rect 10600 4020 10652 4072
rect 10784 4020 10836 4072
rect 11428 4088 11480 4140
rect 12808 4156 12860 4208
rect 13912 4224 13964 4276
rect 12440 4088 12492 4140
rect 7104 3995 7156 4004
rect 7104 3961 7138 3995
rect 7138 3961 7156 3995
rect 7104 3952 7156 3961
rect 7472 3952 7524 4004
rect 4896 3884 4948 3936
rect 6276 3884 6328 3936
rect 8116 3884 8168 3936
rect 9496 3952 9548 4004
rect 12716 4020 12768 4072
rect 13544 4088 13596 4140
rect 13360 4020 13412 4072
rect 13912 4063 13964 4072
rect 13912 4029 13921 4063
rect 13921 4029 13955 4063
rect 13955 4029 13964 4063
rect 13912 4020 13964 4029
rect 11796 3952 11848 4004
rect 15200 4156 15252 4208
rect 14924 4088 14976 4140
rect 9128 3884 9180 3936
rect 9772 3884 9824 3936
rect 9864 3884 9916 3936
rect 10600 3884 10652 3936
rect 11428 3884 11480 3936
rect 12440 3927 12492 3936
rect 12440 3893 12449 3927
rect 12449 3893 12483 3927
rect 12483 3893 12492 3927
rect 12440 3884 12492 3893
rect 12716 3884 12768 3936
rect 12992 3884 13044 3936
rect 13728 3884 13780 3936
rect 14556 3884 14608 3936
rect 15108 3884 15160 3936
rect 5912 3782 5964 3834
rect 5976 3782 6028 3834
rect 6040 3782 6092 3834
rect 6104 3782 6156 3834
rect 10843 3782 10895 3834
rect 10907 3782 10959 3834
rect 10971 3782 11023 3834
rect 11035 3782 11087 3834
rect 3056 3680 3108 3732
rect 3424 3723 3476 3732
rect 3424 3689 3433 3723
rect 3433 3689 3467 3723
rect 3467 3689 3476 3723
rect 3424 3680 3476 3689
rect 4804 3723 4856 3732
rect 4804 3689 4813 3723
rect 4813 3689 4847 3723
rect 4847 3689 4856 3723
rect 4804 3680 4856 3689
rect 5448 3680 5500 3732
rect 6276 3680 6328 3732
rect 6828 3680 6880 3732
rect 1400 3587 1452 3596
rect 1400 3553 1409 3587
rect 1409 3553 1443 3587
rect 1443 3553 1452 3587
rect 1400 3544 1452 3553
rect 2872 3544 2924 3596
rect 2964 3476 3016 3528
rect 4620 3612 4672 3664
rect 5632 3612 5684 3664
rect 5816 3612 5868 3664
rect 7288 3680 7340 3732
rect 7748 3723 7800 3732
rect 7748 3689 7757 3723
rect 7757 3689 7791 3723
rect 7791 3689 7800 3723
rect 7748 3680 7800 3689
rect 7840 3680 7892 3732
rect 3332 3587 3384 3596
rect 3332 3553 3341 3587
rect 3341 3553 3375 3587
rect 3375 3553 3384 3587
rect 3332 3544 3384 3553
rect 4068 3544 4120 3596
rect 4252 3544 4304 3596
rect 8944 3612 8996 3664
rect 9128 3612 9180 3664
rect 9680 3723 9732 3732
rect 9680 3689 9689 3723
rect 9689 3689 9723 3723
rect 9723 3689 9732 3723
rect 9680 3680 9732 3689
rect 9956 3680 10008 3732
rect 10324 3680 10376 3732
rect 10416 3680 10468 3732
rect 11152 3723 11204 3732
rect 11152 3689 11161 3723
rect 11161 3689 11195 3723
rect 11195 3689 11204 3723
rect 11152 3680 11204 3689
rect 11612 3680 11664 3732
rect 11796 3680 11848 3732
rect 12256 3680 12308 3732
rect 12532 3680 12584 3732
rect 12716 3680 12768 3732
rect 12900 3680 12952 3732
rect 13176 3680 13228 3732
rect 13360 3680 13412 3732
rect 14556 3680 14608 3732
rect 14832 3680 14884 3732
rect 9864 3612 9916 3664
rect 3608 3519 3660 3528
rect 3608 3485 3617 3519
rect 3617 3485 3651 3519
rect 3651 3485 3660 3519
rect 3608 3476 3660 3485
rect 4988 3519 5040 3528
rect 4988 3485 4997 3519
rect 4997 3485 5031 3519
rect 5031 3485 5040 3519
rect 4988 3476 5040 3485
rect 5356 3476 5408 3528
rect 5816 3519 5868 3528
rect 3240 3408 3292 3460
rect 4160 3408 4212 3460
rect 5816 3485 5825 3519
rect 5825 3485 5859 3519
rect 5859 3485 5868 3519
rect 5816 3476 5868 3485
rect 6552 3476 6604 3528
rect 7656 3544 7708 3596
rect 204 3340 256 3392
rect 2504 3340 2556 3392
rect 4252 3340 4304 3392
rect 4988 3340 5040 3392
rect 5356 3383 5408 3392
rect 5356 3349 5365 3383
rect 5365 3349 5399 3383
rect 5399 3349 5408 3383
rect 5356 3340 5408 3349
rect 6736 3451 6788 3460
rect 6736 3417 6745 3451
rect 6745 3417 6779 3451
rect 6779 3417 6788 3451
rect 6736 3408 6788 3417
rect 6920 3408 6972 3460
rect 8300 3519 8352 3528
rect 8300 3485 8309 3519
rect 8309 3485 8343 3519
rect 8343 3485 8352 3519
rect 13912 3612 13964 3664
rect 14280 3612 14332 3664
rect 14924 3612 14976 3664
rect 8300 3476 8352 3485
rect 9220 3476 9272 3528
rect 9312 3476 9364 3528
rect 11336 3544 11388 3596
rect 11888 3544 11940 3596
rect 7656 3408 7708 3460
rect 7472 3340 7524 3392
rect 7840 3340 7892 3392
rect 9588 3408 9640 3460
rect 10784 3476 10836 3528
rect 10416 3408 10468 3460
rect 11796 3476 11848 3528
rect 12348 3476 12400 3528
rect 13176 3587 13228 3596
rect 13176 3553 13185 3587
rect 13185 3553 13219 3587
rect 13219 3553 13228 3587
rect 13176 3544 13228 3553
rect 9312 3340 9364 3392
rect 12716 3451 12768 3460
rect 12716 3417 12725 3451
rect 12725 3417 12759 3451
rect 12759 3417 12768 3451
rect 12716 3408 12768 3417
rect 13544 3476 13596 3528
rect 13912 3476 13964 3528
rect 14004 3476 14056 3528
rect 13268 3408 13320 3460
rect 12808 3340 12860 3392
rect 3447 3238 3499 3290
rect 3511 3238 3563 3290
rect 3575 3238 3627 3290
rect 3639 3238 3691 3290
rect 8378 3238 8430 3290
rect 8442 3238 8494 3290
rect 8506 3238 8558 3290
rect 8570 3238 8622 3290
rect 13308 3238 13360 3290
rect 13372 3238 13424 3290
rect 13436 3238 13488 3290
rect 13500 3238 13552 3290
rect 1584 3136 1636 3188
rect 2136 3136 2188 3188
rect 3240 3136 3292 3188
rect 3884 3136 3936 3188
rect 5080 3136 5132 3188
rect 5448 3136 5500 3188
rect 5540 3136 5592 3188
rect 5816 3136 5868 3188
rect 7012 3136 7064 3188
rect 7840 3136 7892 3188
rect 1860 3068 1912 3120
rect 2412 3068 2464 3120
rect 2228 3043 2280 3052
rect 2228 3009 2237 3043
rect 2237 3009 2271 3043
rect 2271 3009 2280 3043
rect 2228 3000 2280 3009
rect 4252 3043 4304 3052
rect 4252 3009 4261 3043
rect 4261 3009 4295 3043
rect 4295 3009 4304 3043
rect 4252 3000 4304 3009
rect 4988 3068 5040 3120
rect 4528 3000 4580 3052
rect 5172 3043 5224 3052
rect 5172 3009 5181 3043
rect 5181 3009 5215 3043
rect 5215 3009 5224 3043
rect 5172 3000 5224 3009
rect 5448 3000 5500 3052
rect 6460 3000 6512 3052
rect 7564 3000 7616 3052
rect 6276 2932 6328 2984
rect 10692 3136 10744 3188
rect 2964 2864 3016 2916
rect 5632 2864 5684 2916
rect 7104 2864 7156 2916
rect 8392 2932 8444 2984
rect 8668 2932 8720 2984
rect 8852 2932 8904 2984
rect 9312 3043 9364 3052
rect 9312 3009 9321 3043
rect 9321 3009 9355 3043
rect 9355 3009 9364 3043
rect 9312 3000 9364 3009
rect 9680 3000 9732 3052
rect 10416 3068 10468 3120
rect 12256 3136 12308 3188
rect 13636 3179 13688 3188
rect 13636 3145 13645 3179
rect 13645 3145 13679 3179
rect 13679 3145 13688 3179
rect 13636 3136 13688 3145
rect 9956 3000 10008 3052
rect 10324 3043 10376 3052
rect 10324 3009 10333 3043
rect 10333 3009 10367 3043
rect 10367 3009 10376 3043
rect 10324 3000 10376 3009
rect 10692 3000 10744 3052
rect 11244 3000 11296 3052
rect 11796 3000 11848 3052
rect 10048 2932 10100 2984
rect 12532 3068 12584 3120
rect 12808 3068 12860 3120
rect 12164 3000 12216 3052
rect 12624 3000 12676 3052
rect 13268 3068 13320 3120
rect 9956 2864 10008 2916
rect 10600 2864 10652 2916
rect 10784 2864 10836 2916
rect 11704 2864 11756 2916
rect 12532 2932 12584 2984
rect 13268 2932 13320 2984
rect 13452 2975 13504 2984
rect 13452 2941 13461 2975
rect 13461 2941 13495 2975
rect 13495 2941 13504 2975
rect 13452 2932 13504 2941
rect 13728 3000 13780 3052
rect 13912 2932 13964 2984
rect 14372 2932 14424 2984
rect 1400 2796 1452 2848
rect 3884 2796 3936 2848
rect 4068 2839 4120 2848
rect 4068 2805 4077 2839
rect 4077 2805 4111 2839
rect 4111 2805 4120 2839
rect 4068 2796 4120 2805
rect 5724 2796 5776 2848
rect 6920 2796 6972 2848
rect 7748 2796 7800 2848
rect 8208 2839 8260 2848
rect 8208 2805 8217 2839
rect 8217 2805 8251 2839
rect 8251 2805 8260 2839
rect 8208 2796 8260 2805
rect 8300 2796 8352 2848
rect 9312 2796 9364 2848
rect 9404 2796 9456 2848
rect 11520 2796 11572 2848
rect 12348 2796 12400 2848
rect 12624 2864 12676 2916
rect 12900 2796 12952 2848
rect 14740 2839 14792 2848
rect 14740 2805 14749 2839
rect 14749 2805 14783 2839
rect 14783 2805 14792 2839
rect 14740 2796 14792 2805
rect 5912 2694 5964 2746
rect 5976 2694 6028 2746
rect 6040 2694 6092 2746
rect 6104 2694 6156 2746
rect 10843 2694 10895 2746
rect 10907 2694 10959 2746
rect 10971 2694 11023 2746
rect 11035 2694 11087 2746
rect 2964 2635 3016 2644
rect 2964 2601 2973 2635
rect 2973 2601 3007 2635
rect 3007 2601 3016 2635
rect 2964 2592 3016 2601
rect 4068 2592 4120 2644
rect 5172 2635 5224 2644
rect 1952 2456 2004 2508
rect 5172 2601 5181 2635
rect 5181 2601 5215 2635
rect 5215 2601 5224 2635
rect 5172 2592 5224 2601
rect 5448 2592 5500 2644
rect 6276 2635 6328 2644
rect 4896 2524 4948 2576
rect 6276 2601 6285 2635
rect 6285 2601 6319 2635
rect 6319 2601 6328 2635
rect 6276 2592 6328 2601
rect 8392 2592 8444 2644
rect 10508 2592 10560 2644
rect 12716 2592 12768 2644
rect 12900 2592 12952 2644
rect 13176 2592 13228 2644
rect 5908 2524 5960 2576
rect 10692 2524 10744 2576
rect 12992 2524 13044 2576
rect 3976 2456 4028 2508
rect 6184 2499 6236 2508
rect 6184 2465 6193 2499
rect 6193 2465 6227 2499
rect 6227 2465 6236 2499
rect 6184 2456 6236 2465
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 2412 2431 2464 2440
rect 2412 2397 2421 2431
rect 2421 2397 2455 2431
rect 2455 2397 2464 2431
rect 2412 2388 2464 2397
rect 3516 2431 3568 2440
rect 3516 2397 3525 2431
rect 3525 2397 3559 2431
rect 3559 2397 3568 2431
rect 3516 2388 3568 2397
rect 3608 2388 3660 2440
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 5448 2388 5500 2397
rect 7840 2456 7892 2508
rect 8024 2456 8076 2508
rect 6644 2388 6696 2440
rect 7932 2388 7984 2440
rect 8944 2388 8996 2440
rect 9128 2499 9180 2508
rect 9128 2465 9137 2499
rect 9137 2465 9171 2499
rect 9171 2465 9180 2499
rect 10140 2499 10192 2508
rect 9128 2456 9180 2465
rect 1032 2320 1084 2372
rect 10140 2465 10149 2499
rect 10149 2465 10183 2499
rect 10183 2465 10192 2499
rect 10140 2456 10192 2465
rect 11796 2499 11848 2508
rect 10416 2431 10468 2440
rect 10416 2397 10425 2431
rect 10425 2397 10459 2431
rect 10459 2397 10468 2431
rect 10416 2388 10468 2397
rect 11152 2388 11204 2440
rect 11796 2465 11805 2499
rect 11805 2465 11839 2499
rect 11839 2465 11848 2499
rect 11796 2456 11848 2465
rect 14924 2524 14976 2576
rect 13176 2499 13228 2508
rect 13176 2465 13185 2499
rect 13185 2465 13219 2499
rect 13219 2465 13228 2499
rect 13176 2456 13228 2465
rect 13084 2388 13136 2440
rect 11428 2320 11480 2372
rect 13452 2320 13504 2372
rect 15292 2456 15344 2508
rect 5356 2252 5408 2304
rect 7104 2295 7156 2304
rect 7104 2261 7113 2295
rect 7113 2261 7147 2295
rect 7147 2261 7156 2295
rect 7104 2252 7156 2261
rect 8116 2295 8168 2304
rect 8116 2261 8125 2295
rect 8125 2261 8159 2295
rect 8159 2261 8168 2295
rect 8116 2252 8168 2261
rect 9772 2295 9824 2304
rect 9772 2261 9781 2295
rect 9781 2261 9815 2295
rect 9815 2261 9824 2295
rect 9772 2252 9824 2261
rect 10600 2252 10652 2304
rect 11980 2295 12032 2304
rect 11980 2261 11989 2295
rect 11989 2261 12023 2295
rect 12023 2261 12032 2295
rect 11980 2252 12032 2261
rect 13912 2295 13964 2304
rect 13912 2261 13921 2295
rect 13921 2261 13955 2295
rect 13955 2261 13964 2295
rect 13912 2252 13964 2261
rect 14464 2295 14516 2304
rect 14464 2261 14473 2295
rect 14473 2261 14507 2295
rect 14507 2261 14516 2295
rect 14464 2252 14516 2261
rect 14556 2252 14608 2304
rect 3447 2150 3499 2202
rect 3511 2150 3563 2202
rect 3575 2150 3627 2202
rect 3639 2150 3691 2202
rect 8378 2150 8430 2202
rect 8442 2150 8494 2202
rect 8506 2150 8558 2202
rect 8570 2150 8622 2202
rect 13308 2150 13360 2202
rect 13372 2150 13424 2202
rect 13436 2150 13488 2202
rect 13500 2150 13552 2202
rect 4068 2048 4120 2100
rect 7288 2048 7340 2100
rect 7380 2048 7432 2100
rect 14464 2048 14516 2100
rect 1768 1980 1820 2032
rect 8208 1980 8260 2032
rect 11704 1980 11756 2032
rect 12624 1980 12676 2032
rect 6552 1912 6604 1964
rect 13912 1912 13964 1964
rect 4436 1844 4488 1896
rect 12900 1844 12952 1896
rect 5448 1776 5500 1828
rect 9404 1776 9456 1828
rect 10140 1776 10192 1828
rect 12440 1776 12492 1828
rect 13360 1776 13412 1828
rect 572 1708 624 1760
rect 11980 1708 12032 1760
rect 3332 1640 3384 1692
rect 8208 1640 8260 1692
rect 14096 1640 14148 1692
rect 6092 1572 6144 1624
rect 11428 1572 11480 1624
rect 5540 1504 5592 1556
rect 9772 1504 9824 1556
rect 2872 1436 2924 1488
rect 10600 1436 10652 1488
rect 3976 1368 4028 1420
rect 7656 1368 7708 1420
rect 7840 1368 7892 1420
rect 14556 1368 14608 1420
rect 7748 1300 7800 1352
rect 13176 1300 13228 1352
rect 7472 1232 7524 1284
rect 14280 1232 14332 1284
rect 9496 1164 9548 1216
rect 10416 1164 10468 1216
rect 15108 1164 15160 1216
rect 9312 1096 9364 1148
rect 12164 1096 12216 1148
rect 12900 892 12952 944
rect 13728 892 13780 944
rect 1860 552 1912 604
rect 11336 552 11388 604
<< metal2 >>
rect 202 17520 258 18000
rect 570 17520 626 18000
rect 1030 17520 1086 18000
rect 1398 17520 1454 18000
rect 1858 17520 1914 18000
rect 2318 17520 2374 18000
rect 2686 17520 2742 18000
rect 3146 17520 3202 18000
rect 3606 17520 3662 18000
rect 3974 17520 4030 18000
rect 4434 17520 4490 18000
rect 4802 17520 4858 18000
rect 5262 17520 5318 18000
rect 5722 17520 5778 18000
rect 6090 17520 6146 18000
rect 6550 17520 6606 18000
rect 7010 17520 7066 18000
rect 7378 17520 7434 18000
rect 7838 17520 7894 18000
rect 8206 17520 8262 18000
rect 8666 17520 8722 18000
rect 9126 17520 9182 18000
rect 9494 17520 9550 18000
rect 9954 17520 10010 18000
rect 10414 17520 10470 18000
rect 10782 17520 10838 18000
rect 11242 17520 11298 18000
rect 11610 17520 11666 18000
rect 12070 17520 12126 18000
rect 12530 17520 12586 18000
rect 12898 17520 12954 18000
rect 13358 17520 13414 18000
rect 13818 17520 13874 18000
rect 14186 17520 14242 18000
rect 14646 17520 14702 18000
rect 15014 17520 15070 18000
rect 15474 17520 15530 18000
rect 15934 17520 15990 18000
rect 16302 17520 16358 18000
rect 16762 17520 16818 18000
rect 216 14618 244 17520
rect 584 15094 612 17520
rect 1044 15978 1072 17520
rect 1032 15972 1084 15978
rect 1032 15914 1084 15920
rect 1412 15162 1440 17520
rect 1400 15156 1452 15162
rect 1400 15098 1452 15104
rect 572 15088 624 15094
rect 572 15030 624 15036
rect 1872 15026 1900 17520
rect 2044 15632 2096 15638
rect 2044 15574 2096 15580
rect 1860 15020 1912 15026
rect 1860 14962 1912 14968
rect 204 14612 256 14618
rect 204 14554 256 14560
rect 1860 14476 1912 14482
rect 1860 14418 1912 14424
rect 1872 13841 1900 14418
rect 1858 13832 1914 13841
rect 1858 13767 1914 13776
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 1584 12640 1636 12646
rect 1584 12582 1636 12588
rect 1492 12096 1544 12102
rect 1492 12038 1544 12044
rect 1504 10062 1532 12038
rect 1596 10130 1624 12582
rect 1688 12073 1716 13262
rect 2056 12730 2084 15574
rect 2332 15065 2360 17520
rect 2700 15434 2728 17520
rect 2962 16280 3018 16289
rect 2962 16215 3018 16224
rect 2780 15496 2832 15502
rect 2780 15438 2832 15444
rect 2688 15428 2740 15434
rect 2688 15370 2740 15376
rect 2318 15056 2374 15065
rect 2318 14991 2374 15000
rect 2792 14958 2820 15438
rect 2870 15192 2926 15201
rect 2870 15127 2926 15136
rect 2228 14952 2280 14958
rect 2226 14920 2228 14929
rect 2780 14952 2832 14958
rect 2280 14920 2282 14929
rect 2780 14894 2832 14900
rect 2226 14855 2282 14864
rect 2780 14272 2832 14278
rect 2780 14214 2832 14220
rect 2792 14006 2820 14214
rect 2780 14000 2832 14006
rect 2502 13968 2558 13977
rect 2228 13932 2280 13938
rect 2780 13942 2832 13948
rect 2502 13903 2558 13912
rect 2228 13874 2280 13880
rect 2136 13864 2188 13870
rect 2136 13806 2188 13812
rect 1964 12702 2084 12730
rect 1964 12322 1992 12702
rect 2044 12640 2096 12646
rect 2044 12582 2096 12588
rect 2056 12442 2084 12582
rect 2044 12436 2096 12442
rect 2044 12378 2096 12384
rect 1780 12294 1992 12322
rect 2042 12336 2098 12345
rect 1674 12064 1730 12073
rect 1674 11999 1730 12008
rect 1676 11552 1728 11558
rect 1676 11494 1728 11500
rect 1584 10124 1636 10130
rect 1584 10066 1636 10072
rect 1492 10056 1544 10062
rect 1492 9998 1544 10004
rect 1504 9586 1532 9998
rect 1492 9580 1544 9586
rect 1492 9522 1544 9528
rect 1688 8498 1716 11494
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1780 8004 1808 12294
rect 2042 12271 2098 12280
rect 2056 11354 2084 12271
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 2044 11076 2096 11082
rect 2044 11018 2096 11024
rect 1858 10976 1914 10985
rect 1858 10911 1914 10920
rect 1872 10198 1900 10911
rect 1950 10704 2006 10713
rect 1950 10639 2006 10648
rect 1964 10606 1992 10639
rect 1952 10600 2004 10606
rect 1952 10542 2004 10548
rect 1860 10192 1912 10198
rect 1860 10134 1912 10140
rect 1858 9888 1914 9897
rect 1858 9823 1914 9832
rect 1872 9110 1900 9823
rect 1860 9104 1912 9110
rect 1860 9046 1912 9052
rect 1596 7976 1808 8004
rect 1308 7744 1360 7750
rect 1308 7686 1360 7692
rect 1320 3641 1348 7686
rect 1400 6112 1452 6118
rect 1400 6054 1452 6060
rect 1412 5914 1440 6054
rect 1400 5908 1452 5914
rect 1400 5850 1452 5856
rect 1398 5808 1454 5817
rect 1398 5743 1400 5752
rect 1452 5743 1454 5752
rect 1400 5714 1452 5720
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 1412 4185 1440 4626
rect 1398 4176 1454 4185
rect 1398 4111 1454 4120
rect 1306 3632 1362 3641
rect 1306 3567 1362 3576
rect 1400 3596 1452 3602
rect 1400 3538 1452 3544
rect 204 3392 256 3398
rect 204 3334 256 3340
rect 216 480 244 3334
rect 1412 2854 1440 3538
rect 1596 3194 1624 7976
rect 1768 7880 1820 7886
rect 1766 7848 1768 7857
rect 1820 7848 1822 7857
rect 1766 7783 1822 7792
rect 1860 7200 1912 7206
rect 1860 7142 1912 7148
rect 1768 6792 1820 6798
rect 1766 6760 1768 6769
rect 1820 6760 1822 6769
rect 1766 6695 1822 6704
rect 1676 6112 1728 6118
rect 1676 6054 1728 6060
rect 1688 3942 1716 6054
rect 1768 5772 1820 5778
rect 1768 5714 1820 5720
rect 1676 3936 1728 3942
rect 1676 3878 1728 3884
rect 1584 3188 1636 3194
rect 1584 3130 1636 3136
rect 1490 3088 1546 3097
rect 1490 3023 1546 3032
rect 1400 2848 1452 2854
rect 1400 2790 1452 2796
rect 1032 2372 1084 2378
rect 1032 2314 1084 2320
rect 572 1760 624 1766
rect 572 1702 624 1708
rect 584 480 612 1702
rect 1044 480 1072 2314
rect 1504 1714 1532 3023
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 1412 1686 1532 1714
rect 1412 480 1440 1686
rect 1688 1465 1716 2382
rect 1780 2038 1808 5714
rect 1872 5216 1900 7142
rect 1952 6860 2004 6866
rect 1952 6802 2004 6808
rect 1964 5642 1992 6802
rect 1952 5636 2004 5642
rect 1952 5578 2004 5584
rect 1872 5188 1992 5216
rect 1858 5128 1914 5137
rect 1858 5063 1914 5072
rect 1872 5030 1900 5063
rect 1860 5024 1912 5030
rect 1860 4966 1912 4972
rect 1858 4720 1914 4729
rect 1858 4655 1914 4664
rect 1872 3126 1900 4655
rect 1964 4570 1992 5188
rect 2056 4729 2084 11018
rect 2148 10470 2176 13806
rect 2136 10464 2188 10470
rect 2136 10406 2188 10412
rect 2136 7948 2188 7954
rect 2136 7890 2188 7896
rect 2148 5370 2176 7890
rect 2240 7857 2268 13874
rect 2516 12374 2544 13903
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2688 13728 2740 13734
rect 2688 13670 2740 13676
rect 2596 12776 2648 12782
rect 2596 12718 2648 12724
rect 2504 12368 2556 12374
rect 2318 12336 2374 12345
rect 2504 12310 2556 12316
rect 2318 12271 2320 12280
rect 2372 12271 2374 12280
rect 2320 12242 2372 12248
rect 2608 12238 2636 12718
rect 2412 12232 2464 12238
rect 2410 12200 2412 12209
rect 2596 12232 2648 12238
rect 2464 12200 2466 12209
rect 2596 12174 2648 12180
rect 2410 12135 2466 12144
rect 2410 11656 2466 11665
rect 2410 11591 2412 11600
rect 2464 11591 2466 11600
rect 2412 11562 2464 11568
rect 2504 11552 2556 11558
rect 2504 11494 2556 11500
rect 2516 11257 2544 11494
rect 2502 11248 2558 11257
rect 2502 11183 2558 11192
rect 2504 11144 2556 11150
rect 2502 11112 2504 11121
rect 2556 11112 2558 11121
rect 2502 11047 2558 11056
rect 2320 10600 2372 10606
rect 2320 10542 2372 10548
rect 2410 10568 2466 10577
rect 2332 10062 2360 10542
rect 2410 10503 2466 10512
rect 2424 10470 2452 10503
rect 2412 10464 2464 10470
rect 2412 10406 2464 10412
rect 2320 10056 2372 10062
rect 2320 9998 2372 10004
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2332 8974 2360 9454
rect 2608 9382 2636 12174
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 2608 9110 2636 9318
rect 2700 9110 2728 13670
rect 2792 13161 2820 13806
rect 2884 13394 2912 15127
rect 2976 15042 3004 16215
rect 3160 15910 3188 17520
rect 3332 15972 3384 15978
rect 3332 15914 3384 15920
rect 3148 15904 3200 15910
rect 3148 15846 3200 15852
rect 3056 15360 3108 15366
rect 3056 15302 3108 15308
rect 3068 15162 3096 15302
rect 3056 15156 3108 15162
rect 3056 15098 3108 15104
rect 3148 15156 3200 15162
rect 3148 15098 3200 15104
rect 3160 15065 3188 15098
rect 3344 15094 3372 15914
rect 3620 15706 3648 17520
rect 3988 17490 4016 17520
rect 3896 17462 4016 17490
rect 3608 15700 3660 15706
rect 3608 15642 3660 15648
rect 3792 15564 3844 15570
rect 3792 15506 3844 15512
rect 3421 15260 3717 15280
rect 3477 15258 3501 15260
rect 3557 15258 3581 15260
rect 3637 15258 3661 15260
rect 3499 15206 3501 15258
rect 3563 15206 3575 15258
rect 3637 15206 3639 15258
rect 3477 15204 3501 15206
rect 3557 15204 3581 15206
rect 3637 15204 3661 15206
rect 3421 15184 3717 15204
rect 3332 15088 3384 15094
rect 3146 15056 3202 15065
rect 2976 15014 3096 15042
rect 2964 14476 3016 14482
rect 2964 14418 3016 14424
rect 2976 14074 3004 14418
rect 2964 14068 3016 14074
rect 2964 14010 3016 14016
rect 3068 13938 3096 15014
rect 3332 15030 3384 15036
rect 3146 14991 3202 15000
rect 3240 14952 3292 14958
rect 3700 14952 3752 14958
rect 3240 14894 3292 14900
rect 3698 14920 3700 14929
rect 3752 14920 3754 14929
rect 3148 14408 3200 14414
rect 3148 14350 3200 14356
rect 3160 14113 3188 14350
rect 3146 14104 3202 14113
rect 3146 14039 3202 14048
rect 3252 13954 3280 14894
rect 3698 14855 3754 14864
rect 3804 14618 3832 15506
rect 3792 14612 3844 14618
rect 3792 14554 3844 14560
rect 3332 14476 3384 14482
rect 3332 14418 3384 14424
rect 3056 13932 3108 13938
rect 3056 13874 3108 13880
rect 3160 13926 3280 13954
rect 3160 13818 3188 13926
rect 3068 13790 3188 13818
rect 3240 13796 3292 13802
rect 3068 13394 3096 13790
rect 3240 13738 3292 13744
rect 2872 13388 2924 13394
rect 2872 13330 2924 13336
rect 3056 13388 3108 13394
rect 3056 13330 3108 13336
rect 2964 13320 3016 13326
rect 2964 13262 3016 13268
rect 2778 13152 2834 13161
rect 2778 13087 2834 13096
rect 2778 12880 2834 12889
rect 2778 12815 2834 12824
rect 2872 12844 2924 12850
rect 2792 10674 2820 12815
rect 2872 12786 2924 12792
rect 2780 10668 2832 10674
rect 2780 10610 2832 10616
rect 2596 9104 2648 9110
rect 2596 9046 2648 9052
rect 2688 9104 2740 9110
rect 2688 9046 2740 9052
rect 2320 8968 2372 8974
rect 2320 8910 2372 8916
rect 2320 8356 2372 8362
rect 2320 8298 2372 8304
rect 2332 7954 2360 8298
rect 2320 7948 2372 7954
rect 2320 7890 2372 7896
rect 2226 7848 2282 7857
rect 2226 7783 2282 7792
rect 2228 7336 2280 7342
rect 2228 7278 2280 7284
rect 2136 5364 2188 5370
rect 2136 5306 2188 5312
rect 2042 4720 2098 4729
rect 2042 4655 2098 4664
rect 1964 4542 2084 4570
rect 1952 4480 2004 4486
rect 1952 4422 2004 4428
rect 1860 3120 1912 3126
rect 1860 3062 1912 3068
rect 1964 2514 1992 4422
rect 2056 3913 2084 4542
rect 2240 4434 2268 7278
rect 2332 6866 2360 7890
rect 2792 7342 2820 10610
rect 2884 9178 2912 12786
rect 2976 11082 3004 13262
rect 3068 12889 3096 13330
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 3054 12880 3110 12889
rect 3160 12850 3188 13126
rect 3054 12815 3110 12824
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 3252 12442 3280 13738
rect 3240 12436 3292 12442
rect 3240 12378 3292 12384
rect 3148 12368 3200 12374
rect 3148 12310 3200 12316
rect 3056 11552 3108 11558
rect 3056 11494 3108 11500
rect 3068 11354 3096 11494
rect 3056 11348 3108 11354
rect 3056 11290 3108 11296
rect 2964 11076 3016 11082
rect 2964 11018 3016 11024
rect 3056 11076 3108 11082
rect 3056 11018 3108 11024
rect 3068 10962 3096 11018
rect 2976 10934 3096 10962
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2870 7440 2926 7449
rect 2870 7375 2926 7384
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 2412 7200 2464 7206
rect 2412 7142 2464 7148
rect 2424 7002 2452 7142
rect 2412 6996 2464 7002
rect 2412 6938 2464 6944
rect 2504 6928 2556 6934
rect 2504 6870 2556 6876
rect 2320 6860 2372 6866
rect 2320 6802 2372 6808
rect 2332 4826 2360 6802
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2320 4820 2372 4826
rect 2320 4762 2372 4768
rect 2320 4684 2372 4690
rect 2320 4626 2372 4632
rect 2148 4406 2268 4434
rect 2148 4078 2176 4406
rect 2228 4276 2280 4282
rect 2228 4218 2280 4224
rect 2136 4072 2188 4078
rect 2136 4014 2188 4020
rect 2136 3936 2188 3942
rect 2042 3904 2098 3913
rect 2136 3878 2188 3884
rect 2042 3839 2098 3848
rect 2148 3194 2176 3878
rect 2136 3188 2188 3194
rect 2136 3130 2188 3136
rect 2240 3058 2268 4218
rect 2332 3505 2360 4626
rect 2318 3496 2374 3505
rect 2318 3431 2374 3440
rect 2424 3346 2452 5510
rect 2516 3398 2544 6870
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 2700 5642 2728 6258
rect 2778 6216 2834 6225
rect 2778 6151 2780 6160
rect 2832 6151 2834 6160
rect 2780 6122 2832 6128
rect 2688 5636 2740 5642
rect 2688 5578 2740 5584
rect 2596 5296 2648 5302
rect 2596 5238 2648 5244
rect 2332 3318 2452 3346
rect 2504 3392 2556 3398
rect 2504 3334 2556 3340
rect 2228 3052 2280 3058
rect 2228 2994 2280 3000
rect 1952 2508 2004 2514
rect 1952 2450 2004 2456
rect 1768 2032 1820 2038
rect 1768 1974 1820 1980
rect 1674 1456 1730 1465
rect 1674 1391 1730 1400
rect 1860 604 1912 610
rect 1860 546 1912 552
rect 1872 480 1900 546
rect 2332 480 2360 3318
rect 2412 3120 2464 3126
rect 2412 3062 2464 3068
rect 2424 2446 2452 3062
rect 2608 2530 2636 5238
rect 2884 5234 2912 7375
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 2780 5092 2832 5098
rect 2780 5034 2832 5040
rect 2792 4865 2820 5034
rect 2778 4856 2834 4865
rect 2688 4820 2740 4826
rect 2778 4791 2834 4800
rect 2688 4762 2740 4768
rect 2700 4078 2728 4762
rect 2884 4690 2912 5170
rect 2976 5030 3004 10934
rect 3056 10464 3108 10470
rect 3054 10432 3056 10441
rect 3108 10432 3110 10441
rect 3054 10367 3110 10376
rect 3056 9444 3108 9450
rect 3160 9432 3188 12310
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 3252 10198 3280 11086
rect 3344 10742 3372 14418
rect 3896 14278 3924 17462
rect 3974 17368 4030 17377
rect 3974 17303 4030 17312
rect 3988 14958 4016 17303
rect 4252 15972 4304 15978
rect 4252 15914 4304 15920
rect 4068 15904 4120 15910
rect 4068 15846 4120 15852
rect 3976 14952 4028 14958
rect 3976 14894 4028 14900
rect 4080 14890 4108 15846
rect 4264 15570 4292 15914
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 4068 14884 4120 14890
rect 4068 14826 4120 14832
rect 4448 14550 4476 17520
rect 4816 14822 4844 17520
rect 5276 15706 5304 17520
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 5632 15496 5684 15502
rect 5632 15438 5684 15444
rect 5448 15428 5500 15434
rect 5448 15370 5500 15376
rect 4988 14952 5040 14958
rect 4988 14894 5040 14900
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 4436 14544 4488 14550
rect 4436 14486 4488 14492
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 3884 14272 3936 14278
rect 3884 14214 3936 14220
rect 4344 14272 4396 14278
rect 4344 14214 4396 14220
rect 3421 14172 3717 14192
rect 3477 14170 3501 14172
rect 3557 14170 3581 14172
rect 3637 14170 3661 14172
rect 3499 14118 3501 14170
rect 3563 14118 3575 14170
rect 3637 14118 3639 14170
rect 3477 14116 3501 14118
rect 3557 14116 3581 14118
rect 3637 14116 3661 14118
rect 3421 14096 3717 14116
rect 4068 14000 4120 14006
rect 4068 13942 4120 13948
rect 3792 13932 3844 13938
rect 3792 13874 3844 13880
rect 3421 13084 3717 13104
rect 3477 13082 3501 13084
rect 3557 13082 3581 13084
rect 3637 13082 3661 13084
rect 3499 13030 3501 13082
rect 3563 13030 3575 13082
rect 3637 13030 3639 13082
rect 3477 13028 3501 13030
rect 3557 13028 3581 13030
rect 3637 13028 3661 13030
rect 3421 13008 3717 13028
rect 3698 12880 3754 12889
rect 3698 12815 3754 12824
rect 3712 12782 3740 12815
rect 3700 12776 3752 12782
rect 3700 12718 3752 12724
rect 3700 12640 3752 12646
rect 3700 12582 3752 12588
rect 3712 12442 3740 12582
rect 3700 12436 3752 12442
rect 3700 12378 3752 12384
rect 3421 11996 3717 12016
rect 3477 11994 3501 11996
rect 3557 11994 3581 11996
rect 3637 11994 3661 11996
rect 3499 11942 3501 11994
rect 3563 11942 3575 11994
rect 3637 11942 3639 11994
rect 3477 11940 3501 11942
rect 3557 11940 3581 11942
rect 3637 11940 3661 11942
rect 3421 11920 3717 11940
rect 3422 11792 3478 11801
rect 3422 11727 3478 11736
rect 3436 11626 3464 11727
rect 3424 11620 3476 11626
rect 3424 11562 3476 11568
rect 3516 11552 3568 11558
rect 3516 11494 3568 11500
rect 3528 11082 3556 11494
rect 3516 11076 3568 11082
rect 3516 11018 3568 11024
rect 3421 10908 3717 10928
rect 3477 10906 3501 10908
rect 3557 10906 3581 10908
rect 3637 10906 3661 10908
rect 3499 10854 3501 10906
rect 3563 10854 3575 10906
rect 3637 10854 3639 10906
rect 3477 10852 3501 10854
rect 3557 10852 3581 10854
rect 3637 10852 3661 10854
rect 3421 10832 3717 10852
rect 3332 10736 3384 10742
rect 3332 10678 3384 10684
rect 3240 10192 3292 10198
rect 3240 10134 3292 10140
rect 3804 10010 3832 13874
rect 3884 13728 3936 13734
rect 3884 13670 3936 13676
rect 3896 12753 3924 13670
rect 3976 13320 4028 13326
rect 3974 13288 3976 13297
rect 4028 13288 4030 13297
rect 3974 13223 4030 13232
rect 3882 12744 3938 12753
rect 3882 12679 3938 12688
rect 3988 12374 4016 13223
rect 4080 12442 4108 13942
rect 4356 13530 4384 14214
rect 4528 13932 4580 13938
rect 4528 13874 4580 13880
rect 4344 13524 4396 13530
rect 4344 13466 4396 13472
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 4436 13184 4488 13190
rect 4436 13126 4488 13132
rect 4172 12850 4200 13126
rect 4160 12844 4212 12850
rect 4160 12786 4212 12792
rect 4448 12782 4476 13126
rect 4436 12776 4488 12782
rect 4436 12718 4488 12724
rect 4252 12708 4304 12714
rect 4252 12650 4304 12656
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 3976 12368 4028 12374
rect 3976 12310 4028 12316
rect 4066 12064 4122 12073
rect 4066 11999 4122 12008
rect 4080 11694 4108 11999
rect 3884 11688 3936 11694
rect 3884 11630 3936 11636
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 3896 10146 3924 11630
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 4080 11354 4108 11494
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 4172 11218 4200 12582
rect 4264 11286 4292 12650
rect 4434 12608 4490 12617
rect 4434 12543 4490 12552
rect 4448 12374 4476 12543
rect 4540 12442 4568 13874
rect 4632 13308 4660 14350
rect 4724 14249 4752 14418
rect 4710 14240 4766 14249
rect 4710 14175 4766 14184
rect 4894 14240 4950 14249
rect 4894 14175 4950 14184
rect 4712 13728 4764 13734
rect 4712 13670 4764 13676
rect 4804 13728 4856 13734
rect 4804 13670 4856 13676
rect 4724 13462 4752 13670
rect 4712 13456 4764 13462
rect 4712 13398 4764 13404
rect 4712 13320 4764 13326
rect 4632 13280 4712 13308
rect 4712 13262 4764 13268
rect 4724 13161 4752 13262
rect 4710 13152 4766 13161
rect 4710 13087 4766 13096
rect 4528 12436 4580 12442
rect 4528 12378 4580 12384
rect 4436 12368 4488 12374
rect 4816 12322 4844 13670
rect 4908 13530 4936 14175
rect 4896 13524 4948 13530
rect 4896 13466 4948 13472
rect 4896 12844 4948 12850
rect 4896 12786 4948 12792
rect 4436 12310 4488 12316
rect 4540 12294 4844 12322
rect 4436 12232 4488 12238
rect 4436 12174 4488 12180
rect 4448 11830 4476 12174
rect 4540 11898 4568 12294
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4528 11892 4580 11898
rect 4528 11834 4580 11840
rect 4436 11824 4488 11830
rect 4436 11766 4488 11772
rect 4252 11280 4304 11286
rect 4252 11222 4304 11228
rect 4448 11218 4476 11766
rect 4724 11558 4752 12174
rect 4816 11762 4844 12174
rect 4804 11756 4856 11762
rect 4804 11698 4856 11704
rect 4908 11694 4936 12786
rect 4896 11688 4948 11694
rect 4896 11630 4948 11636
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 4436 11212 4488 11218
rect 4436 11154 4488 11160
rect 4160 11076 4212 11082
rect 4160 11018 4212 11024
rect 4172 10606 4200 11018
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4160 10600 4212 10606
rect 4160 10542 4212 10548
rect 3896 10118 4108 10146
rect 4172 10130 4200 10542
rect 4632 10470 4660 10746
rect 4804 10736 4856 10742
rect 4908 10724 4936 11630
rect 4856 10696 4936 10724
rect 4804 10678 4856 10684
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 3976 10056 4028 10062
rect 3804 9982 3924 10010
rect 3976 9998 4028 10004
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3421 9820 3717 9840
rect 3477 9818 3501 9820
rect 3557 9818 3581 9820
rect 3637 9818 3661 9820
rect 3499 9766 3501 9818
rect 3563 9766 3575 9818
rect 3637 9766 3639 9818
rect 3477 9764 3501 9766
rect 3557 9764 3581 9766
rect 3637 9764 3661 9766
rect 3421 9744 3717 9764
rect 3804 9450 3832 9862
rect 3896 9625 3924 9982
rect 3882 9616 3938 9625
rect 3882 9551 3938 9560
rect 3108 9404 3188 9432
rect 3792 9444 3844 9450
rect 3056 9386 3108 9392
rect 3792 9386 3844 9392
rect 3421 8732 3717 8752
rect 3477 8730 3501 8732
rect 3557 8730 3581 8732
rect 3637 8730 3661 8732
rect 3499 8678 3501 8730
rect 3563 8678 3575 8730
rect 3637 8678 3639 8730
rect 3477 8676 3501 8678
rect 3557 8676 3581 8678
rect 3637 8676 3661 8678
rect 3421 8656 3717 8676
rect 3698 8392 3754 8401
rect 3332 8356 3384 8362
rect 3698 8327 3754 8336
rect 3332 8298 3384 8304
rect 3344 7886 3372 8298
rect 3712 8090 3740 8327
rect 3896 8294 3924 9551
rect 3988 9178 4016 9998
rect 4080 9178 4108 10118
rect 4160 10124 4212 10130
rect 4160 10066 4212 10072
rect 3976 9172 4028 9178
rect 3976 9114 4028 9120
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 4172 9042 4200 10066
rect 4816 9722 4844 10678
rect 4804 9716 4856 9722
rect 4804 9658 4856 9664
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 4066 8936 4122 8945
rect 4122 8894 4200 8922
rect 4066 8871 4122 8880
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 3700 8084 3752 8090
rect 3700 8026 3752 8032
rect 4172 8022 4200 8894
rect 4160 8016 4212 8022
rect 4160 7958 4212 7964
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3344 7342 3372 7822
rect 3421 7644 3717 7664
rect 3477 7642 3501 7644
rect 3557 7642 3581 7644
rect 3637 7642 3661 7644
rect 3499 7590 3501 7642
rect 3563 7590 3575 7642
rect 3637 7590 3639 7642
rect 3477 7588 3501 7590
rect 3557 7588 3581 7590
rect 3637 7588 3661 7590
rect 3421 7568 3717 7588
rect 3332 7336 3384 7342
rect 3332 7278 3384 7284
rect 3691 7336 3743 7342
rect 3743 7296 3832 7324
rect 3691 7278 3743 7284
rect 3146 7168 3202 7177
rect 3146 7103 3202 7112
rect 3054 6896 3110 6905
rect 3054 6831 3110 6840
rect 3068 6254 3096 6831
rect 3056 6248 3108 6254
rect 3056 6190 3108 6196
rect 3056 6112 3108 6118
rect 3056 6054 3108 6060
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 2872 4684 2924 4690
rect 2872 4626 2924 4632
rect 2962 4584 3018 4593
rect 2962 4519 2964 4528
rect 3016 4519 3018 4528
rect 2964 4490 3016 4496
rect 2962 4448 3018 4457
rect 2962 4383 3018 4392
rect 2688 4072 2740 4078
rect 2688 4014 2740 4020
rect 2780 4004 2832 4010
rect 2780 3946 2832 3952
rect 2608 2502 2728 2530
rect 2412 2440 2464 2446
rect 2412 2382 2464 2388
rect 2700 480 2728 2502
rect 2792 513 2820 3946
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 2884 1494 2912 3538
rect 2976 3534 3004 4383
rect 3068 3738 3096 6054
rect 3160 4622 3188 7103
rect 3344 6322 3372 7278
rect 3421 6556 3717 6576
rect 3477 6554 3501 6556
rect 3557 6554 3581 6556
rect 3637 6554 3661 6556
rect 3499 6502 3501 6554
rect 3563 6502 3575 6554
rect 3637 6502 3639 6554
rect 3477 6500 3501 6502
rect 3557 6500 3581 6502
rect 3637 6500 3661 6502
rect 3421 6480 3717 6500
rect 3332 6316 3384 6322
rect 3804 6304 3832 7296
rect 4068 6792 4120 6798
rect 4066 6760 4068 6769
rect 4120 6760 4122 6769
rect 4066 6695 4122 6704
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 3332 6258 3384 6264
rect 3620 6276 3832 6304
rect 3240 6180 3292 6186
rect 3240 6122 3292 6128
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 3148 4480 3200 4486
rect 3252 4457 3280 6122
rect 3332 5772 3384 5778
rect 3332 5714 3384 5720
rect 3344 5370 3372 5714
rect 3620 5710 3648 6276
rect 3804 6186 3832 6276
rect 3700 6180 3752 6186
rect 3700 6122 3752 6128
rect 3792 6180 3844 6186
rect 3792 6122 3844 6128
rect 3712 6066 3740 6122
rect 3896 6066 3924 6598
rect 3712 6038 3924 6066
rect 3792 5772 3844 5778
rect 3792 5714 3844 5720
rect 3608 5704 3660 5710
rect 3700 5704 3752 5710
rect 3608 5646 3660 5652
rect 3698 5672 3700 5681
rect 3752 5672 3754 5681
rect 3698 5607 3754 5616
rect 3421 5468 3717 5488
rect 3477 5466 3501 5468
rect 3557 5466 3581 5468
rect 3637 5466 3661 5468
rect 3499 5414 3501 5466
rect 3563 5414 3575 5466
rect 3637 5414 3639 5466
rect 3477 5412 3501 5414
rect 3557 5412 3581 5414
rect 3637 5412 3661 5414
rect 3421 5392 3717 5412
rect 3332 5364 3384 5370
rect 3332 5306 3384 5312
rect 3514 5264 3570 5273
rect 3514 5199 3516 5208
rect 3568 5199 3570 5208
rect 3516 5170 3568 5176
rect 3804 5080 3832 5714
rect 3882 5400 3938 5409
rect 3882 5335 3938 5344
rect 3896 5302 3924 5335
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 3712 5052 3832 5080
rect 3332 5024 3384 5030
rect 3384 4984 3648 5012
rect 3332 4966 3384 4972
rect 3620 4622 3648 4984
rect 3712 4690 3740 5052
rect 3884 4752 3936 4758
rect 3884 4694 3936 4700
rect 3700 4684 3752 4690
rect 3700 4626 3752 4632
rect 3608 4616 3660 4622
rect 3608 4558 3660 4564
rect 3792 4480 3844 4486
rect 3148 4422 3200 4428
rect 3238 4448 3294 4457
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 2964 3528 3016 3534
rect 2964 3470 3016 3476
rect 2964 2916 3016 2922
rect 2964 2858 3016 2864
rect 2976 2650 3004 2858
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 2872 1488 2924 1494
rect 2872 1430 2924 1436
rect 2778 504 2834 513
rect 202 0 258 480
rect 570 0 626 480
rect 1030 0 1086 480
rect 1398 0 1454 480
rect 1858 0 1914 480
rect 2318 0 2374 480
rect 2686 0 2742 480
rect 3160 480 3188 4422
rect 3792 4422 3844 4428
rect 3238 4383 3294 4392
rect 3421 4380 3717 4400
rect 3477 4378 3501 4380
rect 3557 4378 3581 4380
rect 3637 4378 3661 4380
rect 3499 4326 3501 4378
rect 3563 4326 3575 4378
rect 3637 4326 3639 4378
rect 3477 4324 3501 4326
rect 3557 4324 3581 4326
rect 3637 4324 3661 4326
rect 3421 4304 3717 4324
rect 3608 4004 3660 4010
rect 3608 3946 3660 3952
rect 3422 3768 3478 3777
rect 3422 3703 3424 3712
rect 3476 3703 3478 3712
rect 3424 3674 3476 3680
rect 3620 3641 3648 3946
rect 3606 3632 3662 3641
rect 3332 3596 3384 3602
rect 3606 3567 3662 3576
rect 3332 3538 3384 3544
rect 3240 3460 3292 3466
rect 3240 3402 3292 3408
rect 3252 3194 3280 3402
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3344 1698 3372 3538
rect 3620 3534 3648 3567
rect 3608 3528 3660 3534
rect 3608 3470 3660 3476
rect 3421 3292 3717 3312
rect 3477 3290 3501 3292
rect 3557 3290 3581 3292
rect 3637 3290 3661 3292
rect 3499 3238 3501 3290
rect 3563 3238 3575 3290
rect 3637 3238 3639 3290
rect 3477 3236 3501 3238
rect 3557 3236 3581 3238
rect 3637 3236 3661 3238
rect 3421 3216 3717 3236
rect 3606 2544 3662 2553
rect 3606 2479 3662 2488
rect 3620 2446 3648 2479
rect 3516 2440 3568 2446
rect 3514 2408 3516 2417
rect 3608 2440 3660 2446
rect 3568 2408 3570 2417
rect 3608 2382 3660 2388
rect 3514 2343 3570 2352
rect 3421 2204 3717 2224
rect 3477 2202 3501 2204
rect 3557 2202 3581 2204
rect 3637 2202 3661 2204
rect 3499 2150 3501 2202
rect 3563 2150 3575 2202
rect 3637 2150 3639 2202
rect 3477 2148 3501 2150
rect 3557 2148 3581 2150
rect 3637 2148 3661 2150
rect 3421 2128 3717 2148
rect 3332 1692 3384 1698
rect 3332 1634 3384 1640
rect 3804 1442 3832 4422
rect 3896 3194 3924 4694
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 3884 2848 3936 2854
rect 3884 2790 3936 2796
rect 3896 2553 3924 2790
rect 3882 2544 3938 2553
rect 3988 2514 4016 6598
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 4080 3602 4108 5714
rect 4172 5574 4200 6394
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4172 5001 4200 5306
rect 4158 4992 4214 5001
rect 4158 4927 4214 4936
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4172 4146 4200 4762
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 4264 3942 4292 9114
rect 5000 9081 5028 14894
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 5080 14340 5132 14346
rect 5080 14282 5132 14288
rect 5092 13938 5120 14282
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 5092 12481 5120 13262
rect 5184 13190 5212 14758
rect 5356 14272 5408 14278
rect 5356 14214 5408 14220
rect 5368 14006 5396 14214
rect 5356 14000 5408 14006
rect 5356 13942 5408 13948
rect 5264 13932 5316 13938
rect 5264 13874 5316 13880
rect 5172 13184 5224 13190
rect 5172 13126 5224 13132
rect 5078 12472 5134 12481
rect 5078 12407 5134 12416
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 5092 11694 5120 12242
rect 5276 11880 5304 13874
rect 5356 13864 5408 13870
rect 5356 13806 5408 13812
rect 5368 13530 5396 13806
rect 5356 13524 5408 13530
rect 5356 13466 5408 13472
rect 5460 12646 5488 15370
rect 5540 15088 5592 15094
rect 5540 15030 5592 15036
rect 5552 14657 5580 15030
rect 5538 14648 5594 14657
rect 5538 14583 5594 14592
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5552 14278 5580 14350
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5552 13394 5580 13670
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5540 13252 5592 13258
rect 5540 13194 5592 13200
rect 5448 12640 5500 12646
rect 5448 12582 5500 12588
rect 5276 11852 5396 11880
rect 5080 11688 5132 11694
rect 5080 11630 5132 11636
rect 5368 11626 5396 11852
rect 5356 11620 5408 11626
rect 5356 11562 5408 11568
rect 5368 11354 5396 11562
rect 5356 11348 5408 11354
rect 5356 11290 5408 11296
rect 5080 10600 5132 10606
rect 5080 10542 5132 10548
rect 5092 10044 5120 10542
rect 5172 10056 5224 10062
rect 5092 10016 5172 10044
rect 5092 9586 5120 10016
rect 5172 9998 5224 10004
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 4986 9072 5042 9081
rect 5092 9042 5120 9522
rect 4986 9007 5042 9016
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5080 8560 5132 8566
rect 5078 8528 5080 8537
rect 5132 8528 5134 8537
rect 5078 8463 5134 8472
rect 4620 8424 4672 8430
rect 4620 8366 4672 8372
rect 4632 7886 4660 8366
rect 4804 8288 4856 8294
rect 4804 8230 4856 8236
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4434 7712 4490 7721
rect 4434 7647 4490 7656
rect 4448 6254 4476 7647
rect 4632 7410 4660 7822
rect 4710 7576 4766 7585
rect 4710 7511 4766 7520
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 4724 7274 4752 7511
rect 4816 7478 4844 8230
rect 4896 8084 4948 8090
rect 4896 8026 4948 8032
rect 4804 7472 4856 7478
rect 4804 7414 4856 7420
rect 4712 7268 4764 7274
rect 4712 7210 4764 7216
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4632 6497 4660 7142
rect 4816 6866 4844 7414
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4618 6488 4674 6497
rect 4618 6423 4674 6432
rect 4528 6384 4580 6390
rect 4528 6326 4580 6332
rect 4618 6352 4674 6361
rect 4436 6248 4488 6254
rect 4436 6190 4488 6196
rect 4344 5636 4396 5642
rect 4344 5578 4396 5584
rect 4356 5098 4384 5578
rect 4434 5536 4490 5545
rect 4434 5471 4490 5480
rect 4448 5302 4476 5471
rect 4436 5296 4488 5302
rect 4436 5238 4488 5244
rect 4344 5092 4396 5098
rect 4344 5034 4396 5040
rect 4436 5024 4488 5030
rect 4436 4966 4488 4972
rect 4342 4312 4398 4321
rect 4342 4247 4398 4256
rect 4356 4214 4384 4247
rect 4344 4208 4396 4214
rect 4344 4150 4396 4156
rect 4342 4040 4398 4049
rect 4342 3975 4398 3984
rect 4160 3936 4212 3942
rect 4160 3878 4212 3884
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 4172 3466 4200 3878
rect 4264 3602 4292 3878
rect 4252 3596 4304 3602
rect 4252 3538 4304 3544
rect 4160 3460 4212 3466
rect 4160 3402 4212 3408
rect 4252 3392 4304 3398
rect 4356 3380 4384 3975
rect 4304 3352 4384 3380
rect 4448 3369 4476 4966
rect 4434 3360 4490 3369
rect 4252 3334 4304 3340
rect 4264 3058 4292 3334
rect 4434 3295 4490 3304
rect 4540 3058 4568 6326
rect 4618 6287 4674 6296
rect 4632 3670 4660 6287
rect 4712 6248 4764 6254
rect 4712 6190 4764 6196
rect 4724 5710 4752 6190
rect 4802 5808 4858 5817
rect 4802 5743 4858 5752
rect 4712 5704 4764 5710
rect 4710 5672 4712 5681
rect 4764 5672 4766 5681
rect 4710 5607 4766 5616
rect 4724 5581 4752 5607
rect 4712 4548 4764 4554
rect 4712 4490 4764 4496
rect 4724 4282 4752 4490
rect 4712 4276 4764 4282
rect 4712 4218 4764 4224
rect 4710 3904 4766 3913
rect 4710 3839 4766 3848
rect 4620 3664 4672 3670
rect 4620 3606 4672 3612
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 4528 3052 4580 3058
rect 4724 3040 4752 3839
rect 4816 3738 4844 5743
rect 4908 4298 4936 8026
rect 5078 7984 5134 7993
rect 5078 7919 5134 7928
rect 5172 7948 5224 7954
rect 5092 7324 5120 7919
rect 5172 7890 5224 7896
rect 5000 7296 5120 7324
rect 5000 4690 5028 7296
rect 5080 7200 5132 7206
rect 5080 7142 5132 7148
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 4986 4312 5042 4321
rect 4908 4270 4986 4298
rect 4986 4247 5042 4256
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4908 3942 4936 4082
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 5000 3534 5028 4247
rect 4988 3528 5040 3534
rect 4988 3470 5040 3476
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 5000 3126 5028 3334
rect 5092 3194 5120 7142
rect 5184 6798 5212 7890
rect 5262 7304 5318 7313
rect 5262 7239 5318 7248
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 5276 5216 5304 7239
rect 5368 6458 5396 8774
rect 5460 8294 5488 12582
rect 5552 10266 5580 13194
rect 5644 11694 5672 15438
rect 5736 14958 5764 17520
rect 6104 15994 6132 17520
rect 6104 15966 6316 15994
rect 5886 15804 6182 15824
rect 5942 15802 5966 15804
rect 6022 15802 6046 15804
rect 6102 15802 6126 15804
rect 5964 15750 5966 15802
rect 6028 15750 6040 15802
rect 6102 15750 6104 15802
rect 5942 15748 5966 15750
rect 6022 15748 6046 15750
rect 6102 15748 6126 15750
rect 5886 15728 6182 15748
rect 6182 15600 6238 15609
rect 5816 15564 5868 15570
rect 6182 15535 6184 15544
rect 5816 15506 5868 15512
rect 6236 15535 6238 15544
rect 6184 15506 6236 15512
rect 5724 14952 5776 14958
rect 5724 14894 5776 14900
rect 5828 14822 5856 15506
rect 6288 15094 6316 15966
rect 6564 15162 6592 17520
rect 7024 16046 7052 17520
rect 7012 16040 7064 16046
rect 7012 15982 7064 15988
rect 6644 15904 6696 15910
rect 6644 15846 6696 15852
rect 6656 15502 6684 15846
rect 6644 15496 6696 15502
rect 6644 15438 6696 15444
rect 7010 15464 7066 15473
rect 7010 15399 7066 15408
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6276 15088 6328 15094
rect 6090 15056 6146 15065
rect 6276 15030 6328 15036
rect 6090 14991 6092 15000
rect 6144 14991 6146 15000
rect 6368 15020 6420 15026
rect 6092 14962 6144 14968
rect 6368 14962 6420 14968
rect 6276 14952 6328 14958
rect 6276 14894 6328 14900
rect 5816 14816 5868 14822
rect 5816 14758 5868 14764
rect 5886 14716 6182 14736
rect 5942 14714 5966 14716
rect 6022 14714 6046 14716
rect 6102 14714 6126 14716
rect 5964 14662 5966 14714
rect 6028 14662 6040 14714
rect 6102 14662 6104 14714
rect 5942 14660 5966 14662
rect 6022 14660 6046 14662
rect 6102 14660 6126 14662
rect 5886 14640 6182 14660
rect 5724 14612 5776 14618
rect 5724 14554 5776 14560
rect 5736 14385 5764 14554
rect 6288 14385 6316 14894
rect 5722 14376 5778 14385
rect 5722 14311 5778 14320
rect 6274 14376 6330 14385
rect 6274 14311 6330 14320
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5724 13796 5776 13802
rect 5724 13738 5776 13744
rect 5736 13433 5764 13738
rect 5722 13424 5778 13433
rect 5722 13359 5778 13368
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 5632 11688 5684 11694
rect 5632 11630 5684 11636
rect 5644 10606 5672 11630
rect 5736 10985 5764 12718
rect 5828 11801 5856 14214
rect 6276 13932 6328 13938
rect 6276 13874 6328 13880
rect 5886 13628 6182 13648
rect 5942 13626 5966 13628
rect 6022 13626 6046 13628
rect 6102 13626 6126 13628
rect 5964 13574 5966 13626
rect 6028 13574 6040 13626
rect 6102 13574 6104 13626
rect 5942 13572 5966 13574
rect 6022 13572 6046 13574
rect 6102 13572 6126 13574
rect 5886 13552 6182 13572
rect 6000 12980 6052 12986
rect 6000 12922 6052 12928
rect 6012 12714 6040 12922
rect 6182 12880 6238 12889
rect 6182 12815 6238 12824
rect 6196 12782 6224 12815
rect 6184 12776 6236 12782
rect 6184 12718 6236 12724
rect 6000 12708 6052 12714
rect 6000 12650 6052 12656
rect 5886 12540 6182 12560
rect 5942 12538 5966 12540
rect 6022 12538 6046 12540
rect 6102 12538 6126 12540
rect 5964 12486 5966 12538
rect 6028 12486 6040 12538
rect 6102 12486 6104 12538
rect 5942 12484 5966 12486
rect 6022 12484 6046 12486
rect 6102 12484 6126 12486
rect 5886 12464 6182 12484
rect 5906 11928 5962 11937
rect 5906 11863 5962 11872
rect 5814 11792 5870 11801
rect 5814 11727 5870 11736
rect 5920 11540 5948 11863
rect 5828 11512 5948 11540
rect 5722 10976 5778 10985
rect 5722 10911 5778 10920
rect 5632 10600 5684 10606
rect 5632 10542 5684 10548
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5828 9738 5856 11512
rect 5886 11452 6182 11472
rect 5942 11450 5966 11452
rect 6022 11450 6046 11452
rect 6102 11450 6126 11452
rect 5964 11398 5966 11450
rect 6028 11398 6040 11450
rect 6102 11398 6104 11450
rect 5942 11396 5966 11398
rect 6022 11396 6046 11398
rect 6102 11396 6126 11398
rect 5886 11376 6182 11396
rect 5886 10364 6182 10384
rect 5942 10362 5966 10364
rect 6022 10362 6046 10364
rect 6102 10362 6126 10364
rect 5964 10310 5966 10362
rect 6028 10310 6040 10362
rect 6102 10310 6104 10362
rect 5942 10308 5966 10310
rect 6022 10308 6046 10310
rect 6102 10308 6126 10310
rect 5886 10288 6182 10308
rect 6288 10198 6316 13874
rect 6380 13569 6408 14962
rect 6460 14952 6512 14958
rect 6460 14894 6512 14900
rect 6366 13560 6422 13569
rect 6366 13495 6422 13504
rect 6380 13297 6408 13495
rect 6366 13288 6422 13297
rect 6366 13223 6422 13232
rect 6368 12844 6420 12850
rect 6368 12786 6420 12792
rect 6380 12374 6408 12786
rect 6368 12368 6420 12374
rect 6368 12310 6420 12316
rect 6368 12096 6420 12102
rect 6368 12038 6420 12044
rect 6380 11354 6408 12038
rect 6368 11348 6420 11354
rect 6368 11290 6420 11296
rect 6276 10192 6328 10198
rect 6276 10134 6328 10140
rect 5644 9710 6132 9738
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5540 8016 5592 8022
rect 5540 7958 5592 7964
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5184 5188 5304 5216
rect 5184 4128 5212 5188
rect 5264 5092 5316 5098
rect 5264 5034 5316 5040
rect 5276 4486 5304 5034
rect 5368 5001 5396 6394
rect 5354 4992 5410 5001
rect 5354 4927 5410 4936
rect 5368 4622 5396 4927
rect 5460 4826 5488 6394
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5448 4548 5500 4554
rect 5448 4490 5500 4496
rect 5264 4480 5316 4486
rect 5264 4422 5316 4428
rect 5460 4282 5488 4490
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 5184 4100 5304 4128
rect 5170 4040 5226 4049
rect 5170 3975 5226 3984
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 4988 3120 5040 3126
rect 4988 3062 5040 3068
rect 5184 3058 5212 3975
rect 5172 3052 5224 3058
rect 4724 3012 4936 3040
rect 4528 2994 4580 3000
rect 4066 2952 4122 2961
rect 4066 2887 4122 2896
rect 4802 2952 4858 2961
rect 4802 2887 4858 2896
rect 4080 2854 4108 2887
rect 4068 2848 4120 2854
rect 4068 2790 4120 2796
rect 4068 2644 4120 2650
rect 4068 2586 4120 2592
rect 3882 2479 3938 2488
rect 3976 2508 4028 2514
rect 3976 2450 4028 2456
rect 4080 2106 4108 2586
rect 4068 2100 4120 2106
rect 4068 2042 4120 2048
rect 4436 1896 4488 1902
rect 4436 1838 4488 1844
rect 3620 1414 3832 1442
rect 3976 1420 4028 1426
rect 3620 480 3648 1414
rect 3976 1362 4028 1368
rect 3988 480 4016 1362
rect 4448 480 4476 1838
rect 4816 480 4844 2887
rect 4908 2582 4936 3012
rect 5172 2994 5224 3000
rect 5170 2680 5226 2689
rect 5170 2615 5172 2624
rect 5224 2615 5226 2624
rect 5172 2586 5224 2592
rect 4896 2576 4948 2582
rect 4896 2518 4948 2524
rect 5276 480 5304 4100
rect 5368 3534 5396 4218
rect 5460 3913 5488 4218
rect 5446 3904 5502 3913
rect 5446 3839 5502 3848
rect 5446 3768 5502 3777
rect 5446 3703 5448 3712
rect 5500 3703 5502 3712
rect 5448 3674 5500 3680
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 5368 2310 5396 3334
rect 5552 3194 5580 7958
rect 5644 7041 5672 9710
rect 6104 9489 6132 9710
rect 6472 9586 6500 14894
rect 6552 14544 6604 14550
rect 6552 14486 6604 14492
rect 6564 13297 6592 14486
rect 6550 13288 6606 13297
rect 6550 13223 6606 13232
rect 6552 13184 6604 13190
rect 6552 13126 6604 13132
rect 6564 12850 6592 13126
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6550 12472 6606 12481
rect 6656 12458 6684 15302
rect 6920 15088 6972 15094
rect 6920 15030 6972 15036
rect 6736 14816 6788 14822
rect 6736 14758 6788 14764
rect 6748 12617 6776 14758
rect 6828 14340 6880 14346
rect 6828 14282 6880 14288
rect 6840 14074 6868 14282
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6932 13462 6960 15030
rect 7024 14657 7052 15399
rect 7104 15360 7156 15366
rect 7104 15302 7156 15308
rect 7196 15360 7248 15366
rect 7196 15302 7248 15308
rect 7010 14648 7066 14657
rect 7116 14618 7144 15302
rect 7010 14583 7066 14592
rect 7104 14612 7156 14618
rect 7024 14482 7052 14583
rect 7104 14554 7156 14560
rect 7012 14476 7064 14482
rect 7012 14418 7064 14424
rect 7104 14340 7156 14346
rect 7104 14282 7156 14288
rect 7010 14104 7066 14113
rect 7010 14039 7012 14048
rect 7064 14039 7066 14048
rect 7012 14010 7064 14016
rect 7116 13705 7144 14282
rect 7208 13802 7236 15302
rect 7392 15178 7420 17520
rect 7472 16176 7524 16182
rect 7472 16118 7524 16124
rect 7484 15570 7512 16118
rect 7472 15564 7524 15570
rect 7472 15506 7524 15512
rect 7484 15337 7512 15506
rect 7470 15328 7526 15337
rect 7470 15263 7526 15272
rect 7392 15150 7696 15178
rect 7288 15020 7340 15026
rect 7288 14962 7340 14968
rect 7196 13796 7248 13802
rect 7196 13738 7248 13744
rect 7300 13734 7328 14962
rect 7668 14958 7696 15150
rect 7380 14952 7432 14958
rect 7380 14894 7432 14900
rect 7656 14952 7708 14958
rect 7656 14894 7708 14900
rect 7392 13977 7420 14894
rect 7656 14816 7708 14822
rect 7656 14758 7708 14764
rect 7564 14612 7616 14618
rect 7564 14554 7616 14560
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 7378 13968 7434 13977
rect 7378 13903 7434 13912
rect 7288 13728 7340 13734
rect 7102 13696 7158 13705
rect 7288 13670 7340 13676
rect 7102 13631 7158 13640
rect 6920 13456 6972 13462
rect 6920 13398 6972 13404
rect 6828 12980 6880 12986
rect 6932 12968 6960 13398
rect 6880 12940 6960 12968
rect 6828 12922 6880 12928
rect 6828 12640 6880 12646
rect 6734 12608 6790 12617
rect 6828 12582 6880 12588
rect 6734 12543 6790 12552
rect 6840 12481 6868 12582
rect 6826 12472 6882 12481
rect 6656 12430 6776 12458
rect 6550 12407 6606 12416
rect 6564 12374 6592 12407
rect 6552 12368 6604 12374
rect 6552 12310 6604 12316
rect 6564 10742 6592 12310
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 6552 10736 6604 10742
rect 6552 10678 6604 10684
rect 6550 10296 6606 10305
rect 6656 10266 6684 11494
rect 6550 10231 6606 10240
rect 6644 10260 6696 10266
rect 6564 9926 6592 10231
rect 6644 10202 6696 10208
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 6460 9580 6512 9586
rect 6460 9522 6512 9528
rect 6090 9480 6146 9489
rect 5724 9444 5776 9450
rect 6090 9415 6146 9424
rect 5724 9386 5776 9392
rect 5736 7721 5764 9386
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 5886 9276 6182 9296
rect 5942 9274 5966 9276
rect 6022 9274 6046 9276
rect 6102 9274 6126 9276
rect 5964 9222 5966 9274
rect 6028 9222 6040 9274
rect 6102 9222 6104 9274
rect 5942 9220 5966 9222
rect 6022 9220 6046 9222
rect 6102 9220 6126 9222
rect 5886 9200 6182 9220
rect 6564 9110 6592 9318
rect 6552 9104 6604 9110
rect 6552 9046 6604 9052
rect 5886 8188 6182 8208
rect 5942 8186 5966 8188
rect 6022 8186 6046 8188
rect 6102 8186 6126 8188
rect 5964 8134 5966 8186
rect 6028 8134 6040 8186
rect 6102 8134 6104 8186
rect 5942 8132 5966 8134
rect 6022 8132 6046 8134
rect 6102 8132 6126 8134
rect 5886 8112 6182 8132
rect 5722 7712 5778 7721
rect 5722 7647 5778 7656
rect 6366 7576 6422 7585
rect 5816 7540 5868 7546
rect 6366 7511 6422 7520
rect 5816 7482 5868 7488
rect 5724 7200 5776 7206
rect 5722 7168 5724 7177
rect 5776 7168 5778 7177
rect 5722 7103 5778 7112
rect 5630 7032 5686 7041
rect 5630 6967 5686 6976
rect 5632 6928 5684 6934
rect 5632 6870 5684 6876
rect 5644 4826 5672 6870
rect 5828 6866 5856 7482
rect 6092 7404 6144 7410
rect 6092 7346 6144 7352
rect 6104 7274 6132 7346
rect 6380 7274 6408 7511
rect 6092 7268 6144 7274
rect 6092 7210 6144 7216
rect 6368 7268 6420 7274
rect 6368 7210 6420 7216
rect 5886 7100 6182 7120
rect 5942 7098 5966 7100
rect 6022 7098 6046 7100
rect 6102 7098 6126 7100
rect 5964 7046 5966 7098
rect 6028 7046 6040 7098
rect 6102 7046 6104 7098
rect 5942 7044 5966 7046
rect 6022 7044 6046 7046
rect 6102 7044 6126 7046
rect 5886 7024 6182 7044
rect 6366 7032 6422 7041
rect 6366 6967 6422 6976
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 5724 6248 5776 6254
rect 5724 6190 5776 6196
rect 5736 5953 5764 6190
rect 5722 5944 5778 5953
rect 5722 5879 5778 5888
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5736 4706 5764 5510
rect 5644 4678 5764 4706
rect 5644 3670 5672 4678
rect 5828 4622 5856 6802
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 6288 6186 6316 6258
rect 6276 6180 6328 6186
rect 6276 6122 6328 6128
rect 6380 6066 6408 6967
rect 6288 6038 6408 6066
rect 5886 6012 6182 6032
rect 5942 6010 5966 6012
rect 6022 6010 6046 6012
rect 6102 6010 6126 6012
rect 5964 5958 5966 6010
rect 6028 5958 6040 6010
rect 6102 5958 6104 6010
rect 5942 5956 5966 5958
rect 6022 5956 6046 5958
rect 6102 5956 6126 5958
rect 5886 5936 6182 5956
rect 5906 5672 5962 5681
rect 5906 5607 5962 5616
rect 5920 5166 5948 5607
rect 6288 5545 6316 6038
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 6368 5568 6420 5574
rect 6274 5536 6330 5545
rect 6368 5510 6420 5516
rect 6274 5471 6330 5480
rect 6380 5166 6408 5510
rect 6472 5302 6500 5714
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 5886 4924 6182 4944
rect 5942 4922 5966 4924
rect 6022 4922 6046 4924
rect 6102 4922 6126 4924
rect 5964 4870 5966 4922
rect 6028 4870 6040 4922
rect 6102 4870 6104 4922
rect 5942 4868 5966 4870
rect 6022 4868 6046 4870
rect 6102 4868 6126 4870
rect 5886 4848 6182 4868
rect 5908 4752 5960 4758
rect 5908 4694 5960 4700
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 5816 4616 5868 4622
rect 5816 4558 5868 4564
rect 5736 4282 5764 4558
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 5920 4214 5948 4694
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 5908 4208 5960 4214
rect 5908 4150 5960 4156
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 5724 4004 5776 4010
rect 5724 3946 5776 3952
rect 5632 3664 5684 3670
rect 5632 3606 5684 3612
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5460 3058 5488 3130
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5736 2938 5764 3946
rect 5828 3670 5856 4082
rect 6012 4060 6040 4422
rect 6288 4264 6316 4966
rect 6380 4758 6408 5102
rect 6458 4856 6514 4865
rect 6458 4791 6514 4800
rect 6368 4752 6420 4758
rect 6368 4694 6420 4700
rect 6368 4276 6420 4282
rect 6288 4236 6368 4264
rect 6368 4218 6420 4224
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6012 4032 6316 4060
rect 6288 3942 6316 4032
rect 6276 3936 6328 3942
rect 6380 3913 6408 4082
rect 6276 3878 6328 3884
rect 6366 3904 6422 3913
rect 5886 3836 6182 3856
rect 6366 3839 6422 3848
rect 5942 3834 5966 3836
rect 6022 3834 6046 3836
rect 6102 3834 6126 3836
rect 5964 3782 5966 3834
rect 6028 3782 6040 3834
rect 6102 3782 6104 3834
rect 5942 3780 5966 3782
rect 6022 3780 6046 3782
rect 6102 3780 6126 3782
rect 5886 3760 6182 3780
rect 6274 3768 6330 3777
rect 6274 3703 6276 3712
rect 6328 3703 6330 3712
rect 6276 3674 6328 3680
rect 5816 3664 5868 3670
rect 5816 3606 5868 3612
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 5828 3194 5856 3470
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 6472 3058 6500 4791
rect 6564 3534 6592 9046
rect 6748 8673 6776 12430
rect 6826 12407 6882 12416
rect 6828 12300 6880 12306
rect 6932 12288 6960 12940
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 6880 12260 6960 12288
rect 6828 12242 6880 12248
rect 6840 11762 6868 12242
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6840 11218 6868 11698
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6840 10674 6868 11154
rect 7024 11082 7052 12922
rect 7300 12730 7328 13670
rect 7116 12702 7328 12730
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 7116 10538 7144 12702
rect 7194 12472 7250 12481
rect 7194 12407 7250 12416
rect 7104 10532 7156 10538
rect 7104 10474 7156 10480
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6840 10198 6868 10406
rect 6828 10192 6880 10198
rect 6828 10134 6880 10140
rect 7208 9654 7236 12407
rect 7392 11744 7420 13903
rect 7484 13530 7512 14214
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7576 12730 7604 14554
rect 7668 13870 7696 14758
rect 7748 14476 7800 14482
rect 7748 14418 7800 14424
rect 7656 13864 7708 13870
rect 7656 13806 7708 13812
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 7484 12702 7604 12730
rect 7484 11937 7512 12702
rect 7562 12608 7618 12617
rect 7562 12543 7618 12552
rect 7470 11928 7526 11937
rect 7470 11863 7526 11872
rect 7392 11716 7512 11744
rect 7380 11620 7432 11626
rect 7380 11562 7432 11568
rect 7392 11354 7420 11562
rect 7484 11529 7512 11716
rect 7576 11642 7604 12543
rect 7668 12481 7696 13330
rect 7654 12472 7710 12481
rect 7654 12407 7710 12416
rect 7576 11614 7696 11642
rect 7564 11552 7616 11558
rect 7470 11520 7526 11529
rect 7564 11494 7616 11500
rect 7470 11455 7526 11464
rect 7380 11348 7432 11354
rect 7576 11336 7604 11494
rect 7380 11290 7432 11296
rect 7484 11308 7604 11336
rect 7484 11234 7512 11308
rect 7668 11268 7696 11614
rect 7392 11218 7512 11234
rect 7380 11212 7512 11218
rect 7432 11206 7512 11212
rect 7576 11240 7696 11268
rect 7380 11154 7432 11160
rect 7392 10826 7420 11154
rect 7576 11014 7604 11240
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 7564 11008 7616 11014
rect 7564 10950 7616 10956
rect 7392 10810 7512 10826
rect 7392 10804 7524 10810
rect 7392 10798 7472 10804
rect 7472 10746 7524 10752
rect 7668 10130 7696 11086
rect 7760 10713 7788 14418
rect 7852 13818 7880 17520
rect 8116 16108 8168 16114
rect 8116 16050 8168 16056
rect 7932 14952 7984 14958
rect 7932 14894 7984 14900
rect 8024 14952 8076 14958
rect 8024 14894 8076 14900
rect 7944 13977 7972 14894
rect 7930 13968 7986 13977
rect 7930 13903 7986 13912
rect 7852 13790 7972 13818
rect 7944 13734 7972 13790
rect 7932 13728 7984 13734
rect 7932 13670 7984 13676
rect 7932 13456 7984 13462
rect 7932 13398 7984 13404
rect 7840 13388 7892 13394
rect 7840 13330 7892 13336
rect 7852 13161 7880 13330
rect 7838 13152 7894 13161
rect 7838 13087 7894 13096
rect 7838 12064 7894 12073
rect 7838 11999 7894 12008
rect 7852 10742 7880 11999
rect 7944 11393 7972 13398
rect 7930 11384 7986 11393
rect 7930 11319 7986 11328
rect 7840 10736 7892 10742
rect 7746 10704 7802 10713
rect 7840 10678 7892 10684
rect 7746 10639 7802 10648
rect 7840 10532 7892 10538
rect 7840 10474 7892 10480
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 7852 9926 7880 10474
rect 8036 10169 8064 14894
rect 8128 14249 8156 16050
rect 8220 15706 8248 17520
rect 8680 16114 8708 17520
rect 9140 16182 9168 17520
rect 9128 16176 9180 16182
rect 9128 16118 9180 16124
rect 8668 16108 8720 16114
rect 8668 16050 8720 16056
rect 9404 16040 9456 16046
rect 9404 15982 9456 15988
rect 9416 15706 9444 15982
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 9404 15700 9456 15706
rect 9404 15642 9456 15648
rect 9036 15564 9088 15570
rect 9036 15506 9088 15512
rect 8668 15496 8720 15502
rect 8666 15464 8668 15473
rect 8760 15496 8812 15502
rect 8720 15464 8722 15473
rect 8760 15438 8812 15444
rect 8666 15399 8722 15408
rect 8352 15260 8648 15280
rect 8408 15258 8432 15260
rect 8488 15258 8512 15260
rect 8568 15258 8592 15260
rect 8430 15206 8432 15258
rect 8494 15206 8506 15258
rect 8568 15206 8570 15258
rect 8408 15204 8432 15206
rect 8488 15204 8512 15206
rect 8568 15204 8592 15206
rect 8352 15184 8648 15204
rect 8680 15026 8708 15399
rect 8668 15020 8720 15026
rect 8668 14962 8720 14968
rect 8772 14906 8800 15438
rect 8496 14878 8800 14906
rect 8850 14920 8906 14929
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8114 14240 8170 14249
rect 8114 14175 8170 14184
rect 8128 13954 8156 14175
rect 8220 14074 8248 14758
rect 8496 14618 8524 14878
rect 8850 14855 8906 14864
rect 8944 14884 8996 14890
rect 8668 14816 8720 14822
rect 8668 14758 8720 14764
rect 8484 14612 8536 14618
rect 8484 14554 8536 14560
rect 8576 14544 8628 14550
rect 8576 14486 8628 14492
rect 8588 14346 8616 14486
rect 8576 14340 8628 14346
rect 8576 14282 8628 14288
rect 8352 14172 8648 14192
rect 8408 14170 8432 14172
rect 8488 14170 8512 14172
rect 8568 14170 8592 14172
rect 8430 14118 8432 14170
rect 8494 14118 8506 14170
rect 8568 14118 8570 14170
rect 8408 14116 8432 14118
rect 8488 14116 8512 14118
rect 8568 14116 8592 14118
rect 8352 14096 8648 14116
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 8680 14006 8708 14758
rect 8864 14618 8892 14855
rect 8944 14826 8996 14832
rect 8956 14618 8984 14826
rect 9048 14822 9076 15506
rect 9312 15428 9364 15434
rect 9312 15370 9364 15376
rect 9324 15065 9352 15370
rect 9310 15056 9366 15065
rect 9310 14991 9366 15000
rect 9036 14816 9088 14822
rect 9036 14758 9088 14764
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 8850 14512 8906 14521
rect 8850 14447 8906 14456
rect 8760 14340 8812 14346
rect 8760 14282 8812 14288
rect 8668 14000 8720 14006
rect 8128 13926 8248 13954
rect 8668 13942 8720 13948
rect 8116 13864 8168 13870
rect 8116 13806 8168 13812
rect 8128 12102 8156 13806
rect 8220 13462 8248 13926
rect 8576 13796 8628 13802
rect 8576 13738 8628 13744
rect 8588 13462 8616 13738
rect 8208 13456 8260 13462
rect 8208 13398 8260 13404
rect 8576 13456 8628 13462
rect 8576 13398 8628 13404
rect 8668 13388 8720 13394
rect 8668 13330 8720 13336
rect 8208 13184 8260 13190
rect 8208 13126 8260 13132
rect 8220 12238 8248 13126
rect 8352 13084 8648 13104
rect 8408 13082 8432 13084
rect 8488 13082 8512 13084
rect 8568 13082 8592 13084
rect 8430 13030 8432 13082
rect 8494 13030 8506 13082
rect 8568 13030 8570 13082
rect 8408 13028 8432 13030
rect 8488 13028 8512 13030
rect 8568 13028 8592 13030
rect 8352 13008 8648 13028
rect 8484 12912 8536 12918
rect 8298 12880 8354 12889
rect 8484 12854 8536 12860
rect 8574 12880 8630 12889
rect 8298 12815 8300 12824
rect 8352 12815 8354 12824
rect 8300 12786 8352 12792
rect 8496 12442 8524 12854
rect 8574 12815 8630 12824
rect 8484 12436 8536 12442
rect 8484 12378 8536 12384
rect 8208 12232 8260 12238
rect 8588 12220 8616 12815
rect 8680 12458 8708 13330
rect 8772 13025 8800 14282
rect 8864 13920 8892 14447
rect 8944 13932 8996 13938
rect 8864 13892 8944 13920
rect 8758 13016 8814 13025
rect 8758 12951 8814 12960
rect 8864 12968 8892 13892
rect 8944 13874 8996 13880
rect 8944 13728 8996 13734
rect 8944 13670 8996 13676
rect 8956 13258 8984 13670
rect 8944 13252 8996 13258
rect 8944 13194 8996 13200
rect 8864 12940 8984 12968
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8772 12617 8800 12718
rect 8956 12714 8984 12940
rect 8944 12708 8996 12714
rect 8944 12650 8996 12656
rect 9048 12617 9076 14758
rect 9324 14113 9352 14991
rect 9508 14600 9536 17520
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 9416 14572 9536 14600
rect 9588 14612 9640 14618
rect 9416 14521 9444 14572
rect 9588 14554 9640 14560
rect 9402 14512 9458 14521
rect 9402 14447 9458 14456
rect 9496 14476 9548 14482
rect 9496 14418 9548 14424
rect 9404 14408 9456 14414
rect 9404 14350 9456 14356
rect 9416 14278 9444 14350
rect 9404 14272 9456 14278
rect 9404 14214 9456 14220
rect 9310 14104 9366 14113
rect 9310 14039 9366 14048
rect 9404 13932 9456 13938
rect 9404 13874 9456 13880
rect 9128 13864 9180 13870
rect 9126 13832 9128 13841
rect 9416 13841 9444 13874
rect 9180 13832 9182 13841
rect 9126 13767 9182 13776
rect 9402 13832 9458 13841
rect 9402 13767 9458 13776
rect 9312 13728 9364 13734
rect 9312 13670 9364 13676
rect 9128 13388 9180 13394
rect 9128 13330 9180 13336
rect 9140 13161 9168 13330
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 9126 13152 9182 13161
rect 9126 13087 9182 13096
rect 9232 12850 9260 13262
rect 9220 12844 9272 12850
rect 9220 12786 9272 12792
rect 9128 12708 9180 12714
rect 9128 12650 9180 12656
rect 8758 12608 8814 12617
rect 8758 12543 8814 12552
rect 9034 12608 9090 12617
rect 9034 12543 9090 12552
rect 9034 12472 9090 12481
rect 8680 12430 8892 12458
rect 8760 12300 8812 12306
rect 8760 12242 8812 12248
rect 8668 12232 8720 12238
rect 8588 12192 8668 12220
rect 8208 12174 8260 12180
rect 8668 12174 8720 12180
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8128 11286 8156 12038
rect 8220 11898 8248 12038
rect 8352 11996 8648 12016
rect 8408 11994 8432 11996
rect 8488 11994 8512 11996
rect 8568 11994 8592 11996
rect 8430 11942 8432 11994
rect 8494 11942 8506 11994
rect 8568 11942 8570 11994
rect 8408 11940 8432 11942
rect 8488 11940 8512 11942
rect 8568 11940 8592 11942
rect 8352 11920 8648 11940
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8116 11280 8168 11286
rect 8116 11222 8168 11228
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 8128 10538 8156 10746
rect 8116 10532 8168 10538
rect 8116 10474 8168 10480
rect 8022 10160 8078 10169
rect 8022 10095 8078 10104
rect 7748 9920 7800 9926
rect 7748 9862 7800 9868
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7196 9648 7248 9654
rect 7196 9590 7248 9596
rect 7380 9648 7432 9654
rect 7380 9590 7432 9596
rect 7654 9616 7710 9625
rect 7104 9580 7156 9586
rect 6932 9540 7104 9568
rect 6734 8664 6790 8673
rect 6932 8634 6960 9540
rect 7104 9522 7156 9528
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 6734 8599 6790 8608
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 6734 8392 6790 8401
rect 6734 8327 6790 8336
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6656 6730 6684 7890
rect 6644 6724 6696 6730
rect 6644 6666 6696 6672
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 6276 2984 6328 2990
rect 5632 2916 5684 2922
rect 5736 2910 5856 2938
rect 6276 2926 6328 2932
rect 5632 2858 5684 2864
rect 5446 2680 5502 2689
rect 5446 2615 5448 2624
rect 5500 2615 5502 2624
rect 5448 2586 5500 2592
rect 5644 2530 5672 2858
rect 5724 2848 5776 2854
rect 5724 2790 5776 2796
rect 5552 2502 5672 2530
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 5356 2304 5408 2310
rect 5356 2246 5408 2252
rect 5460 1834 5488 2382
rect 5448 1828 5500 1834
rect 5448 1770 5500 1776
rect 5552 1562 5580 2502
rect 5540 1556 5592 1562
rect 5540 1498 5592 1504
rect 5736 480 5764 2790
rect 5828 2564 5856 2910
rect 5886 2748 6182 2768
rect 5942 2746 5966 2748
rect 6022 2746 6046 2748
rect 6102 2746 6126 2748
rect 5964 2694 5966 2746
rect 6028 2694 6040 2746
rect 6102 2694 6104 2746
rect 5942 2692 5966 2694
rect 6022 2692 6046 2694
rect 6102 2692 6126 2694
rect 5886 2672 6182 2692
rect 6288 2650 6316 2926
rect 6276 2644 6328 2650
rect 6276 2586 6328 2592
rect 5908 2576 5960 2582
rect 5828 2536 5908 2564
rect 5908 2518 5960 2524
rect 6182 2544 6238 2553
rect 6182 2479 6184 2488
rect 6236 2479 6238 2488
rect 6184 2450 6236 2456
rect 6656 2446 6684 6666
rect 6748 4865 6776 8327
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6840 6934 6868 7278
rect 6828 6928 6880 6934
rect 6828 6870 6880 6876
rect 6840 6322 6868 6870
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6840 5574 6868 6258
rect 6932 5778 6960 8026
rect 7024 6934 7052 8230
rect 7012 6928 7064 6934
rect 7012 6870 7064 6876
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 6840 5234 6868 5510
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 6734 4856 6790 4865
rect 6734 4791 6790 4800
rect 6840 4690 6868 5170
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6736 4208 6788 4214
rect 6736 4150 6788 4156
rect 6748 3466 6776 4150
rect 6840 4146 6868 4626
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6840 3738 6868 4082
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6932 3466 6960 5714
rect 7010 5672 7066 5681
rect 7010 5607 7066 5616
rect 7024 5098 7052 5607
rect 7116 5250 7144 8570
rect 7300 8294 7328 9114
rect 7392 8634 7420 9590
rect 7654 9551 7710 9560
rect 7472 9376 7524 9382
rect 7470 9344 7472 9353
rect 7524 9344 7526 9353
rect 7470 9279 7526 9288
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 7196 7948 7248 7954
rect 7196 7890 7248 7896
rect 7208 6866 7236 7890
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7300 7449 7328 7822
rect 7286 7440 7342 7449
rect 7286 7375 7342 7384
rect 7288 7200 7340 7206
rect 7288 7142 7340 7148
rect 7300 6866 7328 7142
rect 7196 6860 7248 6866
rect 7196 6802 7248 6808
rect 7288 6860 7340 6866
rect 7288 6802 7340 6808
rect 7288 6180 7340 6186
rect 7288 6122 7340 6128
rect 7194 5944 7250 5953
rect 7194 5879 7250 5888
rect 7208 5352 7236 5879
rect 7300 5681 7328 6122
rect 7286 5672 7342 5681
rect 7286 5607 7342 5616
rect 7208 5324 7328 5352
rect 7116 5222 7236 5250
rect 7012 5092 7064 5098
rect 7012 5034 7064 5040
rect 7024 5001 7052 5034
rect 7010 4992 7066 5001
rect 7010 4927 7066 4936
rect 7104 4752 7156 4758
rect 7104 4694 7156 4700
rect 7116 4010 7144 4694
rect 7104 4004 7156 4010
rect 7024 3964 7104 3992
rect 7024 3641 7052 3964
rect 7104 3946 7156 3952
rect 7102 3904 7158 3913
rect 7102 3839 7158 3848
rect 7010 3632 7066 3641
rect 7010 3567 7066 3576
rect 6736 3460 6788 3466
rect 6736 3402 6788 3408
rect 6920 3460 6972 3466
rect 6920 3402 6972 3408
rect 6734 3360 6790 3369
rect 6734 3295 6790 3304
rect 6918 3360 6974 3369
rect 6918 3295 6974 3304
rect 6748 2825 6776 3295
rect 6932 2854 6960 3295
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 6920 2848 6972 2854
rect 6734 2816 6790 2825
rect 6920 2790 6972 2796
rect 6734 2751 6790 2760
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 6552 1964 6604 1970
rect 6552 1906 6604 1912
rect 6092 1624 6144 1630
rect 6092 1566 6144 1572
rect 6104 480 6132 1566
rect 6564 480 6592 1906
rect 7024 480 7052 3130
rect 7116 2922 7144 3839
rect 7208 3233 7236 5222
rect 7300 3738 7328 5324
rect 7392 4078 7420 8570
rect 7484 8498 7512 9279
rect 7564 9172 7616 9178
rect 7564 9114 7616 9120
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7576 8430 7604 9114
rect 7668 9042 7696 9551
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7760 8362 7788 9862
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 8128 9625 8156 9658
rect 8220 9654 8248 11154
rect 8352 10908 8648 10928
rect 8408 10906 8432 10908
rect 8488 10906 8512 10908
rect 8568 10906 8592 10908
rect 8430 10854 8432 10906
rect 8494 10854 8506 10906
rect 8568 10854 8570 10906
rect 8408 10852 8432 10854
rect 8488 10852 8512 10854
rect 8568 10852 8592 10854
rect 8352 10832 8648 10852
rect 8484 10736 8536 10742
rect 8484 10678 8536 10684
rect 8496 10441 8524 10678
rect 8482 10432 8538 10441
rect 8482 10367 8538 10376
rect 8352 9820 8648 9840
rect 8408 9818 8432 9820
rect 8488 9818 8512 9820
rect 8568 9818 8592 9820
rect 8430 9766 8432 9818
rect 8494 9766 8506 9818
rect 8568 9766 8570 9818
rect 8408 9764 8432 9766
rect 8488 9764 8512 9766
rect 8568 9764 8592 9766
rect 8352 9744 8648 9764
rect 8208 9648 8260 9654
rect 8114 9616 8170 9625
rect 8208 9590 8260 9596
rect 8114 9551 8170 9560
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8390 9480 8446 9489
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 7748 8356 7800 8362
rect 7748 8298 7800 8304
rect 7656 7948 7708 7954
rect 7656 7890 7708 7896
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7484 7274 7512 7686
rect 7472 7268 7524 7274
rect 7472 7210 7524 7216
rect 7564 7268 7616 7274
rect 7564 7210 7616 7216
rect 7484 5001 7512 7210
rect 7576 5930 7604 7210
rect 7668 6089 7696 7890
rect 7760 6866 7788 8298
rect 7748 6860 7800 6866
rect 7748 6802 7800 6808
rect 7654 6080 7710 6089
rect 7654 6015 7710 6024
rect 7576 5902 7696 5930
rect 7564 5568 7616 5574
rect 7564 5510 7616 5516
rect 7470 4992 7526 5001
rect 7470 4927 7526 4936
rect 7470 4448 7526 4457
rect 7470 4383 7526 4392
rect 7380 4072 7432 4078
rect 7380 4014 7432 4020
rect 7484 4010 7512 4383
rect 7472 4004 7524 4010
rect 7472 3946 7524 3952
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 7576 3584 7604 5510
rect 7668 4457 7696 5902
rect 7852 5574 7880 8910
rect 7944 8838 7972 9454
rect 8114 9208 8170 9217
rect 8220 9178 8248 9454
rect 8114 9143 8170 9152
rect 8208 9172 8260 9178
rect 7932 8832 7984 8838
rect 7932 8774 7984 8780
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 7944 8022 7972 8434
rect 8024 8424 8076 8430
rect 8128 8412 8156 9143
rect 8208 9114 8260 9120
rect 8312 8820 8340 9454
rect 8390 9415 8392 9424
rect 8444 9415 8446 9424
rect 8392 9386 8444 9392
rect 8220 8792 8340 8820
rect 8220 8634 8248 8792
rect 8352 8732 8648 8752
rect 8408 8730 8432 8732
rect 8488 8730 8512 8732
rect 8568 8730 8592 8732
rect 8430 8678 8432 8730
rect 8494 8678 8506 8730
rect 8568 8678 8570 8730
rect 8408 8676 8432 8678
rect 8488 8676 8512 8678
rect 8568 8676 8592 8678
rect 8352 8656 8648 8676
rect 8680 8634 8708 12174
rect 8772 11937 8800 12242
rect 8864 12102 8892 12430
rect 9034 12407 9090 12416
rect 9048 12238 9076 12407
rect 9036 12232 9088 12238
rect 9036 12174 9088 12180
rect 8852 12096 8904 12102
rect 8852 12038 8904 12044
rect 8758 11928 8814 11937
rect 8758 11863 8814 11872
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 8208 8424 8260 8430
rect 8128 8384 8208 8412
rect 8024 8366 8076 8372
rect 8208 8366 8260 8372
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8036 8294 8064 8366
rect 8024 8288 8076 8294
rect 8024 8230 8076 8236
rect 8208 8084 8260 8090
rect 8208 8026 8260 8032
rect 7932 8016 7984 8022
rect 7932 7958 7984 7964
rect 7944 7410 7972 7958
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 8024 7472 8076 7478
rect 8022 7440 8024 7449
rect 8076 7440 8078 7449
rect 7932 7404 7984 7410
rect 8022 7375 8078 7384
rect 7932 7346 7984 7352
rect 7944 6322 7972 7346
rect 8022 6488 8078 6497
rect 8022 6423 8078 6432
rect 7932 6316 7984 6322
rect 7932 6258 7984 6264
rect 7840 5568 7892 5574
rect 7838 5536 7840 5545
rect 7892 5536 7894 5545
rect 7838 5471 7894 5480
rect 7746 5400 7802 5409
rect 7746 5335 7802 5344
rect 7760 4865 7788 5335
rect 7852 5302 7880 5471
rect 7840 5296 7892 5302
rect 7840 5238 7892 5244
rect 7932 5160 7984 5166
rect 7932 5102 7984 5108
rect 8036 5114 8064 6423
rect 8128 5914 8156 7890
rect 8220 6730 8248 8026
rect 8588 8022 8616 8366
rect 8576 8016 8628 8022
rect 8482 7984 8538 7993
rect 8576 7958 8628 7964
rect 8482 7919 8538 7928
rect 8496 7868 8524 7919
rect 8576 7880 8628 7886
rect 8496 7840 8576 7868
rect 8576 7822 8628 7828
rect 8352 7644 8648 7664
rect 8408 7642 8432 7644
rect 8488 7642 8512 7644
rect 8568 7642 8592 7644
rect 8430 7590 8432 7642
rect 8494 7590 8506 7642
rect 8568 7590 8570 7642
rect 8408 7588 8432 7590
rect 8488 7588 8512 7590
rect 8568 7588 8592 7590
rect 8352 7568 8648 7588
rect 8680 7528 8708 8570
rect 8588 7500 8708 7528
rect 8588 7274 8616 7500
rect 8576 7268 8628 7274
rect 8576 7210 8628 7216
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8208 6724 8260 6730
rect 8208 6666 8260 6672
rect 8352 6556 8648 6576
rect 8408 6554 8432 6556
rect 8488 6554 8512 6556
rect 8568 6554 8592 6556
rect 8430 6502 8432 6554
rect 8494 6502 8506 6554
rect 8568 6502 8570 6554
rect 8408 6500 8432 6502
rect 8488 6500 8512 6502
rect 8568 6500 8592 6502
rect 8352 6480 8648 6500
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 8128 5284 8156 5714
rect 8312 5556 8340 6258
rect 8574 5944 8630 5953
rect 8574 5879 8576 5888
rect 8628 5879 8630 5888
rect 8576 5850 8628 5856
rect 8220 5528 8340 5556
rect 8220 5352 8248 5528
rect 8352 5468 8648 5488
rect 8408 5466 8432 5468
rect 8488 5466 8512 5468
rect 8568 5466 8592 5468
rect 8430 5414 8432 5466
rect 8494 5414 8506 5466
rect 8568 5414 8570 5466
rect 8408 5412 8432 5414
rect 8488 5412 8512 5414
rect 8568 5412 8592 5414
rect 8352 5392 8648 5412
rect 8220 5324 8432 5352
rect 8128 5256 8248 5284
rect 7746 4856 7802 4865
rect 7746 4791 7802 4800
rect 7944 4690 7972 5102
rect 8036 5086 8156 5114
rect 8024 5024 8076 5030
rect 8024 4966 8076 4972
rect 7932 4684 7984 4690
rect 7932 4626 7984 4632
rect 7654 4448 7710 4457
rect 7654 4383 7710 4392
rect 7656 4072 7708 4078
rect 7708 4032 7788 4060
rect 7656 4014 7708 4020
rect 7654 3768 7710 3777
rect 7760 3738 7788 4032
rect 7654 3703 7710 3712
rect 7748 3732 7800 3738
rect 7668 3602 7696 3703
rect 7748 3674 7800 3680
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 7300 3556 7604 3584
rect 7656 3596 7708 3602
rect 7194 3224 7250 3233
rect 7194 3159 7250 3168
rect 7104 2916 7156 2922
rect 7104 2858 7156 2864
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7116 1873 7144 2246
rect 7300 2106 7328 3556
rect 7656 3538 7708 3544
rect 7852 3482 7880 3674
rect 7656 3460 7708 3466
rect 7656 3402 7708 3408
rect 7760 3454 7880 3482
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7288 2100 7340 2106
rect 7288 2042 7340 2048
rect 7380 2100 7432 2106
rect 7380 2042 7432 2048
rect 7102 1864 7158 1873
rect 7102 1799 7158 1808
rect 7392 480 7420 2042
rect 7484 1290 7512 3334
rect 7562 3224 7618 3233
rect 7562 3159 7618 3168
rect 7576 3058 7604 3159
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7668 1426 7696 3402
rect 7760 2854 7788 3454
rect 7840 3392 7892 3398
rect 7840 3334 7892 3340
rect 7852 3194 7880 3334
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 7840 2508 7892 2514
rect 7840 2450 7892 2456
rect 7746 2408 7802 2417
rect 7746 2343 7802 2352
rect 7656 1420 7708 1426
rect 7656 1362 7708 1368
rect 7760 1358 7788 2343
rect 7852 2009 7880 2450
rect 7944 2446 7972 4626
rect 8036 4185 8064 4966
rect 8128 4622 8156 5086
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 8116 4480 8168 4486
rect 8116 4422 8168 4428
rect 8128 4214 8156 4422
rect 8116 4208 8168 4214
rect 8022 4176 8078 4185
rect 8116 4150 8168 4156
rect 8022 4111 8078 4120
rect 8036 2514 8064 4111
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 8128 2553 8156 3878
rect 8220 3516 8248 5256
rect 8404 5234 8432 5324
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8576 4752 8628 4758
rect 8576 4694 8628 4700
rect 8588 4554 8616 4694
rect 8576 4548 8628 4554
rect 8576 4490 8628 4496
rect 8352 4380 8648 4400
rect 8408 4378 8432 4380
rect 8488 4378 8512 4380
rect 8568 4378 8592 4380
rect 8430 4326 8432 4378
rect 8494 4326 8506 4378
rect 8568 4326 8570 4378
rect 8408 4324 8432 4326
rect 8488 4324 8512 4326
rect 8568 4324 8592 4326
rect 8352 4304 8648 4324
rect 8300 3528 8352 3534
rect 8220 3488 8300 3516
rect 8300 3470 8352 3476
rect 8352 3292 8648 3312
rect 8408 3290 8432 3292
rect 8488 3290 8512 3292
rect 8568 3290 8592 3292
rect 8430 3238 8432 3290
rect 8494 3238 8506 3290
rect 8568 3238 8570 3290
rect 8408 3236 8432 3238
rect 8488 3236 8512 3238
rect 8568 3236 8592 3238
rect 8352 3216 8648 3236
rect 8680 2990 8708 7142
rect 8772 5658 8800 11863
rect 8850 11520 8906 11529
rect 8850 11455 8906 11464
rect 8864 11286 8892 11455
rect 8852 11280 8904 11286
rect 8852 11222 8904 11228
rect 8852 11144 8904 11150
rect 8850 11112 8852 11121
rect 8904 11112 8906 11121
rect 8850 11047 8906 11056
rect 8852 11008 8904 11014
rect 8850 10976 8852 10985
rect 8904 10976 8906 10985
rect 8850 10911 8906 10920
rect 9048 10674 9076 12174
rect 9140 11354 9168 12650
rect 9218 11928 9274 11937
rect 9218 11863 9274 11872
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 8944 10464 8996 10470
rect 8944 10406 8996 10412
rect 8850 9752 8906 9761
rect 8850 9687 8906 9696
rect 8864 9450 8892 9687
rect 8852 9444 8904 9450
rect 8852 9386 8904 9392
rect 8850 8664 8906 8673
rect 8850 8599 8852 8608
rect 8904 8599 8906 8608
rect 8852 8570 8904 8576
rect 8956 8090 8984 10406
rect 9048 9722 9076 10610
rect 9140 10198 9168 11290
rect 9232 11150 9260 11863
rect 9220 11144 9272 11150
rect 9324 11121 9352 13670
rect 9508 12986 9536 14418
rect 9600 14278 9628 14554
rect 9770 14512 9826 14521
rect 9876 14482 9904 15846
rect 9968 15502 9996 17520
rect 10048 15564 10100 15570
rect 10048 15506 10100 15512
rect 9956 15496 10008 15502
rect 9956 15438 10008 15444
rect 9770 14447 9772 14456
rect 9824 14447 9826 14456
rect 9864 14476 9916 14482
rect 9772 14418 9824 14424
rect 9864 14418 9916 14424
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9588 14272 9640 14278
rect 9588 14214 9640 14220
rect 9586 14104 9642 14113
rect 9586 14039 9642 14048
rect 9600 14006 9628 14039
rect 9588 14000 9640 14006
rect 9588 13942 9640 13948
rect 9588 13864 9640 13870
rect 9588 13806 9640 13812
rect 9496 12980 9548 12986
rect 9496 12922 9548 12928
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 9508 12646 9536 12786
rect 9600 12714 9628 13806
rect 9588 12708 9640 12714
rect 9588 12650 9640 12656
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9586 12608 9642 12617
rect 9402 12472 9458 12481
rect 9402 12407 9404 12416
rect 9456 12407 9458 12416
rect 9404 12378 9456 12384
rect 9402 12200 9458 12209
rect 9402 12135 9458 12144
rect 9220 11086 9272 11092
rect 9310 11112 9366 11121
rect 9128 10192 9180 10198
rect 9128 10134 9180 10140
rect 9232 10062 9260 11086
rect 9310 11047 9366 11056
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9036 9716 9088 9722
rect 9036 9658 9088 9664
rect 9312 9376 9364 9382
rect 9312 9318 9364 9324
rect 9324 9217 9352 9318
rect 9310 9208 9366 9217
rect 9310 9143 9366 9152
rect 9220 9036 9272 9042
rect 9220 8978 9272 8984
rect 9128 8832 9180 8838
rect 9126 8800 9128 8809
rect 9180 8800 9182 8809
rect 9126 8735 9182 8744
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 9034 8256 9090 8265
rect 9034 8191 9090 8200
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8850 7984 8906 7993
rect 8850 7919 8906 7928
rect 8864 7002 8892 7919
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8956 7585 8984 7686
rect 8942 7576 8998 7585
rect 8942 7511 8998 7520
rect 8956 7274 8984 7511
rect 8944 7268 8996 7274
rect 8944 7210 8996 7216
rect 9048 7002 9076 8191
rect 8852 6996 8904 7002
rect 8852 6938 8904 6944
rect 9036 6996 9088 7002
rect 9036 6938 9088 6944
rect 8864 5778 8892 6938
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 8956 5914 8984 6802
rect 9034 6624 9090 6633
rect 9034 6559 9090 6568
rect 9048 6186 9076 6559
rect 9036 6180 9088 6186
rect 9036 6122 9088 6128
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 8772 5630 8984 5658
rect 8760 5568 8812 5574
rect 8760 5510 8812 5516
rect 8772 4146 8800 5510
rect 8852 5092 8904 5098
rect 8852 5034 8904 5040
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 8758 3224 8814 3233
rect 8758 3159 8814 3168
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 8668 2984 8720 2990
rect 8668 2926 8720 2932
rect 8208 2848 8260 2854
rect 8208 2790 8260 2796
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 8220 2689 8248 2790
rect 8206 2680 8262 2689
rect 8206 2615 8262 2624
rect 8312 2564 8340 2790
rect 8404 2650 8432 2926
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 8114 2544 8170 2553
rect 8024 2508 8076 2514
rect 8114 2479 8170 2488
rect 8220 2536 8340 2564
rect 8024 2450 8076 2456
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 8114 2408 8170 2417
rect 8114 2343 8170 2352
rect 8128 2310 8156 2343
rect 8116 2304 8168 2310
rect 8116 2246 8168 2252
rect 8220 2038 8248 2536
rect 8352 2204 8648 2224
rect 8408 2202 8432 2204
rect 8488 2202 8512 2204
rect 8568 2202 8592 2204
rect 8430 2150 8432 2202
rect 8494 2150 8506 2202
rect 8568 2150 8570 2202
rect 8408 2148 8432 2150
rect 8488 2148 8512 2150
rect 8568 2148 8592 2150
rect 8352 2128 8648 2148
rect 8208 2032 8260 2038
rect 7838 2000 7894 2009
rect 8208 1974 8260 1980
rect 7838 1935 7894 1944
rect 8208 1692 8260 1698
rect 8208 1634 8260 1640
rect 7840 1420 7892 1426
rect 7840 1362 7892 1368
rect 7748 1352 7800 1358
rect 7748 1294 7800 1300
rect 7472 1284 7524 1290
rect 7472 1226 7524 1232
rect 7852 480 7880 1362
rect 8220 480 8248 1634
rect 8680 480 8708 2926
rect 8772 2689 8800 3159
rect 8864 2990 8892 5034
rect 8956 4282 8984 5630
rect 8944 4276 8996 4282
rect 8944 4218 8996 4224
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 8956 3670 8984 4082
rect 8944 3664 8996 3670
rect 8944 3606 8996 3612
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 8956 2836 8984 3606
rect 8864 2808 8984 2836
rect 8758 2680 8814 2689
rect 8758 2615 8814 2624
rect 8864 2122 8892 2808
rect 8944 2440 8996 2446
rect 9048 2428 9076 6122
rect 9140 5098 9168 8570
rect 9232 8498 9260 8978
rect 9324 8838 9352 9143
rect 9312 8832 9364 8838
rect 9312 8774 9364 8780
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 9220 8356 9272 8362
rect 9220 8298 9272 8304
rect 9232 7834 9260 8298
rect 9232 7806 9352 7834
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 9232 7546 9260 7686
rect 9220 7540 9272 7546
rect 9220 7482 9272 7488
rect 9324 7426 9352 7806
rect 9232 7398 9352 7426
rect 9232 5710 9260 7398
rect 9310 7032 9366 7041
rect 9310 6967 9366 6976
rect 9324 6934 9352 6967
rect 9312 6928 9364 6934
rect 9312 6870 9364 6876
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9324 5710 9352 5850
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9232 5098 9260 5646
rect 9128 5092 9180 5098
rect 9128 5034 9180 5040
rect 9220 5092 9272 5098
rect 9220 5034 9272 5040
rect 9324 5001 9352 5646
rect 9416 5216 9444 12135
rect 9508 11898 9536 12582
rect 9586 12543 9642 12552
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9496 11620 9548 11626
rect 9496 11562 9548 11568
rect 9508 11014 9536 11562
rect 9496 11008 9548 11014
rect 9496 10950 9548 10956
rect 9508 10674 9536 10950
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9508 10130 9536 10610
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9496 9648 9548 9654
rect 9496 9590 9548 9596
rect 9508 9450 9536 9590
rect 9496 9444 9548 9450
rect 9496 9386 9548 9392
rect 9508 5778 9536 9386
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9600 5681 9628 12543
rect 9692 5794 9720 14350
rect 9772 14340 9824 14346
rect 9772 14282 9824 14288
rect 9784 14249 9812 14282
rect 9770 14240 9826 14249
rect 9770 14175 9826 14184
rect 9772 14000 9824 14006
rect 9772 13942 9824 13948
rect 9784 12073 9812 13942
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9876 13258 9904 13806
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 9864 13252 9916 13258
rect 9864 13194 9916 13200
rect 9862 13152 9918 13161
rect 9862 13087 9918 13096
rect 9876 12481 9904 13087
rect 9862 12472 9918 12481
rect 9862 12407 9918 12416
rect 9770 12064 9826 12073
rect 9770 11999 9826 12008
rect 9772 11620 9824 11626
rect 9772 11562 9824 11568
rect 9784 10538 9812 11562
rect 9772 10532 9824 10538
rect 9772 10474 9824 10480
rect 9784 10266 9812 10474
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 9876 10146 9904 12407
rect 9968 12306 9996 13466
rect 10060 13462 10088 15506
rect 10230 15464 10286 15473
rect 10428 15434 10456 17520
rect 10796 16017 10824 17520
rect 10782 16008 10838 16017
rect 10782 15943 10838 15952
rect 10817 15804 11113 15824
rect 10873 15802 10897 15804
rect 10953 15802 10977 15804
rect 11033 15802 11057 15804
rect 10895 15750 10897 15802
rect 10959 15750 10971 15802
rect 11033 15750 11035 15802
rect 10873 15748 10897 15750
rect 10953 15748 10977 15750
rect 11033 15748 11057 15750
rect 10817 15728 11113 15748
rect 11152 15564 11204 15570
rect 11152 15506 11204 15512
rect 10230 15399 10286 15408
rect 10416 15428 10468 15434
rect 10244 14890 10272 15399
rect 10416 15370 10468 15376
rect 10324 15360 10376 15366
rect 10324 15302 10376 15308
rect 10232 14884 10284 14890
rect 10232 14826 10284 14832
rect 10232 14476 10284 14482
rect 10152 14436 10232 14464
rect 10048 13456 10100 13462
rect 10048 13398 10100 13404
rect 10048 13320 10100 13326
rect 10048 13262 10100 13268
rect 10060 12986 10088 13262
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 9954 12200 10010 12209
rect 9954 12135 10010 12144
rect 9968 11218 9996 12135
rect 10060 12073 10088 12786
rect 10046 12064 10102 12073
rect 10046 11999 10102 12008
rect 9956 11212 10008 11218
rect 9956 11154 10008 11160
rect 9968 10266 9996 11154
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 9784 10118 9904 10146
rect 9784 5896 9812 10118
rect 10152 9110 10180 14436
rect 10232 14418 10284 14424
rect 10230 13152 10286 13161
rect 10230 13087 10286 13096
rect 10244 12918 10272 13087
rect 10232 12912 10284 12918
rect 10232 12854 10284 12860
rect 10336 12646 10364 15302
rect 10508 15020 10560 15026
rect 10508 14962 10560 14968
rect 10520 14414 10548 14962
rect 10600 14952 10652 14958
rect 10784 14952 10836 14958
rect 10600 14894 10652 14900
rect 10704 14912 10784 14940
rect 10612 14793 10640 14894
rect 10598 14784 10654 14793
rect 10598 14719 10654 14728
rect 10704 14600 10732 14912
rect 10784 14894 10836 14900
rect 10817 14716 11113 14736
rect 10873 14714 10897 14716
rect 10953 14714 10977 14716
rect 11033 14714 11057 14716
rect 10895 14662 10897 14714
rect 10959 14662 10971 14714
rect 11033 14662 11035 14714
rect 10873 14660 10897 14662
rect 10953 14660 10977 14662
rect 11033 14660 11057 14662
rect 10817 14640 11113 14660
rect 10704 14572 10824 14600
rect 10600 14544 10652 14550
rect 10600 14486 10652 14492
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 10416 14340 10468 14346
rect 10416 14282 10468 14288
rect 10428 13938 10456 14282
rect 10416 13932 10468 13938
rect 10416 13874 10468 13880
rect 10414 13832 10470 13841
rect 10414 13767 10470 13776
rect 10428 13326 10456 13767
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10324 12640 10376 12646
rect 10324 12582 10376 12588
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 10244 11218 10272 11630
rect 10232 11212 10284 11218
rect 10232 11154 10284 11160
rect 10230 9752 10286 9761
rect 10230 9687 10286 9696
rect 10244 9625 10272 9687
rect 10230 9616 10286 9625
rect 10230 9551 10286 9560
rect 10244 9450 10272 9551
rect 10232 9444 10284 9450
rect 10232 9386 10284 9392
rect 9956 9104 10008 9110
rect 9876 9064 9956 9092
rect 9876 6746 9904 9064
rect 9956 9046 10008 9052
rect 10140 9104 10192 9110
rect 10140 9046 10192 9052
rect 10046 8528 10102 8537
rect 10046 8463 10102 8472
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 9968 7954 9996 8230
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 9968 7449 9996 7890
rect 9954 7440 10010 7449
rect 9954 7375 10010 7384
rect 9954 7032 10010 7041
rect 9954 6967 10010 6976
rect 9968 6866 9996 6967
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 9876 6718 9996 6746
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 9876 6458 9904 6598
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9968 6338 9996 6718
rect 10060 6458 10088 8463
rect 10140 8424 10192 8430
rect 10140 8366 10192 8372
rect 10152 8022 10180 8366
rect 10230 8120 10286 8129
rect 10230 8055 10286 8064
rect 10140 8016 10192 8022
rect 10140 7958 10192 7964
rect 10152 7410 10180 7958
rect 10244 7721 10272 8055
rect 10336 8004 10364 12582
rect 10414 12472 10470 12481
rect 10414 12407 10470 12416
rect 10428 12209 10456 12407
rect 10520 12322 10548 14350
rect 10612 14249 10640 14486
rect 10692 14476 10744 14482
rect 10692 14418 10744 14424
rect 10598 14240 10654 14249
rect 10598 14175 10654 14184
rect 10704 13682 10732 14418
rect 10796 13802 10824 14572
rect 10784 13796 10836 13802
rect 10784 13738 10836 13744
rect 10612 13654 10732 13682
rect 10612 13444 10640 13654
rect 10817 13628 11113 13648
rect 10873 13626 10897 13628
rect 10953 13626 10977 13628
rect 11033 13626 11057 13628
rect 10895 13574 10897 13626
rect 10959 13574 10971 13626
rect 11033 13574 11035 13626
rect 10873 13572 10897 13574
rect 10953 13572 10977 13574
rect 11033 13572 11057 13574
rect 10817 13552 11113 13572
rect 10876 13456 10928 13462
rect 10612 13416 10732 13444
rect 10704 12850 10732 13416
rect 10876 13398 10928 13404
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 10796 12889 10824 13126
rect 10782 12880 10838 12889
rect 10692 12844 10744 12850
rect 10782 12815 10838 12824
rect 10692 12786 10744 12792
rect 10888 12696 10916 13398
rect 10968 13252 11020 13258
rect 10968 13194 11020 13200
rect 11060 13252 11112 13258
rect 11060 13194 11112 13200
rect 10980 12832 11008 13194
rect 11072 12986 11100 13194
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 11060 12844 11112 12850
rect 10980 12804 11060 12832
rect 11060 12786 11112 12792
rect 10968 12708 11020 12714
rect 10888 12668 10968 12696
rect 10968 12650 11020 12656
rect 10817 12540 11113 12560
rect 10873 12538 10897 12540
rect 10953 12538 10977 12540
rect 11033 12538 11057 12540
rect 10895 12486 10897 12538
rect 10959 12486 10971 12538
rect 11033 12486 11035 12538
rect 10873 12484 10897 12486
rect 10953 12484 10977 12486
rect 11033 12484 11057 12486
rect 10817 12464 11113 12484
rect 10520 12306 10640 12322
rect 10520 12300 10652 12306
rect 10520 12294 10600 12300
rect 10600 12242 10652 12248
rect 10692 12300 10744 12306
rect 10692 12242 10744 12248
rect 10508 12232 10560 12238
rect 10414 12200 10470 12209
rect 10508 12174 10560 12180
rect 10414 12135 10470 12144
rect 10520 12073 10548 12174
rect 10506 12064 10562 12073
rect 10506 11999 10562 12008
rect 10520 11898 10548 11999
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 10414 11792 10470 11801
rect 10612 11778 10640 12242
rect 10414 11727 10470 11736
rect 10520 11750 10640 11778
rect 10428 11626 10456 11727
rect 10416 11620 10468 11626
rect 10416 11562 10468 11568
rect 10414 11384 10470 11393
rect 10414 11319 10416 11328
rect 10468 11319 10470 11328
rect 10416 11290 10468 11296
rect 10428 10282 10456 11290
rect 10520 10441 10548 11750
rect 10704 11676 10732 12242
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 11058 12200 11114 12209
rect 10888 11801 10916 12174
rect 10980 12102 11008 12174
rect 11058 12135 11114 12144
rect 11072 12102 11100 12135
rect 10968 12096 11020 12102
rect 10966 12064 10968 12073
rect 11060 12096 11112 12102
rect 11020 12064 11022 12073
rect 11060 12038 11112 12044
rect 10966 11999 11022 12008
rect 10980 11973 11008 11999
rect 11058 11928 11114 11937
rect 11058 11863 11114 11872
rect 10874 11792 10930 11801
rect 10874 11727 10930 11736
rect 10612 11648 10732 11676
rect 10612 11354 10640 11648
rect 11072 11626 11100 11863
rect 11060 11620 11112 11626
rect 11060 11562 11112 11568
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10704 10742 10732 11494
rect 10817 11452 11113 11472
rect 10873 11450 10897 11452
rect 10953 11450 10977 11452
rect 11033 11450 11057 11452
rect 10895 11398 10897 11450
rect 10959 11398 10971 11450
rect 11033 11398 11035 11450
rect 10873 11396 10897 11398
rect 10953 11396 10977 11398
rect 11033 11396 11057 11398
rect 10817 11376 11113 11396
rect 11164 11286 11192 15506
rect 11256 14906 11284 17520
rect 11256 14878 11376 14906
rect 11348 14822 11376 14878
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 11256 12782 11284 14758
rect 11348 13870 11376 14758
rect 11426 13968 11482 13977
rect 11624 13954 11652 17520
rect 11796 15972 11848 15978
rect 11796 15914 11848 15920
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 11426 13903 11482 13912
rect 11532 13926 11652 13954
rect 11336 13864 11388 13870
rect 11336 13806 11388 13812
rect 11334 13696 11390 13705
rect 11334 13631 11390 13640
rect 11348 13530 11376 13631
rect 11336 13524 11388 13530
rect 11336 13466 11388 13472
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 11348 13161 11376 13262
rect 11440 13258 11468 13903
rect 11428 13252 11480 13258
rect 11428 13194 11480 13200
rect 11532 13190 11560 13926
rect 11716 13852 11744 14418
rect 11624 13824 11744 13852
rect 11808 13841 11836 15914
rect 11888 14816 11940 14822
rect 11888 14758 11940 14764
rect 11794 13832 11850 13841
rect 11624 13734 11652 13824
rect 11794 13767 11850 13776
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 11520 13184 11572 13190
rect 11334 13152 11390 13161
rect 11520 13126 11572 13132
rect 11334 13087 11390 13096
rect 11244 12776 11296 12782
rect 11244 12718 11296 12724
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 11256 12306 11284 12582
rect 11348 12481 11376 13087
rect 11518 12880 11574 12889
rect 11518 12815 11574 12824
rect 11428 12708 11480 12714
rect 11428 12650 11480 12656
rect 11440 12617 11468 12650
rect 11426 12608 11482 12617
rect 11426 12543 11482 12552
rect 11334 12472 11390 12481
rect 11334 12407 11390 12416
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11244 12300 11296 12306
rect 11244 12242 11296 12248
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 11348 11880 11376 12174
rect 11256 11852 11376 11880
rect 11152 11280 11204 11286
rect 11152 11222 11204 11228
rect 11256 11014 11284 11852
rect 11336 11756 11388 11762
rect 11336 11698 11388 11704
rect 11348 11218 11376 11698
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11060 11008 11112 11014
rect 11060 10950 11112 10956
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 11072 10810 11100 10950
rect 11150 10840 11206 10849
rect 11060 10804 11112 10810
rect 11150 10775 11206 10784
rect 11060 10746 11112 10752
rect 10692 10736 10744 10742
rect 10692 10678 10744 10684
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10612 10470 10640 10610
rect 10600 10464 10652 10470
rect 10506 10432 10562 10441
rect 10600 10406 10652 10412
rect 10506 10367 10562 10376
rect 10817 10364 11113 10384
rect 10873 10362 10897 10364
rect 10953 10362 10977 10364
rect 11033 10362 11057 10364
rect 10895 10310 10897 10362
rect 10959 10310 10971 10362
rect 11033 10310 11035 10362
rect 10873 10308 10897 10310
rect 10953 10308 10977 10310
rect 11033 10308 11057 10310
rect 10598 10296 10654 10305
rect 10428 10254 10548 10282
rect 10416 10192 10468 10198
rect 10416 10134 10468 10140
rect 10428 8129 10456 10134
rect 10520 9160 10548 10254
rect 10817 10288 11113 10308
rect 10598 10231 10654 10240
rect 10612 9976 10640 10231
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 10692 9988 10744 9994
rect 10612 9948 10692 9976
rect 10692 9930 10744 9936
rect 10966 9752 11022 9761
rect 10966 9687 10968 9696
rect 11020 9687 11022 9696
rect 10968 9658 11020 9664
rect 11072 9489 11100 10066
rect 11058 9480 11114 9489
rect 11058 9415 11114 9424
rect 10817 9276 11113 9296
rect 10873 9274 10897 9276
rect 10953 9274 10977 9276
rect 11033 9274 11057 9276
rect 10895 9222 10897 9274
rect 10959 9222 10971 9274
rect 11033 9222 11035 9274
rect 10873 9220 10897 9222
rect 10953 9220 10977 9222
rect 11033 9220 11057 9222
rect 10817 9200 11113 9220
rect 10520 9132 10916 9160
rect 10782 8936 10838 8945
rect 10782 8871 10838 8880
rect 10692 8560 10744 8566
rect 10690 8528 10692 8537
rect 10744 8528 10746 8537
rect 10690 8463 10746 8472
rect 10796 8430 10824 8871
rect 10888 8537 10916 9132
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 11072 8838 11100 8978
rect 11164 8974 11192 10775
rect 11256 10606 11284 10950
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 11244 10192 11296 10198
rect 11244 10134 11296 10140
rect 11256 9518 11284 10134
rect 11348 10062 11376 11154
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11348 9586 11376 9998
rect 11440 9654 11468 12378
rect 11532 11354 11560 12815
rect 11520 11348 11572 11354
rect 11520 11290 11572 11296
rect 11518 10840 11574 10849
rect 11518 10775 11574 10784
rect 11428 9648 11480 9654
rect 11428 9590 11480 9596
rect 11336 9580 11388 9586
rect 11336 9522 11388 9528
rect 11244 9512 11296 9518
rect 11244 9454 11296 9460
rect 11256 9382 11284 9454
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11242 9208 11298 9217
rect 11348 9178 11376 9522
rect 11426 9480 11482 9489
rect 11426 9415 11482 9424
rect 11242 9143 11244 9152
rect 11296 9143 11298 9152
rect 11336 9172 11388 9178
rect 11244 9114 11296 9120
rect 11336 9114 11388 9120
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 10874 8528 10930 8537
rect 10874 8463 10930 8472
rect 10600 8424 10652 8430
rect 10520 8384 10600 8412
rect 10414 8120 10470 8129
rect 10520 8090 10548 8384
rect 10600 8366 10652 8372
rect 10784 8424 10836 8430
rect 10980 8378 11008 8570
rect 10784 8366 10836 8372
rect 10888 8350 11008 8378
rect 10888 8276 10916 8350
rect 10612 8248 10916 8276
rect 10414 8055 10470 8064
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 10336 7976 10456 8004
rect 10230 7712 10286 7721
rect 10230 7647 10286 7656
rect 10428 7460 10456 7976
rect 10506 7576 10562 7585
rect 10506 7511 10562 7520
rect 10336 7432 10456 7460
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 10152 7002 10180 7346
rect 10336 7206 10364 7432
rect 10324 7200 10376 7206
rect 10324 7142 10376 7148
rect 10414 7168 10470 7177
rect 10230 7032 10286 7041
rect 10140 6996 10192 7002
rect 10230 6967 10286 6976
rect 10140 6938 10192 6944
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 9876 6310 9996 6338
rect 10152 6322 10180 6938
rect 10140 6316 10192 6322
rect 9876 6118 9904 6310
rect 10140 6258 10192 6264
rect 10244 6118 10272 6967
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9956 6112 10008 6118
rect 10232 6112 10284 6118
rect 9956 6054 10008 6060
rect 10060 6072 10232 6100
rect 9784 5868 9904 5896
rect 9692 5766 9812 5794
rect 9586 5672 9642 5681
rect 9586 5607 9642 5616
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9416 5188 9536 5216
rect 9508 5098 9536 5188
rect 9404 5092 9456 5098
rect 9404 5034 9456 5040
rect 9496 5092 9548 5098
rect 9496 5034 9548 5040
rect 9310 4992 9366 5001
rect 9310 4927 9366 4936
rect 9128 4752 9180 4758
rect 9128 4694 9180 4700
rect 9140 4321 9168 4694
rect 9324 4622 9352 4927
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 9220 4548 9272 4554
rect 9220 4490 9272 4496
rect 9126 4312 9182 4321
rect 9126 4247 9182 4256
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9140 3670 9168 3878
rect 9128 3664 9180 3670
rect 9128 3606 9180 3612
rect 9232 3534 9260 4490
rect 9310 4448 9366 4457
rect 9310 4383 9366 4392
rect 9324 3534 9352 4383
rect 9220 3528 9272 3534
rect 9126 3496 9182 3505
rect 9220 3470 9272 3476
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9126 3431 9182 3440
rect 9140 2961 9168 3431
rect 9126 2952 9182 2961
rect 9126 2887 9182 2896
rect 9128 2508 9180 2514
rect 9232 2496 9260 3470
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9324 3058 9352 3334
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 9416 2854 9444 5034
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9496 4276 9548 4282
rect 9496 4218 9548 4224
rect 9508 4185 9536 4218
rect 9494 4176 9550 4185
rect 9600 4146 9628 4966
rect 9692 4826 9720 5510
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 9784 4706 9812 5766
rect 9876 4826 9904 5868
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 9692 4678 9812 4706
rect 9494 4111 9550 4120
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9496 4004 9548 4010
rect 9496 3946 9548 3952
rect 9312 2848 9364 2854
rect 9312 2790 9364 2796
rect 9404 2848 9456 2854
rect 9404 2790 9456 2796
rect 9180 2468 9260 2496
rect 9128 2450 9180 2456
rect 8996 2400 9076 2428
rect 8944 2382 8996 2388
rect 9140 2281 9168 2450
rect 9126 2272 9182 2281
rect 9126 2207 9182 2216
rect 8864 2094 9168 2122
rect 9140 480 9168 2094
rect 9324 1154 9352 2790
rect 9416 1834 9444 2790
rect 9508 1986 9536 3946
rect 9692 3738 9720 4678
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9784 4282 9812 4558
rect 9876 4321 9904 4762
rect 9968 4690 9996 6054
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 9862 4312 9918 4321
rect 9772 4276 9824 4282
rect 9862 4247 9918 4256
rect 9772 4218 9824 4224
rect 9770 4176 9826 4185
rect 9770 4111 9826 4120
rect 9784 4078 9812 4111
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9784 3516 9812 3878
rect 9876 3670 9904 3878
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 9864 3664 9916 3670
rect 9864 3606 9916 3612
rect 9968 3516 9996 3674
rect 9784 3488 9996 3516
rect 9588 3460 9640 3466
rect 9640 3420 9720 3448
rect 9588 3402 9640 3408
rect 9692 3380 9720 3420
rect 9692 3352 9904 3380
rect 9678 3224 9734 3233
rect 9678 3159 9734 3168
rect 9692 3058 9720 3159
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9772 2304 9824 2310
rect 9772 2246 9824 2252
rect 9678 2000 9734 2009
rect 9508 1958 9678 1986
rect 9678 1935 9734 1944
rect 9404 1828 9456 1834
rect 9404 1770 9456 1776
rect 9784 1562 9812 2246
rect 9876 1737 9904 3352
rect 9954 3224 10010 3233
rect 9954 3159 10010 3168
rect 9968 3058 9996 3159
rect 9956 3052 10008 3058
rect 9956 2994 10008 3000
rect 10060 2990 10088 6072
rect 10232 6054 10284 6060
rect 10232 5908 10284 5914
rect 10152 5868 10232 5896
rect 10152 4146 10180 5868
rect 10232 5850 10284 5856
rect 10230 5808 10286 5817
rect 10230 5743 10286 5752
rect 10244 5642 10272 5743
rect 10232 5636 10284 5642
rect 10232 5578 10284 5584
rect 10232 5092 10284 5098
rect 10232 5034 10284 5040
rect 10244 4672 10272 5034
rect 10336 4826 10364 7142
rect 10414 7103 10470 7112
rect 10428 5114 10456 7103
rect 10520 5302 10548 7511
rect 10612 5914 10640 8248
rect 11256 8242 11284 9114
rect 11348 9042 11376 9114
rect 11336 9036 11388 9042
rect 11336 8978 11388 8984
rect 11440 8922 11468 9415
rect 11348 8906 11468 8922
rect 11336 8900 11468 8906
rect 11388 8894 11468 8900
rect 11336 8842 11388 8848
rect 11532 8566 11560 10775
rect 11624 8820 11652 13670
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11716 13433 11744 13466
rect 11702 13424 11758 13433
rect 11702 13359 11758 13368
rect 11702 13288 11758 13297
rect 11702 13223 11758 13232
rect 11716 13002 11744 13223
rect 11716 12974 11836 13002
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11716 10810 11744 12786
rect 11808 11642 11836 12974
rect 11900 12050 11928 14758
rect 12084 14657 12112 17520
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 12070 14648 12126 14657
rect 12070 14583 12126 14592
rect 11978 14512 12034 14521
rect 11978 14447 12034 14456
rect 11992 13433 12020 14447
rect 12176 13530 12204 15098
rect 12346 14376 12402 14385
rect 12346 14311 12402 14320
rect 12256 14272 12308 14278
rect 12256 14214 12308 14220
rect 12164 13524 12216 13530
rect 12164 13466 12216 13472
rect 11978 13424 12034 13433
rect 11978 13359 12034 13368
rect 12164 13320 12216 13326
rect 12162 13288 12164 13297
rect 12216 13288 12218 13297
rect 12162 13223 12218 13232
rect 12176 12986 12204 13223
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 11992 12442 12020 12718
rect 12084 12442 12112 12854
rect 12164 12844 12216 12850
rect 12164 12786 12216 12792
rect 12176 12646 12204 12786
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 12072 12436 12124 12442
rect 12072 12378 12124 12384
rect 11900 12022 12204 12050
rect 12070 11928 12126 11937
rect 12070 11863 12126 11872
rect 11980 11824 12032 11830
rect 11980 11766 12032 11772
rect 11808 11614 11928 11642
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11808 10606 11836 11494
rect 11900 11354 11928 11614
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 11888 11144 11940 11150
rect 11992 11132 12020 11766
rect 11940 11104 12020 11132
rect 11888 11086 11940 11092
rect 11900 10674 11928 11086
rect 11980 10736 12032 10742
rect 11978 10704 11980 10713
rect 12032 10704 12034 10713
rect 11888 10668 11940 10674
rect 11978 10639 12034 10648
rect 11888 10610 11940 10616
rect 11796 10600 11848 10606
rect 11796 10542 11848 10548
rect 11704 10464 11756 10470
rect 11702 10432 11704 10441
rect 11756 10432 11758 10441
rect 11702 10367 11758 10376
rect 11900 10130 11928 10610
rect 11888 10124 11940 10130
rect 11888 10066 11940 10072
rect 12084 9976 12112 11863
rect 12176 11642 12204 12022
rect 12268 11762 12296 14214
rect 12360 14074 12388 14311
rect 12348 14068 12400 14074
rect 12348 14010 12400 14016
rect 12440 14000 12492 14006
rect 12440 13942 12492 13948
rect 12348 13932 12400 13938
rect 12348 13874 12400 13880
rect 12360 13705 12388 13874
rect 12452 13841 12480 13942
rect 12438 13832 12494 13841
rect 12438 13767 12494 13776
rect 12440 13728 12492 13734
rect 12346 13696 12402 13705
rect 12440 13670 12492 13676
rect 12346 13631 12402 13640
rect 12360 13433 12388 13631
rect 12346 13424 12402 13433
rect 12452 13410 12480 13670
rect 12544 13512 12572 17520
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 12714 14240 12770 14249
rect 12714 14175 12770 14184
rect 12728 13870 12756 14175
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 12544 13484 12664 13512
rect 12452 13382 12572 13410
rect 12346 13359 12402 13368
rect 12348 13252 12400 13258
rect 12348 13194 12400 13200
rect 12360 12322 12388 13194
rect 12440 12912 12492 12918
rect 12440 12854 12492 12860
rect 12452 12753 12480 12854
rect 12438 12744 12494 12753
rect 12438 12679 12494 12688
rect 12360 12294 12480 12322
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 12256 11756 12308 11762
rect 12256 11698 12308 11704
rect 12360 11694 12388 12174
rect 12452 11830 12480 12294
rect 12544 12186 12572 13382
rect 12636 12288 12664 13484
rect 12728 12458 12756 13806
rect 12820 12646 12848 14554
rect 12912 13462 12940 17520
rect 13372 15473 13400 17520
rect 13358 15464 13414 15473
rect 13358 15399 13414 15408
rect 13832 15366 13860 17520
rect 13912 15428 13964 15434
rect 13912 15370 13964 15376
rect 13820 15360 13872 15366
rect 13820 15302 13872 15308
rect 13282 15260 13578 15280
rect 13338 15258 13362 15260
rect 13418 15258 13442 15260
rect 13498 15258 13522 15260
rect 13360 15206 13362 15258
rect 13424 15206 13436 15258
rect 13498 15206 13500 15258
rect 13338 15204 13362 15206
rect 13418 15204 13442 15206
rect 13498 15204 13522 15206
rect 13282 15184 13578 15204
rect 12992 14952 13044 14958
rect 12992 14894 13044 14900
rect 12900 13456 12952 13462
rect 12900 13398 12952 13404
rect 12912 12889 12940 13398
rect 12898 12880 12954 12889
rect 12898 12815 12954 12824
rect 12900 12776 12952 12782
rect 12900 12718 12952 12724
rect 12808 12640 12860 12646
rect 12912 12617 12940 12718
rect 12808 12582 12860 12588
rect 12898 12608 12954 12617
rect 12898 12543 12954 12552
rect 12898 12472 12954 12481
rect 12728 12430 12848 12458
rect 12636 12260 12756 12288
rect 12728 12209 12756 12260
rect 12714 12200 12770 12209
rect 12544 12158 12664 12186
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12440 11824 12492 11830
rect 12440 11766 12492 11772
rect 12348 11688 12400 11694
rect 12176 11614 12296 11642
rect 12348 11630 12400 11636
rect 12164 11008 12216 11014
rect 12164 10950 12216 10956
rect 12176 10198 12204 10950
rect 12164 10192 12216 10198
rect 12164 10134 12216 10140
rect 12268 10112 12296 11614
rect 12544 11286 12572 12038
rect 12636 11694 12664 12158
rect 12714 12135 12770 12144
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 12624 11552 12676 11558
rect 12624 11494 12676 11500
rect 12636 11354 12664 11494
rect 12728 11393 12756 12038
rect 12714 11384 12770 11393
rect 12624 11348 12676 11354
rect 12714 11319 12770 11328
rect 12624 11290 12676 11296
rect 12440 11280 12492 11286
rect 12440 11222 12492 11228
rect 12532 11280 12584 11286
rect 12820 11234 12848 12430
rect 12898 12407 12954 12416
rect 12912 12238 12940 12407
rect 12900 12232 12952 12238
rect 12900 12174 12952 12180
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12912 11937 12940 12038
rect 12898 11928 12954 11937
rect 12898 11863 12954 11872
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12532 11222 12584 11228
rect 12452 10248 12480 11222
rect 12636 11206 12848 11234
rect 12636 10470 12664 11206
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12806 10976 12862 10985
rect 12624 10464 12676 10470
rect 12624 10406 12676 10412
rect 12452 10220 12664 10248
rect 12348 10124 12400 10130
rect 12268 10084 12348 10112
rect 12348 10066 12400 10072
rect 12084 9948 12204 9976
rect 12070 9888 12126 9897
rect 12070 9823 12126 9832
rect 11704 9648 11756 9654
rect 11704 9590 11756 9596
rect 11716 9217 11744 9590
rect 11980 9512 12032 9518
rect 11980 9454 12032 9460
rect 11886 9344 11942 9353
rect 11886 9279 11942 9288
rect 11702 9208 11758 9217
rect 11702 9143 11758 9152
rect 11796 9104 11848 9110
rect 11796 9046 11848 9052
rect 11808 8945 11836 9046
rect 11900 9042 11928 9279
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11794 8936 11850 8945
rect 11794 8871 11850 8880
rect 11624 8792 11928 8820
rect 11520 8560 11572 8566
rect 11520 8502 11572 8508
rect 11796 8560 11848 8566
rect 11796 8502 11848 8508
rect 11428 8492 11480 8498
rect 11428 8434 11480 8440
rect 11164 8214 11284 8242
rect 10817 8188 11113 8208
rect 10873 8186 10897 8188
rect 10953 8186 10977 8188
rect 11033 8186 11057 8188
rect 10895 8134 10897 8186
rect 10959 8134 10971 8186
rect 11033 8134 11035 8186
rect 10873 8132 10897 8134
rect 10953 8132 10977 8134
rect 11033 8132 11057 8134
rect 10817 8112 11113 8132
rect 11164 7834 11192 8214
rect 11242 8120 11298 8129
rect 11242 8055 11298 8064
rect 11072 7806 11192 7834
rect 10782 7576 10838 7585
rect 10782 7511 10838 7520
rect 10690 7440 10746 7449
rect 10690 7375 10746 7384
rect 10704 6798 10732 7375
rect 10796 7313 10824 7511
rect 11072 7449 11100 7806
rect 11152 7744 11204 7750
rect 11256 7732 11284 8055
rect 11204 7704 11284 7732
rect 11152 7686 11204 7692
rect 11058 7440 11114 7449
rect 11058 7375 11114 7384
rect 10968 7336 11020 7342
rect 10782 7304 10838 7313
rect 10782 7239 10838 7248
rect 10966 7304 10968 7313
rect 11020 7304 11022 7313
rect 11164 7274 11192 7686
rect 11334 7576 11390 7585
rect 11334 7511 11390 7520
rect 11348 7478 11376 7511
rect 11336 7472 11388 7478
rect 11336 7414 11388 7420
rect 11440 7410 11468 8434
rect 11520 8424 11572 8430
rect 11520 8366 11572 8372
rect 11428 7404 11480 7410
rect 11428 7346 11480 7352
rect 11256 7274 11468 7290
rect 10966 7239 11022 7248
rect 11152 7268 11204 7274
rect 11152 7210 11204 7216
rect 11256 7268 11480 7274
rect 11256 7262 11428 7268
rect 10817 7100 11113 7120
rect 10873 7098 10897 7100
rect 10953 7098 10977 7100
rect 11033 7098 11057 7100
rect 10895 7046 10897 7098
rect 10959 7046 10971 7098
rect 11033 7046 11035 7098
rect 10873 7044 10897 7046
rect 10953 7044 10977 7046
rect 11033 7044 11057 7046
rect 10817 7024 11113 7044
rect 10784 6860 10836 6866
rect 10784 6802 10836 6808
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10796 6644 10824 6802
rect 10704 6616 10824 6644
rect 10600 5908 10652 5914
rect 10600 5850 10652 5856
rect 10704 5846 10732 6616
rect 11256 6474 11284 7262
rect 11428 7210 11480 7216
rect 11336 7200 11388 7206
rect 11334 7168 11336 7177
rect 11388 7168 11390 7177
rect 11334 7103 11390 7112
rect 11336 6996 11388 7002
rect 11336 6938 11388 6944
rect 11164 6446 11284 6474
rect 11348 6458 11376 6938
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 11336 6452 11388 6458
rect 10817 6012 11113 6032
rect 10873 6010 10897 6012
rect 10953 6010 10977 6012
rect 11033 6010 11057 6012
rect 10895 5958 10897 6010
rect 10959 5958 10971 6010
rect 11033 5958 11035 6010
rect 10873 5956 10897 5958
rect 10953 5956 10977 5958
rect 11033 5956 11057 5958
rect 10817 5936 11113 5956
rect 10692 5840 10744 5846
rect 10692 5782 10744 5788
rect 10968 5840 11020 5846
rect 11164 5828 11192 6446
rect 11336 6394 11388 6400
rect 11244 6384 11296 6390
rect 11244 6326 11296 6332
rect 11256 5914 11284 6326
rect 11336 6180 11388 6186
rect 11336 6122 11388 6128
rect 11244 5908 11296 5914
rect 11244 5850 11296 5856
rect 11020 5800 11192 5828
rect 10968 5782 11020 5788
rect 10784 5704 10836 5710
rect 11060 5704 11112 5710
rect 10784 5646 10836 5652
rect 11058 5672 11060 5681
rect 11112 5672 11114 5681
rect 10796 5574 10824 5646
rect 11058 5607 11114 5616
rect 11242 5672 11298 5681
rect 11242 5607 11298 5616
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10508 5296 10560 5302
rect 10508 5238 10560 5244
rect 10428 5098 10640 5114
rect 10428 5092 10652 5098
rect 10428 5086 10600 5092
rect 10600 5034 10652 5040
rect 10416 5024 10468 5030
rect 10416 4966 10468 4972
rect 10324 4820 10376 4826
rect 10324 4762 10376 4768
rect 10428 4758 10456 4966
rect 10508 4820 10560 4826
rect 10704 4808 10732 5510
rect 10796 5358 11008 5386
rect 10796 5098 10824 5358
rect 10876 5296 10928 5302
rect 10876 5238 10928 5244
rect 10784 5092 10836 5098
rect 10784 5034 10836 5040
rect 10888 5012 10916 5238
rect 10980 5234 11008 5358
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 11256 5098 11284 5607
rect 11244 5092 11296 5098
rect 11244 5034 11296 5040
rect 10888 4984 11192 5012
rect 10817 4924 11113 4944
rect 10873 4922 10897 4924
rect 10953 4922 10977 4924
rect 11033 4922 11057 4924
rect 10895 4870 10897 4922
rect 10959 4870 10971 4922
rect 11033 4870 11035 4922
rect 10873 4868 10897 4870
rect 10953 4868 10977 4870
rect 11033 4868 11057 4870
rect 10817 4848 11113 4868
rect 10704 4780 10824 4808
rect 10508 4762 10560 4768
rect 10416 4752 10468 4758
rect 10416 4694 10468 4700
rect 10235 4644 10272 4672
rect 10235 4536 10263 4644
rect 10520 4604 10548 4762
rect 10336 4576 10548 4604
rect 10600 4616 10652 4622
rect 10235 4508 10272 4536
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 10244 4026 10272 4508
rect 10336 4214 10364 4576
rect 10600 4558 10652 4564
rect 10414 4448 10470 4457
rect 10414 4383 10470 4392
rect 10419 4264 10447 4383
rect 10419 4236 10456 4264
rect 10324 4208 10376 4214
rect 10324 4150 10376 4156
rect 10152 3998 10272 4026
rect 10324 4072 10376 4078
rect 10324 4014 10376 4020
rect 10048 2984 10100 2990
rect 10048 2926 10100 2932
rect 9956 2916 10008 2922
rect 9956 2858 10008 2864
rect 9968 2145 9996 2858
rect 10152 2514 10180 3998
rect 10230 3768 10286 3777
rect 10336 3738 10364 4014
rect 10428 3738 10456 4236
rect 10508 4208 10560 4214
rect 10508 4150 10560 4156
rect 10230 3703 10286 3712
rect 10324 3732 10376 3738
rect 10244 3040 10272 3703
rect 10324 3674 10376 3680
rect 10416 3732 10468 3738
rect 10416 3674 10468 3680
rect 10416 3460 10468 3466
rect 10416 3402 10468 3408
rect 10428 3126 10456 3402
rect 10416 3120 10468 3126
rect 10416 3062 10468 3068
rect 10324 3052 10376 3058
rect 10244 3012 10324 3040
rect 10324 2994 10376 3000
rect 10414 2680 10470 2689
rect 10520 2650 10548 4150
rect 10612 4078 10640 4558
rect 10796 4162 10824 4780
rect 10968 4752 11020 4758
rect 11020 4712 11100 4740
rect 10968 4694 11020 4700
rect 10876 4684 10928 4690
rect 10876 4626 10928 4632
rect 10704 4134 10824 4162
rect 10600 4072 10652 4078
rect 10600 4014 10652 4020
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10612 2922 10640 3878
rect 10704 3194 10732 4134
rect 10784 4072 10836 4078
rect 10782 4040 10784 4049
rect 10888 4060 10916 4626
rect 11072 4486 11100 4712
rect 10968 4480 11020 4486
rect 10968 4422 11020 4428
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 10980 4282 11008 4422
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 11060 4208 11112 4214
rect 11164 4196 11192 4984
rect 11348 4826 11376 6122
rect 11440 5710 11468 6734
rect 11532 6186 11560 8366
rect 11704 8016 11756 8022
rect 11704 7958 11756 7964
rect 11610 7440 11666 7449
rect 11610 7375 11666 7384
rect 11520 6180 11572 6186
rect 11520 6122 11572 6128
rect 11518 6080 11574 6089
rect 11518 6015 11574 6024
rect 11532 5846 11560 6015
rect 11520 5840 11572 5846
rect 11520 5782 11572 5788
rect 11428 5704 11480 5710
rect 11428 5646 11480 5652
rect 11520 5704 11572 5710
rect 11520 5646 11572 5652
rect 11532 5080 11560 5646
rect 11440 5052 11560 5080
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11244 4752 11296 4758
rect 11244 4694 11296 4700
rect 11112 4168 11192 4196
rect 11060 4150 11112 4156
rect 11256 4060 11284 4694
rect 11336 4616 11388 4622
rect 11336 4558 11388 4564
rect 11348 4486 11376 4558
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 11336 4208 11388 4214
rect 11336 4150 11388 4156
rect 10836 4040 10838 4049
rect 10888 4032 11284 4060
rect 10782 3975 10838 3984
rect 10817 3836 11113 3856
rect 10873 3834 10897 3836
rect 10953 3834 10977 3836
rect 11033 3834 11057 3836
rect 10895 3782 10897 3834
rect 10959 3782 10971 3834
rect 11033 3782 11035 3834
rect 10873 3780 10897 3782
rect 10953 3780 10977 3782
rect 11033 3780 11057 3782
rect 10817 3760 11113 3780
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 10692 3188 10744 3194
rect 10692 3130 10744 3136
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10704 2961 10732 2994
rect 10690 2952 10746 2961
rect 10600 2916 10652 2922
rect 10796 2922 10824 3470
rect 10690 2887 10746 2896
rect 10784 2916 10836 2922
rect 10600 2858 10652 2864
rect 10784 2858 10836 2864
rect 10817 2748 11113 2768
rect 10873 2746 10897 2748
rect 10953 2746 10977 2748
rect 11033 2746 11057 2748
rect 10895 2694 10897 2746
rect 10959 2694 10971 2746
rect 11033 2694 11035 2746
rect 10873 2692 10897 2694
rect 10953 2692 10977 2694
rect 11033 2692 11057 2694
rect 10817 2672 11113 2692
rect 10414 2615 10470 2624
rect 10508 2644 10560 2650
rect 10140 2508 10192 2514
rect 10140 2450 10192 2456
rect 9954 2136 10010 2145
rect 9954 2071 10010 2080
rect 9862 1728 9918 1737
rect 9862 1663 9918 1672
rect 9772 1556 9824 1562
rect 9772 1498 9824 1504
rect 9496 1216 9548 1222
rect 9496 1158 9548 1164
rect 9312 1148 9364 1154
rect 9312 1090 9364 1096
rect 9508 480 9536 1158
rect 9968 480 9996 2071
rect 10152 1834 10180 2450
rect 10428 2446 10456 2615
rect 11164 2632 11192 3674
rect 11348 3602 11376 4150
rect 11440 4146 11468 5052
rect 11518 4992 11574 5001
rect 11518 4927 11574 4936
rect 11428 4140 11480 4146
rect 11428 4082 11480 4088
rect 11428 3936 11480 3942
rect 11532 3913 11560 4927
rect 11624 4554 11652 7375
rect 11716 6662 11744 7958
rect 11808 6934 11836 8502
rect 11900 7002 11928 8792
rect 11888 6996 11940 7002
rect 11888 6938 11940 6944
rect 11796 6928 11848 6934
rect 11796 6870 11848 6876
rect 11992 6798 12020 9454
rect 12084 7478 12112 9823
rect 12176 9450 12204 9948
rect 12164 9444 12216 9450
rect 12164 9386 12216 9392
rect 12164 9172 12216 9178
rect 12164 9114 12216 9120
rect 12072 7472 12124 7478
rect 12176 7449 12204 9114
rect 12360 8566 12388 10066
rect 12440 9444 12492 9450
rect 12440 9386 12492 9392
rect 12452 8838 12480 9386
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12636 8634 12664 10220
rect 12728 9926 12756 10950
rect 12806 10911 12862 10920
rect 12820 10588 12848 10911
rect 12912 10742 12940 11494
rect 13004 11286 13032 14894
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 13282 14172 13578 14192
rect 13338 14170 13362 14172
rect 13418 14170 13442 14172
rect 13498 14170 13522 14172
rect 13360 14118 13362 14170
rect 13424 14118 13436 14170
rect 13498 14118 13500 14170
rect 13338 14116 13362 14118
rect 13418 14116 13442 14118
rect 13498 14116 13522 14118
rect 13282 14096 13578 14116
rect 13084 13388 13136 13394
rect 13084 13330 13136 13336
rect 13096 12986 13124 13330
rect 13176 13320 13228 13326
rect 13176 13262 13228 13268
rect 13452 13320 13504 13326
rect 13504 13280 13676 13308
rect 13452 13262 13504 13268
rect 13084 12980 13136 12986
rect 13084 12922 13136 12928
rect 13188 12889 13216 13262
rect 13282 13084 13578 13104
rect 13338 13082 13362 13084
rect 13418 13082 13442 13084
rect 13498 13082 13522 13084
rect 13360 13030 13362 13082
rect 13424 13030 13436 13082
rect 13498 13030 13500 13082
rect 13338 13028 13362 13030
rect 13418 13028 13442 13030
rect 13498 13028 13522 13030
rect 13282 13008 13578 13028
rect 13174 12880 13230 12889
rect 13174 12815 13230 12824
rect 13268 12844 13320 12850
rect 13268 12786 13320 12792
rect 13174 12744 13230 12753
rect 13174 12679 13230 12688
rect 13188 12442 13216 12679
rect 13176 12436 13228 12442
rect 13176 12378 13228 12384
rect 13188 12306 13216 12378
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 13084 12164 13136 12170
rect 13084 12106 13136 12112
rect 12992 11280 13044 11286
rect 12992 11222 13044 11228
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 12900 10736 12952 10742
rect 12900 10678 12952 10684
rect 12820 10560 12940 10588
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12820 10180 12848 10406
rect 12912 10282 12940 10560
rect 13004 10538 13032 11086
rect 13096 10792 13124 12106
rect 13280 12084 13308 12786
rect 13452 12640 13504 12646
rect 13452 12582 13504 12588
rect 13464 12442 13492 12582
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 13188 12056 13308 12084
rect 13188 11257 13216 12056
rect 13282 11996 13578 12016
rect 13338 11994 13362 11996
rect 13418 11994 13442 11996
rect 13498 11994 13522 11996
rect 13360 11942 13362 11994
rect 13424 11942 13436 11994
rect 13498 11942 13500 11994
rect 13338 11940 13362 11942
rect 13418 11940 13442 11942
rect 13498 11940 13522 11942
rect 13282 11920 13578 11940
rect 13360 11824 13412 11830
rect 13266 11792 13322 11801
rect 13360 11766 13412 11772
rect 13544 11824 13596 11830
rect 13544 11766 13596 11772
rect 13266 11727 13322 11736
rect 13174 11248 13230 11257
rect 13174 11183 13230 11192
rect 13280 11132 13308 11727
rect 13372 11354 13400 11766
rect 13450 11656 13506 11665
rect 13450 11591 13506 11600
rect 13464 11558 13492 11591
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 13556 11257 13584 11766
rect 13542 11248 13598 11257
rect 13542 11183 13598 11192
rect 13648 11200 13676 13280
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13740 12646 13768 13126
rect 13832 12918 13860 14418
rect 13820 12912 13872 12918
rect 13820 12854 13872 12860
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13924 12424 13952 15370
rect 14200 15094 14228 17520
rect 14660 15178 14688 17520
rect 14660 15150 14872 15178
rect 14188 15088 14240 15094
rect 14002 15056 14058 15065
rect 14188 15030 14240 15036
rect 14740 15088 14792 15094
rect 14740 15030 14792 15036
rect 14002 14991 14058 15000
rect 14016 13462 14044 14991
rect 14278 14920 14334 14929
rect 14278 14855 14334 14864
rect 14188 14272 14240 14278
rect 14188 14214 14240 14220
rect 14004 13456 14056 13462
rect 14004 13398 14056 13404
rect 14200 12782 14228 14214
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 14188 12436 14240 12442
rect 13924 12396 14044 12424
rect 13818 12336 13874 12345
rect 13818 12271 13874 12280
rect 13912 12300 13964 12306
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13740 11762 13768 12174
rect 13832 11898 13860 12271
rect 14016 12288 14044 12396
rect 14188 12378 14240 12384
rect 14016 12260 14136 12288
rect 13912 12242 13964 12248
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13728 11756 13780 11762
rect 13728 11698 13780 11704
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13648 11172 13768 11200
rect 13360 11144 13412 11150
rect 13280 11104 13360 11132
rect 13360 11086 13412 11092
rect 13634 11112 13690 11121
rect 13634 11047 13690 11056
rect 13282 10908 13578 10928
rect 13338 10906 13362 10908
rect 13418 10906 13442 10908
rect 13498 10906 13522 10908
rect 13360 10854 13362 10906
rect 13424 10854 13436 10906
rect 13498 10854 13500 10906
rect 13338 10852 13362 10854
rect 13418 10852 13442 10854
rect 13498 10852 13522 10854
rect 13282 10832 13578 10852
rect 13096 10764 13400 10792
rect 13372 10674 13400 10764
rect 13542 10704 13598 10713
rect 13360 10668 13412 10674
rect 13542 10639 13598 10648
rect 13360 10610 13412 10616
rect 12992 10532 13044 10538
rect 12992 10474 13044 10480
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 13174 10432 13230 10441
rect 12912 10266 13032 10282
rect 12912 10260 13044 10266
rect 12912 10254 12992 10260
rect 12992 10202 13044 10208
rect 12820 10152 12940 10180
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12808 9444 12860 9450
rect 12808 9386 12860 9392
rect 12716 9104 12768 9110
rect 12716 9046 12768 9052
rect 12728 8838 12756 9046
rect 12716 8832 12768 8838
rect 12716 8774 12768 8780
rect 12820 8673 12848 9386
rect 12806 8664 12862 8673
rect 12624 8628 12676 8634
rect 12806 8599 12862 8608
rect 12624 8570 12676 8576
rect 12348 8560 12400 8566
rect 12348 8502 12400 8508
rect 12530 8528 12586 8537
rect 12530 8463 12586 8472
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 12452 7954 12480 8366
rect 12544 8090 12572 8463
rect 12912 8265 12940 10152
rect 12992 9512 13044 9518
rect 12992 9454 13044 9460
rect 12898 8256 12954 8265
rect 12898 8191 12954 8200
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 12440 7948 12492 7954
rect 12440 7890 12492 7896
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 12072 7414 12124 7420
rect 12162 7440 12218 7449
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 11716 6322 11744 6598
rect 11794 6352 11850 6361
rect 11704 6316 11756 6322
rect 11794 6287 11850 6296
rect 11704 6258 11756 6264
rect 11716 5234 11744 6258
rect 11808 5914 11836 6287
rect 11900 6254 11928 6598
rect 11888 6248 11940 6254
rect 11888 6190 11940 6196
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 11796 5908 11848 5914
rect 11796 5850 11848 5856
rect 11900 5760 11928 6054
rect 11992 5846 12020 6734
rect 12084 6361 12112 7414
rect 12360 7410 12388 7822
rect 12532 7472 12584 7478
rect 12438 7440 12494 7449
rect 12162 7375 12218 7384
rect 12348 7404 12400 7410
rect 12532 7414 12584 7420
rect 12438 7375 12494 7384
rect 12348 7346 12400 7352
rect 12254 7304 12310 7313
rect 12254 7239 12310 7248
rect 12348 7268 12400 7274
rect 12162 7032 12218 7041
rect 12162 6967 12218 6976
rect 12176 6934 12204 6967
rect 12164 6928 12216 6934
rect 12164 6870 12216 6876
rect 12268 6440 12296 7239
rect 12348 7210 12400 7216
rect 12360 7002 12388 7210
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 12360 6633 12388 6802
rect 12346 6624 12402 6633
rect 12346 6559 12402 6568
rect 12176 6412 12296 6440
rect 12070 6352 12126 6361
rect 12070 6287 12126 6296
rect 12072 6248 12124 6254
rect 12072 6190 12124 6196
rect 11980 5840 12032 5846
rect 11980 5782 12032 5788
rect 11808 5732 11928 5760
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 11808 5114 11836 5732
rect 11980 5704 12032 5710
rect 11900 5664 11980 5692
rect 11900 5234 11928 5664
rect 11980 5646 12032 5652
rect 11978 5536 12034 5545
rect 11978 5471 12034 5480
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 11808 5086 11928 5114
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11702 4856 11758 4865
rect 11702 4791 11704 4800
rect 11756 4791 11758 4800
rect 11704 4762 11756 4768
rect 11612 4548 11664 4554
rect 11612 4490 11664 4496
rect 11624 4214 11652 4490
rect 11808 4457 11836 4966
rect 11794 4448 11850 4457
rect 11794 4383 11850 4392
rect 11794 4312 11850 4321
rect 11716 4270 11794 4298
rect 11612 4208 11664 4214
rect 11612 4150 11664 4156
rect 11716 3992 11744 4270
rect 11794 4247 11850 4256
rect 11604 3964 11744 3992
rect 11796 4004 11848 4010
rect 11428 3878 11480 3884
rect 11518 3904 11574 3913
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 10508 2586 10560 2592
rect 10796 2604 11192 2632
rect 10692 2576 10744 2582
rect 10692 2518 10744 2524
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 10600 2304 10652 2310
rect 10600 2246 10652 2252
rect 10140 1828 10192 1834
rect 10140 1770 10192 1776
rect 10612 1494 10640 2246
rect 10704 1601 10732 2518
rect 10690 1592 10746 1601
rect 10690 1527 10746 1536
rect 10600 1488 10652 1494
rect 10600 1430 10652 1436
rect 10416 1216 10468 1222
rect 10416 1158 10468 1164
rect 10428 480 10456 1158
rect 10796 480 10824 2604
rect 11152 2440 11204 2446
rect 11256 2428 11284 2994
rect 11440 2496 11468 3878
rect 11518 3839 11574 3848
rect 11604 3754 11632 3964
rect 11796 3946 11848 3952
rect 11702 3904 11758 3913
rect 11702 3839 11758 3848
rect 11604 3738 11652 3754
rect 11604 3732 11664 3738
rect 11604 3726 11612 3732
rect 11612 3674 11664 3680
rect 11716 3516 11744 3839
rect 11808 3738 11836 3946
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 11900 3602 11928 5086
rect 11992 5001 12020 5471
rect 11978 4992 12034 5001
rect 11978 4927 12034 4936
rect 12084 4865 12112 6190
rect 12070 4856 12126 4865
rect 12070 4791 12126 4800
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 11992 3777 12020 4626
rect 12084 4282 12112 4791
rect 12072 4276 12124 4282
rect 12072 4218 12124 4224
rect 11978 3768 12034 3777
rect 12176 3754 12204 6412
rect 12348 6384 12400 6390
rect 12254 6352 12310 6361
rect 12348 6326 12400 6332
rect 12254 6287 12310 6296
rect 12268 6089 12296 6287
rect 12254 6080 12310 6089
rect 12254 6015 12310 6024
rect 12256 5364 12308 5370
rect 12256 5306 12308 5312
rect 12268 4758 12296 5306
rect 12360 5302 12388 6326
rect 12452 6254 12480 7375
rect 12544 6905 12572 7414
rect 12636 7342 12664 7958
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 12898 7712 12954 7721
rect 12624 7336 12676 7342
rect 12622 7304 12624 7313
rect 12676 7304 12678 7313
rect 12622 7239 12678 7248
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12530 6896 12586 6905
rect 12530 6831 12586 6840
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12530 6080 12586 6089
rect 12452 5914 12480 6054
rect 12530 6015 12586 6024
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12438 5672 12494 5681
rect 12438 5607 12440 5616
rect 12492 5607 12494 5616
rect 12440 5578 12492 5584
rect 12544 5352 12572 6015
rect 12636 5692 12664 7142
rect 12728 7041 12756 7686
rect 12714 7032 12770 7041
rect 12714 6967 12770 6976
rect 12714 6896 12770 6905
rect 12714 6831 12770 6840
rect 12728 6798 12756 6831
rect 12716 6792 12768 6798
rect 12716 6734 12768 6740
rect 12716 6656 12768 6662
rect 12716 6598 12768 6604
rect 12728 6458 12756 6598
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12716 6248 12768 6254
rect 12820 6225 12848 7686
rect 12898 7647 12954 7656
rect 12912 7206 12940 7647
rect 12900 7200 12952 7206
rect 13004 7177 13032 9454
rect 13096 8294 13124 10406
rect 13174 10367 13230 10376
rect 13188 9518 13216 10367
rect 13556 10146 13584 10639
rect 13648 10266 13676 11047
rect 13740 10985 13768 11172
rect 13726 10976 13782 10985
rect 13726 10911 13782 10920
rect 13832 10826 13860 11494
rect 13740 10798 13860 10826
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13556 10118 13676 10146
rect 13282 9820 13578 9840
rect 13338 9818 13362 9820
rect 13418 9818 13442 9820
rect 13498 9818 13522 9820
rect 13360 9766 13362 9818
rect 13424 9766 13436 9818
rect 13498 9766 13500 9818
rect 13338 9764 13362 9766
rect 13418 9764 13442 9766
rect 13498 9764 13522 9766
rect 13282 9744 13578 9764
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 13268 9376 13320 9382
rect 13266 9344 13268 9353
rect 13320 9344 13322 9353
rect 13266 9279 13322 9288
rect 13464 9217 13492 9522
rect 13648 9489 13676 10118
rect 13634 9480 13690 9489
rect 13634 9415 13690 9424
rect 13450 9208 13506 9217
rect 13450 9143 13506 9152
rect 13740 9110 13768 10798
rect 13818 10568 13874 10577
rect 13818 10503 13820 10512
rect 13872 10503 13874 10512
rect 13820 10474 13872 10480
rect 13818 9616 13874 9625
rect 13818 9551 13874 9560
rect 13728 9104 13780 9110
rect 13728 9046 13780 9052
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 13282 8732 13578 8752
rect 13338 8730 13362 8732
rect 13418 8730 13442 8732
rect 13498 8730 13522 8732
rect 13360 8678 13362 8730
rect 13424 8678 13436 8730
rect 13498 8678 13500 8730
rect 13338 8676 13362 8678
rect 13418 8676 13442 8678
rect 13498 8676 13522 8678
rect 13282 8656 13578 8676
rect 13452 8560 13504 8566
rect 13452 8502 13504 8508
rect 13084 8288 13136 8294
rect 13084 8230 13136 8236
rect 13464 7993 13492 8502
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 13082 7984 13138 7993
rect 13450 7984 13506 7993
rect 13082 7919 13138 7928
rect 13176 7948 13228 7954
rect 13096 7410 13124 7919
rect 13450 7919 13506 7928
rect 13176 7890 13228 7896
rect 13084 7404 13136 7410
rect 13084 7346 13136 7352
rect 12900 7142 12952 7148
rect 12990 7168 13046 7177
rect 12912 7002 12940 7142
rect 12990 7103 13046 7112
rect 12990 7032 13046 7041
rect 12900 6996 12952 7002
rect 12990 6967 13046 6976
rect 12900 6938 12952 6944
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 12912 6390 12940 6734
rect 12900 6384 12952 6390
rect 12900 6326 12952 6332
rect 12716 6190 12768 6196
rect 12806 6216 12862 6225
rect 12728 6066 12756 6190
rect 12806 6151 12862 6160
rect 12728 6038 12940 6066
rect 12806 5944 12862 5953
rect 12806 5879 12862 5888
rect 12820 5846 12848 5879
rect 12808 5840 12860 5846
rect 12912 5817 12940 6038
rect 12808 5782 12860 5788
rect 12898 5808 12954 5817
rect 12898 5743 12954 5752
rect 12912 5710 12940 5743
rect 12900 5704 12952 5710
rect 12636 5664 12848 5692
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 12452 5324 12572 5352
rect 12622 5400 12678 5409
rect 12622 5335 12678 5344
rect 12348 5296 12400 5302
rect 12348 5238 12400 5244
rect 12256 4752 12308 4758
rect 12256 4694 12308 4700
rect 12254 4448 12310 4457
rect 12254 4383 12310 4392
rect 12268 3913 12296 4383
rect 12452 4146 12480 5324
rect 12636 5250 12664 5335
rect 12544 5234 12664 5250
rect 12532 5228 12664 5234
rect 12584 5222 12664 5228
rect 12532 5170 12584 5176
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 12532 5024 12584 5030
rect 12532 4966 12584 4972
rect 12544 4826 12572 4966
rect 12636 4826 12664 5102
rect 12532 4820 12584 4826
rect 12532 4762 12584 4768
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12624 4480 12676 4486
rect 12624 4422 12676 4428
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 12544 4049 12572 4422
rect 12530 4040 12586 4049
rect 12530 3975 12586 3984
rect 12440 3936 12492 3942
rect 12254 3904 12310 3913
rect 12440 3878 12492 3884
rect 12254 3839 12310 3848
rect 12176 3738 12296 3754
rect 12176 3732 12308 3738
rect 12176 3726 12256 3732
rect 11978 3703 12034 3712
rect 12256 3674 12308 3680
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 11796 3528 11848 3534
rect 11716 3488 11796 3516
rect 11796 3470 11848 3476
rect 11610 3088 11666 3097
rect 11808 3058 11836 3470
rect 12268 3369 12296 3674
rect 12452 3641 12480 3878
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 12438 3632 12494 3641
rect 12438 3567 12494 3576
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 11886 3360 11942 3369
rect 11886 3295 11942 3304
rect 12254 3360 12310 3369
rect 12254 3295 12310 3304
rect 11900 3097 11928 3295
rect 12256 3188 12308 3194
rect 12256 3130 12308 3136
rect 11886 3088 11942 3097
rect 11610 3023 11666 3032
rect 11796 3052 11848 3058
rect 11520 2848 11572 2854
rect 11520 2790 11572 2796
rect 11532 2689 11560 2790
rect 11518 2680 11574 2689
rect 11518 2615 11574 2624
rect 11204 2400 11284 2428
rect 11348 2468 11468 2496
rect 11152 2382 11204 2388
rect 11242 1456 11298 1465
rect 11242 1391 11298 1400
rect 11256 480 11284 1391
rect 11348 610 11376 2468
rect 11428 2372 11480 2378
rect 11428 2314 11480 2320
rect 11440 1630 11468 2314
rect 11428 1624 11480 1630
rect 11428 1566 11480 1572
rect 11336 604 11388 610
rect 11336 546 11388 552
rect 11624 480 11652 3023
rect 11886 3023 11942 3032
rect 12164 3052 12216 3058
rect 11796 2994 11848 3000
rect 12164 2994 12216 3000
rect 11704 2916 11756 2922
rect 11704 2858 11756 2864
rect 11716 2038 11744 2858
rect 11794 2544 11850 2553
rect 11794 2479 11796 2488
rect 11848 2479 11850 2488
rect 11796 2450 11848 2456
rect 11980 2304 12032 2310
rect 11980 2246 12032 2252
rect 11704 2032 11756 2038
rect 11704 1974 11756 1980
rect 11992 1766 12020 2246
rect 12070 2136 12126 2145
rect 12070 2071 12126 2080
rect 11980 1760 12032 1766
rect 11980 1702 12032 1708
rect 12084 480 12112 2071
rect 12176 1154 12204 2994
rect 12268 2961 12296 3130
rect 12254 2952 12310 2961
rect 12254 2887 12310 2896
rect 12360 2854 12388 3470
rect 12438 3360 12494 3369
rect 12438 3295 12494 3304
rect 12348 2848 12400 2854
rect 12348 2790 12400 2796
rect 12452 1834 12480 3295
rect 12544 3126 12572 3674
rect 12532 3120 12584 3126
rect 12532 3062 12584 3068
rect 12636 3058 12664 4422
rect 12728 4078 12756 5510
rect 12820 4214 12848 5664
rect 12900 5646 12952 5652
rect 12898 5536 12954 5545
rect 12898 5471 12954 5480
rect 12912 5302 12940 5471
rect 13004 5409 13032 6967
rect 13188 6866 13216 7890
rect 13282 7644 13578 7664
rect 13338 7642 13362 7644
rect 13418 7642 13442 7644
rect 13498 7642 13522 7644
rect 13360 7590 13362 7642
rect 13424 7590 13436 7642
rect 13498 7590 13500 7642
rect 13338 7588 13362 7590
rect 13418 7588 13442 7590
rect 13498 7588 13522 7590
rect 13282 7568 13578 7588
rect 13360 7268 13412 7274
rect 13360 7210 13412 7216
rect 13372 7177 13400 7210
rect 13452 7200 13504 7206
rect 13358 7168 13414 7177
rect 13452 7142 13504 7148
rect 13358 7103 13414 7112
rect 13084 6860 13136 6866
rect 13084 6802 13136 6808
rect 13176 6860 13228 6866
rect 13176 6802 13228 6808
rect 13096 6322 13124 6802
rect 13464 6730 13492 7142
rect 13176 6724 13228 6730
rect 13176 6666 13228 6672
rect 13452 6724 13504 6730
rect 13452 6666 13504 6672
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 13188 6254 13216 6666
rect 13282 6556 13578 6576
rect 13338 6554 13362 6556
rect 13418 6554 13442 6556
rect 13498 6554 13522 6556
rect 13360 6502 13362 6554
rect 13424 6502 13436 6554
rect 13498 6502 13500 6554
rect 13338 6500 13362 6502
rect 13418 6500 13442 6502
rect 13498 6500 13522 6502
rect 13282 6480 13578 6500
rect 13648 6458 13676 8434
rect 13740 8401 13768 8774
rect 13832 8634 13860 9551
rect 13924 9466 13952 12242
rect 14108 11642 14136 12260
rect 14016 11614 14136 11642
rect 14016 10130 14044 11614
rect 14096 11552 14148 11558
rect 14096 11494 14148 11500
rect 14108 11121 14136 11494
rect 14200 11218 14228 12378
rect 14188 11212 14240 11218
rect 14188 11154 14240 11160
rect 14094 11112 14150 11121
rect 14094 11047 14150 11056
rect 14200 10996 14228 11154
rect 14108 10968 14228 10996
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 13924 9438 14044 9466
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13726 8392 13782 8401
rect 13726 8327 13782 8336
rect 13728 8288 13780 8294
rect 13728 8230 13780 8236
rect 13636 6452 13688 6458
rect 13636 6394 13688 6400
rect 13740 6338 13768 8230
rect 13820 7812 13872 7818
rect 13820 7754 13872 7760
rect 13648 6310 13768 6338
rect 13176 6248 13228 6254
rect 13176 6190 13228 6196
rect 13268 6248 13320 6254
rect 13268 6190 13320 6196
rect 13450 6216 13506 6225
rect 13280 5710 13308 6190
rect 13450 6151 13506 6160
rect 13464 6118 13492 6151
rect 13452 6112 13504 6118
rect 13452 6054 13504 6060
rect 13464 5710 13492 6054
rect 13268 5704 13320 5710
rect 13188 5664 13268 5692
rect 12990 5400 13046 5409
rect 12990 5335 13046 5344
rect 12900 5296 12952 5302
rect 12900 5238 12952 5244
rect 12898 5128 12954 5137
rect 12898 5063 12954 5072
rect 13084 5092 13136 5098
rect 12912 4690 12940 5063
rect 13084 5034 13136 5040
rect 12900 4684 12952 4690
rect 12900 4626 12952 4632
rect 12992 4616 13044 4622
rect 12990 4584 12992 4593
rect 13044 4584 13046 4593
rect 12900 4548 12952 4554
rect 12990 4519 13046 4528
rect 12900 4490 12952 4496
rect 12912 4457 12940 4490
rect 12898 4448 12954 4457
rect 12898 4383 12954 4392
rect 12808 4208 12860 4214
rect 12808 4150 12860 4156
rect 12716 4072 12768 4078
rect 12716 4014 12768 4020
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 12728 3738 12756 3878
rect 12716 3732 12768 3738
rect 12716 3674 12768 3680
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 12716 3460 12768 3466
rect 12716 3402 12768 3408
rect 12624 3052 12676 3058
rect 12624 2994 12676 3000
rect 12532 2984 12584 2990
rect 12532 2926 12584 2932
rect 12440 1828 12492 1834
rect 12440 1770 12492 1776
rect 12164 1148 12216 1154
rect 12164 1090 12216 1096
rect 12544 480 12572 2926
rect 12624 2916 12676 2922
rect 12624 2858 12676 2864
rect 12636 2038 12664 2858
rect 12728 2650 12756 3402
rect 12808 3392 12860 3398
rect 12808 3334 12860 3340
rect 12820 3126 12848 3334
rect 12808 3120 12860 3126
rect 12808 3062 12860 3068
rect 12912 2854 12940 3674
rect 12900 2848 12952 2854
rect 12900 2790 12952 2796
rect 12716 2644 12768 2650
rect 12716 2586 12768 2592
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 12624 2032 12676 2038
rect 12624 1974 12676 1980
rect 12912 1902 12940 2586
rect 13004 2582 13032 3878
rect 12992 2576 13044 2582
rect 12992 2518 13044 2524
rect 13096 2446 13124 5034
rect 13188 4758 13216 5664
rect 13268 5646 13320 5652
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 13282 5468 13578 5488
rect 13338 5466 13362 5468
rect 13418 5466 13442 5468
rect 13498 5466 13522 5468
rect 13360 5414 13362 5466
rect 13424 5414 13436 5466
rect 13498 5414 13500 5466
rect 13338 5412 13362 5414
rect 13418 5412 13442 5414
rect 13498 5412 13522 5414
rect 13282 5392 13578 5412
rect 13268 5024 13320 5030
rect 13268 4966 13320 4972
rect 13176 4752 13228 4758
rect 13176 4694 13228 4700
rect 13280 4468 13308 4966
rect 13542 4720 13598 4729
rect 13542 4655 13544 4664
rect 13596 4655 13598 4664
rect 13544 4626 13596 4632
rect 13188 4440 13308 4468
rect 13188 3738 13216 4440
rect 13282 4380 13578 4400
rect 13338 4378 13362 4380
rect 13418 4378 13442 4380
rect 13498 4378 13522 4380
rect 13360 4326 13362 4378
rect 13424 4326 13436 4378
rect 13498 4326 13500 4378
rect 13338 4324 13362 4326
rect 13418 4324 13442 4326
rect 13498 4324 13522 4326
rect 13282 4304 13578 4324
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 13360 4072 13412 4078
rect 13360 4014 13412 4020
rect 13266 3768 13322 3777
rect 13176 3732 13228 3738
rect 13372 3738 13400 4014
rect 13266 3703 13322 3712
rect 13360 3732 13412 3738
rect 13176 3674 13228 3680
rect 13174 3632 13230 3641
rect 13174 3567 13176 3576
rect 13228 3567 13230 3576
rect 13176 3538 13228 3544
rect 13188 2650 13216 3538
rect 13280 3466 13308 3703
rect 13360 3674 13412 3680
rect 13556 3534 13584 4082
rect 13648 3652 13676 6310
rect 13832 6254 13860 7754
rect 13924 6934 13952 9318
rect 14016 8838 14044 9438
rect 14108 8906 14136 10968
rect 14200 10062 14228 10093
rect 14188 10056 14240 10062
rect 14186 10024 14188 10033
rect 14240 10024 14242 10033
rect 14186 9959 14242 9968
rect 14096 8900 14148 8906
rect 14096 8842 14148 8848
rect 14004 8832 14056 8838
rect 14004 8774 14056 8780
rect 14096 8560 14148 8566
rect 14096 8502 14148 8508
rect 14108 8401 14136 8502
rect 14094 8392 14150 8401
rect 14004 8356 14056 8362
rect 14094 8327 14150 8336
rect 14004 8298 14056 8304
rect 14016 7818 14044 8298
rect 14200 8242 14228 9959
rect 14292 9654 14320 14855
rect 14556 14544 14608 14550
rect 14556 14486 14608 14492
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 14372 12912 14424 12918
rect 14372 12854 14424 12860
rect 14384 11150 14412 12854
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14476 10810 14504 14350
rect 14464 10804 14516 10810
rect 14464 10746 14516 10752
rect 14372 10532 14424 10538
rect 14372 10474 14424 10480
rect 14280 9648 14332 9654
rect 14280 9590 14332 9596
rect 14280 8900 14332 8906
rect 14280 8842 14332 8848
rect 14108 8214 14228 8242
rect 14004 7812 14056 7818
rect 14004 7754 14056 7760
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 13912 6928 13964 6934
rect 13912 6870 13964 6876
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 13910 6216 13966 6225
rect 13910 6151 13912 6160
rect 13964 6151 13966 6160
rect 13912 6122 13964 6128
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13740 5302 13768 5850
rect 13832 5681 13860 6054
rect 13818 5672 13874 5681
rect 13818 5607 13874 5616
rect 13728 5296 13780 5302
rect 13728 5238 13780 5244
rect 13924 5234 13952 6122
rect 14016 5778 14044 7482
rect 14108 7478 14136 8214
rect 14292 7970 14320 8842
rect 14200 7942 14320 7970
rect 14096 7472 14148 7478
rect 14096 7414 14148 7420
rect 14096 7268 14148 7274
rect 14096 7210 14148 7216
rect 14108 7002 14136 7210
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 14200 6866 14228 7942
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14292 7410 14320 7822
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14280 7268 14332 7274
rect 14280 7210 14332 7216
rect 14188 6860 14240 6866
rect 14188 6802 14240 6808
rect 14188 6656 14240 6662
rect 14188 6598 14240 6604
rect 14094 6352 14150 6361
rect 14094 6287 14150 6296
rect 14108 5914 14136 6287
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 14004 5772 14056 5778
rect 14004 5714 14056 5720
rect 14096 5704 14148 5710
rect 14096 5646 14148 5652
rect 14004 5568 14056 5574
rect 14004 5510 14056 5516
rect 13820 5228 13872 5234
rect 13820 5170 13872 5176
rect 13912 5228 13964 5234
rect 13912 5170 13964 5176
rect 13832 5030 13860 5170
rect 14016 5098 14044 5510
rect 14004 5092 14056 5098
rect 14004 5034 14056 5040
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 13912 5024 13964 5030
rect 13912 4966 13964 4972
rect 14002 4992 14058 5001
rect 13726 4856 13782 4865
rect 13726 4791 13782 4800
rect 13740 4622 13768 4791
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13728 3936 13780 3942
rect 13726 3904 13728 3913
rect 13780 3904 13782 3913
rect 13726 3839 13782 3848
rect 13648 3624 13768 3652
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13634 3496 13690 3505
rect 13268 3460 13320 3466
rect 13634 3431 13690 3440
rect 13268 3402 13320 3408
rect 13282 3292 13578 3312
rect 13338 3290 13362 3292
rect 13418 3290 13442 3292
rect 13498 3290 13522 3292
rect 13360 3238 13362 3290
rect 13424 3238 13436 3290
rect 13498 3238 13500 3290
rect 13338 3236 13362 3238
rect 13418 3236 13442 3238
rect 13498 3236 13522 3238
rect 13282 3216 13578 3236
rect 13648 3194 13676 3431
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 13268 3120 13320 3126
rect 13266 3088 13268 3097
rect 13320 3088 13322 3097
rect 13266 3023 13322 3032
rect 13450 3088 13506 3097
rect 13740 3058 13768 3624
rect 13450 3023 13506 3032
rect 13728 3052 13780 3058
rect 13464 2990 13492 3023
rect 13728 2994 13780 3000
rect 13268 2984 13320 2990
rect 13268 2926 13320 2932
rect 13452 2984 13504 2990
rect 13832 2938 13860 4966
rect 13924 4282 13952 4966
rect 14002 4927 14058 4936
rect 13912 4276 13964 4282
rect 13912 4218 13964 4224
rect 13912 4072 13964 4078
rect 13910 4040 13912 4049
rect 13964 4040 13966 4049
rect 13910 3975 13966 3984
rect 13924 3670 13952 3975
rect 13912 3664 13964 3670
rect 13912 3606 13964 3612
rect 14016 3534 14044 4927
rect 13912 3528 13964 3534
rect 13912 3470 13964 3476
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 13924 2990 13952 3470
rect 14108 3380 14136 5646
rect 14016 3352 14136 3380
rect 13452 2926 13504 2932
rect 13176 2644 13228 2650
rect 13176 2586 13228 2592
rect 13174 2544 13230 2553
rect 13174 2479 13176 2488
rect 13228 2479 13230 2488
rect 13176 2450 13228 2456
rect 13084 2440 13136 2446
rect 13280 2394 13308 2926
rect 13740 2910 13860 2938
rect 13912 2984 13964 2990
rect 13912 2926 13964 2932
rect 13450 2680 13506 2689
rect 13450 2615 13506 2624
rect 13084 2382 13136 2388
rect 13188 2366 13308 2394
rect 13464 2378 13492 2615
rect 13452 2372 13504 2378
rect 12900 1896 12952 1902
rect 12900 1838 12952 1844
rect 13188 1358 13216 2366
rect 13452 2314 13504 2320
rect 13282 2204 13578 2224
rect 13338 2202 13362 2204
rect 13418 2202 13442 2204
rect 13498 2202 13522 2204
rect 13360 2150 13362 2202
rect 13424 2150 13436 2202
rect 13498 2150 13500 2202
rect 13338 2148 13362 2150
rect 13418 2148 13442 2150
rect 13498 2148 13522 2150
rect 13282 2128 13578 2148
rect 13360 1828 13412 1834
rect 13360 1770 13412 1776
rect 13176 1352 13228 1358
rect 13176 1294 13228 1300
rect 12900 944 12952 950
rect 12900 886 12952 892
rect 12912 480 12940 886
rect 13372 480 13400 1770
rect 13740 950 13768 2910
rect 14016 2836 14044 3352
rect 14200 3108 14228 6598
rect 14292 3670 14320 7210
rect 14280 3664 14332 3670
rect 14280 3606 14332 3612
rect 13832 2808 14044 2836
rect 14108 3080 14228 3108
rect 13728 944 13780 950
rect 13728 886 13780 892
rect 13832 480 13860 2808
rect 13912 2304 13964 2310
rect 13912 2246 13964 2252
rect 13924 1970 13952 2246
rect 13912 1964 13964 1970
rect 13912 1906 13964 1912
rect 14108 1698 14136 3080
rect 14186 2952 14242 2961
rect 14186 2887 14242 2896
rect 14096 1692 14148 1698
rect 14096 1634 14148 1640
rect 14200 480 14228 2887
rect 14292 1290 14320 3606
rect 14384 2990 14412 10474
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14476 10169 14504 10406
rect 14462 10160 14518 10169
rect 14462 10095 14518 10104
rect 14464 9920 14516 9926
rect 14464 9862 14516 9868
rect 14476 7698 14504 9862
rect 14568 9178 14596 14486
rect 14752 12186 14780 15030
rect 14660 12158 14780 12186
rect 14660 10538 14688 12158
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14752 11354 14780 12038
rect 14844 11694 14872 15150
rect 14924 12640 14976 12646
rect 14924 12582 14976 12588
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 14830 11520 14886 11529
rect 14830 11455 14886 11464
rect 14740 11348 14792 11354
rect 14740 11290 14792 11296
rect 14740 10804 14792 10810
rect 14740 10746 14792 10752
rect 14648 10532 14700 10538
rect 14648 10474 14700 10480
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14752 8922 14780 10746
rect 14660 8894 14780 8922
rect 14554 8392 14610 8401
rect 14554 8327 14556 8336
rect 14608 8327 14610 8336
rect 14556 8298 14608 8304
rect 14660 8022 14688 8894
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14648 8016 14700 8022
rect 14648 7958 14700 7964
rect 14476 7670 14596 7698
rect 14464 7472 14516 7478
rect 14464 7414 14516 7420
rect 14476 7154 14504 7414
rect 14568 7342 14596 7670
rect 14752 7426 14780 8774
rect 14660 7398 14780 7426
rect 14556 7336 14608 7342
rect 14556 7278 14608 7284
rect 14476 7126 14596 7154
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 14476 5370 14504 6802
rect 14464 5364 14516 5370
rect 14464 5306 14516 5312
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 14476 3777 14504 4966
rect 14568 3942 14596 7126
rect 14660 6118 14688 7398
rect 14844 7290 14872 11455
rect 14752 7262 14872 7290
rect 14752 6390 14780 7262
rect 14832 7200 14884 7206
rect 14832 7142 14884 7148
rect 14740 6384 14792 6390
rect 14740 6326 14792 6332
rect 14740 6248 14792 6254
rect 14740 6190 14792 6196
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14660 5030 14688 6054
rect 14752 5914 14780 6190
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 14648 5024 14700 5030
rect 14700 4984 14780 5012
rect 14648 4966 14700 4972
rect 14646 4856 14702 4865
rect 14646 4791 14702 4800
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14462 3768 14518 3777
rect 14462 3703 14518 3712
rect 14556 3732 14608 3738
rect 14556 3674 14608 3680
rect 14372 2984 14424 2990
rect 14372 2926 14424 2932
rect 14568 2417 14596 3674
rect 14554 2408 14610 2417
rect 14554 2343 14610 2352
rect 14464 2304 14516 2310
rect 14464 2246 14516 2252
rect 14556 2304 14608 2310
rect 14556 2246 14608 2252
rect 14476 2106 14504 2246
rect 14464 2100 14516 2106
rect 14464 2042 14516 2048
rect 14568 1426 14596 2246
rect 14556 1420 14608 1426
rect 14556 1362 14608 1368
rect 14280 1284 14332 1290
rect 14280 1226 14332 1232
rect 14660 480 14688 4791
rect 14752 3516 14780 4984
rect 14844 3738 14872 7142
rect 14936 6458 14964 12582
rect 15028 11744 15056 17520
rect 15488 14414 15516 17520
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15948 14006 15976 17520
rect 15936 14000 15988 14006
rect 15936 13942 15988 13948
rect 15290 13288 15346 13297
rect 15290 13223 15346 13232
rect 15304 11762 15332 13223
rect 15384 12708 15436 12714
rect 15384 12650 15436 12656
rect 15292 11756 15344 11762
rect 15028 11716 15240 11744
rect 15016 11620 15068 11626
rect 15016 11562 15068 11568
rect 15028 10810 15056 11562
rect 15016 10804 15068 10810
rect 15016 10746 15068 10752
rect 15016 10668 15068 10674
rect 15016 10610 15068 10616
rect 15028 9722 15056 10610
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 15016 9716 15068 9722
rect 15016 9658 15068 9664
rect 15014 9616 15070 9625
rect 15120 9586 15148 10542
rect 15212 10441 15240 11716
rect 15292 11698 15344 11704
rect 15292 11620 15344 11626
rect 15292 11562 15344 11568
rect 15198 10432 15254 10441
rect 15198 10367 15254 10376
rect 15014 9551 15070 9560
rect 15108 9580 15160 9586
rect 15028 7410 15056 9551
rect 15108 9522 15160 9528
rect 15108 8288 15160 8294
rect 15108 8230 15160 8236
rect 15120 7857 15148 8230
rect 15106 7848 15162 7857
rect 15106 7783 15162 7792
rect 15016 7404 15068 7410
rect 15016 7346 15068 7352
rect 15028 6798 15056 7346
rect 15108 7336 15160 7342
rect 15108 7278 15160 7284
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 14924 6452 14976 6458
rect 14924 6394 14976 6400
rect 15120 6338 15148 7278
rect 15198 6896 15254 6905
rect 15198 6831 15200 6840
rect 15252 6831 15254 6840
rect 15200 6802 15252 6808
rect 15016 6316 15068 6322
rect 15120 6310 15240 6338
rect 15016 6258 15068 6264
rect 15028 6225 15056 6258
rect 15014 6216 15070 6225
rect 15014 6151 15070 6160
rect 14924 5228 14976 5234
rect 14924 5170 14976 5176
rect 14936 4622 14964 5170
rect 15016 5092 15068 5098
rect 15016 5034 15068 5040
rect 14924 4616 14976 4622
rect 14924 4558 14976 4564
rect 15028 4185 15056 5034
rect 15212 4214 15240 6310
rect 15304 4826 15332 11562
rect 15396 10470 15424 12650
rect 16316 11830 16344 17520
rect 16776 12442 16804 17520
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 16304 11824 16356 11830
rect 16304 11766 16356 11772
rect 15476 11008 15528 11014
rect 15476 10950 15528 10956
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15488 9081 15516 10950
rect 15936 10464 15988 10470
rect 15936 10406 15988 10412
rect 15474 9072 15530 9081
rect 15474 9007 15530 9016
rect 15382 8936 15438 8945
rect 15382 8871 15438 8880
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 15200 4208 15252 4214
rect 15014 4176 15070 4185
rect 14924 4140 14976 4146
rect 15200 4150 15252 4156
rect 15014 4111 15070 4120
rect 14924 4082 14976 4088
rect 14832 3732 14884 3738
rect 14832 3674 14884 3680
rect 14936 3670 14964 4082
rect 15108 3936 15160 3942
rect 15014 3904 15070 3913
rect 15108 3878 15160 3884
rect 15014 3839 15070 3848
rect 14924 3664 14976 3670
rect 14924 3606 14976 3612
rect 14752 3488 14964 3516
rect 14740 2848 14792 2854
rect 14740 2790 14792 2796
rect 14752 1737 14780 2790
rect 14936 2582 14964 3488
rect 14924 2576 14976 2582
rect 14924 2518 14976 2524
rect 15028 2009 15056 3839
rect 15014 2000 15070 2009
rect 15014 1935 15070 1944
rect 14738 1728 14794 1737
rect 14738 1663 14794 1672
rect 15028 480 15056 1935
rect 15120 1222 15148 3878
rect 15304 2514 15332 4762
rect 15396 3097 15424 8871
rect 15476 6180 15528 6186
rect 15476 6122 15528 6128
rect 15382 3088 15438 3097
rect 15382 3023 15438 3032
rect 15292 2508 15344 2514
rect 15292 2450 15344 2456
rect 15108 1216 15160 1222
rect 15108 1158 15160 1164
rect 15488 480 15516 6122
rect 15948 2825 15976 10406
rect 16764 5296 16816 5302
rect 16764 5238 16816 5244
rect 16304 5092 16356 5098
rect 16304 5034 16356 5040
rect 15934 2816 15990 2825
rect 15934 2751 15990 2760
rect 15948 480 15976 2751
rect 16316 480 16344 5034
rect 16776 480 16804 5238
rect 2778 439 2834 448
rect 3146 0 3202 480
rect 3606 0 3662 480
rect 3974 0 4030 480
rect 4434 0 4490 480
rect 4802 0 4858 480
rect 5262 0 5318 480
rect 5722 0 5778 480
rect 6090 0 6146 480
rect 6550 0 6606 480
rect 7010 0 7066 480
rect 7378 0 7434 480
rect 7838 0 7894 480
rect 8206 0 8262 480
rect 8666 0 8722 480
rect 9126 0 9182 480
rect 9494 0 9550 480
rect 9954 0 10010 480
rect 10414 0 10470 480
rect 10782 0 10838 480
rect 11242 0 11298 480
rect 11610 0 11666 480
rect 12070 0 12126 480
rect 12530 0 12586 480
rect 12898 0 12954 480
rect 13358 0 13414 480
rect 13818 0 13874 480
rect 14186 0 14242 480
rect 14646 0 14702 480
rect 15014 0 15070 480
rect 15474 0 15530 480
rect 15934 0 15990 480
rect 16302 0 16358 480
rect 16762 0 16818 480
<< via2 >>
rect 1858 13776 1914 13832
rect 2962 16224 3018 16280
rect 2318 15000 2374 15056
rect 2870 15136 2926 15192
rect 2226 14900 2228 14920
rect 2228 14900 2280 14920
rect 2280 14900 2282 14920
rect 2226 14864 2282 14900
rect 2502 13912 2558 13968
rect 1674 12008 1730 12064
rect 2042 12280 2098 12336
rect 1858 10920 1914 10976
rect 1950 10648 2006 10704
rect 1858 9832 1914 9888
rect 1398 5772 1454 5808
rect 1398 5752 1400 5772
rect 1400 5752 1452 5772
rect 1452 5752 1454 5772
rect 1398 4120 1454 4176
rect 1306 3576 1362 3632
rect 1766 7828 1768 7848
rect 1768 7828 1820 7848
rect 1820 7828 1822 7848
rect 1766 7792 1822 7828
rect 1766 6740 1768 6760
rect 1768 6740 1820 6760
rect 1820 6740 1822 6760
rect 1766 6704 1822 6740
rect 1490 3032 1546 3088
rect 1858 5072 1914 5128
rect 1858 4664 1914 4720
rect 2318 12300 2374 12336
rect 2318 12280 2320 12300
rect 2320 12280 2372 12300
rect 2372 12280 2374 12300
rect 2410 12180 2412 12200
rect 2412 12180 2464 12200
rect 2464 12180 2466 12200
rect 2410 12144 2466 12180
rect 2410 11620 2466 11656
rect 2410 11600 2412 11620
rect 2412 11600 2464 11620
rect 2464 11600 2466 11620
rect 2502 11192 2558 11248
rect 2502 11092 2504 11112
rect 2504 11092 2556 11112
rect 2556 11092 2558 11112
rect 2502 11056 2558 11092
rect 2410 10512 2466 10568
rect 3421 15258 3477 15260
rect 3501 15258 3557 15260
rect 3581 15258 3637 15260
rect 3661 15258 3717 15260
rect 3421 15206 3447 15258
rect 3447 15206 3477 15258
rect 3501 15206 3511 15258
rect 3511 15206 3557 15258
rect 3581 15206 3627 15258
rect 3627 15206 3637 15258
rect 3661 15206 3691 15258
rect 3691 15206 3717 15258
rect 3421 15204 3477 15206
rect 3501 15204 3557 15206
rect 3581 15204 3637 15206
rect 3661 15204 3717 15206
rect 3146 15000 3202 15056
rect 3698 14900 3700 14920
rect 3700 14900 3752 14920
rect 3752 14900 3754 14920
rect 3146 14048 3202 14104
rect 3698 14864 3754 14900
rect 2778 13096 2834 13152
rect 2778 12824 2834 12880
rect 2226 7792 2282 7848
rect 2042 4664 2098 4720
rect 3054 12824 3110 12880
rect 2870 7384 2926 7440
rect 2042 3848 2098 3904
rect 2318 3440 2374 3496
rect 2778 6180 2834 6216
rect 2778 6160 2780 6180
rect 2780 6160 2832 6180
rect 2832 6160 2834 6180
rect 1674 1400 1730 1456
rect 2778 4800 2834 4856
rect 3054 10412 3056 10432
rect 3056 10412 3108 10432
rect 3108 10412 3110 10432
rect 3054 10376 3110 10412
rect 3974 17312 4030 17368
rect 3421 14170 3477 14172
rect 3501 14170 3557 14172
rect 3581 14170 3637 14172
rect 3661 14170 3717 14172
rect 3421 14118 3447 14170
rect 3447 14118 3477 14170
rect 3501 14118 3511 14170
rect 3511 14118 3557 14170
rect 3581 14118 3627 14170
rect 3627 14118 3637 14170
rect 3661 14118 3691 14170
rect 3691 14118 3717 14170
rect 3421 14116 3477 14118
rect 3501 14116 3557 14118
rect 3581 14116 3637 14118
rect 3661 14116 3717 14118
rect 3421 13082 3477 13084
rect 3501 13082 3557 13084
rect 3581 13082 3637 13084
rect 3661 13082 3717 13084
rect 3421 13030 3447 13082
rect 3447 13030 3477 13082
rect 3501 13030 3511 13082
rect 3511 13030 3557 13082
rect 3581 13030 3627 13082
rect 3627 13030 3637 13082
rect 3661 13030 3691 13082
rect 3691 13030 3717 13082
rect 3421 13028 3477 13030
rect 3501 13028 3557 13030
rect 3581 13028 3637 13030
rect 3661 13028 3717 13030
rect 3698 12824 3754 12880
rect 3421 11994 3477 11996
rect 3501 11994 3557 11996
rect 3581 11994 3637 11996
rect 3661 11994 3717 11996
rect 3421 11942 3447 11994
rect 3447 11942 3477 11994
rect 3501 11942 3511 11994
rect 3511 11942 3557 11994
rect 3581 11942 3627 11994
rect 3627 11942 3637 11994
rect 3661 11942 3691 11994
rect 3691 11942 3717 11994
rect 3421 11940 3477 11942
rect 3501 11940 3557 11942
rect 3581 11940 3637 11942
rect 3661 11940 3717 11942
rect 3422 11736 3478 11792
rect 3421 10906 3477 10908
rect 3501 10906 3557 10908
rect 3581 10906 3637 10908
rect 3661 10906 3717 10908
rect 3421 10854 3447 10906
rect 3447 10854 3477 10906
rect 3501 10854 3511 10906
rect 3511 10854 3557 10906
rect 3581 10854 3627 10906
rect 3627 10854 3637 10906
rect 3661 10854 3691 10906
rect 3691 10854 3717 10906
rect 3421 10852 3477 10854
rect 3501 10852 3557 10854
rect 3581 10852 3637 10854
rect 3661 10852 3717 10854
rect 3974 13268 3976 13288
rect 3976 13268 4028 13288
rect 4028 13268 4030 13288
rect 3974 13232 4030 13268
rect 3882 12688 3938 12744
rect 4066 12008 4122 12064
rect 4434 12552 4490 12608
rect 4710 14184 4766 14240
rect 4894 14184 4950 14240
rect 4710 13096 4766 13152
rect 3421 9818 3477 9820
rect 3501 9818 3557 9820
rect 3581 9818 3637 9820
rect 3661 9818 3717 9820
rect 3421 9766 3447 9818
rect 3447 9766 3477 9818
rect 3501 9766 3511 9818
rect 3511 9766 3557 9818
rect 3581 9766 3627 9818
rect 3627 9766 3637 9818
rect 3661 9766 3691 9818
rect 3691 9766 3717 9818
rect 3421 9764 3477 9766
rect 3501 9764 3557 9766
rect 3581 9764 3637 9766
rect 3661 9764 3717 9766
rect 3882 9560 3938 9616
rect 3421 8730 3477 8732
rect 3501 8730 3557 8732
rect 3581 8730 3637 8732
rect 3661 8730 3717 8732
rect 3421 8678 3447 8730
rect 3447 8678 3477 8730
rect 3501 8678 3511 8730
rect 3511 8678 3557 8730
rect 3581 8678 3627 8730
rect 3627 8678 3637 8730
rect 3661 8678 3691 8730
rect 3691 8678 3717 8730
rect 3421 8676 3477 8678
rect 3501 8676 3557 8678
rect 3581 8676 3637 8678
rect 3661 8676 3717 8678
rect 3698 8336 3754 8392
rect 4066 8880 4122 8936
rect 3421 7642 3477 7644
rect 3501 7642 3557 7644
rect 3581 7642 3637 7644
rect 3661 7642 3717 7644
rect 3421 7590 3447 7642
rect 3447 7590 3477 7642
rect 3501 7590 3511 7642
rect 3511 7590 3557 7642
rect 3581 7590 3627 7642
rect 3627 7590 3637 7642
rect 3661 7590 3691 7642
rect 3691 7590 3717 7642
rect 3421 7588 3477 7590
rect 3501 7588 3557 7590
rect 3581 7588 3637 7590
rect 3661 7588 3717 7590
rect 3146 7112 3202 7168
rect 3054 6840 3110 6896
rect 2962 4548 3018 4584
rect 2962 4528 2964 4548
rect 2964 4528 3016 4548
rect 3016 4528 3018 4548
rect 2962 4392 3018 4448
rect 3421 6554 3477 6556
rect 3501 6554 3557 6556
rect 3581 6554 3637 6556
rect 3661 6554 3717 6556
rect 3421 6502 3447 6554
rect 3447 6502 3477 6554
rect 3501 6502 3511 6554
rect 3511 6502 3557 6554
rect 3581 6502 3627 6554
rect 3627 6502 3637 6554
rect 3661 6502 3691 6554
rect 3691 6502 3717 6554
rect 3421 6500 3477 6502
rect 3501 6500 3557 6502
rect 3581 6500 3637 6502
rect 3661 6500 3717 6502
rect 4066 6740 4068 6760
rect 4068 6740 4120 6760
rect 4120 6740 4122 6760
rect 4066 6704 4122 6740
rect 3698 5652 3700 5672
rect 3700 5652 3752 5672
rect 3752 5652 3754 5672
rect 3698 5616 3754 5652
rect 3421 5466 3477 5468
rect 3501 5466 3557 5468
rect 3581 5466 3637 5468
rect 3661 5466 3717 5468
rect 3421 5414 3447 5466
rect 3447 5414 3477 5466
rect 3501 5414 3511 5466
rect 3511 5414 3557 5466
rect 3581 5414 3627 5466
rect 3627 5414 3637 5466
rect 3661 5414 3691 5466
rect 3691 5414 3717 5466
rect 3421 5412 3477 5414
rect 3501 5412 3557 5414
rect 3581 5412 3637 5414
rect 3661 5412 3717 5414
rect 3514 5228 3570 5264
rect 3514 5208 3516 5228
rect 3516 5208 3568 5228
rect 3568 5208 3570 5228
rect 3882 5344 3938 5400
rect 2778 448 2834 504
rect 3238 4392 3294 4448
rect 3421 4378 3477 4380
rect 3501 4378 3557 4380
rect 3581 4378 3637 4380
rect 3661 4378 3717 4380
rect 3421 4326 3447 4378
rect 3447 4326 3477 4378
rect 3501 4326 3511 4378
rect 3511 4326 3557 4378
rect 3581 4326 3627 4378
rect 3627 4326 3637 4378
rect 3661 4326 3691 4378
rect 3691 4326 3717 4378
rect 3421 4324 3477 4326
rect 3501 4324 3557 4326
rect 3581 4324 3637 4326
rect 3661 4324 3717 4326
rect 3422 3732 3478 3768
rect 3422 3712 3424 3732
rect 3424 3712 3476 3732
rect 3476 3712 3478 3732
rect 3606 3576 3662 3632
rect 3421 3290 3477 3292
rect 3501 3290 3557 3292
rect 3581 3290 3637 3292
rect 3661 3290 3717 3292
rect 3421 3238 3447 3290
rect 3447 3238 3477 3290
rect 3501 3238 3511 3290
rect 3511 3238 3557 3290
rect 3581 3238 3627 3290
rect 3627 3238 3637 3290
rect 3661 3238 3691 3290
rect 3691 3238 3717 3290
rect 3421 3236 3477 3238
rect 3501 3236 3557 3238
rect 3581 3236 3637 3238
rect 3661 3236 3717 3238
rect 3606 2488 3662 2544
rect 3514 2388 3516 2408
rect 3516 2388 3568 2408
rect 3568 2388 3570 2408
rect 3514 2352 3570 2388
rect 3421 2202 3477 2204
rect 3501 2202 3557 2204
rect 3581 2202 3637 2204
rect 3661 2202 3717 2204
rect 3421 2150 3447 2202
rect 3447 2150 3477 2202
rect 3501 2150 3511 2202
rect 3511 2150 3557 2202
rect 3581 2150 3627 2202
rect 3627 2150 3637 2202
rect 3661 2150 3691 2202
rect 3691 2150 3717 2202
rect 3421 2148 3477 2150
rect 3501 2148 3557 2150
rect 3581 2148 3637 2150
rect 3661 2148 3717 2150
rect 3882 2488 3938 2544
rect 4158 4936 4214 4992
rect 5078 12416 5134 12472
rect 5538 14592 5594 14648
rect 4986 9016 5042 9072
rect 5078 8508 5080 8528
rect 5080 8508 5132 8528
rect 5132 8508 5134 8528
rect 5078 8472 5134 8508
rect 4434 7656 4490 7712
rect 4710 7520 4766 7576
rect 4618 6432 4674 6488
rect 4434 5480 4490 5536
rect 4342 4256 4398 4312
rect 4342 3984 4398 4040
rect 4434 3304 4490 3360
rect 4618 6296 4674 6352
rect 4802 5752 4858 5808
rect 4710 5652 4712 5672
rect 4712 5652 4764 5672
rect 4764 5652 4766 5672
rect 4710 5616 4766 5652
rect 4710 3848 4766 3904
rect 5078 7928 5134 7984
rect 4986 4256 5042 4312
rect 5262 7248 5318 7304
rect 5886 15802 5942 15804
rect 5966 15802 6022 15804
rect 6046 15802 6102 15804
rect 6126 15802 6182 15804
rect 5886 15750 5912 15802
rect 5912 15750 5942 15802
rect 5966 15750 5976 15802
rect 5976 15750 6022 15802
rect 6046 15750 6092 15802
rect 6092 15750 6102 15802
rect 6126 15750 6156 15802
rect 6156 15750 6182 15802
rect 5886 15748 5942 15750
rect 5966 15748 6022 15750
rect 6046 15748 6102 15750
rect 6126 15748 6182 15750
rect 6182 15564 6238 15600
rect 6182 15544 6184 15564
rect 6184 15544 6236 15564
rect 6236 15544 6238 15564
rect 7010 15408 7066 15464
rect 6090 15020 6146 15056
rect 6090 15000 6092 15020
rect 6092 15000 6144 15020
rect 6144 15000 6146 15020
rect 5886 14714 5942 14716
rect 5966 14714 6022 14716
rect 6046 14714 6102 14716
rect 6126 14714 6182 14716
rect 5886 14662 5912 14714
rect 5912 14662 5942 14714
rect 5966 14662 5976 14714
rect 5976 14662 6022 14714
rect 6046 14662 6092 14714
rect 6092 14662 6102 14714
rect 6126 14662 6156 14714
rect 6156 14662 6182 14714
rect 5886 14660 5942 14662
rect 5966 14660 6022 14662
rect 6046 14660 6102 14662
rect 6126 14660 6182 14662
rect 5722 14320 5778 14376
rect 6274 14320 6330 14376
rect 5722 13368 5778 13424
rect 5886 13626 5942 13628
rect 5966 13626 6022 13628
rect 6046 13626 6102 13628
rect 6126 13626 6182 13628
rect 5886 13574 5912 13626
rect 5912 13574 5942 13626
rect 5966 13574 5976 13626
rect 5976 13574 6022 13626
rect 6046 13574 6092 13626
rect 6092 13574 6102 13626
rect 6126 13574 6156 13626
rect 6156 13574 6182 13626
rect 5886 13572 5942 13574
rect 5966 13572 6022 13574
rect 6046 13572 6102 13574
rect 6126 13572 6182 13574
rect 6182 12824 6238 12880
rect 5886 12538 5942 12540
rect 5966 12538 6022 12540
rect 6046 12538 6102 12540
rect 6126 12538 6182 12540
rect 5886 12486 5912 12538
rect 5912 12486 5942 12538
rect 5966 12486 5976 12538
rect 5976 12486 6022 12538
rect 6046 12486 6092 12538
rect 6092 12486 6102 12538
rect 6126 12486 6156 12538
rect 6156 12486 6182 12538
rect 5886 12484 5942 12486
rect 5966 12484 6022 12486
rect 6046 12484 6102 12486
rect 6126 12484 6182 12486
rect 5906 11872 5962 11928
rect 5814 11736 5870 11792
rect 5722 10920 5778 10976
rect 5886 11450 5942 11452
rect 5966 11450 6022 11452
rect 6046 11450 6102 11452
rect 6126 11450 6182 11452
rect 5886 11398 5912 11450
rect 5912 11398 5942 11450
rect 5966 11398 5976 11450
rect 5976 11398 6022 11450
rect 6046 11398 6092 11450
rect 6092 11398 6102 11450
rect 6126 11398 6156 11450
rect 6156 11398 6182 11450
rect 5886 11396 5942 11398
rect 5966 11396 6022 11398
rect 6046 11396 6102 11398
rect 6126 11396 6182 11398
rect 5886 10362 5942 10364
rect 5966 10362 6022 10364
rect 6046 10362 6102 10364
rect 6126 10362 6182 10364
rect 5886 10310 5912 10362
rect 5912 10310 5942 10362
rect 5966 10310 5976 10362
rect 5976 10310 6022 10362
rect 6046 10310 6092 10362
rect 6092 10310 6102 10362
rect 6126 10310 6156 10362
rect 6156 10310 6182 10362
rect 5886 10308 5942 10310
rect 5966 10308 6022 10310
rect 6046 10308 6102 10310
rect 6126 10308 6182 10310
rect 6366 13504 6422 13560
rect 6366 13232 6422 13288
rect 5354 4936 5410 4992
rect 5170 3984 5226 4040
rect 4066 2896 4122 2952
rect 4802 2896 4858 2952
rect 5170 2644 5226 2680
rect 5170 2624 5172 2644
rect 5172 2624 5224 2644
rect 5224 2624 5226 2644
rect 5446 3848 5502 3904
rect 5446 3732 5502 3768
rect 5446 3712 5448 3732
rect 5448 3712 5500 3732
rect 5500 3712 5502 3732
rect 6550 13232 6606 13288
rect 6550 12416 6606 12472
rect 7010 14592 7066 14648
rect 7010 14068 7066 14104
rect 7010 14048 7012 14068
rect 7012 14048 7064 14068
rect 7064 14048 7066 14068
rect 7470 15272 7526 15328
rect 7378 13912 7434 13968
rect 7102 13640 7158 13696
rect 6734 12552 6790 12608
rect 6550 10240 6606 10296
rect 6090 9424 6146 9480
rect 5886 9274 5942 9276
rect 5966 9274 6022 9276
rect 6046 9274 6102 9276
rect 6126 9274 6182 9276
rect 5886 9222 5912 9274
rect 5912 9222 5942 9274
rect 5966 9222 5976 9274
rect 5976 9222 6022 9274
rect 6046 9222 6092 9274
rect 6092 9222 6102 9274
rect 6126 9222 6156 9274
rect 6156 9222 6182 9274
rect 5886 9220 5942 9222
rect 5966 9220 6022 9222
rect 6046 9220 6102 9222
rect 6126 9220 6182 9222
rect 5886 8186 5942 8188
rect 5966 8186 6022 8188
rect 6046 8186 6102 8188
rect 6126 8186 6182 8188
rect 5886 8134 5912 8186
rect 5912 8134 5942 8186
rect 5966 8134 5976 8186
rect 5976 8134 6022 8186
rect 6046 8134 6092 8186
rect 6092 8134 6102 8186
rect 6126 8134 6156 8186
rect 6156 8134 6182 8186
rect 5886 8132 5942 8134
rect 5966 8132 6022 8134
rect 6046 8132 6102 8134
rect 6126 8132 6182 8134
rect 5722 7656 5778 7712
rect 6366 7520 6422 7576
rect 5722 7148 5724 7168
rect 5724 7148 5776 7168
rect 5776 7148 5778 7168
rect 5722 7112 5778 7148
rect 5630 6976 5686 7032
rect 5886 7098 5942 7100
rect 5966 7098 6022 7100
rect 6046 7098 6102 7100
rect 6126 7098 6182 7100
rect 5886 7046 5912 7098
rect 5912 7046 5942 7098
rect 5966 7046 5976 7098
rect 5976 7046 6022 7098
rect 6046 7046 6092 7098
rect 6092 7046 6102 7098
rect 6126 7046 6156 7098
rect 6156 7046 6182 7098
rect 5886 7044 5942 7046
rect 5966 7044 6022 7046
rect 6046 7044 6102 7046
rect 6126 7044 6182 7046
rect 6366 6976 6422 7032
rect 5722 5888 5778 5944
rect 5886 6010 5942 6012
rect 5966 6010 6022 6012
rect 6046 6010 6102 6012
rect 6126 6010 6182 6012
rect 5886 5958 5912 6010
rect 5912 5958 5942 6010
rect 5966 5958 5976 6010
rect 5976 5958 6022 6010
rect 6046 5958 6092 6010
rect 6092 5958 6102 6010
rect 6126 5958 6156 6010
rect 6156 5958 6182 6010
rect 5886 5956 5942 5958
rect 5966 5956 6022 5958
rect 6046 5956 6102 5958
rect 6126 5956 6182 5958
rect 5906 5616 5962 5672
rect 6274 5480 6330 5536
rect 5886 4922 5942 4924
rect 5966 4922 6022 4924
rect 6046 4922 6102 4924
rect 6126 4922 6182 4924
rect 5886 4870 5912 4922
rect 5912 4870 5942 4922
rect 5966 4870 5976 4922
rect 5976 4870 6022 4922
rect 6046 4870 6092 4922
rect 6092 4870 6102 4922
rect 6126 4870 6156 4922
rect 6156 4870 6182 4922
rect 5886 4868 5942 4870
rect 5966 4868 6022 4870
rect 6046 4868 6102 4870
rect 6126 4868 6182 4870
rect 6458 4800 6514 4856
rect 6366 3848 6422 3904
rect 5886 3834 5942 3836
rect 5966 3834 6022 3836
rect 6046 3834 6102 3836
rect 6126 3834 6182 3836
rect 5886 3782 5912 3834
rect 5912 3782 5942 3834
rect 5966 3782 5976 3834
rect 5976 3782 6022 3834
rect 6046 3782 6092 3834
rect 6092 3782 6102 3834
rect 6126 3782 6156 3834
rect 6156 3782 6182 3834
rect 5886 3780 5942 3782
rect 5966 3780 6022 3782
rect 6046 3780 6102 3782
rect 6126 3780 6182 3782
rect 6274 3732 6330 3768
rect 6274 3712 6276 3732
rect 6276 3712 6328 3732
rect 6328 3712 6330 3732
rect 6826 12416 6882 12472
rect 7194 12416 7250 12472
rect 7562 12552 7618 12608
rect 7470 11872 7526 11928
rect 7654 12416 7710 12472
rect 7470 11464 7526 11520
rect 7930 13912 7986 13968
rect 7838 13096 7894 13152
rect 7838 12008 7894 12064
rect 7930 11328 7986 11384
rect 7746 10648 7802 10704
rect 8666 15444 8668 15464
rect 8668 15444 8720 15464
rect 8720 15444 8722 15464
rect 8666 15408 8722 15444
rect 8352 15258 8408 15260
rect 8432 15258 8488 15260
rect 8512 15258 8568 15260
rect 8592 15258 8648 15260
rect 8352 15206 8378 15258
rect 8378 15206 8408 15258
rect 8432 15206 8442 15258
rect 8442 15206 8488 15258
rect 8512 15206 8558 15258
rect 8558 15206 8568 15258
rect 8592 15206 8622 15258
rect 8622 15206 8648 15258
rect 8352 15204 8408 15206
rect 8432 15204 8488 15206
rect 8512 15204 8568 15206
rect 8592 15204 8648 15206
rect 8114 14184 8170 14240
rect 8850 14864 8906 14920
rect 8352 14170 8408 14172
rect 8432 14170 8488 14172
rect 8512 14170 8568 14172
rect 8592 14170 8648 14172
rect 8352 14118 8378 14170
rect 8378 14118 8408 14170
rect 8432 14118 8442 14170
rect 8442 14118 8488 14170
rect 8512 14118 8558 14170
rect 8558 14118 8568 14170
rect 8592 14118 8622 14170
rect 8622 14118 8648 14170
rect 8352 14116 8408 14118
rect 8432 14116 8488 14118
rect 8512 14116 8568 14118
rect 8592 14116 8648 14118
rect 9310 15000 9366 15056
rect 8850 14456 8906 14512
rect 8352 13082 8408 13084
rect 8432 13082 8488 13084
rect 8512 13082 8568 13084
rect 8592 13082 8648 13084
rect 8352 13030 8378 13082
rect 8378 13030 8408 13082
rect 8432 13030 8442 13082
rect 8442 13030 8488 13082
rect 8512 13030 8558 13082
rect 8558 13030 8568 13082
rect 8592 13030 8622 13082
rect 8622 13030 8648 13082
rect 8352 13028 8408 13030
rect 8432 13028 8488 13030
rect 8512 13028 8568 13030
rect 8592 13028 8648 13030
rect 8298 12844 8354 12880
rect 8298 12824 8300 12844
rect 8300 12824 8352 12844
rect 8352 12824 8354 12844
rect 8574 12824 8630 12880
rect 8758 12960 8814 13016
rect 9402 14456 9458 14512
rect 9310 14048 9366 14104
rect 9126 13812 9128 13832
rect 9128 13812 9180 13832
rect 9180 13812 9182 13832
rect 9126 13776 9182 13812
rect 9402 13776 9458 13832
rect 9126 13096 9182 13152
rect 8758 12552 8814 12608
rect 9034 12552 9090 12608
rect 8352 11994 8408 11996
rect 8432 11994 8488 11996
rect 8512 11994 8568 11996
rect 8592 11994 8648 11996
rect 8352 11942 8378 11994
rect 8378 11942 8408 11994
rect 8432 11942 8442 11994
rect 8442 11942 8488 11994
rect 8512 11942 8558 11994
rect 8558 11942 8568 11994
rect 8592 11942 8622 11994
rect 8622 11942 8648 11994
rect 8352 11940 8408 11942
rect 8432 11940 8488 11942
rect 8512 11940 8568 11942
rect 8592 11940 8648 11942
rect 8022 10104 8078 10160
rect 6734 8608 6790 8664
rect 6734 8336 6790 8392
rect 5446 2644 5502 2680
rect 5446 2624 5448 2644
rect 5448 2624 5500 2644
rect 5500 2624 5502 2644
rect 5886 2746 5942 2748
rect 5966 2746 6022 2748
rect 6046 2746 6102 2748
rect 6126 2746 6182 2748
rect 5886 2694 5912 2746
rect 5912 2694 5942 2746
rect 5966 2694 5976 2746
rect 5976 2694 6022 2746
rect 6046 2694 6092 2746
rect 6092 2694 6102 2746
rect 6126 2694 6156 2746
rect 6156 2694 6182 2746
rect 5886 2692 5942 2694
rect 5966 2692 6022 2694
rect 6046 2692 6102 2694
rect 6126 2692 6182 2694
rect 6182 2508 6238 2544
rect 6182 2488 6184 2508
rect 6184 2488 6236 2508
rect 6236 2488 6238 2508
rect 6734 4800 6790 4856
rect 7010 5616 7066 5672
rect 7654 9560 7710 9616
rect 7470 9324 7472 9344
rect 7472 9324 7524 9344
rect 7524 9324 7526 9344
rect 7470 9288 7526 9324
rect 7286 7384 7342 7440
rect 7194 5888 7250 5944
rect 7286 5616 7342 5672
rect 7010 4936 7066 4992
rect 7102 3848 7158 3904
rect 7010 3576 7066 3632
rect 6734 3304 6790 3360
rect 6918 3304 6974 3360
rect 6734 2760 6790 2816
rect 8352 10906 8408 10908
rect 8432 10906 8488 10908
rect 8512 10906 8568 10908
rect 8592 10906 8648 10908
rect 8352 10854 8378 10906
rect 8378 10854 8408 10906
rect 8432 10854 8442 10906
rect 8442 10854 8488 10906
rect 8512 10854 8558 10906
rect 8558 10854 8568 10906
rect 8592 10854 8622 10906
rect 8622 10854 8648 10906
rect 8352 10852 8408 10854
rect 8432 10852 8488 10854
rect 8512 10852 8568 10854
rect 8592 10852 8648 10854
rect 8482 10376 8538 10432
rect 8352 9818 8408 9820
rect 8432 9818 8488 9820
rect 8512 9818 8568 9820
rect 8592 9818 8648 9820
rect 8352 9766 8378 9818
rect 8378 9766 8408 9818
rect 8432 9766 8442 9818
rect 8442 9766 8488 9818
rect 8512 9766 8558 9818
rect 8558 9766 8568 9818
rect 8592 9766 8622 9818
rect 8622 9766 8648 9818
rect 8352 9764 8408 9766
rect 8432 9764 8488 9766
rect 8512 9764 8568 9766
rect 8592 9764 8648 9766
rect 8114 9560 8170 9616
rect 7654 6024 7710 6080
rect 7470 4936 7526 4992
rect 7470 4392 7526 4448
rect 8114 9152 8170 9208
rect 8390 9444 8446 9480
rect 8390 9424 8392 9444
rect 8392 9424 8444 9444
rect 8444 9424 8446 9444
rect 8352 8730 8408 8732
rect 8432 8730 8488 8732
rect 8512 8730 8568 8732
rect 8592 8730 8648 8732
rect 8352 8678 8378 8730
rect 8378 8678 8408 8730
rect 8432 8678 8442 8730
rect 8442 8678 8488 8730
rect 8512 8678 8558 8730
rect 8558 8678 8568 8730
rect 8592 8678 8622 8730
rect 8622 8678 8648 8730
rect 8352 8676 8408 8678
rect 8432 8676 8488 8678
rect 8512 8676 8568 8678
rect 8592 8676 8648 8678
rect 9034 12416 9090 12472
rect 8758 11872 8814 11928
rect 8022 7420 8024 7440
rect 8024 7420 8076 7440
rect 8076 7420 8078 7440
rect 8022 7384 8078 7420
rect 8022 6432 8078 6488
rect 7838 5516 7840 5536
rect 7840 5516 7892 5536
rect 7892 5516 7894 5536
rect 7838 5480 7894 5516
rect 7746 5344 7802 5400
rect 8482 7928 8538 7984
rect 8352 7642 8408 7644
rect 8432 7642 8488 7644
rect 8512 7642 8568 7644
rect 8592 7642 8648 7644
rect 8352 7590 8378 7642
rect 8378 7590 8408 7642
rect 8432 7590 8442 7642
rect 8442 7590 8488 7642
rect 8512 7590 8558 7642
rect 8558 7590 8568 7642
rect 8592 7590 8622 7642
rect 8622 7590 8648 7642
rect 8352 7588 8408 7590
rect 8432 7588 8488 7590
rect 8512 7588 8568 7590
rect 8592 7588 8648 7590
rect 8352 6554 8408 6556
rect 8432 6554 8488 6556
rect 8512 6554 8568 6556
rect 8592 6554 8648 6556
rect 8352 6502 8378 6554
rect 8378 6502 8408 6554
rect 8432 6502 8442 6554
rect 8442 6502 8488 6554
rect 8512 6502 8558 6554
rect 8558 6502 8568 6554
rect 8592 6502 8622 6554
rect 8622 6502 8648 6554
rect 8352 6500 8408 6502
rect 8432 6500 8488 6502
rect 8512 6500 8568 6502
rect 8592 6500 8648 6502
rect 8574 5908 8630 5944
rect 8574 5888 8576 5908
rect 8576 5888 8628 5908
rect 8628 5888 8630 5908
rect 8352 5466 8408 5468
rect 8432 5466 8488 5468
rect 8512 5466 8568 5468
rect 8592 5466 8648 5468
rect 8352 5414 8378 5466
rect 8378 5414 8408 5466
rect 8432 5414 8442 5466
rect 8442 5414 8488 5466
rect 8512 5414 8558 5466
rect 8558 5414 8568 5466
rect 8592 5414 8622 5466
rect 8622 5414 8648 5466
rect 8352 5412 8408 5414
rect 8432 5412 8488 5414
rect 8512 5412 8568 5414
rect 8592 5412 8648 5414
rect 7746 4800 7802 4856
rect 7654 4392 7710 4448
rect 7654 3712 7710 3768
rect 7194 3168 7250 3224
rect 7102 1808 7158 1864
rect 7562 3168 7618 3224
rect 7746 2352 7802 2408
rect 8022 4120 8078 4176
rect 8352 4378 8408 4380
rect 8432 4378 8488 4380
rect 8512 4378 8568 4380
rect 8592 4378 8648 4380
rect 8352 4326 8378 4378
rect 8378 4326 8408 4378
rect 8432 4326 8442 4378
rect 8442 4326 8488 4378
rect 8512 4326 8558 4378
rect 8558 4326 8568 4378
rect 8592 4326 8622 4378
rect 8622 4326 8648 4378
rect 8352 4324 8408 4326
rect 8432 4324 8488 4326
rect 8512 4324 8568 4326
rect 8592 4324 8648 4326
rect 8352 3290 8408 3292
rect 8432 3290 8488 3292
rect 8512 3290 8568 3292
rect 8592 3290 8648 3292
rect 8352 3238 8378 3290
rect 8378 3238 8408 3290
rect 8432 3238 8442 3290
rect 8442 3238 8488 3290
rect 8512 3238 8558 3290
rect 8558 3238 8568 3290
rect 8592 3238 8622 3290
rect 8622 3238 8648 3290
rect 8352 3236 8408 3238
rect 8432 3236 8488 3238
rect 8512 3236 8568 3238
rect 8592 3236 8648 3238
rect 8850 11464 8906 11520
rect 8850 11092 8852 11112
rect 8852 11092 8904 11112
rect 8904 11092 8906 11112
rect 8850 11056 8906 11092
rect 8850 10956 8852 10976
rect 8852 10956 8904 10976
rect 8904 10956 8906 10976
rect 8850 10920 8906 10956
rect 9218 11872 9274 11928
rect 8850 9696 8906 9752
rect 8850 8628 8906 8664
rect 8850 8608 8852 8628
rect 8852 8608 8904 8628
rect 8904 8608 8906 8628
rect 9770 14476 9826 14512
rect 9770 14456 9772 14476
rect 9772 14456 9824 14476
rect 9824 14456 9826 14476
rect 9586 14048 9642 14104
rect 9402 12436 9458 12472
rect 9402 12416 9404 12436
rect 9404 12416 9456 12436
rect 9456 12416 9458 12436
rect 9402 12144 9458 12200
rect 9310 11056 9366 11112
rect 9310 9152 9366 9208
rect 9126 8780 9128 8800
rect 9128 8780 9180 8800
rect 9180 8780 9182 8800
rect 9126 8744 9182 8780
rect 9034 8200 9090 8256
rect 8850 7928 8906 7984
rect 8942 7520 8998 7576
rect 9034 6568 9090 6624
rect 8758 3168 8814 3224
rect 8206 2624 8262 2680
rect 8114 2488 8170 2544
rect 8114 2352 8170 2408
rect 8352 2202 8408 2204
rect 8432 2202 8488 2204
rect 8512 2202 8568 2204
rect 8592 2202 8648 2204
rect 8352 2150 8378 2202
rect 8378 2150 8408 2202
rect 8432 2150 8442 2202
rect 8442 2150 8488 2202
rect 8512 2150 8558 2202
rect 8558 2150 8568 2202
rect 8592 2150 8622 2202
rect 8622 2150 8648 2202
rect 8352 2148 8408 2150
rect 8432 2148 8488 2150
rect 8512 2148 8568 2150
rect 8592 2148 8648 2150
rect 7838 1944 7894 2000
rect 8758 2624 8814 2680
rect 9310 6976 9366 7032
rect 9586 12552 9642 12608
rect 9770 14184 9826 14240
rect 9862 13096 9918 13152
rect 9862 12416 9918 12472
rect 9770 12008 9826 12064
rect 10230 15408 10286 15464
rect 10782 15952 10838 16008
rect 10817 15802 10873 15804
rect 10897 15802 10953 15804
rect 10977 15802 11033 15804
rect 11057 15802 11113 15804
rect 10817 15750 10843 15802
rect 10843 15750 10873 15802
rect 10897 15750 10907 15802
rect 10907 15750 10953 15802
rect 10977 15750 11023 15802
rect 11023 15750 11033 15802
rect 11057 15750 11087 15802
rect 11087 15750 11113 15802
rect 10817 15748 10873 15750
rect 10897 15748 10953 15750
rect 10977 15748 11033 15750
rect 11057 15748 11113 15750
rect 9954 12144 10010 12200
rect 10046 12008 10102 12064
rect 10230 13096 10286 13152
rect 10598 14728 10654 14784
rect 10817 14714 10873 14716
rect 10897 14714 10953 14716
rect 10977 14714 11033 14716
rect 11057 14714 11113 14716
rect 10817 14662 10843 14714
rect 10843 14662 10873 14714
rect 10897 14662 10907 14714
rect 10907 14662 10953 14714
rect 10977 14662 11023 14714
rect 11023 14662 11033 14714
rect 11057 14662 11087 14714
rect 11087 14662 11113 14714
rect 10817 14660 10873 14662
rect 10897 14660 10953 14662
rect 10977 14660 11033 14662
rect 11057 14660 11113 14662
rect 10414 13776 10470 13832
rect 10230 9696 10286 9752
rect 10230 9560 10286 9616
rect 10046 8472 10102 8528
rect 9954 7384 10010 7440
rect 9954 6976 10010 7032
rect 10230 8064 10286 8120
rect 10414 12416 10470 12472
rect 10598 14184 10654 14240
rect 10817 13626 10873 13628
rect 10897 13626 10953 13628
rect 10977 13626 11033 13628
rect 11057 13626 11113 13628
rect 10817 13574 10843 13626
rect 10843 13574 10873 13626
rect 10897 13574 10907 13626
rect 10907 13574 10953 13626
rect 10977 13574 11023 13626
rect 11023 13574 11033 13626
rect 11057 13574 11087 13626
rect 11087 13574 11113 13626
rect 10817 13572 10873 13574
rect 10897 13572 10953 13574
rect 10977 13572 11033 13574
rect 11057 13572 11113 13574
rect 10782 12824 10838 12880
rect 10817 12538 10873 12540
rect 10897 12538 10953 12540
rect 10977 12538 11033 12540
rect 11057 12538 11113 12540
rect 10817 12486 10843 12538
rect 10843 12486 10873 12538
rect 10897 12486 10907 12538
rect 10907 12486 10953 12538
rect 10977 12486 11023 12538
rect 11023 12486 11033 12538
rect 11057 12486 11087 12538
rect 11087 12486 11113 12538
rect 10817 12484 10873 12486
rect 10897 12484 10953 12486
rect 10977 12484 11033 12486
rect 11057 12484 11113 12486
rect 10414 12144 10470 12200
rect 10506 12008 10562 12064
rect 10414 11736 10470 11792
rect 10414 11348 10470 11384
rect 10414 11328 10416 11348
rect 10416 11328 10468 11348
rect 10468 11328 10470 11348
rect 11058 12144 11114 12200
rect 10966 12044 10968 12064
rect 10968 12044 11020 12064
rect 11020 12044 11022 12064
rect 10966 12008 11022 12044
rect 11058 11872 11114 11928
rect 10874 11736 10930 11792
rect 10817 11450 10873 11452
rect 10897 11450 10953 11452
rect 10977 11450 11033 11452
rect 11057 11450 11113 11452
rect 10817 11398 10843 11450
rect 10843 11398 10873 11450
rect 10897 11398 10907 11450
rect 10907 11398 10953 11450
rect 10977 11398 11023 11450
rect 11023 11398 11033 11450
rect 11057 11398 11087 11450
rect 11087 11398 11113 11450
rect 10817 11396 10873 11398
rect 10897 11396 10953 11398
rect 10977 11396 11033 11398
rect 11057 11396 11113 11398
rect 11426 13912 11482 13968
rect 11334 13640 11390 13696
rect 11794 13776 11850 13832
rect 11334 13096 11390 13152
rect 11518 12824 11574 12880
rect 11426 12552 11482 12608
rect 11334 12416 11390 12472
rect 11150 10784 11206 10840
rect 10506 10376 10562 10432
rect 10817 10362 10873 10364
rect 10897 10362 10953 10364
rect 10977 10362 11033 10364
rect 11057 10362 11113 10364
rect 10817 10310 10843 10362
rect 10843 10310 10873 10362
rect 10897 10310 10907 10362
rect 10907 10310 10953 10362
rect 10977 10310 11023 10362
rect 11023 10310 11033 10362
rect 11057 10310 11087 10362
rect 11087 10310 11113 10362
rect 10817 10308 10873 10310
rect 10897 10308 10953 10310
rect 10977 10308 11033 10310
rect 11057 10308 11113 10310
rect 10598 10240 10654 10296
rect 10966 9716 11022 9752
rect 10966 9696 10968 9716
rect 10968 9696 11020 9716
rect 11020 9696 11022 9716
rect 11058 9424 11114 9480
rect 10817 9274 10873 9276
rect 10897 9274 10953 9276
rect 10977 9274 11033 9276
rect 11057 9274 11113 9276
rect 10817 9222 10843 9274
rect 10843 9222 10873 9274
rect 10897 9222 10907 9274
rect 10907 9222 10953 9274
rect 10977 9222 11023 9274
rect 11023 9222 11033 9274
rect 11057 9222 11087 9274
rect 11087 9222 11113 9274
rect 10817 9220 10873 9222
rect 10897 9220 10953 9222
rect 10977 9220 11033 9222
rect 11057 9220 11113 9222
rect 10782 8880 10838 8936
rect 10690 8508 10692 8528
rect 10692 8508 10744 8528
rect 10744 8508 10746 8528
rect 10690 8472 10746 8508
rect 11518 10784 11574 10840
rect 11242 9172 11298 9208
rect 11426 9424 11482 9480
rect 11242 9152 11244 9172
rect 11244 9152 11296 9172
rect 11296 9152 11298 9172
rect 10874 8472 10930 8528
rect 10414 8064 10470 8120
rect 10230 7656 10286 7712
rect 10506 7520 10562 7576
rect 10230 6976 10286 7032
rect 9586 5616 9642 5672
rect 9310 4936 9366 4992
rect 9126 4256 9182 4312
rect 9310 4392 9366 4448
rect 9126 3440 9182 3496
rect 9126 2896 9182 2952
rect 9494 4120 9550 4176
rect 9126 2216 9182 2272
rect 9862 4256 9918 4312
rect 9770 4120 9826 4176
rect 9678 3168 9734 3224
rect 9678 1944 9734 2000
rect 9954 3168 10010 3224
rect 10230 5752 10286 5808
rect 10414 7112 10470 7168
rect 11702 13368 11758 13424
rect 11702 13232 11758 13288
rect 12070 14592 12126 14648
rect 11978 14456 12034 14512
rect 12346 14320 12402 14376
rect 11978 13368 12034 13424
rect 12162 13268 12164 13288
rect 12164 13268 12216 13288
rect 12216 13268 12218 13288
rect 12162 13232 12218 13268
rect 12070 11872 12126 11928
rect 11978 10684 11980 10704
rect 11980 10684 12032 10704
rect 12032 10684 12034 10704
rect 11978 10648 12034 10684
rect 11702 10412 11704 10432
rect 11704 10412 11756 10432
rect 11756 10412 11758 10432
rect 11702 10376 11758 10412
rect 12438 13776 12494 13832
rect 12346 13640 12402 13696
rect 12346 13368 12402 13424
rect 12714 14184 12770 14240
rect 12438 12688 12494 12744
rect 13358 15408 13414 15464
rect 13282 15258 13338 15260
rect 13362 15258 13418 15260
rect 13442 15258 13498 15260
rect 13522 15258 13578 15260
rect 13282 15206 13308 15258
rect 13308 15206 13338 15258
rect 13362 15206 13372 15258
rect 13372 15206 13418 15258
rect 13442 15206 13488 15258
rect 13488 15206 13498 15258
rect 13522 15206 13552 15258
rect 13552 15206 13578 15258
rect 13282 15204 13338 15206
rect 13362 15204 13418 15206
rect 13442 15204 13498 15206
rect 13522 15204 13578 15206
rect 12898 12824 12954 12880
rect 12898 12552 12954 12608
rect 12714 12144 12770 12200
rect 12714 11328 12770 11384
rect 12898 12416 12954 12472
rect 12898 11872 12954 11928
rect 12070 9832 12126 9888
rect 11886 9288 11942 9344
rect 11702 9152 11758 9208
rect 11794 8880 11850 8936
rect 10817 8186 10873 8188
rect 10897 8186 10953 8188
rect 10977 8186 11033 8188
rect 11057 8186 11113 8188
rect 10817 8134 10843 8186
rect 10843 8134 10873 8186
rect 10897 8134 10907 8186
rect 10907 8134 10953 8186
rect 10977 8134 11023 8186
rect 11023 8134 11033 8186
rect 11057 8134 11087 8186
rect 11087 8134 11113 8186
rect 10817 8132 10873 8134
rect 10897 8132 10953 8134
rect 10977 8132 11033 8134
rect 11057 8132 11113 8134
rect 11242 8064 11298 8120
rect 10782 7520 10838 7576
rect 10690 7384 10746 7440
rect 11058 7384 11114 7440
rect 10782 7248 10838 7304
rect 10966 7284 10968 7304
rect 10968 7284 11020 7304
rect 11020 7284 11022 7304
rect 10966 7248 11022 7284
rect 11334 7520 11390 7576
rect 10817 7098 10873 7100
rect 10897 7098 10953 7100
rect 10977 7098 11033 7100
rect 11057 7098 11113 7100
rect 10817 7046 10843 7098
rect 10843 7046 10873 7098
rect 10897 7046 10907 7098
rect 10907 7046 10953 7098
rect 10977 7046 11023 7098
rect 11023 7046 11033 7098
rect 11057 7046 11087 7098
rect 11087 7046 11113 7098
rect 10817 7044 10873 7046
rect 10897 7044 10953 7046
rect 10977 7044 11033 7046
rect 11057 7044 11113 7046
rect 11334 7148 11336 7168
rect 11336 7148 11388 7168
rect 11388 7148 11390 7168
rect 11334 7112 11390 7148
rect 10817 6010 10873 6012
rect 10897 6010 10953 6012
rect 10977 6010 11033 6012
rect 11057 6010 11113 6012
rect 10817 5958 10843 6010
rect 10843 5958 10873 6010
rect 10897 5958 10907 6010
rect 10907 5958 10953 6010
rect 10977 5958 11023 6010
rect 11023 5958 11033 6010
rect 11057 5958 11087 6010
rect 11087 5958 11113 6010
rect 10817 5956 10873 5958
rect 10897 5956 10953 5958
rect 10977 5956 11033 5958
rect 11057 5956 11113 5958
rect 11058 5652 11060 5672
rect 11060 5652 11112 5672
rect 11112 5652 11114 5672
rect 11058 5616 11114 5652
rect 11242 5616 11298 5672
rect 10817 4922 10873 4924
rect 10897 4922 10953 4924
rect 10977 4922 11033 4924
rect 11057 4922 11113 4924
rect 10817 4870 10843 4922
rect 10843 4870 10873 4922
rect 10897 4870 10907 4922
rect 10907 4870 10953 4922
rect 10977 4870 11023 4922
rect 11023 4870 11033 4922
rect 11057 4870 11087 4922
rect 11087 4870 11113 4922
rect 10817 4868 10873 4870
rect 10897 4868 10953 4870
rect 10977 4868 11033 4870
rect 11057 4868 11113 4870
rect 10414 4392 10470 4448
rect 10230 3712 10286 3768
rect 10414 2624 10470 2680
rect 11610 7384 11666 7440
rect 11518 6024 11574 6080
rect 10782 4020 10784 4040
rect 10784 4020 10836 4040
rect 10836 4020 10838 4040
rect 10782 3984 10838 4020
rect 10817 3834 10873 3836
rect 10897 3834 10953 3836
rect 10977 3834 11033 3836
rect 11057 3834 11113 3836
rect 10817 3782 10843 3834
rect 10843 3782 10873 3834
rect 10897 3782 10907 3834
rect 10907 3782 10953 3834
rect 10977 3782 11023 3834
rect 11023 3782 11033 3834
rect 11057 3782 11087 3834
rect 11087 3782 11113 3834
rect 10817 3780 10873 3782
rect 10897 3780 10953 3782
rect 10977 3780 11033 3782
rect 11057 3780 11113 3782
rect 10690 2896 10746 2952
rect 10817 2746 10873 2748
rect 10897 2746 10953 2748
rect 10977 2746 11033 2748
rect 11057 2746 11113 2748
rect 10817 2694 10843 2746
rect 10843 2694 10873 2746
rect 10897 2694 10907 2746
rect 10907 2694 10953 2746
rect 10977 2694 11023 2746
rect 11023 2694 11033 2746
rect 11057 2694 11087 2746
rect 11087 2694 11113 2746
rect 10817 2692 10873 2694
rect 10897 2692 10953 2694
rect 10977 2692 11033 2694
rect 11057 2692 11113 2694
rect 9954 2080 10010 2136
rect 9862 1672 9918 1728
rect 11518 4936 11574 4992
rect 12806 10920 12862 10976
rect 13282 14170 13338 14172
rect 13362 14170 13418 14172
rect 13442 14170 13498 14172
rect 13522 14170 13578 14172
rect 13282 14118 13308 14170
rect 13308 14118 13338 14170
rect 13362 14118 13372 14170
rect 13372 14118 13418 14170
rect 13442 14118 13488 14170
rect 13488 14118 13498 14170
rect 13522 14118 13552 14170
rect 13552 14118 13578 14170
rect 13282 14116 13338 14118
rect 13362 14116 13418 14118
rect 13442 14116 13498 14118
rect 13522 14116 13578 14118
rect 13282 13082 13338 13084
rect 13362 13082 13418 13084
rect 13442 13082 13498 13084
rect 13522 13082 13578 13084
rect 13282 13030 13308 13082
rect 13308 13030 13338 13082
rect 13362 13030 13372 13082
rect 13372 13030 13418 13082
rect 13442 13030 13488 13082
rect 13488 13030 13498 13082
rect 13522 13030 13552 13082
rect 13552 13030 13578 13082
rect 13282 13028 13338 13030
rect 13362 13028 13418 13030
rect 13442 13028 13498 13030
rect 13522 13028 13578 13030
rect 13174 12824 13230 12880
rect 13174 12688 13230 12744
rect 13282 11994 13338 11996
rect 13362 11994 13418 11996
rect 13442 11994 13498 11996
rect 13522 11994 13578 11996
rect 13282 11942 13308 11994
rect 13308 11942 13338 11994
rect 13362 11942 13372 11994
rect 13372 11942 13418 11994
rect 13442 11942 13488 11994
rect 13488 11942 13498 11994
rect 13522 11942 13552 11994
rect 13552 11942 13578 11994
rect 13282 11940 13338 11942
rect 13362 11940 13418 11942
rect 13442 11940 13498 11942
rect 13522 11940 13578 11942
rect 13266 11736 13322 11792
rect 13174 11192 13230 11248
rect 13450 11600 13506 11656
rect 13542 11192 13598 11248
rect 14002 15000 14058 15056
rect 14278 14864 14334 14920
rect 13818 12280 13874 12336
rect 13634 11056 13690 11112
rect 13282 10906 13338 10908
rect 13362 10906 13418 10908
rect 13442 10906 13498 10908
rect 13522 10906 13578 10908
rect 13282 10854 13308 10906
rect 13308 10854 13338 10906
rect 13362 10854 13372 10906
rect 13372 10854 13418 10906
rect 13442 10854 13488 10906
rect 13488 10854 13498 10906
rect 13522 10854 13552 10906
rect 13552 10854 13578 10906
rect 13282 10852 13338 10854
rect 13362 10852 13418 10854
rect 13442 10852 13498 10854
rect 13522 10852 13578 10854
rect 13542 10648 13598 10704
rect 12806 8608 12862 8664
rect 12530 8472 12586 8528
rect 12898 8200 12954 8256
rect 11794 6296 11850 6352
rect 12162 7384 12218 7440
rect 12438 7384 12494 7440
rect 12254 7248 12310 7304
rect 12162 6976 12218 7032
rect 12346 6568 12402 6624
rect 12070 6296 12126 6352
rect 11978 5480 12034 5536
rect 11702 4820 11758 4856
rect 11702 4800 11704 4820
rect 11704 4800 11756 4820
rect 11756 4800 11758 4820
rect 11794 4392 11850 4448
rect 11794 4256 11850 4312
rect 10690 1536 10746 1592
rect 11518 3848 11574 3904
rect 11702 3848 11758 3904
rect 11978 4936 12034 4992
rect 12070 4800 12126 4856
rect 11978 3712 12034 3768
rect 12254 6296 12310 6352
rect 12254 6024 12310 6080
rect 12622 7284 12624 7304
rect 12624 7284 12676 7304
rect 12676 7284 12678 7304
rect 12622 7248 12678 7284
rect 12530 6840 12586 6896
rect 12530 6024 12586 6080
rect 12438 5636 12494 5672
rect 12438 5616 12440 5636
rect 12440 5616 12492 5636
rect 12492 5616 12494 5636
rect 12714 6976 12770 7032
rect 12714 6840 12770 6896
rect 12898 7656 12954 7712
rect 13174 10376 13230 10432
rect 13726 10920 13782 10976
rect 13282 9818 13338 9820
rect 13362 9818 13418 9820
rect 13442 9818 13498 9820
rect 13522 9818 13578 9820
rect 13282 9766 13308 9818
rect 13308 9766 13338 9818
rect 13362 9766 13372 9818
rect 13372 9766 13418 9818
rect 13442 9766 13488 9818
rect 13488 9766 13498 9818
rect 13522 9766 13552 9818
rect 13552 9766 13578 9818
rect 13282 9764 13338 9766
rect 13362 9764 13418 9766
rect 13442 9764 13498 9766
rect 13522 9764 13578 9766
rect 13266 9324 13268 9344
rect 13268 9324 13320 9344
rect 13320 9324 13322 9344
rect 13266 9288 13322 9324
rect 13634 9424 13690 9480
rect 13450 9152 13506 9208
rect 13818 10532 13874 10568
rect 13818 10512 13820 10532
rect 13820 10512 13872 10532
rect 13872 10512 13874 10532
rect 13818 9560 13874 9616
rect 13282 8730 13338 8732
rect 13362 8730 13418 8732
rect 13442 8730 13498 8732
rect 13522 8730 13578 8732
rect 13282 8678 13308 8730
rect 13308 8678 13338 8730
rect 13362 8678 13372 8730
rect 13372 8678 13418 8730
rect 13442 8678 13488 8730
rect 13488 8678 13498 8730
rect 13522 8678 13552 8730
rect 13552 8678 13578 8730
rect 13282 8676 13338 8678
rect 13362 8676 13418 8678
rect 13442 8676 13498 8678
rect 13522 8676 13578 8678
rect 13082 7928 13138 7984
rect 13450 7928 13506 7984
rect 12990 7112 13046 7168
rect 12990 6976 13046 7032
rect 12806 6160 12862 6216
rect 12806 5888 12862 5944
rect 12898 5752 12954 5808
rect 12622 5344 12678 5400
rect 12254 4392 12310 4448
rect 12530 3984 12586 4040
rect 12254 3848 12310 3904
rect 11610 3032 11666 3088
rect 12438 3576 12494 3632
rect 11886 3304 11942 3360
rect 12254 3304 12310 3360
rect 11518 2624 11574 2680
rect 11242 1400 11298 1456
rect 11886 3032 11942 3088
rect 11794 2508 11850 2544
rect 11794 2488 11796 2508
rect 11796 2488 11848 2508
rect 11848 2488 11850 2508
rect 12070 2080 12126 2136
rect 12254 2896 12310 2952
rect 12438 3304 12494 3360
rect 12898 5480 12954 5536
rect 13282 7642 13338 7644
rect 13362 7642 13418 7644
rect 13442 7642 13498 7644
rect 13522 7642 13578 7644
rect 13282 7590 13308 7642
rect 13308 7590 13338 7642
rect 13362 7590 13372 7642
rect 13372 7590 13418 7642
rect 13442 7590 13488 7642
rect 13488 7590 13498 7642
rect 13522 7590 13552 7642
rect 13552 7590 13578 7642
rect 13282 7588 13338 7590
rect 13362 7588 13418 7590
rect 13442 7588 13498 7590
rect 13522 7588 13578 7590
rect 13358 7112 13414 7168
rect 13282 6554 13338 6556
rect 13362 6554 13418 6556
rect 13442 6554 13498 6556
rect 13522 6554 13578 6556
rect 13282 6502 13308 6554
rect 13308 6502 13338 6554
rect 13362 6502 13372 6554
rect 13372 6502 13418 6554
rect 13442 6502 13488 6554
rect 13488 6502 13498 6554
rect 13522 6502 13552 6554
rect 13552 6502 13578 6554
rect 13282 6500 13338 6502
rect 13362 6500 13418 6502
rect 13442 6500 13498 6502
rect 13522 6500 13578 6502
rect 14094 11056 14150 11112
rect 13726 8336 13782 8392
rect 13450 6160 13506 6216
rect 12990 5344 13046 5400
rect 12898 5072 12954 5128
rect 12990 4564 12992 4584
rect 12992 4564 13044 4584
rect 13044 4564 13046 4584
rect 12990 4528 13046 4564
rect 12898 4392 12954 4448
rect 13282 5466 13338 5468
rect 13362 5466 13418 5468
rect 13442 5466 13498 5468
rect 13522 5466 13578 5468
rect 13282 5414 13308 5466
rect 13308 5414 13338 5466
rect 13362 5414 13372 5466
rect 13372 5414 13418 5466
rect 13442 5414 13488 5466
rect 13488 5414 13498 5466
rect 13522 5414 13552 5466
rect 13552 5414 13578 5466
rect 13282 5412 13338 5414
rect 13362 5412 13418 5414
rect 13442 5412 13498 5414
rect 13522 5412 13578 5414
rect 13542 4684 13598 4720
rect 13542 4664 13544 4684
rect 13544 4664 13596 4684
rect 13596 4664 13598 4684
rect 13282 4378 13338 4380
rect 13362 4378 13418 4380
rect 13442 4378 13498 4380
rect 13522 4378 13578 4380
rect 13282 4326 13308 4378
rect 13308 4326 13338 4378
rect 13362 4326 13372 4378
rect 13372 4326 13418 4378
rect 13442 4326 13488 4378
rect 13488 4326 13498 4378
rect 13522 4326 13552 4378
rect 13552 4326 13578 4378
rect 13282 4324 13338 4326
rect 13362 4324 13418 4326
rect 13442 4324 13498 4326
rect 13522 4324 13578 4326
rect 13266 3712 13322 3768
rect 13174 3596 13230 3632
rect 13174 3576 13176 3596
rect 13176 3576 13228 3596
rect 13228 3576 13230 3596
rect 14186 10004 14188 10024
rect 14188 10004 14240 10024
rect 14240 10004 14242 10024
rect 14186 9968 14242 10004
rect 14094 8336 14150 8392
rect 13910 6180 13966 6216
rect 13910 6160 13912 6180
rect 13912 6160 13964 6180
rect 13964 6160 13966 6180
rect 13818 5616 13874 5672
rect 14094 6296 14150 6352
rect 13726 4800 13782 4856
rect 13726 3884 13728 3904
rect 13728 3884 13780 3904
rect 13780 3884 13782 3904
rect 13726 3848 13782 3884
rect 13634 3440 13690 3496
rect 13282 3290 13338 3292
rect 13362 3290 13418 3292
rect 13442 3290 13498 3292
rect 13522 3290 13578 3292
rect 13282 3238 13308 3290
rect 13308 3238 13338 3290
rect 13362 3238 13372 3290
rect 13372 3238 13418 3290
rect 13442 3238 13488 3290
rect 13488 3238 13498 3290
rect 13522 3238 13552 3290
rect 13552 3238 13578 3290
rect 13282 3236 13338 3238
rect 13362 3236 13418 3238
rect 13442 3236 13498 3238
rect 13522 3236 13578 3238
rect 13266 3068 13268 3088
rect 13268 3068 13320 3088
rect 13320 3068 13322 3088
rect 13266 3032 13322 3068
rect 13450 3032 13506 3088
rect 14002 4936 14058 4992
rect 13910 4020 13912 4040
rect 13912 4020 13964 4040
rect 13964 4020 13966 4040
rect 13910 3984 13966 4020
rect 13174 2508 13230 2544
rect 13174 2488 13176 2508
rect 13176 2488 13228 2508
rect 13228 2488 13230 2508
rect 13450 2624 13506 2680
rect 13282 2202 13338 2204
rect 13362 2202 13418 2204
rect 13442 2202 13498 2204
rect 13522 2202 13578 2204
rect 13282 2150 13308 2202
rect 13308 2150 13338 2202
rect 13362 2150 13372 2202
rect 13372 2150 13418 2202
rect 13442 2150 13488 2202
rect 13488 2150 13498 2202
rect 13522 2150 13552 2202
rect 13552 2150 13578 2202
rect 13282 2148 13338 2150
rect 13362 2148 13418 2150
rect 13442 2148 13498 2150
rect 13522 2148 13578 2150
rect 14186 2896 14242 2952
rect 14462 10104 14518 10160
rect 14830 11464 14886 11520
rect 14554 8356 14610 8392
rect 14554 8336 14556 8356
rect 14556 8336 14608 8356
rect 14608 8336 14610 8356
rect 14646 4800 14702 4856
rect 14462 3712 14518 3768
rect 14554 2352 14610 2408
rect 15290 13232 15346 13288
rect 15014 9560 15070 9616
rect 15198 10376 15254 10432
rect 15106 7792 15162 7848
rect 15198 6860 15254 6896
rect 15198 6840 15200 6860
rect 15200 6840 15252 6860
rect 15252 6840 15254 6860
rect 15014 6160 15070 6216
rect 15474 9016 15530 9072
rect 15382 8880 15438 8936
rect 15014 4120 15070 4176
rect 15014 3848 15070 3904
rect 15014 1944 15070 2000
rect 14738 1672 14794 1728
rect 15382 3032 15438 3088
rect 15934 2760 15990 2816
<< metal3 >>
rect 0 17370 480 17400
rect 3969 17370 4035 17373
rect 0 17368 4035 17370
rect 0 17312 3974 17368
rect 4030 17312 4035 17368
rect 0 17310 4035 17312
rect 0 17280 480 17310
rect 3969 17307 4035 17310
rect 0 16282 480 16312
rect 2957 16282 3023 16285
rect 0 16280 3023 16282
rect 0 16224 2962 16280
rect 3018 16224 3023 16280
rect 0 16222 3023 16224
rect 0 16192 480 16222
rect 2957 16219 3023 16222
rect 10174 15948 10180 16012
rect 10244 16010 10250 16012
rect 10777 16010 10843 16013
rect 10244 16008 10843 16010
rect 10244 15952 10782 16008
rect 10838 15952 10843 16008
rect 10244 15950 10843 15952
rect 10244 15948 10250 15950
rect 10777 15947 10843 15950
rect 5874 15808 6194 15809
rect 5874 15744 5882 15808
rect 5946 15744 5962 15808
rect 6026 15744 6042 15808
rect 6106 15744 6122 15808
rect 6186 15744 6194 15808
rect 5874 15743 6194 15744
rect 10805 15808 11125 15809
rect 10805 15744 10813 15808
rect 10877 15744 10893 15808
rect 10957 15744 10973 15808
rect 11037 15744 11053 15808
rect 11117 15744 11125 15808
rect 10805 15743 11125 15744
rect 6177 15602 6243 15605
rect 12566 15602 12572 15604
rect 6177 15600 12572 15602
rect 6177 15544 6182 15600
rect 6238 15544 12572 15600
rect 6177 15542 12572 15544
rect 6177 15539 6243 15542
rect 12566 15540 12572 15542
rect 12636 15540 12642 15604
rect 7005 15466 7071 15469
rect 8661 15466 8727 15469
rect 7005 15464 8727 15466
rect 7005 15408 7010 15464
rect 7066 15408 8666 15464
rect 8722 15408 8727 15464
rect 7005 15406 8727 15408
rect 7005 15403 7071 15406
rect 8661 15403 8727 15406
rect 10225 15466 10291 15469
rect 12934 15466 12940 15468
rect 10225 15464 12940 15466
rect 10225 15408 10230 15464
rect 10286 15408 12940 15464
rect 10225 15406 12940 15408
rect 10225 15403 10291 15406
rect 12934 15404 12940 15406
rect 13004 15466 13010 15468
rect 13353 15466 13419 15469
rect 13004 15464 13419 15466
rect 13004 15408 13358 15464
rect 13414 15408 13419 15464
rect 13004 15406 13419 15408
rect 13004 15404 13010 15406
rect 13353 15403 13419 15406
rect 7465 15332 7531 15333
rect 7414 15330 7420 15332
rect 7374 15270 7420 15330
rect 7484 15328 7531 15332
rect 7526 15272 7531 15328
rect 7414 15268 7420 15270
rect 7484 15268 7531 15272
rect 7465 15267 7531 15268
rect 3409 15264 3729 15265
rect 0 15194 480 15224
rect 3409 15200 3417 15264
rect 3481 15200 3497 15264
rect 3561 15200 3577 15264
rect 3641 15200 3657 15264
rect 3721 15200 3729 15264
rect 3409 15199 3729 15200
rect 8340 15264 8660 15265
rect 8340 15200 8348 15264
rect 8412 15200 8428 15264
rect 8492 15200 8508 15264
rect 8572 15200 8588 15264
rect 8652 15200 8660 15264
rect 8340 15199 8660 15200
rect 13270 15264 13590 15265
rect 13270 15200 13278 15264
rect 13342 15200 13358 15264
rect 13422 15200 13438 15264
rect 13502 15200 13518 15264
rect 13582 15200 13590 15264
rect 13270 15199 13590 15200
rect 2865 15194 2931 15197
rect 0 15192 2931 15194
rect 0 15136 2870 15192
rect 2926 15136 2931 15192
rect 0 15134 2931 15136
rect 0 15104 480 15134
rect 2865 15131 2931 15134
rect 3926 15134 6562 15194
rect 2313 15058 2379 15061
rect 3141 15058 3207 15061
rect 3926 15058 3986 15134
rect 2313 15056 3207 15058
rect 2313 15000 2318 15056
rect 2374 15000 3146 15056
rect 3202 15000 3207 15056
rect 2313 14998 3207 15000
rect 2313 14995 2379 14998
rect 3141 14995 3207 14998
rect 3558 14998 3986 15058
rect 6085 15058 6151 15061
rect 6310 15058 6316 15060
rect 6085 15056 6316 15058
rect 6085 15000 6090 15056
rect 6146 15000 6316 15056
rect 6085 14998 6316 15000
rect 2221 14922 2287 14925
rect 3558 14922 3618 14998
rect 6085 14995 6151 14998
rect 6310 14996 6316 14998
rect 6380 14996 6386 15060
rect 6502 15058 6562 15134
rect 9305 15058 9371 15061
rect 6502 15056 9371 15058
rect 6502 15000 9310 15056
rect 9366 15000 9371 15056
rect 6502 14998 9371 15000
rect 9305 14995 9371 14998
rect 13997 15058 14063 15061
rect 16520 15058 17000 15088
rect 13997 15056 17000 15058
rect 13997 15000 14002 15056
rect 14058 15000 17000 15056
rect 13997 14998 17000 15000
rect 13997 14995 14063 14998
rect 16520 14968 17000 14998
rect 2221 14920 3618 14922
rect 2221 14864 2226 14920
rect 2282 14864 3618 14920
rect 2221 14862 3618 14864
rect 3693 14922 3759 14925
rect 8845 14922 8911 14925
rect 14273 14922 14339 14925
rect 3693 14920 8770 14922
rect 3693 14864 3698 14920
rect 3754 14864 8770 14920
rect 3693 14862 8770 14864
rect 2221 14859 2287 14862
rect 3693 14859 3759 14862
rect 5874 14720 6194 14721
rect 5874 14656 5882 14720
rect 5946 14656 5962 14720
rect 6026 14656 6042 14720
rect 6106 14656 6122 14720
rect 6186 14656 6194 14720
rect 5874 14655 6194 14656
rect 3182 14588 3188 14652
rect 3252 14650 3258 14652
rect 5533 14650 5599 14653
rect 3252 14648 5780 14650
rect 3252 14592 5538 14648
rect 5594 14592 5780 14648
rect 3252 14590 5780 14592
rect 3252 14588 3258 14590
rect 5533 14587 5599 14590
rect 5720 14514 5780 14590
rect 6678 14588 6684 14652
rect 6748 14650 6754 14652
rect 7005 14650 7071 14653
rect 6748 14648 7071 14650
rect 6748 14592 7010 14648
rect 7066 14592 7071 14648
rect 6748 14590 7071 14592
rect 8710 14650 8770 14862
rect 8845 14920 14339 14922
rect 8845 14864 8850 14920
rect 8906 14864 14278 14920
rect 14334 14864 14339 14920
rect 8845 14862 14339 14864
rect 8845 14859 8911 14862
rect 14273 14859 14339 14862
rect 9070 14724 9076 14788
rect 9140 14786 9146 14788
rect 10593 14786 10659 14789
rect 9140 14784 10659 14786
rect 9140 14728 10598 14784
rect 10654 14728 10659 14784
rect 9140 14726 10659 14728
rect 9140 14724 9146 14726
rect 10593 14723 10659 14726
rect 10805 14720 11125 14721
rect 10805 14656 10813 14720
rect 10877 14656 10893 14720
rect 10957 14656 10973 14720
rect 11037 14656 11053 14720
rect 11117 14656 11125 14720
rect 10805 14655 11125 14656
rect 8710 14590 10610 14650
rect 6748 14588 6754 14590
rect 7005 14587 7071 14590
rect 8845 14514 8911 14517
rect 9397 14514 9463 14517
rect 9765 14516 9831 14517
rect 9765 14514 9812 14516
rect 5720 14512 9463 14514
rect 5720 14456 8850 14512
rect 8906 14456 9402 14512
rect 9458 14456 9463 14512
rect 5720 14454 9463 14456
rect 9720 14512 9812 14514
rect 9720 14456 9770 14512
rect 9720 14454 9812 14456
rect 8845 14451 8911 14454
rect 9397 14451 9463 14454
rect 9765 14452 9812 14454
rect 9876 14452 9882 14516
rect 10550 14514 10610 14590
rect 11462 14588 11468 14652
rect 11532 14650 11538 14652
rect 12065 14650 12131 14653
rect 11532 14648 12131 14650
rect 11532 14592 12070 14648
rect 12126 14592 12131 14648
rect 11532 14590 12131 14592
rect 11532 14588 11538 14590
rect 12065 14587 12131 14590
rect 11973 14514 12039 14517
rect 10550 14512 12039 14514
rect 10550 14456 11978 14512
rect 12034 14456 12039 14512
rect 10550 14454 12039 14456
rect 9765 14451 9831 14452
rect 11973 14451 12039 14454
rect 5574 14316 5580 14380
rect 5644 14378 5650 14380
rect 5717 14378 5783 14381
rect 5644 14376 5783 14378
rect 5644 14320 5722 14376
rect 5778 14320 5783 14376
rect 5644 14318 5783 14320
rect 5644 14316 5650 14318
rect 5717 14315 5783 14318
rect 6269 14378 6335 14381
rect 12341 14378 12407 14381
rect 6269 14376 12407 14378
rect 6269 14320 6274 14376
rect 6330 14320 12346 14376
rect 12402 14320 12407 14376
rect 6269 14318 12407 14320
rect 6269 14315 6335 14318
rect 12341 14315 12407 14318
rect 4705 14242 4771 14245
rect 4889 14242 4955 14245
rect 8109 14242 8175 14245
rect 4705 14240 8175 14242
rect 4705 14184 4710 14240
rect 4766 14184 4894 14240
rect 4950 14184 8114 14240
rect 8170 14184 8175 14240
rect 4705 14182 8175 14184
rect 4705 14179 4771 14182
rect 4889 14179 4955 14182
rect 8109 14179 8175 14182
rect 9622 14180 9628 14244
rect 9692 14242 9698 14244
rect 9765 14242 9831 14245
rect 9692 14240 9831 14242
rect 9692 14184 9770 14240
rect 9826 14184 9831 14240
rect 9692 14182 9831 14184
rect 9692 14180 9698 14182
rect 9765 14179 9831 14182
rect 10593 14242 10659 14245
rect 12709 14242 12775 14245
rect 10593 14240 12775 14242
rect 10593 14184 10598 14240
rect 10654 14184 12714 14240
rect 12770 14184 12775 14240
rect 10593 14182 12775 14184
rect 10593 14179 10659 14182
rect 12709 14179 12775 14182
rect 3409 14176 3729 14177
rect 0 14106 480 14136
rect 3409 14112 3417 14176
rect 3481 14112 3497 14176
rect 3561 14112 3577 14176
rect 3641 14112 3657 14176
rect 3721 14112 3729 14176
rect 3409 14111 3729 14112
rect 8340 14176 8660 14177
rect 8340 14112 8348 14176
rect 8412 14112 8428 14176
rect 8492 14112 8508 14176
rect 8572 14112 8588 14176
rect 8652 14112 8660 14176
rect 8340 14111 8660 14112
rect 13270 14176 13590 14177
rect 13270 14112 13278 14176
rect 13342 14112 13358 14176
rect 13422 14112 13438 14176
rect 13502 14112 13518 14176
rect 13582 14112 13590 14176
rect 13270 14111 13590 14112
rect 3141 14106 3207 14109
rect 0 14104 3207 14106
rect 0 14048 3146 14104
rect 3202 14048 3207 14104
rect 0 14046 3207 14048
rect 0 14016 480 14046
rect 3141 14043 3207 14046
rect 4470 14044 4476 14108
rect 4540 14106 4546 14108
rect 7005 14106 7071 14109
rect 9305 14108 9371 14109
rect 4540 14104 7071 14106
rect 4540 14048 7010 14104
rect 7066 14048 7071 14104
rect 4540 14046 7071 14048
rect 4540 14044 4546 14046
rect 7005 14043 7071 14046
rect 9254 14044 9260 14108
rect 9324 14106 9371 14108
rect 9581 14106 9647 14109
rect 10358 14106 10364 14108
rect 9324 14104 9416 14106
rect 9366 14048 9416 14104
rect 9324 14046 9416 14048
rect 9581 14104 10364 14106
rect 9581 14048 9586 14104
rect 9642 14048 10364 14104
rect 9581 14046 10364 14048
rect 9324 14044 9371 14046
rect 9305 14043 9371 14044
rect 9581 14043 9647 14046
rect 10358 14044 10364 14046
rect 10428 14044 10434 14108
rect 10542 14044 10548 14108
rect 10612 14106 10618 14108
rect 10612 14046 11668 14106
rect 10612 14044 10618 14046
rect 2497 13970 2563 13973
rect 7373 13970 7439 13973
rect 2497 13968 7439 13970
rect 2497 13912 2502 13968
rect 2558 13912 7378 13968
rect 7434 13912 7439 13968
rect 2497 13910 7439 13912
rect 2497 13907 2563 13910
rect 7373 13907 7439 13910
rect 7925 13970 7991 13973
rect 11421 13970 11487 13973
rect 7925 13968 11487 13970
rect 7925 13912 7930 13968
rect 7986 13912 11426 13968
rect 11482 13912 11487 13968
rect 7925 13910 11487 13912
rect 7925 13907 7991 13910
rect 11421 13907 11487 13910
rect 1853 13834 1919 13837
rect 9121 13834 9187 13837
rect 1853 13832 9187 13834
rect 1853 13776 1858 13832
rect 1914 13776 9126 13832
rect 9182 13776 9187 13832
rect 1853 13774 9187 13776
rect 1853 13771 1919 13774
rect 9121 13771 9187 13774
rect 9397 13834 9463 13837
rect 10409 13834 10475 13837
rect 9397 13832 10475 13834
rect 9397 13776 9402 13832
rect 9458 13776 10414 13832
rect 10470 13776 10475 13832
rect 9397 13774 10475 13776
rect 9397 13771 9463 13774
rect 10409 13771 10475 13774
rect 10550 13774 11346 13834
rect 6494 13636 6500 13700
rect 6564 13698 6570 13700
rect 7097 13698 7163 13701
rect 6564 13696 7163 13698
rect 6564 13640 7102 13696
rect 7158 13640 7163 13696
rect 6564 13638 7163 13640
rect 9124 13698 9184 13771
rect 10550 13698 10610 13774
rect 9124 13638 10610 13698
rect 11286 13701 11346 13774
rect 11286 13698 11395 13701
rect 11608 13698 11668 14046
rect 11789 13836 11855 13837
rect 12433 13836 12499 13837
rect 11789 13832 11836 13836
rect 11900 13834 11906 13836
rect 12382 13834 12388 13836
rect 11789 13776 11794 13832
rect 11789 13772 11836 13776
rect 11900 13774 11946 13834
rect 12342 13774 12388 13834
rect 12452 13832 12499 13836
rect 12494 13776 12499 13832
rect 11900 13772 11906 13774
rect 12382 13772 12388 13774
rect 12452 13772 12499 13776
rect 11789 13771 11855 13772
rect 12433 13771 12499 13772
rect 12341 13698 12407 13701
rect 11286 13696 11530 13698
rect 11286 13640 11334 13696
rect 11390 13640 11530 13696
rect 11286 13638 11530 13640
rect 11608 13696 12407 13698
rect 11608 13640 12346 13696
rect 12402 13640 12407 13696
rect 11608 13638 12407 13640
rect 6564 13636 6570 13638
rect 7097 13635 7163 13638
rect 11329 13635 11395 13638
rect 5874 13632 6194 13633
rect 5874 13568 5882 13632
rect 5946 13568 5962 13632
rect 6026 13568 6042 13632
rect 6106 13568 6122 13632
rect 6186 13568 6194 13632
rect 5874 13567 6194 13568
rect 10805 13632 11125 13633
rect 10805 13568 10813 13632
rect 10877 13568 10893 13632
rect 10957 13568 10973 13632
rect 11037 13568 11053 13632
rect 11117 13568 11125 13632
rect 10805 13567 11125 13568
rect 6361 13562 6427 13565
rect 10542 13562 10548 13564
rect 6361 13560 10548 13562
rect 6361 13504 6366 13560
rect 6422 13504 10548 13560
rect 6361 13502 10548 13504
rect 6361 13499 6427 13502
rect 10542 13500 10548 13502
rect 10612 13500 10618 13564
rect 11470 13562 11530 13638
rect 12341 13635 12407 13638
rect 12198 13562 12204 13564
rect 11470 13502 12204 13562
rect 12198 13500 12204 13502
rect 12268 13500 12274 13564
rect 5717 13426 5783 13429
rect 11697 13426 11763 13429
rect 11973 13426 12039 13429
rect 5717 13424 11763 13426
rect 5717 13368 5722 13424
rect 5778 13368 11702 13424
rect 11758 13368 11763 13424
rect 5717 13366 11763 13368
rect 5717 13363 5783 13366
rect 11697 13363 11763 13366
rect 11838 13424 12039 13426
rect 11838 13368 11978 13424
rect 12034 13368 12039 13424
rect 11838 13366 12039 13368
rect 3969 13290 4035 13293
rect 6361 13290 6427 13293
rect 3969 13288 6427 13290
rect 3969 13232 3974 13288
rect 4030 13232 6366 13288
rect 6422 13232 6427 13288
rect 3969 13230 6427 13232
rect 3969 13227 4035 13230
rect 6361 13227 6427 13230
rect 6545 13290 6611 13293
rect 11697 13290 11763 13293
rect 11838 13290 11898 13366
rect 11973 13363 12039 13366
rect 12341 13426 12407 13429
rect 12341 13424 12818 13426
rect 12341 13368 12346 13424
rect 12402 13368 12818 13424
rect 12341 13366 12818 13368
rect 12341 13363 12407 13366
rect 6545 13288 11530 13290
rect 6545 13232 6550 13288
rect 6606 13232 11530 13288
rect 6545 13230 11530 13232
rect 6545 13227 6611 13230
rect 0 13154 480 13184
rect 2773 13154 2839 13157
rect 0 13152 2839 13154
rect 0 13096 2778 13152
rect 2834 13096 2839 13152
rect 0 13094 2839 13096
rect 0 13064 480 13094
rect 2773 13091 2839 13094
rect 4705 13154 4771 13157
rect 7833 13154 7899 13157
rect 4705 13152 7899 13154
rect 4705 13096 4710 13152
rect 4766 13096 7838 13152
rect 7894 13096 7899 13152
rect 4705 13094 7899 13096
rect 4705 13091 4771 13094
rect 7833 13091 7899 13094
rect 9121 13154 9187 13157
rect 9857 13154 9923 13157
rect 9121 13152 9923 13154
rect 9121 13096 9126 13152
rect 9182 13096 9862 13152
rect 9918 13096 9923 13152
rect 9121 13094 9923 13096
rect 9121 13091 9187 13094
rect 9857 13091 9923 13094
rect 10225 13154 10291 13157
rect 11329 13154 11395 13157
rect 10225 13152 11395 13154
rect 10225 13096 10230 13152
rect 10286 13096 11334 13152
rect 11390 13096 11395 13152
rect 10225 13094 11395 13096
rect 10225 13091 10291 13094
rect 11329 13091 11395 13094
rect 3409 13088 3729 13089
rect 3409 13024 3417 13088
rect 3481 13024 3497 13088
rect 3561 13024 3577 13088
rect 3641 13024 3657 13088
rect 3721 13024 3729 13088
rect 3409 13023 3729 13024
rect 8340 13088 8660 13089
rect 8340 13024 8348 13088
rect 8412 13024 8428 13088
rect 8492 13024 8508 13088
rect 8572 13024 8588 13088
rect 8652 13024 8660 13088
rect 8340 13023 8660 13024
rect 8753 13018 8819 13021
rect 9438 13018 9444 13020
rect 3926 12958 7666 13018
rect 2773 12882 2839 12885
rect 3049 12882 3115 12885
rect 3693 12882 3759 12885
rect 3926 12882 3986 12958
rect 2773 12880 3986 12882
rect 2773 12824 2778 12880
rect 2834 12824 3054 12880
rect 3110 12824 3698 12880
rect 3754 12824 3986 12880
rect 2773 12822 3986 12824
rect 6177 12882 6243 12885
rect 7230 12882 7236 12884
rect 6177 12880 7236 12882
rect 6177 12824 6182 12880
rect 6238 12824 7236 12880
rect 6177 12822 7236 12824
rect 2773 12819 2839 12822
rect 3049 12819 3115 12822
rect 3693 12819 3759 12822
rect 6177 12819 6243 12822
rect 7230 12820 7236 12822
rect 7300 12820 7306 12884
rect 7606 12882 7666 12958
rect 8753 13016 9444 13018
rect 8753 12960 8758 13016
rect 8814 12960 9444 13016
rect 8753 12958 9444 12960
rect 8753 12955 8819 12958
rect 9438 12956 9444 12958
rect 9508 12956 9514 13020
rect 11470 12885 11530 13230
rect 11697 13288 11898 13290
rect 11697 13232 11702 13288
rect 11758 13232 11898 13288
rect 11697 13230 11898 13232
rect 11697 13227 11763 13230
rect 12014 13228 12020 13292
rect 12084 13290 12090 13292
rect 12157 13290 12223 13293
rect 12084 13288 12223 13290
rect 12084 13232 12162 13288
rect 12218 13232 12223 13288
rect 12084 13230 12223 13232
rect 12758 13290 12818 13366
rect 15285 13290 15351 13293
rect 12758 13288 15351 13290
rect 12758 13232 15290 13288
rect 15346 13232 15351 13288
rect 12758 13230 15351 13232
rect 12084 13228 12090 13230
rect 12157 13227 12223 13230
rect 15285 13227 15351 13230
rect 13270 13088 13590 13089
rect 13270 13024 13278 13088
rect 13342 13024 13358 13088
rect 13422 13024 13438 13088
rect 13502 13024 13518 13088
rect 13582 13024 13590 13088
rect 13270 13023 13590 13024
rect 8293 12882 8359 12885
rect 7606 12880 8359 12882
rect 7606 12824 8298 12880
rect 8354 12824 8359 12880
rect 7606 12822 8359 12824
rect 8293 12819 8359 12822
rect 8569 12882 8635 12885
rect 10777 12882 10843 12885
rect 8569 12880 10843 12882
rect 8569 12824 8574 12880
rect 8630 12824 10782 12880
rect 10838 12824 10843 12880
rect 8569 12822 10843 12824
rect 11470 12880 11579 12885
rect 11470 12824 11518 12880
rect 11574 12824 11579 12880
rect 11470 12822 11579 12824
rect 8569 12819 8635 12822
rect 10777 12819 10843 12822
rect 11513 12819 11579 12822
rect 12893 12880 12959 12885
rect 13169 12884 13235 12885
rect 13118 12882 13124 12884
rect 12893 12824 12898 12880
rect 12954 12824 12959 12880
rect 12893 12819 12959 12824
rect 13078 12822 13124 12882
rect 13188 12880 13235 12884
rect 13230 12824 13235 12880
rect 13118 12820 13124 12822
rect 13188 12820 13235 12824
rect 13169 12819 13235 12820
rect 3877 12746 3943 12749
rect 12433 12746 12499 12749
rect 3877 12744 12499 12746
rect 3877 12688 3882 12744
rect 3938 12688 12438 12744
rect 12494 12688 12499 12744
rect 3877 12686 12499 12688
rect 12896 12746 12956 12819
rect 13169 12746 13235 12749
rect 12896 12744 13235 12746
rect 12896 12688 13174 12744
rect 13230 12688 13235 12744
rect 12896 12686 13235 12688
rect 3877 12683 3943 12686
rect 12433 12683 12499 12686
rect 13169 12683 13235 12686
rect 4429 12612 4495 12613
rect 4429 12610 4476 12612
rect 4384 12608 4476 12610
rect 4384 12552 4434 12608
rect 4384 12550 4476 12552
rect 4429 12548 4476 12550
rect 4540 12548 4546 12612
rect 6729 12610 6795 12613
rect 7557 12610 7623 12613
rect 6729 12608 7623 12610
rect 6729 12552 6734 12608
rect 6790 12552 7562 12608
rect 7618 12552 7623 12608
rect 6729 12550 7623 12552
rect 4429 12547 4495 12548
rect 6729 12547 6795 12550
rect 7557 12547 7623 12550
rect 8753 12610 8819 12613
rect 8886 12610 8892 12612
rect 8753 12608 8892 12610
rect 8753 12552 8758 12608
rect 8814 12552 8892 12608
rect 8753 12550 8892 12552
rect 8753 12547 8819 12550
rect 8886 12548 8892 12550
rect 8956 12548 8962 12612
rect 9029 12610 9095 12613
rect 9581 12610 9647 12613
rect 9029 12608 9647 12610
rect 9029 12552 9034 12608
rect 9090 12552 9586 12608
rect 9642 12552 9647 12608
rect 9029 12550 9647 12552
rect 9029 12547 9095 12550
rect 9581 12547 9647 12550
rect 11421 12610 11487 12613
rect 11646 12610 11652 12612
rect 11421 12608 11652 12610
rect 11421 12552 11426 12608
rect 11482 12552 11652 12608
rect 11421 12550 11652 12552
rect 11421 12547 11487 12550
rect 11646 12548 11652 12550
rect 11716 12548 11722 12612
rect 12750 12548 12756 12612
rect 12820 12610 12826 12612
rect 12893 12610 12959 12613
rect 12820 12608 12959 12610
rect 12820 12552 12898 12608
rect 12954 12552 12959 12608
rect 12820 12550 12959 12552
rect 12820 12548 12826 12550
rect 12893 12547 12959 12550
rect 5874 12544 6194 12545
rect 5874 12480 5882 12544
rect 5946 12480 5962 12544
rect 6026 12480 6042 12544
rect 6106 12480 6122 12544
rect 6186 12480 6194 12544
rect 5874 12479 6194 12480
rect 10805 12544 11125 12545
rect 10805 12480 10813 12544
rect 10877 12480 10893 12544
rect 10957 12480 10973 12544
rect 11037 12480 11053 12544
rect 11117 12480 11125 12544
rect 10805 12479 11125 12480
rect 5073 12474 5139 12477
rect 2086 12472 5139 12474
rect 2086 12416 5078 12472
rect 5134 12416 5139 12472
rect 2086 12414 5139 12416
rect 2086 12341 2146 12414
rect 5073 12411 5139 12414
rect 6545 12474 6611 12477
rect 6678 12474 6684 12476
rect 6545 12472 6684 12474
rect 6545 12416 6550 12472
rect 6606 12416 6684 12472
rect 6545 12414 6684 12416
rect 6545 12411 6611 12414
rect 6678 12412 6684 12414
rect 6748 12412 6754 12476
rect 6821 12474 6887 12477
rect 7189 12474 7255 12477
rect 6821 12472 7255 12474
rect 6821 12416 6826 12472
rect 6882 12416 7194 12472
rect 7250 12416 7255 12472
rect 6821 12414 7255 12416
rect 6821 12411 6887 12414
rect 7189 12411 7255 12414
rect 7649 12474 7715 12477
rect 9029 12474 9095 12477
rect 9397 12476 9463 12477
rect 9397 12474 9444 12476
rect 7649 12472 9095 12474
rect 7649 12416 7654 12472
rect 7710 12416 9034 12472
rect 9090 12416 9095 12472
rect 7649 12414 9095 12416
rect 9352 12472 9444 12474
rect 9352 12416 9402 12472
rect 9352 12414 9444 12416
rect 7649 12411 7715 12414
rect 9029 12411 9095 12414
rect 9397 12412 9444 12414
rect 9508 12412 9514 12476
rect 9857 12474 9923 12477
rect 10409 12474 10475 12477
rect 9857 12472 10475 12474
rect 9857 12416 9862 12472
rect 9918 12416 10414 12472
rect 10470 12416 10475 12472
rect 9857 12414 10475 12416
rect 9397 12411 9463 12412
rect 9857 12411 9923 12414
rect 10409 12411 10475 12414
rect 11329 12474 11395 12477
rect 12893 12474 12959 12477
rect 11329 12472 12959 12474
rect 11329 12416 11334 12472
rect 11390 12416 12898 12472
rect 12954 12416 12959 12472
rect 11329 12414 12959 12416
rect 11329 12411 11395 12414
rect 12893 12411 12959 12414
rect 2037 12336 2146 12341
rect 2037 12280 2042 12336
rect 2098 12280 2146 12336
rect 2037 12278 2146 12280
rect 2313 12338 2379 12341
rect 13813 12338 13879 12341
rect 2313 12336 13879 12338
rect 2313 12280 2318 12336
rect 2374 12280 13818 12336
rect 13874 12280 13879 12336
rect 2313 12278 13879 12280
rect 2037 12275 2103 12278
rect 2313 12275 2379 12278
rect 13813 12275 13879 12278
rect 2405 12202 2471 12205
rect 2405 12200 8954 12202
rect 2405 12144 2410 12200
rect 2466 12144 8954 12200
rect 2405 12142 8954 12144
rect 2405 12139 2471 12142
rect 0 12066 480 12096
rect 1669 12066 1735 12069
rect 0 12064 1735 12066
rect 0 12008 1674 12064
rect 1730 12008 1735 12064
rect 0 12006 1735 12008
rect 0 11976 480 12006
rect 1669 12003 1735 12006
rect 4061 12066 4127 12069
rect 5574 12066 5580 12068
rect 4061 12064 5580 12066
rect 4061 12008 4066 12064
rect 4122 12008 5580 12064
rect 4061 12006 5580 12008
rect 4061 12003 4127 12006
rect 5574 12004 5580 12006
rect 5644 12066 5650 12068
rect 7833 12066 7899 12069
rect 5644 12064 7899 12066
rect 5644 12008 7838 12064
rect 7894 12008 7899 12064
rect 5644 12006 7899 12008
rect 8894 12066 8954 12142
rect 9254 12140 9260 12204
rect 9324 12202 9330 12204
rect 9397 12202 9463 12205
rect 9324 12200 9463 12202
rect 9324 12144 9402 12200
rect 9458 12144 9463 12200
rect 9324 12142 9463 12144
rect 9324 12140 9330 12142
rect 9397 12139 9463 12142
rect 9806 12140 9812 12204
rect 9876 12202 9882 12204
rect 9949 12202 10015 12205
rect 9876 12200 10015 12202
rect 9876 12144 9954 12200
rect 10010 12144 10015 12200
rect 9876 12142 10015 12144
rect 9876 12140 9882 12142
rect 9949 12139 10015 12142
rect 10409 12202 10475 12205
rect 11053 12202 11119 12205
rect 10409 12200 11119 12202
rect 10409 12144 10414 12200
rect 10470 12144 11058 12200
rect 11114 12144 11119 12200
rect 10409 12142 11119 12144
rect 10409 12139 10475 12142
rect 11053 12139 11119 12142
rect 12709 12202 12775 12205
rect 14406 12202 14412 12204
rect 12709 12200 14412 12202
rect 12709 12144 12714 12200
rect 12770 12144 14412 12200
rect 12709 12142 14412 12144
rect 12709 12139 12775 12142
rect 14406 12140 14412 12142
rect 14476 12140 14482 12204
rect 9765 12066 9831 12069
rect 8894 12064 9831 12066
rect 8894 12008 9770 12064
rect 9826 12008 9831 12064
rect 8894 12006 9831 12008
rect 5644 12004 5650 12006
rect 7833 12003 7899 12006
rect 9765 12003 9831 12006
rect 10041 12066 10107 12069
rect 10501 12066 10567 12069
rect 10041 12064 10567 12066
rect 10041 12008 10046 12064
rect 10102 12008 10506 12064
rect 10562 12008 10567 12064
rect 10041 12006 10567 12008
rect 10041 12003 10107 12006
rect 10501 12003 10567 12006
rect 10961 12066 11027 12069
rect 11278 12066 11284 12068
rect 10961 12064 11284 12066
rect 10961 12008 10966 12064
rect 11022 12008 11284 12064
rect 10961 12006 11284 12008
rect 10961 12003 11027 12006
rect 11278 12004 11284 12006
rect 11348 12004 11354 12068
rect 3409 12000 3729 12001
rect 3409 11936 3417 12000
rect 3481 11936 3497 12000
rect 3561 11936 3577 12000
rect 3641 11936 3657 12000
rect 3721 11936 3729 12000
rect 3409 11935 3729 11936
rect 8340 12000 8660 12001
rect 8340 11936 8348 12000
rect 8412 11936 8428 12000
rect 8492 11936 8508 12000
rect 8572 11936 8588 12000
rect 8652 11936 8660 12000
rect 8340 11935 8660 11936
rect 13270 12000 13590 12001
rect 13270 11936 13278 12000
rect 13342 11936 13358 12000
rect 13422 11936 13438 12000
rect 13502 11936 13518 12000
rect 13582 11936 13590 12000
rect 13270 11935 13590 11936
rect 5901 11930 5967 11933
rect 7465 11930 7531 11933
rect 5214 11928 7531 11930
rect 5214 11872 5906 11928
rect 5962 11872 7470 11928
rect 7526 11872 7531 11928
rect 5214 11870 7531 11872
rect 3417 11794 3483 11797
rect 5214 11794 5274 11870
rect 5901 11867 5967 11870
rect 7465 11867 7531 11870
rect 8753 11930 8819 11933
rect 9070 11930 9076 11932
rect 8753 11928 9076 11930
rect 8753 11872 8758 11928
rect 8814 11872 9076 11928
rect 8753 11870 9076 11872
rect 8753 11867 8819 11870
rect 9070 11868 9076 11870
rect 9140 11868 9146 11932
rect 9213 11930 9279 11933
rect 9622 11930 9628 11932
rect 9213 11928 9628 11930
rect 9213 11872 9218 11928
rect 9274 11872 9628 11928
rect 9213 11870 9628 11872
rect 9213 11867 9279 11870
rect 9622 11868 9628 11870
rect 9692 11868 9698 11932
rect 10358 11868 10364 11932
rect 10428 11930 10434 11932
rect 11053 11930 11119 11933
rect 10428 11928 11119 11930
rect 10428 11872 11058 11928
rect 11114 11872 11119 11928
rect 10428 11870 11119 11872
rect 10428 11868 10434 11870
rect 11053 11867 11119 11870
rect 12065 11930 12131 11933
rect 12893 11930 12959 11933
rect 12065 11928 12959 11930
rect 12065 11872 12070 11928
rect 12126 11872 12898 11928
rect 12954 11872 12959 11928
rect 12065 11870 12959 11872
rect 12065 11867 12131 11870
rect 12893 11867 12959 11870
rect 3417 11792 5274 11794
rect 3417 11736 3422 11792
rect 3478 11736 5274 11792
rect 3417 11734 5274 11736
rect 5809 11794 5875 11797
rect 10409 11796 10475 11797
rect 9990 11794 9996 11796
rect 5809 11792 9996 11794
rect 5809 11736 5814 11792
rect 5870 11736 9996 11792
rect 5809 11734 9996 11736
rect 3417 11731 3483 11734
rect 5809 11731 5875 11734
rect 9990 11732 9996 11734
rect 10060 11732 10066 11796
rect 10358 11794 10364 11796
rect 10318 11734 10364 11794
rect 10428 11792 10475 11796
rect 10470 11736 10475 11792
rect 10358 11732 10364 11734
rect 10428 11732 10475 11736
rect 10409 11731 10475 11732
rect 10869 11794 10935 11797
rect 13261 11794 13327 11797
rect 10869 11792 13327 11794
rect 10869 11736 10874 11792
rect 10930 11736 13266 11792
rect 13322 11736 13327 11792
rect 10869 11734 13327 11736
rect 10869 11731 10935 11734
rect 13261 11731 13327 11734
rect 2405 11658 2471 11661
rect 13445 11658 13511 11661
rect 2405 11656 13511 11658
rect 2405 11600 2410 11656
rect 2466 11600 13450 11656
rect 13506 11600 13511 11656
rect 2405 11598 13511 11600
rect 2405 11595 2471 11598
rect 13445 11595 13511 11598
rect 7465 11522 7531 11525
rect 8845 11522 8911 11525
rect 7465 11520 8911 11522
rect 7465 11464 7470 11520
rect 7526 11464 8850 11520
rect 8906 11464 8911 11520
rect 7465 11462 8911 11464
rect 7465 11459 7531 11462
rect 8845 11459 8911 11462
rect 11646 11460 11652 11524
rect 11716 11522 11722 11524
rect 14825 11522 14891 11525
rect 11716 11520 14891 11522
rect 11716 11464 14830 11520
rect 14886 11464 14891 11520
rect 11716 11462 14891 11464
rect 11716 11460 11722 11462
rect 14825 11459 14891 11462
rect 5874 11456 6194 11457
rect 5874 11392 5882 11456
rect 5946 11392 5962 11456
rect 6026 11392 6042 11456
rect 6106 11392 6122 11456
rect 6186 11392 6194 11456
rect 5874 11391 6194 11392
rect 10805 11456 11125 11457
rect 10805 11392 10813 11456
rect 10877 11392 10893 11456
rect 10957 11392 10973 11456
rect 11037 11392 11053 11456
rect 11117 11392 11125 11456
rect 10805 11391 11125 11392
rect 7782 11324 7788 11388
rect 7852 11386 7858 11388
rect 7925 11386 7991 11389
rect 10409 11386 10475 11389
rect 12709 11386 12775 11389
rect 7852 11384 10475 11386
rect 7852 11328 7930 11384
rect 7986 11328 10414 11384
rect 10470 11328 10475 11384
rect 7852 11326 10475 11328
rect 7852 11324 7858 11326
rect 7925 11323 7991 11326
rect 10409 11323 10475 11326
rect 11286 11384 12775 11386
rect 11286 11328 12714 11384
rect 12770 11328 12775 11384
rect 11286 11326 12775 11328
rect 2497 11250 2563 11253
rect 11286 11250 11346 11326
rect 12709 11323 12775 11326
rect 2497 11248 11346 11250
rect 2497 11192 2502 11248
rect 2558 11192 11346 11248
rect 2497 11190 11346 11192
rect 2497 11187 2563 11190
rect 11646 11188 11652 11252
rect 11716 11250 11722 11252
rect 13169 11250 13235 11253
rect 11716 11248 13235 11250
rect 11716 11192 13174 11248
rect 13230 11192 13235 11248
rect 11716 11190 13235 11192
rect 11716 11188 11722 11190
rect 13169 11187 13235 11190
rect 13537 11250 13603 11253
rect 14958 11250 14964 11252
rect 13537 11248 14964 11250
rect 13537 11192 13542 11248
rect 13598 11192 14964 11248
rect 13537 11190 14964 11192
rect 13537 11187 13603 11190
rect 14958 11188 14964 11190
rect 15028 11188 15034 11252
rect 2497 11114 2563 11117
rect 8845 11114 8911 11117
rect 2497 11112 8911 11114
rect 2497 11056 2502 11112
rect 2558 11056 8850 11112
rect 8906 11056 8911 11112
rect 2497 11054 8911 11056
rect 2497 11051 2563 11054
rect 8845 11051 8911 11054
rect 9305 11114 9371 11117
rect 13629 11114 13695 11117
rect 14089 11116 14155 11117
rect 14038 11114 14044 11116
rect 9305 11112 13695 11114
rect 9305 11056 9310 11112
rect 9366 11056 13634 11112
rect 13690 11056 13695 11112
rect 9305 11054 13695 11056
rect 13998 11054 14044 11114
rect 14108 11112 14155 11116
rect 14150 11056 14155 11112
rect 9305 11051 9371 11054
rect 13629 11051 13695 11054
rect 14038 11052 14044 11054
rect 14108 11052 14155 11056
rect 14089 11051 14155 11052
rect 0 10978 480 11008
rect 1853 10978 1919 10981
rect 0 10976 1919 10978
rect 0 10920 1858 10976
rect 1914 10920 1919 10976
rect 0 10918 1919 10920
rect 0 10888 480 10918
rect 1853 10915 1919 10918
rect 5717 10978 5783 10981
rect 7414 10978 7420 10980
rect 5717 10976 7420 10978
rect 5717 10920 5722 10976
rect 5778 10920 7420 10976
rect 5717 10918 7420 10920
rect 5717 10915 5783 10918
rect 7414 10916 7420 10918
rect 7484 10916 7490 10980
rect 8845 10978 8911 10981
rect 9622 10978 9628 10980
rect 8845 10976 9628 10978
rect 8845 10920 8850 10976
rect 8906 10920 9628 10976
rect 8845 10918 9628 10920
rect 8845 10915 8911 10918
rect 9622 10916 9628 10918
rect 9692 10978 9698 10980
rect 12801 10978 12867 10981
rect 9692 10976 12867 10978
rect 9692 10920 12806 10976
rect 12862 10920 12867 10976
rect 9692 10918 12867 10920
rect 9692 10916 9698 10918
rect 12801 10915 12867 10918
rect 13721 10976 13787 10981
rect 13721 10920 13726 10976
rect 13782 10920 13787 10976
rect 13721 10915 13787 10920
rect 3409 10912 3729 10913
rect 3409 10848 3417 10912
rect 3481 10848 3497 10912
rect 3561 10848 3577 10912
rect 3641 10848 3657 10912
rect 3721 10848 3729 10912
rect 3409 10847 3729 10848
rect 8340 10912 8660 10913
rect 8340 10848 8348 10912
rect 8412 10848 8428 10912
rect 8492 10848 8508 10912
rect 8572 10848 8588 10912
rect 8652 10848 8660 10912
rect 8340 10847 8660 10848
rect 13270 10912 13590 10913
rect 13270 10848 13278 10912
rect 13342 10848 13358 10912
rect 13422 10848 13438 10912
rect 13502 10848 13518 10912
rect 13582 10848 13590 10912
rect 13270 10847 13590 10848
rect 9990 10780 9996 10844
rect 10060 10842 10066 10844
rect 11145 10842 11211 10845
rect 10060 10840 11211 10842
rect 10060 10784 11150 10840
rect 11206 10784 11211 10840
rect 10060 10782 11211 10784
rect 10060 10780 10066 10782
rect 11145 10779 11211 10782
rect 11513 10842 11579 10845
rect 12014 10842 12020 10844
rect 11513 10840 12020 10842
rect 11513 10784 11518 10840
rect 11574 10784 12020 10840
rect 11513 10782 12020 10784
rect 11513 10779 11579 10782
rect 12014 10780 12020 10782
rect 12084 10780 12090 10844
rect 1945 10706 2011 10709
rect 6494 10706 6500 10708
rect 1945 10704 6500 10706
rect 1945 10648 1950 10704
rect 2006 10648 6500 10704
rect 1945 10646 6500 10648
rect 1945 10643 2011 10646
rect 6494 10644 6500 10646
rect 6564 10644 6570 10708
rect 7741 10706 7807 10709
rect 11973 10706 12039 10709
rect 7741 10704 12039 10706
rect 7741 10648 7746 10704
rect 7802 10648 11978 10704
rect 12034 10648 12039 10704
rect 7741 10646 12039 10648
rect 7741 10643 7807 10646
rect 11973 10643 12039 10646
rect 13537 10706 13603 10709
rect 13724 10706 13784 10915
rect 13537 10704 13784 10706
rect 13537 10648 13542 10704
rect 13598 10648 13784 10704
rect 13537 10646 13784 10648
rect 13537 10643 13603 10646
rect 2405 10570 2471 10573
rect 13813 10570 13879 10573
rect 2405 10568 13879 10570
rect 2405 10512 2410 10568
rect 2466 10512 13818 10568
rect 13874 10512 13879 10568
rect 2405 10510 13879 10512
rect 2405 10507 2471 10510
rect 13813 10507 13879 10510
rect 3049 10434 3115 10437
rect 3182 10434 3188 10436
rect 3049 10432 3188 10434
rect 3049 10376 3054 10432
rect 3110 10376 3188 10432
rect 3049 10374 3188 10376
rect 3049 10371 3115 10374
rect 3182 10372 3188 10374
rect 3252 10372 3258 10436
rect 7230 10372 7236 10436
rect 7300 10434 7306 10436
rect 8477 10434 8543 10437
rect 7300 10432 8543 10434
rect 7300 10376 8482 10432
rect 8538 10376 8543 10432
rect 7300 10374 8543 10376
rect 7300 10372 7306 10374
rect 8477 10371 8543 10374
rect 10174 10372 10180 10436
rect 10244 10434 10250 10436
rect 10501 10434 10567 10437
rect 10244 10432 10567 10434
rect 10244 10376 10506 10432
rect 10562 10376 10567 10432
rect 10244 10374 10567 10376
rect 10244 10372 10250 10374
rect 10501 10371 10567 10374
rect 11697 10434 11763 10437
rect 13169 10434 13235 10437
rect 15193 10434 15259 10437
rect 11697 10432 15259 10434
rect 11697 10376 11702 10432
rect 11758 10376 13174 10432
rect 13230 10376 15198 10432
rect 15254 10376 15259 10432
rect 11697 10374 15259 10376
rect 11697 10371 11763 10374
rect 13169 10371 13235 10374
rect 15193 10371 15259 10374
rect 5874 10368 6194 10369
rect 5874 10304 5882 10368
rect 5946 10304 5962 10368
rect 6026 10304 6042 10368
rect 6106 10304 6122 10368
rect 6186 10304 6194 10368
rect 5874 10303 6194 10304
rect 10805 10368 11125 10369
rect 10805 10304 10813 10368
rect 10877 10304 10893 10368
rect 10957 10304 10973 10368
rect 11037 10304 11053 10368
rect 11117 10304 11125 10368
rect 10805 10303 11125 10304
rect 6545 10298 6611 10301
rect 8886 10298 8892 10300
rect 6545 10296 8892 10298
rect 6545 10240 6550 10296
rect 6606 10240 8892 10296
rect 6545 10238 8892 10240
rect 6545 10235 6611 10238
rect 8886 10236 8892 10238
rect 8956 10298 8962 10300
rect 10593 10298 10659 10301
rect 8956 10296 10659 10298
rect 8956 10240 10598 10296
rect 10654 10240 10659 10296
rect 8956 10238 10659 10240
rect 8956 10236 8962 10238
rect 10593 10235 10659 10238
rect 12022 10238 13048 10298
rect 8017 10162 8083 10165
rect 12022 10162 12082 10238
rect 8017 10160 12082 10162
rect 8017 10104 8022 10160
rect 8078 10104 12082 10160
rect 8017 10102 12082 10104
rect 12988 10162 13048 10238
rect 14457 10162 14523 10165
rect 12988 10160 14523 10162
rect 12988 10104 14462 10160
rect 14518 10104 14523 10160
rect 12988 10102 14523 10104
rect 8017 10099 8083 10102
rect 14457 10099 14523 10102
rect 6310 9964 6316 10028
rect 6380 10026 6386 10028
rect 14181 10026 14247 10029
rect 6380 9992 12818 10026
rect 12988 10024 14247 10026
rect 12988 9992 14186 10024
rect 6380 9968 14186 9992
rect 14242 9968 14247 10024
rect 6380 9966 14247 9968
rect 6380 9964 6386 9966
rect 12758 9932 13048 9966
rect 14181 9963 14247 9966
rect 0 9890 480 9920
rect 1853 9890 1919 9893
rect 11646 9890 11652 9892
rect 0 9888 1919 9890
rect 0 9832 1858 9888
rect 1914 9832 1919 9888
rect 0 9830 1919 9832
rect 0 9800 480 9830
rect 1853 9827 1919 9830
rect 9262 9830 11652 9890
rect 3409 9824 3729 9825
rect 3409 9760 3417 9824
rect 3481 9760 3497 9824
rect 3561 9760 3577 9824
rect 3641 9760 3657 9824
rect 3721 9760 3729 9824
rect 3409 9759 3729 9760
rect 8340 9824 8660 9825
rect 8340 9760 8348 9824
rect 8412 9760 8428 9824
rect 8492 9760 8508 9824
rect 8572 9760 8588 9824
rect 8652 9760 8660 9824
rect 8340 9759 8660 9760
rect 8845 9754 8911 9757
rect 9262 9754 9322 9830
rect 11646 9828 11652 9830
rect 11716 9828 11722 9892
rect 11830 9828 11836 9892
rect 11900 9890 11906 9892
rect 12065 9890 12131 9893
rect 11900 9888 12131 9890
rect 11900 9832 12070 9888
rect 12126 9832 12131 9888
rect 11900 9830 12131 9832
rect 11900 9828 11906 9830
rect 12065 9827 12131 9830
rect 13270 9824 13590 9825
rect 13270 9760 13278 9824
rect 13342 9760 13358 9824
rect 13422 9760 13438 9824
rect 13502 9760 13518 9824
rect 13582 9760 13590 9824
rect 13270 9759 13590 9760
rect 8845 9752 9322 9754
rect 8845 9696 8850 9752
rect 8906 9696 9322 9752
rect 8845 9694 9322 9696
rect 10225 9754 10291 9757
rect 10961 9754 11027 9757
rect 10225 9752 11027 9754
rect 10225 9696 10230 9752
rect 10286 9696 10966 9752
rect 11022 9696 11027 9752
rect 10225 9694 11027 9696
rect 8845 9691 8911 9694
rect 10225 9691 10291 9694
rect 10961 9691 11027 9694
rect 3877 9618 3943 9621
rect 7649 9618 7715 9621
rect 3877 9616 7715 9618
rect 3877 9560 3882 9616
rect 3938 9560 7654 9616
rect 7710 9560 7715 9616
rect 3877 9558 7715 9560
rect 3877 9555 3943 9558
rect 7649 9555 7715 9558
rect 8109 9618 8175 9621
rect 10225 9618 10291 9621
rect 8109 9616 10291 9618
rect 8109 9560 8114 9616
rect 8170 9560 10230 9616
rect 10286 9560 10291 9616
rect 8109 9558 10291 9560
rect 8109 9555 8175 9558
rect 10225 9555 10291 9558
rect 10358 9556 10364 9620
rect 10428 9618 10434 9620
rect 13813 9618 13879 9621
rect 15009 9620 15075 9621
rect 10428 9616 13879 9618
rect 10428 9560 13818 9616
rect 13874 9560 13879 9616
rect 10428 9558 13879 9560
rect 10428 9556 10434 9558
rect 13813 9555 13879 9558
rect 14958 9556 14964 9620
rect 15028 9618 15075 9620
rect 15028 9616 15120 9618
rect 15070 9560 15120 9616
rect 15028 9558 15120 9560
rect 15028 9556 15075 9558
rect 15009 9555 15075 9556
rect 6085 9482 6151 9485
rect 8385 9482 8451 9485
rect 11053 9482 11119 9485
rect 6085 9480 7528 9482
rect 6085 9424 6090 9480
rect 6146 9424 7528 9480
rect 6085 9422 7528 9424
rect 6085 9419 6151 9422
rect 7468 9349 7528 9422
rect 8385 9480 11119 9482
rect 8385 9424 8390 9480
rect 8446 9424 11058 9480
rect 11114 9424 11119 9480
rect 8385 9422 11119 9424
rect 8385 9419 8451 9422
rect 11053 9419 11119 9422
rect 11421 9482 11487 9485
rect 13629 9482 13695 9485
rect 11421 9480 13695 9482
rect 11421 9424 11426 9480
rect 11482 9424 13634 9480
rect 13690 9424 13695 9480
rect 11421 9422 13695 9424
rect 11421 9419 11487 9422
rect 13629 9419 13695 9422
rect 7465 9346 7531 9349
rect 9438 9346 9444 9348
rect 7465 9344 9444 9346
rect 7465 9288 7470 9344
rect 7526 9288 9444 9344
rect 7465 9286 9444 9288
rect 7465 9283 7531 9286
rect 9438 9284 9444 9286
rect 9508 9284 9514 9348
rect 11646 9346 11652 9348
rect 11240 9286 11652 9346
rect 5874 9280 6194 9281
rect 5874 9216 5882 9280
rect 5946 9216 5962 9280
rect 6026 9216 6042 9280
rect 6106 9216 6122 9280
rect 6186 9216 6194 9280
rect 5874 9215 6194 9216
rect 10805 9280 11125 9281
rect 10805 9216 10813 9280
rect 10877 9216 10893 9280
rect 10957 9216 10973 9280
rect 11037 9216 11053 9280
rect 11117 9216 11125 9280
rect 10805 9215 11125 9216
rect 11240 9213 11300 9286
rect 11646 9284 11652 9286
rect 11716 9284 11722 9348
rect 11881 9346 11947 9349
rect 13261 9346 13327 9349
rect 11881 9344 13327 9346
rect 11881 9288 11886 9344
rect 11942 9288 13266 9344
rect 13322 9288 13327 9344
rect 11881 9286 13327 9288
rect 11881 9283 11947 9286
rect 13261 9283 13327 9286
rect 8109 9210 8175 9213
rect 9305 9210 9371 9213
rect 8109 9208 9371 9210
rect 8109 9152 8114 9208
rect 8170 9152 9310 9208
rect 9366 9152 9371 9208
rect 8109 9150 9371 9152
rect 8109 9147 8175 9150
rect 9305 9147 9371 9150
rect 11237 9208 11303 9213
rect 11237 9152 11242 9208
rect 11298 9152 11303 9208
rect 11237 9147 11303 9152
rect 11697 9210 11763 9213
rect 13445 9210 13511 9213
rect 11697 9208 13511 9210
rect 11697 9152 11702 9208
rect 11758 9152 13450 9208
rect 13506 9152 13511 9208
rect 11697 9150 13511 9152
rect 11697 9147 11763 9150
rect 13445 9147 13511 9150
rect 4981 9074 5047 9077
rect 12014 9074 12020 9076
rect 4981 9072 12020 9074
rect 4981 9016 4986 9072
rect 5042 9016 12020 9072
rect 4981 9014 12020 9016
rect 4981 9011 5047 9014
rect 12014 9012 12020 9014
rect 12084 9012 12090 9076
rect 15469 9074 15535 9077
rect 16520 9074 17000 9104
rect 15469 9072 17000 9074
rect 15469 9016 15474 9072
rect 15530 9016 17000 9072
rect 15469 9014 17000 9016
rect 15469 9011 15535 9014
rect 16520 8984 17000 9014
rect 0 8938 480 8968
rect 4061 8938 4127 8941
rect 0 8936 4127 8938
rect 0 8880 4066 8936
rect 4122 8880 4127 8936
rect 0 8878 4127 8880
rect 0 8848 480 8878
rect 4061 8875 4127 8878
rect 9806 8876 9812 8940
rect 9876 8938 9882 8940
rect 10777 8938 10843 8941
rect 9876 8936 10843 8938
rect 9876 8880 10782 8936
rect 10838 8880 10843 8936
rect 9876 8878 10843 8880
rect 9876 8876 9882 8878
rect 10777 8875 10843 8878
rect 11789 8938 11855 8941
rect 15377 8938 15443 8941
rect 11789 8936 15443 8938
rect 11789 8880 11794 8936
rect 11850 8880 15382 8936
rect 15438 8880 15443 8936
rect 11789 8878 15443 8880
rect 11789 8875 11855 8878
rect 15377 8875 15443 8878
rect 9121 8802 9187 8805
rect 11646 8802 11652 8804
rect 9121 8800 11652 8802
rect 9121 8744 9126 8800
rect 9182 8744 11652 8800
rect 9121 8742 11652 8744
rect 9121 8739 9187 8742
rect 11646 8740 11652 8742
rect 11716 8740 11722 8804
rect 3409 8736 3729 8737
rect 3409 8672 3417 8736
rect 3481 8672 3497 8736
rect 3561 8672 3577 8736
rect 3641 8672 3657 8736
rect 3721 8672 3729 8736
rect 3409 8671 3729 8672
rect 8340 8736 8660 8737
rect 8340 8672 8348 8736
rect 8412 8672 8428 8736
rect 8492 8672 8508 8736
rect 8572 8672 8588 8736
rect 8652 8672 8660 8736
rect 8340 8671 8660 8672
rect 13270 8736 13590 8737
rect 13270 8672 13278 8736
rect 13342 8672 13358 8736
rect 13422 8672 13438 8736
rect 13502 8672 13518 8736
rect 13582 8672 13590 8736
rect 13270 8671 13590 8672
rect 6729 8666 6795 8669
rect 8150 8666 8156 8668
rect 6729 8664 8156 8666
rect 6729 8608 6734 8664
rect 6790 8608 8156 8664
rect 6729 8606 8156 8608
rect 6729 8603 6795 8606
rect 8150 8604 8156 8606
rect 8220 8604 8226 8668
rect 8845 8666 8911 8669
rect 12801 8666 12867 8669
rect 8845 8664 12867 8666
rect 8845 8608 8850 8664
rect 8906 8608 12806 8664
rect 12862 8608 12867 8664
rect 8845 8606 12867 8608
rect 8845 8603 8911 8606
rect 12801 8603 12867 8606
rect 5073 8530 5139 8533
rect 10041 8530 10107 8533
rect 10685 8530 10751 8533
rect 5073 8528 10751 8530
rect 5073 8472 5078 8528
rect 5134 8472 10046 8528
rect 10102 8472 10690 8528
rect 10746 8472 10751 8528
rect 5073 8470 10751 8472
rect 5073 8467 5139 8470
rect 10041 8467 10107 8470
rect 10685 8467 10751 8470
rect 10869 8530 10935 8533
rect 12525 8530 12591 8533
rect 10869 8528 12591 8530
rect 10869 8472 10874 8528
rect 10930 8472 12530 8528
rect 12586 8472 12591 8528
rect 10869 8470 12591 8472
rect 10869 8467 10935 8470
rect 12525 8467 12591 8470
rect 3693 8394 3759 8397
rect 6729 8394 6795 8397
rect 13721 8394 13787 8397
rect 3693 8392 13787 8394
rect 3693 8336 3698 8392
rect 3754 8336 6734 8392
rect 6790 8336 13726 8392
rect 13782 8336 13787 8392
rect 3693 8334 13787 8336
rect 3693 8331 3759 8334
rect 6729 8331 6795 8334
rect 13721 8331 13787 8334
rect 13854 8332 13860 8396
rect 13924 8394 13930 8396
rect 14089 8394 14155 8397
rect 13924 8392 14155 8394
rect 13924 8336 14094 8392
rect 14150 8336 14155 8392
rect 13924 8334 14155 8336
rect 13924 8332 13930 8334
rect 14089 8331 14155 8334
rect 14222 8332 14228 8396
rect 14292 8394 14298 8396
rect 14549 8394 14615 8397
rect 14292 8392 14615 8394
rect 14292 8336 14554 8392
rect 14610 8336 14615 8392
rect 14292 8334 14615 8336
rect 14292 8332 14298 8334
rect 14549 8331 14615 8334
rect 7414 8196 7420 8260
rect 7484 8258 7490 8260
rect 9029 8258 9095 8261
rect 7484 8256 9095 8258
rect 7484 8200 9034 8256
rect 9090 8200 9095 8256
rect 7484 8198 9095 8200
rect 7484 8196 7490 8198
rect 9029 8195 9095 8198
rect 12893 8258 12959 8261
rect 14958 8258 14964 8260
rect 12893 8256 14964 8258
rect 12893 8200 12898 8256
rect 12954 8200 14964 8256
rect 12893 8198 14964 8200
rect 12893 8195 12959 8198
rect 14958 8196 14964 8198
rect 15028 8196 15034 8260
rect 5874 8192 6194 8193
rect 5874 8128 5882 8192
rect 5946 8128 5962 8192
rect 6026 8128 6042 8192
rect 6106 8128 6122 8192
rect 6186 8128 6194 8192
rect 5874 8127 6194 8128
rect 10805 8192 11125 8193
rect 10805 8128 10813 8192
rect 10877 8128 10893 8192
rect 10957 8128 10973 8192
rect 11037 8128 11053 8192
rect 11117 8128 11125 8192
rect 10805 8127 11125 8128
rect 10225 8122 10291 8125
rect 6870 8120 10291 8122
rect 6870 8064 10230 8120
rect 10286 8064 10291 8120
rect 6870 8062 10291 8064
rect 5073 7986 5139 7989
rect 6870 7986 6930 8062
rect 10225 8059 10291 8062
rect 10409 8122 10475 8125
rect 11237 8124 11303 8125
rect 10542 8122 10548 8124
rect 10409 8120 10548 8122
rect 10409 8064 10414 8120
rect 10470 8064 10548 8120
rect 10409 8062 10548 8064
rect 10409 8059 10475 8062
rect 10542 8060 10548 8062
rect 10612 8060 10618 8124
rect 11237 8120 11284 8124
rect 11348 8122 11354 8124
rect 11237 8064 11242 8120
rect 11237 8060 11284 8064
rect 11348 8062 11394 8122
rect 11348 8060 11354 8062
rect 11237 8059 11303 8060
rect 5073 7984 6930 7986
rect 5073 7928 5078 7984
rect 5134 7928 6930 7984
rect 5073 7926 6930 7928
rect 5073 7923 5139 7926
rect 7046 7924 7052 7988
rect 7116 7986 7122 7988
rect 8477 7986 8543 7989
rect 7116 7984 8543 7986
rect 7116 7928 8482 7984
rect 8538 7928 8543 7984
rect 7116 7926 8543 7928
rect 7116 7924 7122 7926
rect 8477 7923 8543 7926
rect 8845 7986 8911 7989
rect 13077 7986 13143 7989
rect 8845 7984 13143 7986
rect 8845 7928 8850 7984
rect 8906 7928 13082 7984
rect 13138 7928 13143 7984
rect 8845 7926 13143 7928
rect 8845 7923 8911 7926
rect 13077 7923 13143 7926
rect 13445 7986 13511 7989
rect 13670 7986 13676 7988
rect 13445 7984 13676 7986
rect 13445 7928 13450 7984
rect 13506 7928 13676 7984
rect 13445 7926 13676 7928
rect 13445 7923 13511 7926
rect 13670 7924 13676 7926
rect 13740 7924 13746 7988
rect 0 7850 480 7880
rect 1761 7850 1827 7853
rect 0 7848 1827 7850
rect 0 7792 1766 7848
rect 1822 7792 1827 7848
rect 0 7790 1827 7792
rect 0 7760 480 7790
rect 1761 7787 1827 7790
rect 2221 7850 2287 7853
rect 9070 7850 9076 7852
rect 2221 7848 9076 7850
rect 2221 7792 2226 7848
rect 2282 7792 9076 7848
rect 2221 7790 9076 7792
rect 2221 7787 2287 7790
rect 9070 7788 9076 7790
rect 9140 7788 9146 7852
rect 15101 7850 15167 7853
rect 10044 7848 15167 7850
rect 10044 7792 15106 7848
rect 15162 7792 15167 7848
rect 10044 7790 15167 7792
rect 4429 7714 4495 7717
rect 5717 7714 5783 7717
rect 4429 7712 7666 7714
rect 4429 7656 4434 7712
rect 4490 7656 5722 7712
rect 5778 7656 7666 7712
rect 4429 7654 7666 7656
rect 4429 7651 4495 7654
rect 5717 7651 5783 7654
rect 3409 7648 3729 7649
rect 3409 7584 3417 7648
rect 3481 7584 3497 7648
rect 3561 7584 3577 7648
rect 3641 7584 3657 7648
rect 3721 7584 3729 7648
rect 3409 7583 3729 7584
rect 4705 7578 4771 7581
rect 6361 7578 6427 7581
rect 4705 7576 6427 7578
rect 4705 7520 4710 7576
rect 4766 7520 6366 7576
rect 6422 7520 6427 7576
rect 4705 7518 6427 7520
rect 4705 7515 4771 7518
rect 6361 7515 6427 7518
rect 2865 7442 2931 7445
rect 7281 7442 7347 7445
rect 7606 7444 7666 7654
rect 8340 7648 8660 7649
rect 8340 7584 8348 7648
rect 8412 7584 8428 7648
rect 8492 7584 8508 7648
rect 8572 7584 8588 7648
rect 8652 7584 8660 7648
rect 8340 7583 8660 7584
rect 8937 7580 9003 7581
rect 8886 7578 8892 7580
rect 8846 7518 8892 7578
rect 8956 7576 9003 7580
rect 8998 7520 9003 7576
rect 8886 7516 8892 7518
rect 8956 7516 9003 7520
rect 10044 7578 10104 7790
rect 15101 7787 15167 7790
rect 10225 7714 10291 7717
rect 11462 7714 11468 7716
rect 10225 7712 11468 7714
rect 10225 7656 10230 7712
rect 10286 7656 11468 7712
rect 10225 7654 11468 7656
rect 10225 7651 10291 7654
rect 11462 7652 11468 7654
rect 11532 7714 11538 7716
rect 12893 7714 12959 7717
rect 11532 7712 12959 7714
rect 11532 7656 12898 7712
rect 12954 7656 12959 7712
rect 11532 7654 12959 7656
rect 11532 7652 11538 7654
rect 12893 7651 12959 7654
rect 13270 7648 13590 7649
rect 13270 7584 13278 7648
rect 13342 7584 13358 7648
rect 13422 7584 13438 7648
rect 13502 7584 13518 7648
rect 13582 7584 13590 7648
rect 13270 7583 13590 7584
rect 10501 7578 10567 7581
rect 10044 7576 10567 7578
rect 10044 7520 10506 7576
rect 10562 7520 10567 7576
rect 10044 7518 10567 7520
rect 8937 7515 9003 7516
rect 10501 7515 10567 7518
rect 10777 7578 10843 7581
rect 11329 7578 11395 7581
rect 10777 7576 11395 7578
rect 10777 7520 10782 7576
rect 10838 7520 11334 7576
rect 11390 7520 11395 7576
rect 10777 7518 11395 7520
rect 10777 7515 10843 7518
rect 11329 7515 11395 7518
rect 2865 7440 7347 7442
rect 2865 7384 2870 7440
rect 2926 7384 7286 7440
rect 7342 7384 7347 7440
rect 2865 7382 7347 7384
rect 2865 7379 2931 7382
rect 7281 7379 7347 7382
rect 7598 7380 7604 7444
rect 7668 7442 7674 7444
rect 8017 7442 8083 7445
rect 7668 7440 8083 7442
rect 7668 7384 8022 7440
rect 8078 7384 8083 7440
rect 7668 7382 8083 7384
rect 7668 7380 7674 7382
rect 8017 7379 8083 7382
rect 9949 7442 10015 7445
rect 10685 7442 10751 7445
rect 9949 7440 10751 7442
rect 9949 7384 9954 7440
rect 10010 7384 10690 7440
rect 10746 7384 10751 7440
rect 9949 7382 10751 7384
rect 9949 7379 10015 7382
rect 10685 7379 10751 7382
rect 11053 7442 11119 7445
rect 11278 7442 11284 7444
rect 11053 7440 11284 7442
rect 11053 7384 11058 7440
rect 11114 7384 11284 7440
rect 11053 7382 11284 7384
rect 11053 7379 11119 7382
rect 11278 7380 11284 7382
rect 11348 7380 11354 7444
rect 11605 7442 11671 7445
rect 12157 7442 12223 7445
rect 11605 7440 12223 7442
rect 11605 7384 11610 7440
rect 11666 7384 12162 7440
rect 12218 7384 12223 7440
rect 11605 7382 12223 7384
rect 11605 7379 11671 7382
rect 12157 7379 12223 7382
rect 12433 7442 12499 7445
rect 12934 7442 12940 7444
rect 12433 7440 12940 7442
rect 12433 7384 12438 7440
rect 12494 7384 12940 7440
rect 12433 7382 12940 7384
rect 12433 7379 12499 7382
rect 12934 7380 12940 7382
rect 13004 7380 13010 7444
rect 5257 7306 5323 7309
rect 10777 7306 10843 7309
rect 5257 7304 10843 7306
rect 5257 7248 5262 7304
rect 5318 7248 10782 7304
rect 10838 7248 10843 7304
rect 5257 7246 10843 7248
rect 5257 7243 5323 7246
rect 10777 7243 10843 7246
rect 10961 7306 11027 7309
rect 11608 7306 11668 7379
rect 10961 7304 11668 7306
rect 10961 7248 10966 7304
rect 11022 7248 11668 7304
rect 10961 7246 11668 7248
rect 12249 7306 12315 7309
rect 12382 7306 12388 7308
rect 12249 7304 12388 7306
rect 12249 7248 12254 7304
rect 12310 7248 12388 7304
rect 12249 7246 12388 7248
rect 10961 7243 11027 7246
rect 12249 7243 12315 7246
rect 12382 7244 12388 7246
rect 12452 7244 12458 7308
rect 12617 7306 12683 7309
rect 12934 7306 12940 7308
rect 12617 7304 12940 7306
rect 12617 7248 12622 7304
rect 12678 7248 12940 7304
rect 12617 7246 12940 7248
rect 12617 7243 12683 7246
rect 12934 7244 12940 7246
rect 13004 7244 13010 7308
rect 3141 7170 3207 7173
rect 5717 7170 5783 7173
rect 3141 7168 5783 7170
rect 3141 7112 3146 7168
rect 3202 7112 5722 7168
rect 5778 7112 5783 7168
rect 3141 7110 5783 7112
rect 3141 7107 3207 7110
rect 5717 7107 5783 7110
rect 10409 7170 10475 7173
rect 10542 7170 10548 7172
rect 10409 7168 10548 7170
rect 10409 7112 10414 7168
rect 10470 7112 10548 7168
rect 10409 7110 10548 7112
rect 10409 7107 10475 7110
rect 10542 7108 10548 7110
rect 10612 7108 10618 7172
rect 11329 7170 11395 7173
rect 11462 7170 11468 7172
rect 11329 7168 11468 7170
rect 11329 7112 11334 7168
rect 11390 7112 11468 7168
rect 11329 7110 11468 7112
rect 11329 7107 11395 7110
rect 11462 7108 11468 7110
rect 11532 7108 11538 7172
rect 12382 7108 12388 7172
rect 12452 7170 12458 7172
rect 12985 7170 13051 7173
rect 12452 7168 13051 7170
rect 12452 7112 12990 7168
rect 13046 7112 13051 7168
rect 12452 7110 13051 7112
rect 12452 7108 12458 7110
rect 12985 7107 13051 7110
rect 13353 7170 13419 7173
rect 14774 7170 14780 7172
rect 13353 7168 14780 7170
rect 13353 7112 13358 7168
rect 13414 7112 14780 7168
rect 13353 7110 14780 7112
rect 13353 7107 13419 7110
rect 14774 7108 14780 7110
rect 14844 7108 14850 7172
rect 5874 7104 6194 7105
rect 5874 7040 5882 7104
rect 5946 7040 5962 7104
rect 6026 7040 6042 7104
rect 6106 7040 6122 7104
rect 6186 7040 6194 7104
rect 5874 7039 6194 7040
rect 10805 7104 11125 7105
rect 10805 7040 10813 7104
rect 10877 7040 10893 7104
rect 10957 7040 10973 7104
rect 11037 7040 11053 7104
rect 11117 7040 11125 7104
rect 10805 7039 11125 7040
rect 5206 6972 5212 7036
rect 5276 7034 5282 7036
rect 5625 7034 5691 7037
rect 5276 7032 5691 7034
rect 5276 6976 5630 7032
rect 5686 6976 5691 7032
rect 5276 6974 5691 6976
rect 5276 6972 5282 6974
rect 5625 6971 5691 6974
rect 6361 7034 6427 7037
rect 9305 7034 9371 7037
rect 6361 7032 9371 7034
rect 6361 6976 6366 7032
rect 6422 6976 9310 7032
rect 9366 6976 9371 7032
rect 6361 6974 9371 6976
rect 6361 6971 6427 6974
rect 9305 6971 9371 6974
rect 9949 7034 10015 7037
rect 10225 7034 10291 7037
rect 9949 7032 10291 7034
rect 9949 6976 9954 7032
rect 10010 6976 10230 7032
rect 10286 6976 10291 7032
rect 9949 6974 10291 6976
rect 9949 6971 10015 6974
rect 10225 6971 10291 6974
rect 11830 6972 11836 7036
rect 11900 7034 11906 7036
rect 12157 7034 12223 7037
rect 11900 7032 12223 7034
rect 11900 6976 12162 7032
rect 12218 6976 12223 7032
rect 11900 6974 12223 6976
rect 11900 6972 11906 6974
rect 12157 6971 12223 6974
rect 12709 7034 12775 7037
rect 12985 7034 13051 7037
rect 12709 7032 13051 7034
rect 12709 6976 12714 7032
rect 12770 6976 12990 7032
rect 13046 6976 13051 7032
rect 12709 6974 13051 6976
rect 12709 6971 12775 6974
rect 12985 6971 13051 6974
rect 3049 6898 3115 6901
rect 12525 6898 12591 6901
rect 3049 6896 12591 6898
rect 3049 6840 3054 6896
rect 3110 6840 12530 6896
rect 12586 6840 12591 6896
rect 3049 6838 12591 6840
rect 3049 6835 3115 6838
rect 12525 6835 12591 6838
rect 12709 6898 12775 6901
rect 15193 6898 15259 6901
rect 12709 6896 15259 6898
rect 12709 6840 12714 6896
rect 12770 6840 15198 6896
rect 15254 6840 15259 6896
rect 12709 6838 15259 6840
rect 12709 6835 12775 6838
rect 15193 6835 15259 6838
rect 0 6762 480 6792
rect 1761 6762 1827 6765
rect 0 6760 1827 6762
rect 0 6704 1766 6760
rect 1822 6704 1827 6760
rect 0 6702 1827 6704
rect 0 6672 480 6702
rect 1761 6699 1827 6702
rect 4061 6762 4127 6765
rect 14038 6762 14044 6764
rect 4061 6760 14044 6762
rect 4061 6704 4066 6760
rect 4122 6704 14044 6760
rect 4061 6702 14044 6704
rect 4061 6699 4127 6702
rect 14038 6700 14044 6702
rect 14108 6700 14114 6764
rect 9029 6626 9095 6629
rect 10174 6626 10180 6628
rect 9029 6624 10180 6626
rect 9029 6568 9034 6624
rect 9090 6568 10180 6624
rect 9029 6566 10180 6568
rect 9029 6563 9095 6566
rect 10174 6564 10180 6566
rect 10244 6626 10250 6628
rect 11462 6626 11468 6628
rect 10244 6566 11468 6626
rect 10244 6564 10250 6566
rect 11462 6564 11468 6566
rect 11532 6564 11538 6628
rect 11830 6564 11836 6628
rect 11900 6626 11906 6628
rect 12341 6626 12407 6629
rect 11900 6624 12407 6626
rect 11900 6568 12346 6624
rect 12402 6568 12407 6624
rect 11900 6566 12407 6568
rect 11900 6564 11906 6566
rect 12341 6563 12407 6566
rect 3409 6560 3729 6561
rect 3409 6496 3417 6560
rect 3481 6496 3497 6560
rect 3561 6496 3577 6560
rect 3641 6496 3657 6560
rect 3721 6496 3729 6560
rect 3409 6495 3729 6496
rect 8340 6560 8660 6561
rect 8340 6496 8348 6560
rect 8412 6496 8428 6560
rect 8492 6496 8508 6560
rect 8572 6496 8588 6560
rect 8652 6496 8660 6560
rect 8340 6495 8660 6496
rect 13270 6560 13590 6561
rect 13270 6496 13278 6560
rect 13342 6496 13358 6560
rect 13422 6496 13438 6560
rect 13502 6496 13518 6560
rect 13582 6496 13590 6560
rect 13270 6495 13590 6496
rect 4613 6490 4679 6493
rect 8017 6490 8083 6493
rect 4613 6488 8083 6490
rect 4613 6432 4618 6488
rect 4674 6432 8022 6488
rect 8078 6432 8083 6488
rect 4613 6430 8083 6432
rect 4613 6427 4679 6430
rect 8017 6427 8083 6430
rect 9990 6428 9996 6492
rect 10060 6490 10066 6492
rect 10060 6430 13186 6490
rect 10060 6428 10066 6430
rect 4613 6354 4679 6357
rect 11789 6354 11855 6357
rect 4613 6352 11855 6354
rect 4613 6296 4618 6352
rect 4674 6296 11794 6352
rect 11850 6296 11855 6352
rect 4613 6294 11855 6296
rect 4613 6291 4679 6294
rect 11789 6291 11855 6294
rect 12065 6354 12131 6357
rect 12249 6354 12315 6357
rect 12065 6352 12315 6354
rect 12065 6296 12070 6352
rect 12126 6296 12254 6352
rect 12310 6296 12315 6352
rect 12065 6294 12315 6296
rect 13126 6354 13186 6430
rect 14089 6354 14155 6357
rect 13126 6352 14155 6354
rect 13126 6296 14094 6352
rect 14150 6296 14155 6352
rect 13126 6294 14155 6296
rect 12065 6291 12131 6294
rect 12249 6291 12315 6294
rect 14089 6291 14155 6294
rect 2773 6218 2839 6221
rect 12801 6218 12867 6221
rect 2773 6216 12867 6218
rect 2773 6160 2778 6216
rect 2834 6160 12806 6216
rect 12862 6160 12867 6216
rect 2773 6158 12867 6160
rect 2773 6155 2839 6158
rect 12801 6155 12867 6158
rect 13445 6218 13511 6221
rect 13670 6218 13676 6220
rect 13445 6216 13676 6218
rect 13445 6160 13450 6216
rect 13506 6160 13676 6216
rect 13445 6158 13676 6160
rect 13445 6155 13511 6158
rect 13670 6156 13676 6158
rect 13740 6156 13746 6220
rect 13905 6218 13971 6221
rect 15009 6218 15075 6221
rect 13905 6216 15075 6218
rect 13905 6160 13910 6216
rect 13966 6160 15014 6216
rect 15070 6160 15075 6216
rect 13905 6158 15075 6160
rect 13905 6155 13971 6158
rect 15009 6155 15075 6158
rect 7649 6082 7715 6085
rect 11513 6084 11579 6085
rect 11462 6082 11468 6084
rect 7649 6080 10656 6082
rect 7649 6024 7654 6080
rect 7710 6024 10656 6080
rect 7649 6022 10656 6024
rect 11386 6022 11468 6082
rect 11532 6082 11579 6084
rect 12249 6082 12315 6085
rect 12525 6084 12591 6085
rect 12525 6082 12572 6084
rect 11532 6080 12315 6082
rect 11574 6024 12254 6080
rect 12310 6024 12315 6080
rect 7649 6019 7715 6022
rect 5874 6016 6194 6017
rect 5874 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6122 6016
rect 6186 5952 6194 6016
rect 5874 5951 6194 5952
rect 4470 5884 4476 5948
rect 4540 5946 4546 5948
rect 5717 5946 5783 5949
rect 4540 5944 5783 5946
rect 4540 5888 5722 5944
rect 5778 5888 5783 5944
rect 4540 5886 5783 5888
rect 4540 5884 4546 5886
rect 5717 5883 5783 5886
rect 7189 5946 7255 5949
rect 7414 5946 7420 5948
rect 7189 5944 7420 5946
rect 7189 5888 7194 5944
rect 7250 5888 7420 5944
rect 7189 5886 7420 5888
rect 7189 5883 7255 5886
rect 7414 5884 7420 5886
rect 7484 5946 7490 5948
rect 8569 5946 8635 5949
rect 9254 5946 9260 5948
rect 7484 5944 9260 5946
rect 7484 5888 8574 5944
rect 8630 5888 9260 5944
rect 7484 5886 9260 5888
rect 7484 5884 7490 5886
rect 8569 5883 8635 5886
rect 9254 5884 9260 5886
rect 9324 5884 9330 5948
rect 1393 5810 1459 5813
rect 4102 5810 4108 5812
rect 1393 5808 4108 5810
rect 1393 5752 1398 5808
rect 1454 5752 4108 5808
rect 1393 5750 4108 5752
rect 1393 5747 1459 5750
rect 4102 5748 4108 5750
rect 4172 5748 4178 5812
rect 4797 5810 4863 5813
rect 10225 5810 10291 5813
rect 4797 5808 10291 5810
rect 4797 5752 4802 5808
rect 4858 5752 10230 5808
rect 10286 5752 10291 5808
rect 4797 5750 10291 5752
rect 10596 5810 10656 6022
rect 11462 6020 11468 6022
rect 11532 6022 12315 6024
rect 12480 6080 12572 6082
rect 12480 6024 12530 6080
rect 12480 6022 12572 6024
rect 11532 6020 11579 6022
rect 11513 6019 11579 6020
rect 12249 6019 12315 6022
rect 12525 6020 12572 6022
rect 12636 6020 12642 6084
rect 12525 6019 12591 6020
rect 10805 6016 11125 6017
rect 10805 5952 10813 6016
rect 10877 5952 10893 6016
rect 10957 5952 10973 6016
rect 11037 5952 11053 6016
rect 11117 5952 11125 6016
rect 10805 5951 11125 5952
rect 12801 5946 12867 5949
rect 11240 5944 12867 5946
rect 11240 5888 12806 5944
rect 12862 5888 12867 5944
rect 11240 5886 12867 5888
rect 11240 5810 11300 5886
rect 12801 5883 12867 5886
rect 12382 5810 12388 5812
rect 10596 5750 11300 5810
rect 11470 5750 12388 5810
rect 4797 5747 4863 5750
rect 10225 5747 10291 5750
rect 0 5674 480 5704
rect 3693 5674 3759 5677
rect 0 5672 3759 5674
rect 0 5616 3698 5672
rect 3754 5616 3759 5672
rect 0 5614 3759 5616
rect 0 5584 480 5614
rect 3693 5611 3759 5614
rect 4705 5674 4771 5677
rect 5901 5674 5967 5677
rect 7005 5676 7071 5677
rect 7005 5674 7052 5676
rect 4705 5672 5967 5674
rect 4705 5616 4710 5672
rect 4766 5616 5906 5672
rect 5962 5616 5967 5672
rect 4705 5614 5967 5616
rect 6960 5672 7052 5674
rect 6960 5616 7010 5672
rect 6960 5614 7052 5616
rect 4705 5611 4771 5614
rect 5901 5611 5967 5614
rect 7005 5612 7052 5614
rect 7116 5612 7122 5676
rect 7281 5674 7347 5677
rect 9581 5674 9647 5677
rect 11053 5674 11119 5677
rect 7281 5672 8908 5674
rect 7281 5616 7286 5672
rect 7342 5616 8908 5672
rect 7281 5614 8908 5616
rect 7005 5611 7071 5612
rect 7281 5611 7347 5614
rect 4429 5538 4495 5541
rect 6269 5538 6335 5541
rect 4429 5536 6335 5538
rect 4429 5480 4434 5536
rect 4490 5480 6274 5536
rect 6330 5480 6335 5536
rect 4429 5478 6335 5480
rect 4429 5475 4495 5478
rect 6269 5475 6335 5478
rect 6494 5476 6500 5540
rect 6564 5538 6570 5540
rect 7833 5538 7899 5541
rect 6564 5536 7899 5538
rect 6564 5480 7838 5536
rect 7894 5480 7899 5536
rect 6564 5478 7899 5480
rect 8848 5538 8908 5614
rect 9581 5672 11119 5674
rect 9581 5616 9586 5672
rect 9642 5616 11058 5672
rect 11114 5616 11119 5672
rect 9581 5614 11119 5616
rect 9581 5611 9647 5614
rect 11053 5611 11119 5614
rect 11237 5674 11303 5677
rect 11470 5674 11530 5750
rect 12382 5748 12388 5750
rect 12452 5748 12458 5812
rect 12893 5810 12959 5813
rect 13670 5810 13676 5812
rect 12893 5808 13676 5810
rect 12893 5752 12898 5808
rect 12954 5752 13676 5808
rect 12893 5750 13676 5752
rect 12893 5747 12959 5750
rect 13670 5748 13676 5750
rect 13740 5748 13746 5812
rect 11237 5672 11530 5674
rect 11237 5616 11242 5672
rect 11298 5616 11530 5672
rect 11237 5614 11530 5616
rect 11237 5611 11303 5614
rect 12014 5612 12020 5676
rect 12084 5674 12090 5676
rect 12433 5674 12499 5677
rect 12084 5672 12499 5674
rect 12084 5616 12438 5672
rect 12494 5616 12499 5672
rect 12084 5614 12499 5616
rect 12084 5612 12090 5614
rect 12433 5611 12499 5614
rect 12566 5612 12572 5676
rect 12636 5674 12642 5676
rect 13813 5674 13879 5677
rect 12636 5672 13879 5674
rect 12636 5616 13818 5672
rect 13874 5616 13879 5672
rect 12636 5614 13879 5616
rect 12636 5612 12642 5614
rect 13813 5611 13879 5614
rect 11973 5538 12039 5541
rect 8848 5536 12039 5538
rect 8848 5480 11978 5536
rect 12034 5480 12039 5536
rect 8848 5478 12039 5480
rect 6564 5476 6570 5478
rect 7833 5475 7899 5478
rect 11973 5475 12039 5478
rect 12198 5476 12204 5540
rect 12268 5538 12274 5540
rect 12893 5538 12959 5541
rect 12268 5536 12959 5538
rect 12268 5480 12898 5536
rect 12954 5480 12959 5536
rect 12268 5478 12959 5480
rect 12268 5476 12274 5478
rect 12893 5475 12959 5478
rect 3409 5472 3729 5473
rect 3409 5408 3417 5472
rect 3481 5408 3497 5472
rect 3561 5408 3577 5472
rect 3641 5408 3657 5472
rect 3721 5408 3729 5472
rect 3409 5407 3729 5408
rect 8340 5472 8660 5473
rect 8340 5408 8348 5472
rect 8412 5408 8428 5472
rect 8492 5408 8508 5472
rect 8572 5408 8588 5472
rect 8652 5408 8660 5472
rect 8340 5407 8660 5408
rect 13270 5472 13590 5473
rect 13270 5408 13278 5472
rect 13342 5408 13358 5472
rect 13422 5408 13438 5472
rect 13502 5408 13518 5472
rect 13582 5408 13590 5472
rect 13270 5407 13590 5408
rect 3877 5402 3943 5405
rect 7741 5402 7807 5405
rect 3877 5400 7807 5402
rect 3877 5344 3882 5400
rect 3938 5344 7746 5400
rect 7802 5344 7807 5400
rect 3877 5342 7807 5344
rect 3877 5339 3943 5342
rect 7741 5339 7807 5342
rect 8886 5340 8892 5404
rect 8956 5402 8962 5404
rect 12617 5402 12683 5405
rect 12985 5402 13051 5405
rect 8956 5400 13051 5402
rect 8956 5344 12622 5400
rect 12678 5344 12990 5400
rect 13046 5344 13051 5400
rect 8956 5342 13051 5344
rect 8956 5340 8962 5342
rect 12617 5339 12683 5342
rect 12985 5339 13051 5342
rect 3509 5266 3575 5269
rect 13854 5266 13860 5268
rect 3509 5264 13860 5266
rect 3509 5208 3514 5264
rect 3570 5208 13860 5264
rect 3509 5206 13860 5208
rect 3509 5203 3575 5206
rect 13854 5204 13860 5206
rect 13924 5204 13930 5268
rect 1853 5130 1919 5133
rect 12893 5130 12959 5133
rect 1853 5128 12959 5130
rect 1853 5072 1858 5128
rect 1914 5072 12898 5128
rect 12954 5072 12959 5128
rect 1853 5070 12959 5072
rect 1853 5067 1919 5070
rect 12893 5067 12959 5070
rect 4153 4994 4219 4997
rect 5349 4994 5415 4997
rect 4153 4992 5415 4994
rect 4153 4936 4158 4992
rect 4214 4936 5354 4992
rect 5410 4936 5415 4992
rect 4153 4934 5415 4936
rect 4153 4931 4219 4934
rect 5349 4931 5415 4934
rect 6678 4932 6684 4996
rect 6748 4994 6754 4996
rect 7005 4994 7071 4997
rect 6748 4992 7071 4994
rect 6748 4936 7010 4992
rect 7066 4936 7071 4992
rect 6748 4934 7071 4936
rect 6748 4932 6754 4934
rect 7005 4931 7071 4934
rect 7465 4994 7531 4997
rect 9305 4994 9371 4997
rect 7465 4992 9371 4994
rect 7465 4936 7470 4992
rect 7526 4936 9310 4992
rect 9366 4936 9371 4992
rect 7465 4934 9371 4936
rect 7465 4931 7531 4934
rect 9305 4931 9371 4934
rect 11513 4994 11579 4997
rect 11830 4994 11836 4996
rect 11513 4992 11836 4994
rect 11513 4936 11518 4992
rect 11574 4936 11836 4992
rect 11513 4934 11836 4936
rect 11513 4931 11579 4934
rect 11830 4932 11836 4934
rect 11900 4932 11906 4996
rect 11973 4994 12039 4997
rect 13997 4994 14063 4997
rect 11973 4992 14063 4994
rect 11973 4936 11978 4992
rect 12034 4936 14002 4992
rect 14058 4936 14063 4992
rect 11973 4934 14063 4936
rect 11973 4931 12039 4934
rect 13997 4931 14063 4934
rect 5874 4928 6194 4929
rect 5874 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6122 4928
rect 6186 4864 6194 4928
rect 5874 4863 6194 4864
rect 10805 4928 11125 4929
rect 10805 4864 10813 4928
rect 10877 4864 10893 4928
rect 10957 4864 10973 4928
rect 11037 4864 11053 4928
rect 11117 4864 11125 4928
rect 10805 4863 11125 4864
rect 2773 4858 2839 4861
rect 5206 4858 5212 4860
rect 2773 4856 5212 4858
rect 2773 4800 2778 4856
rect 2834 4800 5212 4856
rect 2773 4798 5212 4800
rect 2773 4795 2839 4798
rect 5206 4796 5212 4798
rect 5276 4796 5282 4860
rect 6453 4858 6519 4861
rect 6729 4858 6795 4861
rect 6453 4856 6795 4858
rect 6453 4800 6458 4856
rect 6514 4800 6734 4856
rect 6790 4800 6795 4856
rect 6453 4798 6795 4800
rect 6453 4795 6519 4798
rect 6729 4795 6795 4798
rect 7741 4858 7807 4861
rect 10358 4858 10364 4860
rect 7741 4856 10364 4858
rect 7741 4800 7746 4856
rect 7802 4800 10364 4856
rect 7741 4798 10364 4800
rect 7741 4795 7807 4798
rect 10358 4796 10364 4798
rect 10428 4796 10434 4860
rect 11697 4858 11763 4861
rect 11830 4858 11836 4860
rect 11697 4856 11836 4858
rect 11697 4800 11702 4856
rect 11758 4800 11836 4856
rect 11697 4798 11836 4800
rect 11697 4795 11763 4798
rect 11830 4796 11836 4798
rect 11900 4796 11906 4860
rect 12065 4858 12131 4861
rect 13721 4858 13787 4861
rect 12065 4856 13787 4858
rect 12065 4800 12070 4856
rect 12126 4800 13726 4856
rect 13782 4800 13787 4856
rect 12065 4798 13787 4800
rect 12065 4795 12131 4798
rect 13721 4795 13787 4798
rect 14641 4858 14707 4861
rect 14774 4858 14780 4860
rect 14641 4856 14780 4858
rect 14641 4800 14646 4856
rect 14702 4800 14780 4856
rect 14641 4798 14780 4800
rect 14641 4795 14707 4798
rect 14774 4796 14780 4798
rect 14844 4796 14850 4860
rect 0 4722 480 4752
rect 1853 4722 1919 4725
rect 0 4720 1919 4722
rect 0 4664 1858 4720
rect 1914 4664 1919 4720
rect 0 4662 1919 4664
rect 0 4632 480 4662
rect 1853 4659 1919 4662
rect 2037 4722 2103 4725
rect 13537 4722 13603 4725
rect 2037 4720 13603 4722
rect 2037 4664 2042 4720
rect 2098 4664 13542 4720
rect 13598 4664 13603 4720
rect 2037 4662 13603 4664
rect 2037 4659 2103 4662
rect 13537 4659 13603 4662
rect 2957 4586 3023 4589
rect 12985 4586 13051 4589
rect 2957 4584 13051 4586
rect 2957 4528 2962 4584
rect 3018 4528 12990 4584
rect 13046 4528 13051 4584
rect 2957 4526 13051 4528
rect 2957 4523 3023 4526
rect 12985 4523 13051 4526
rect 2957 4450 3023 4453
rect 3233 4450 3299 4453
rect 7465 4450 7531 4453
rect 7649 4450 7715 4453
rect 2957 4448 3299 4450
rect 2957 4392 2962 4448
rect 3018 4392 3238 4448
rect 3294 4392 3299 4448
rect 2957 4390 3299 4392
rect 2957 4387 3023 4390
rect 3233 4387 3299 4390
rect 4156 4448 7715 4450
rect 4156 4392 7470 4448
rect 7526 4392 7654 4448
rect 7710 4392 7715 4448
rect 4156 4390 7715 4392
rect 3409 4384 3729 4385
rect 3409 4320 3417 4384
rect 3481 4320 3497 4384
rect 3561 4320 3577 4384
rect 3641 4320 3657 4384
rect 3721 4320 3729 4384
rect 3409 4319 3729 4320
rect 1393 4178 1459 4181
rect 4156 4178 4216 4390
rect 7465 4387 7531 4390
rect 7649 4387 7715 4390
rect 9070 4388 9076 4452
rect 9140 4450 9146 4452
rect 9305 4450 9371 4453
rect 9140 4448 9371 4450
rect 9140 4392 9310 4448
rect 9366 4392 9371 4448
rect 9140 4390 9371 4392
rect 9140 4388 9146 4390
rect 9305 4387 9371 4390
rect 9622 4388 9628 4452
rect 9692 4388 9698 4452
rect 9990 4388 9996 4452
rect 10060 4450 10066 4452
rect 10409 4450 10475 4453
rect 10060 4448 10475 4450
rect 10060 4392 10414 4448
rect 10470 4392 10475 4448
rect 10060 4390 10475 4392
rect 10060 4388 10066 4390
rect 8340 4384 8660 4385
rect 8340 4320 8348 4384
rect 8412 4320 8428 4384
rect 8492 4320 8508 4384
rect 8572 4320 8588 4384
rect 8652 4320 8660 4384
rect 8340 4319 8660 4320
rect 4337 4314 4403 4317
rect 4470 4314 4476 4316
rect 4337 4312 4476 4314
rect 4337 4256 4342 4312
rect 4398 4256 4476 4312
rect 4337 4254 4476 4256
rect 4337 4251 4403 4254
rect 4470 4252 4476 4254
rect 4540 4252 4546 4316
rect 4981 4314 5047 4317
rect 9121 4316 9187 4317
rect 4981 4312 8218 4314
rect 4981 4256 4986 4312
rect 5042 4256 8218 4312
rect 4981 4254 8218 4256
rect 4981 4251 5047 4254
rect 8017 4178 8083 4181
rect 1393 4176 4216 4178
rect 1393 4120 1398 4176
rect 1454 4120 4216 4176
rect 1393 4118 4216 4120
rect 4340 4176 8083 4178
rect 4340 4120 8022 4176
rect 8078 4120 8083 4176
rect 4340 4118 8083 4120
rect 8158 4178 8218 4254
rect 9070 4252 9076 4316
rect 9140 4314 9187 4316
rect 9630 4314 9690 4388
rect 10409 4387 10475 4390
rect 10542 4388 10548 4452
rect 10612 4450 10618 4452
rect 11789 4450 11855 4453
rect 10612 4448 11855 4450
rect 10612 4392 11794 4448
rect 11850 4392 11855 4448
rect 10612 4390 11855 4392
rect 10612 4388 10618 4390
rect 11789 4387 11855 4390
rect 12249 4450 12315 4453
rect 12893 4450 12959 4453
rect 12249 4448 12959 4450
rect 12249 4392 12254 4448
rect 12310 4392 12898 4448
rect 12954 4392 12959 4448
rect 12249 4390 12959 4392
rect 12249 4387 12315 4390
rect 12893 4387 12959 4390
rect 13270 4384 13590 4385
rect 13270 4320 13278 4384
rect 13342 4320 13358 4384
rect 13422 4320 13438 4384
rect 13502 4320 13518 4384
rect 13582 4320 13590 4384
rect 13270 4319 13590 4320
rect 9140 4312 9690 4314
rect 9182 4256 9690 4312
rect 9140 4254 9690 4256
rect 9857 4314 9923 4317
rect 11789 4314 11855 4317
rect 12014 4314 12020 4316
rect 9857 4312 11668 4314
rect 9857 4256 9862 4312
rect 9918 4256 11668 4312
rect 9857 4254 11668 4256
rect 9140 4252 9187 4254
rect 9121 4251 9187 4252
rect 9857 4251 9923 4254
rect 9489 4180 9555 4181
rect 8886 4178 8892 4180
rect 8158 4118 8892 4178
rect 1393 4115 1459 4118
rect 4340 4045 4400 4118
rect 8017 4115 8083 4118
rect 8886 4116 8892 4118
rect 8956 4116 8962 4180
rect 9438 4116 9444 4180
rect 9508 4178 9555 4180
rect 9765 4180 9831 4181
rect 9765 4178 9812 4180
rect 9508 4176 9600 4178
rect 9550 4120 9600 4176
rect 9508 4118 9600 4120
rect 9720 4176 9812 4178
rect 9720 4120 9770 4176
rect 9720 4118 9812 4120
rect 9508 4116 9555 4118
rect 9489 4115 9555 4116
rect 9765 4116 9812 4118
rect 9876 4116 9882 4180
rect 11608 4178 11668 4254
rect 11789 4312 12020 4314
rect 11789 4256 11794 4312
rect 11850 4256 12020 4312
rect 11789 4254 12020 4256
rect 11789 4251 11855 4254
rect 12014 4252 12020 4254
rect 12084 4252 12090 4316
rect 15009 4178 15075 4181
rect 10182 4118 11530 4178
rect 11608 4176 15075 4178
rect 11608 4120 15014 4176
rect 15070 4120 15075 4176
rect 11608 4118 15075 4120
rect 9765 4115 9831 4116
rect 4337 4040 4403 4045
rect 4337 3984 4342 4040
rect 4398 3984 4403 4040
rect 4337 3979 4403 3984
rect 5165 4042 5231 4045
rect 10182 4042 10242 4118
rect 5165 4040 10242 4042
rect 5165 3984 5170 4040
rect 5226 3984 10242 4040
rect 5165 3982 10242 3984
rect 5165 3979 5231 3982
rect 10358 3980 10364 4044
rect 10428 4042 10434 4044
rect 10777 4042 10843 4045
rect 11470 4042 11530 4118
rect 15009 4115 15075 4118
rect 12525 4042 12591 4045
rect 10428 4040 11392 4042
rect 10428 3984 10782 4040
rect 10838 3984 11392 4040
rect 10428 3982 11392 3984
rect 11470 4040 12591 4042
rect 11470 3984 12530 4040
rect 12586 3984 12591 4040
rect 11470 3982 12591 3984
rect 10428 3980 10434 3982
rect 10777 3979 10843 3982
rect 2037 3906 2103 3909
rect 4705 3906 4771 3909
rect 5441 3908 5507 3909
rect 5390 3906 5396 3908
rect 2037 3904 4771 3906
rect 2037 3848 2042 3904
rect 2098 3848 4710 3904
rect 4766 3848 4771 3904
rect 2037 3846 4771 3848
rect 5350 3846 5396 3906
rect 5460 3904 5507 3908
rect 5502 3848 5507 3904
rect 2037 3843 2103 3846
rect 4705 3843 4771 3846
rect 5390 3844 5396 3846
rect 5460 3844 5507 3848
rect 5441 3843 5507 3844
rect 6361 3906 6427 3909
rect 6494 3906 6500 3908
rect 6361 3904 6500 3906
rect 6361 3848 6366 3904
rect 6422 3848 6500 3904
rect 6361 3846 6500 3848
rect 6361 3843 6427 3846
rect 6494 3844 6500 3846
rect 6564 3844 6570 3908
rect 7097 3906 7163 3909
rect 10542 3906 10548 3908
rect 7097 3904 10548 3906
rect 7097 3848 7102 3904
rect 7158 3848 10548 3904
rect 7097 3846 10548 3848
rect 7097 3843 7163 3846
rect 10542 3844 10548 3846
rect 10612 3844 10618 3908
rect 11332 3906 11392 3982
rect 12525 3979 12591 3982
rect 13905 4042 13971 4045
rect 14406 4042 14412 4044
rect 13905 4040 14412 4042
rect 13905 3984 13910 4040
rect 13966 3984 14412 4040
rect 13905 3982 14412 3984
rect 13905 3979 13971 3982
rect 14406 3980 14412 3982
rect 14476 3980 14482 4044
rect 11513 3906 11579 3909
rect 11332 3904 11579 3906
rect 11332 3848 11518 3904
rect 11574 3848 11579 3904
rect 11332 3846 11579 3848
rect 11513 3843 11579 3846
rect 11697 3906 11763 3909
rect 12249 3906 12315 3909
rect 11697 3904 12315 3906
rect 11697 3848 11702 3904
rect 11758 3848 12254 3904
rect 12310 3848 12315 3904
rect 11697 3846 12315 3848
rect 11697 3843 11763 3846
rect 12249 3843 12315 3846
rect 13721 3906 13787 3909
rect 15009 3906 15075 3909
rect 13721 3904 15075 3906
rect 13721 3848 13726 3904
rect 13782 3848 15014 3904
rect 15070 3848 15075 3904
rect 13721 3846 15075 3848
rect 13721 3843 13787 3846
rect 15009 3843 15075 3846
rect 5874 3840 6194 3841
rect 5874 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6122 3840
rect 6186 3776 6194 3840
rect 5874 3775 6194 3776
rect 10805 3840 11125 3841
rect 10805 3776 10813 3840
rect 10877 3776 10893 3840
rect 10957 3776 10973 3840
rect 11037 3776 11053 3840
rect 11117 3776 11125 3840
rect 10805 3775 11125 3776
rect 3182 3708 3188 3772
rect 3252 3770 3258 3772
rect 3417 3770 3483 3773
rect 5441 3770 5507 3773
rect 3252 3768 5507 3770
rect 3252 3712 3422 3768
rect 3478 3712 5446 3768
rect 5502 3712 5507 3768
rect 3252 3710 5507 3712
rect 3252 3708 3258 3710
rect 3417 3707 3483 3710
rect 5441 3707 5507 3710
rect 6269 3770 6335 3773
rect 7649 3770 7715 3773
rect 6269 3768 7715 3770
rect 6269 3712 6274 3768
rect 6330 3712 7654 3768
rect 7710 3712 7715 3768
rect 6269 3710 7715 3712
rect 6269 3707 6335 3710
rect 7649 3707 7715 3710
rect 8150 3708 8156 3772
rect 8220 3770 8226 3772
rect 10225 3770 10291 3773
rect 11973 3772 12039 3773
rect 11973 3770 12020 3772
rect 8220 3768 10291 3770
rect 8220 3712 10230 3768
rect 10286 3712 10291 3768
rect 8220 3710 10291 3712
rect 11928 3768 12020 3770
rect 11928 3712 11978 3768
rect 11928 3710 12020 3712
rect 8220 3708 8226 3710
rect 10225 3707 10291 3710
rect 11973 3708 12020 3710
rect 12084 3708 12090 3772
rect 12382 3708 12388 3772
rect 12452 3770 12458 3772
rect 13261 3770 13327 3773
rect 14457 3770 14523 3773
rect 12452 3710 13186 3770
rect 12452 3708 12458 3710
rect 11973 3707 12039 3708
rect 0 3634 480 3664
rect 13126 3637 13186 3710
rect 13261 3768 14523 3770
rect 13261 3712 13266 3768
rect 13322 3712 14462 3768
rect 14518 3712 14523 3768
rect 13261 3710 14523 3712
rect 13261 3707 13327 3710
rect 14457 3707 14523 3710
rect 1301 3634 1367 3637
rect 0 3632 1367 3634
rect 0 3576 1306 3632
rect 1362 3576 1367 3632
rect 0 3574 1367 3576
rect 0 3544 480 3574
rect 1301 3571 1367 3574
rect 3601 3634 3667 3637
rect 7005 3634 7071 3637
rect 12433 3634 12499 3637
rect 3601 3632 7071 3634
rect 3601 3576 3606 3632
rect 3662 3576 7010 3632
rect 7066 3576 7071 3632
rect 3601 3574 7071 3576
rect 3601 3571 3667 3574
rect 7005 3571 7071 3574
rect 7560 3632 12499 3634
rect 7560 3576 12438 3632
rect 12494 3576 12499 3632
rect 7560 3574 12499 3576
rect 13126 3632 13235 3637
rect 13126 3576 13174 3632
rect 13230 3576 13235 3632
rect 13126 3574 13235 3576
rect 2313 3498 2379 3501
rect 7560 3498 7620 3574
rect 12433 3571 12499 3574
rect 13169 3571 13235 3574
rect 9121 3498 9187 3501
rect 13629 3498 13695 3501
rect 2313 3496 7620 3498
rect 2313 3440 2318 3496
rect 2374 3440 7620 3496
rect 2313 3438 7620 3440
rect 7790 3438 8954 3498
rect 2313 3435 2379 3438
rect 4429 3362 4495 3365
rect 6729 3362 6795 3365
rect 4429 3360 6795 3362
rect 4429 3304 4434 3360
rect 4490 3304 6734 3360
rect 6790 3304 6795 3360
rect 4429 3302 6795 3304
rect 4429 3299 4495 3302
rect 6729 3299 6795 3302
rect 6913 3362 6979 3365
rect 7790 3362 7850 3438
rect 6913 3360 7850 3362
rect 6913 3304 6918 3360
rect 6974 3304 7850 3360
rect 6913 3302 7850 3304
rect 8894 3362 8954 3438
rect 9121 3496 13695 3498
rect 9121 3440 9126 3496
rect 9182 3440 13634 3496
rect 13690 3440 13695 3496
rect 9121 3438 13695 3440
rect 9121 3435 9187 3438
rect 13629 3435 13695 3438
rect 11881 3362 11947 3365
rect 12249 3364 12315 3365
rect 8894 3360 11947 3362
rect 8894 3304 11886 3360
rect 11942 3304 11947 3360
rect 8894 3302 11947 3304
rect 6913 3299 6979 3302
rect 11881 3299 11947 3302
rect 12198 3300 12204 3364
rect 12268 3362 12315 3364
rect 12433 3362 12499 3365
rect 12566 3362 12572 3364
rect 12268 3360 12360 3362
rect 12310 3304 12360 3360
rect 12268 3302 12360 3304
rect 12433 3360 12572 3362
rect 12433 3304 12438 3360
rect 12494 3304 12572 3360
rect 12433 3302 12572 3304
rect 12268 3300 12315 3302
rect 12249 3299 12315 3300
rect 12433 3299 12499 3302
rect 12566 3300 12572 3302
rect 12636 3300 12642 3364
rect 3409 3296 3729 3297
rect 3409 3232 3417 3296
rect 3481 3232 3497 3296
rect 3561 3232 3577 3296
rect 3641 3232 3657 3296
rect 3721 3232 3729 3296
rect 3409 3231 3729 3232
rect 8340 3296 8660 3297
rect 8340 3232 8348 3296
rect 8412 3232 8428 3296
rect 8492 3232 8508 3296
rect 8572 3232 8588 3296
rect 8652 3232 8660 3296
rect 8340 3231 8660 3232
rect 13270 3296 13590 3297
rect 13270 3232 13278 3296
rect 13342 3232 13358 3296
rect 13422 3232 13438 3296
rect 13502 3232 13518 3296
rect 13582 3232 13590 3296
rect 13270 3231 13590 3232
rect 7189 3226 7255 3229
rect 3926 3224 7255 3226
rect 3926 3168 7194 3224
rect 7250 3168 7255 3224
rect 3926 3166 7255 3168
rect 1485 3090 1551 3093
rect 3926 3090 3986 3166
rect 7189 3163 7255 3166
rect 7557 3228 7623 3229
rect 7557 3224 7604 3228
rect 7668 3226 7674 3228
rect 8753 3226 8819 3229
rect 9673 3226 9739 3229
rect 7557 3168 7562 3224
rect 7557 3164 7604 3168
rect 7668 3166 7714 3226
rect 8753 3224 9739 3226
rect 8753 3168 8758 3224
rect 8814 3168 9678 3224
rect 9734 3168 9739 3224
rect 8753 3166 9739 3168
rect 7668 3164 7674 3166
rect 7557 3163 7623 3164
rect 8753 3163 8819 3166
rect 9673 3163 9739 3166
rect 9949 3226 10015 3229
rect 13118 3226 13124 3228
rect 9949 3224 13124 3226
rect 9949 3168 9954 3224
rect 10010 3168 13124 3224
rect 9949 3166 13124 3168
rect 9949 3163 10015 3166
rect 13118 3164 13124 3166
rect 13188 3164 13194 3228
rect 11605 3092 11671 3093
rect 1485 3088 3986 3090
rect 1485 3032 1490 3088
rect 1546 3032 3986 3088
rect 1485 3030 3986 3032
rect 4662 3030 11530 3090
rect 1485 3027 1551 3030
rect 4061 2954 4127 2957
rect 4662 2954 4722 3030
rect 4061 2952 4722 2954
rect 4061 2896 4066 2952
rect 4122 2896 4722 2952
rect 4061 2894 4722 2896
rect 4797 2954 4863 2957
rect 9121 2954 9187 2957
rect 4797 2952 9187 2954
rect 4797 2896 4802 2952
rect 4858 2896 9126 2952
rect 9182 2896 9187 2952
rect 4797 2894 9187 2896
rect 4061 2891 4127 2894
rect 4797 2891 4863 2894
rect 9121 2891 9187 2894
rect 10685 2954 10751 2957
rect 11278 2954 11284 2956
rect 10685 2952 11284 2954
rect 10685 2896 10690 2952
rect 10746 2896 11284 2952
rect 10685 2894 11284 2896
rect 10685 2891 10751 2894
rect 11278 2892 11284 2894
rect 11348 2892 11354 2956
rect 11470 2954 11530 3030
rect 11605 3088 11652 3092
rect 11716 3090 11722 3092
rect 11881 3090 11947 3093
rect 13261 3090 13327 3093
rect 11605 3032 11610 3088
rect 11605 3028 11652 3032
rect 11716 3030 11762 3090
rect 11881 3088 13327 3090
rect 11881 3032 11886 3088
rect 11942 3032 13266 3088
rect 13322 3032 13327 3088
rect 11881 3030 13327 3032
rect 11716 3028 11722 3030
rect 11605 3027 11671 3028
rect 11881 3027 11947 3030
rect 13261 3027 13327 3030
rect 13445 3090 13511 3093
rect 13670 3090 13676 3092
rect 13445 3088 13676 3090
rect 13445 3032 13450 3088
rect 13506 3032 13676 3088
rect 13445 3030 13676 3032
rect 13445 3027 13511 3030
rect 13670 3028 13676 3030
rect 13740 3028 13746 3092
rect 15377 3090 15443 3093
rect 16520 3090 17000 3120
rect 15377 3088 17000 3090
rect 15377 3032 15382 3088
rect 15438 3032 17000 3088
rect 15377 3030 17000 3032
rect 15377 3027 15443 3030
rect 16520 3000 17000 3030
rect 12249 2954 12315 2957
rect 11470 2952 12315 2954
rect 11470 2896 12254 2952
rect 12310 2896 12315 2952
rect 11470 2894 12315 2896
rect 12249 2891 12315 2894
rect 14181 2954 14247 2957
rect 14958 2954 14964 2956
rect 14181 2952 14964 2954
rect 14181 2896 14186 2952
rect 14242 2896 14964 2952
rect 14181 2894 14964 2896
rect 14181 2891 14247 2894
rect 14958 2892 14964 2894
rect 15028 2892 15034 2956
rect 6729 2818 6795 2821
rect 9438 2818 9444 2820
rect 6729 2816 9444 2818
rect 6729 2760 6734 2816
rect 6790 2760 9444 2816
rect 6729 2758 9444 2760
rect 6729 2755 6795 2758
rect 9438 2756 9444 2758
rect 9508 2756 9514 2820
rect 15929 2818 15995 2821
rect 11792 2816 15995 2818
rect 11792 2760 15934 2816
rect 15990 2760 15995 2816
rect 11792 2758 15995 2760
rect 5874 2752 6194 2753
rect 5874 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6122 2752
rect 6186 2688 6194 2752
rect 5874 2687 6194 2688
rect 10805 2752 11125 2753
rect 10805 2688 10813 2752
rect 10877 2688 10893 2752
rect 10957 2688 10973 2752
rect 11037 2688 11053 2752
rect 11117 2688 11125 2752
rect 10805 2687 11125 2688
rect 5165 2684 5231 2685
rect 5441 2684 5507 2685
rect 5165 2682 5212 2684
rect 5120 2680 5212 2682
rect 5120 2624 5170 2680
rect 5120 2622 5212 2624
rect 5165 2620 5212 2622
rect 5276 2620 5282 2684
rect 5390 2620 5396 2684
rect 5460 2682 5507 2684
rect 5460 2680 5552 2682
rect 5502 2624 5552 2680
rect 5460 2622 5552 2624
rect 5460 2620 5507 2622
rect 7782 2620 7788 2684
rect 7852 2682 7858 2684
rect 8201 2682 8267 2685
rect 8753 2682 8819 2685
rect 7852 2680 8267 2682
rect 7852 2624 8206 2680
rect 8262 2624 8267 2680
rect 7852 2622 8267 2624
rect 7852 2620 7858 2622
rect 5165 2619 5231 2620
rect 5441 2619 5507 2620
rect 0 2546 480 2576
rect 3601 2546 3667 2549
rect 0 2544 3667 2546
rect 0 2488 3606 2544
rect 3662 2488 3667 2544
rect 0 2486 3667 2488
rect 0 2456 480 2486
rect 3601 2483 3667 2486
rect 3877 2546 3943 2549
rect 6177 2546 6243 2549
rect 7790 2546 7850 2620
rect 8201 2619 8267 2622
rect 8388 2680 8819 2682
rect 8388 2624 8758 2680
rect 8814 2624 8819 2680
rect 8388 2622 8819 2624
rect 3877 2544 7850 2546
rect 3877 2488 3882 2544
rect 3938 2488 6182 2544
rect 6238 2488 7850 2544
rect 3877 2486 7850 2488
rect 8109 2546 8175 2549
rect 8388 2546 8448 2622
rect 8753 2619 8819 2622
rect 8886 2620 8892 2684
rect 8956 2682 8962 2684
rect 10409 2682 10475 2685
rect 8956 2680 10475 2682
rect 8956 2624 10414 2680
rect 10470 2624 10475 2680
rect 8956 2622 10475 2624
rect 8956 2620 8962 2622
rect 10409 2619 10475 2622
rect 11513 2682 11579 2685
rect 11792 2682 11852 2758
rect 15929 2755 15995 2758
rect 11513 2680 11852 2682
rect 11513 2624 11518 2680
rect 11574 2624 11852 2680
rect 11513 2622 11852 2624
rect 11513 2619 11579 2622
rect 12198 2620 12204 2684
rect 12268 2682 12274 2684
rect 13445 2682 13511 2685
rect 12268 2680 13511 2682
rect 12268 2624 13450 2680
rect 13506 2624 13511 2680
rect 12268 2622 13511 2624
rect 12268 2620 12274 2622
rect 13445 2619 13511 2622
rect 8109 2544 8448 2546
rect 8109 2488 8114 2544
rect 8170 2488 8448 2544
rect 8109 2486 8448 2488
rect 3877 2483 3943 2486
rect 6177 2483 6243 2486
rect 8109 2483 8175 2486
rect 9254 2484 9260 2548
rect 9324 2546 9330 2548
rect 11789 2546 11855 2549
rect 12014 2546 12020 2548
rect 9324 2544 12020 2546
rect 9324 2488 11794 2544
rect 11850 2488 12020 2544
rect 9324 2486 12020 2488
rect 9324 2484 9330 2486
rect 11789 2483 11855 2486
rect 12014 2484 12020 2486
rect 12084 2484 12090 2548
rect 12934 2484 12940 2548
rect 13004 2546 13010 2548
rect 13169 2546 13235 2549
rect 13004 2544 13235 2546
rect 13004 2488 13174 2544
rect 13230 2488 13235 2544
rect 13004 2486 13235 2488
rect 13004 2484 13010 2486
rect 13169 2483 13235 2486
rect 3509 2410 3575 2413
rect 6678 2410 6684 2412
rect 3509 2408 6684 2410
rect 3509 2352 3514 2408
rect 3570 2352 6684 2408
rect 3509 2350 6684 2352
rect 3509 2347 3575 2350
rect 6678 2348 6684 2350
rect 6748 2410 6754 2412
rect 7741 2410 7807 2413
rect 6748 2408 7807 2410
rect 6748 2352 7746 2408
rect 7802 2352 7807 2408
rect 6748 2350 7807 2352
rect 6748 2348 6754 2350
rect 7741 2347 7807 2350
rect 8109 2410 8175 2413
rect 12750 2410 12756 2412
rect 8109 2408 12756 2410
rect 8109 2352 8114 2408
rect 8170 2352 12756 2408
rect 8109 2350 12756 2352
rect 8109 2347 8175 2350
rect 12750 2348 12756 2350
rect 12820 2348 12826 2412
rect 14549 2410 14615 2413
rect 12896 2408 14615 2410
rect 12896 2352 14554 2408
rect 14610 2352 14615 2408
rect 12896 2350 14615 2352
rect 9121 2274 9187 2277
rect 12896 2274 12956 2350
rect 14549 2347 14615 2350
rect 9121 2272 12956 2274
rect 9121 2216 9126 2272
rect 9182 2216 12956 2272
rect 9121 2214 12956 2216
rect 9121 2211 9187 2214
rect 3409 2208 3729 2209
rect 3409 2144 3417 2208
rect 3481 2144 3497 2208
rect 3561 2144 3577 2208
rect 3641 2144 3657 2208
rect 3721 2144 3729 2208
rect 3409 2143 3729 2144
rect 8340 2208 8660 2209
rect 8340 2144 8348 2208
rect 8412 2144 8428 2208
rect 8492 2144 8508 2208
rect 8572 2144 8588 2208
rect 8652 2144 8660 2208
rect 8340 2143 8660 2144
rect 13270 2208 13590 2209
rect 13270 2144 13278 2208
rect 13342 2144 13358 2208
rect 13422 2144 13438 2208
rect 13502 2144 13518 2208
rect 13582 2144 13590 2208
rect 13270 2143 13590 2144
rect 9949 2138 10015 2141
rect 9492 2136 10015 2138
rect 9492 2080 9954 2136
rect 10010 2080 10015 2136
rect 9492 2078 10015 2080
rect 7833 2002 7899 2005
rect 9492 2002 9552 2078
rect 9949 2075 10015 2078
rect 11462 2076 11468 2140
rect 11532 2138 11538 2140
rect 12065 2138 12131 2141
rect 11532 2136 12131 2138
rect 11532 2080 12070 2136
rect 12126 2080 12131 2136
rect 11532 2078 12131 2080
rect 11532 2076 11538 2078
rect 12065 2075 12131 2078
rect 7833 2000 9552 2002
rect 7833 1944 7838 2000
rect 7894 1944 9552 2000
rect 7833 1942 9552 1944
rect 9673 2002 9739 2005
rect 15009 2002 15075 2005
rect 9673 2000 15075 2002
rect 9673 1944 9678 2000
rect 9734 1944 15014 2000
rect 15070 1944 15075 2000
rect 9673 1942 15075 1944
rect 7833 1939 7899 1942
rect 9673 1939 9739 1942
rect 15009 1939 15075 1942
rect 7097 1866 7163 1869
rect 14222 1866 14228 1868
rect 7097 1864 14228 1866
rect 7097 1808 7102 1864
rect 7158 1808 14228 1864
rect 7097 1806 14228 1808
rect 7097 1803 7163 1806
rect 14222 1804 14228 1806
rect 14292 1804 14298 1868
rect 9857 1730 9923 1733
rect 14733 1730 14799 1733
rect 9857 1728 14799 1730
rect 9857 1672 9862 1728
rect 9918 1672 14738 1728
rect 14794 1672 14799 1728
rect 9857 1670 14799 1672
rect 9857 1667 9923 1670
rect 14733 1667 14799 1670
rect 10685 1594 10751 1597
rect 11830 1594 11836 1596
rect 10685 1592 11836 1594
rect 10685 1536 10690 1592
rect 10746 1536 11836 1592
rect 10685 1534 11836 1536
rect 10685 1531 10751 1534
rect 11830 1532 11836 1534
rect 11900 1532 11906 1596
rect 0 1458 480 1488
rect 1669 1458 1735 1461
rect 0 1456 1735 1458
rect 0 1400 1674 1456
rect 1730 1400 1735 1456
rect 0 1398 1735 1400
rect 0 1368 480 1398
rect 1669 1395 1735 1398
rect 9070 1396 9076 1460
rect 9140 1458 9146 1460
rect 11237 1458 11303 1461
rect 9140 1456 11303 1458
rect 9140 1400 11242 1456
rect 11298 1400 11303 1456
rect 9140 1398 11303 1400
rect 9140 1396 9146 1398
rect 11237 1395 11303 1398
rect 0 506 480 536
rect 2773 506 2839 509
rect 0 504 2839 506
rect 0 448 2778 504
rect 2834 448 2839 504
rect 0 446 2839 448
rect 0 416 480 446
rect 2773 443 2839 446
<< via3 >>
rect 10180 15948 10244 16012
rect 5882 15804 5946 15808
rect 5882 15748 5886 15804
rect 5886 15748 5942 15804
rect 5942 15748 5946 15804
rect 5882 15744 5946 15748
rect 5962 15804 6026 15808
rect 5962 15748 5966 15804
rect 5966 15748 6022 15804
rect 6022 15748 6026 15804
rect 5962 15744 6026 15748
rect 6042 15804 6106 15808
rect 6042 15748 6046 15804
rect 6046 15748 6102 15804
rect 6102 15748 6106 15804
rect 6042 15744 6106 15748
rect 6122 15804 6186 15808
rect 6122 15748 6126 15804
rect 6126 15748 6182 15804
rect 6182 15748 6186 15804
rect 6122 15744 6186 15748
rect 10813 15804 10877 15808
rect 10813 15748 10817 15804
rect 10817 15748 10873 15804
rect 10873 15748 10877 15804
rect 10813 15744 10877 15748
rect 10893 15804 10957 15808
rect 10893 15748 10897 15804
rect 10897 15748 10953 15804
rect 10953 15748 10957 15804
rect 10893 15744 10957 15748
rect 10973 15804 11037 15808
rect 10973 15748 10977 15804
rect 10977 15748 11033 15804
rect 11033 15748 11037 15804
rect 10973 15744 11037 15748
rect 11053 15804 11117 15808
rect 11053 15748 11057 15804
rect 11057 15748 11113 15804
rect 11113 15748 11117 15804
rect 11053 15744 11117 15748
rect 12572 15540 12636 15604
rect 12940 15404 13004 15468
rect 7420 15328 7484 15332
rect 7420 15272 7470 15328
rect 7470 15272 7484 15328
rect 7420 15268 7484 15272
rect 3417 15260 3481 15264
rect 3417 15204 3421 15260
rect 3421 15204 3477 15260
rect 3477 15204 3481 15260
rect 3417 15200 3481 15204
rect 3497 15260 3561 15264
rect 3497 15204 3501 15260
rect 3501 15204 3557 15260
rect 3557 15204 3561 15260
rect 3497 15200 3561 15204
rect 3577 15260 3641 15264
rect 3577 15204 3581 15260
rect 3581 15204 3637 15260
rect 3637 15204 3641 15260
rect 3577 15200 3641 15204
rect 3657 15260 3721 15264
rect 3657 15204 3661 15260
rect 3661 15204 3717 15260
rect 3717 15204 3721 15260
rect 3657 15200 3721 15204
rect 8348 15260 8412 15264
rect 8348 15204 8352 15260
rect 8352 15204 8408 15260
rect 8408 15204 8412 15260
rect 8348 15200 8412 15204
rect 8428 15260 8492 15264
rect 8428 15204 8432 15260
rect 8432 15204 8488 15260
rect 8488 15204 8492 15260
rect 8428 15200 8492 15204
rect 8508 15260 8572 15264
rect 8508 15204 8512 15260
rect 8512 15204 8568 15260
rect 8568 15204 8572 15260
rect 8508 15200 8572 15204
rect 8588 15260 8652 15264
rect 8588 15204 8592 15260
rect 8592 15204 8648 15260
rect 8648 15204 8652 15260
rect 8588 15200 8652 15204
rect 13278 15260 13342 15264
rect 13278 15204 13282 15260
rect 13282 15204 13338 15260
rect 13338 15204 13342 15260
rect 13278 15200 13342 15204
rect 13358 15260 13422 15264
rect 13358 15204 13362 15260
rect 13362 15204 13418 15260
rect 13418 15204 13422 15260
rect 13358 15200 13422 15204
rect 13438 15260 13502 15264
rect 13438 15204 13442 15260
rect 13442 15204 13498 15260
rect 13498 15204 13502 15260
rect 13438 15200 13502 15204
rect 13518 15260 13582 15264
rect 13518 15204 13522 15260
rect 13522 15204 13578 15260
rect 13578 15204 13582 15260
rect 13518 15200 13582 15204
rect 6316 14996 6380 15060
rect 5882 14716 5946 14720
rect 5882 14660 5886 14716
rect 5886 14660 5942 14716
rect 5942 14660 5946 14716
rect 5882 14656 5946 14660
rect 5962 14716 6026 14720
rect 5962 14660 5966 14716
rect 5966 14660 6022 14716
rect 6022 14660 6026 14716
rect 5962 14656 6026 14660
rect 6042 14716 6106 14720
rect 6042 14660 6046 14716
rect 6046 14660 6102 14716
rect 6102 14660 6106 14716
rect 6042 14656 6106 14660
rect 6122 14716 6186 14720
rect 6122 14660 6126 14716
rect 6126 14660 6182 14716
rect 6182 14660 6186 14716
rect 6122 14656 6186 14660
rect 3188 14588 3252 14652
rect 6684 14588 6748 14652
rect 9076 14724 9140 14788
rect 10813 14716 10877 14720
rect 10813 14660 10817 14716
rect 10817 14660 10873 14716
rect 10873 14660 10877 14716
rect 10813 14656 10877 14660
rect 10893 14716 10957 14720
rect 10893 14660 10897 14716
rect 10897 14660 10953 14716
rect 10953 14660 10957 14716
rect 10893 14656 10957 14660
rect 10973 14716 11037 14720
rect 10973 14660 10977 14716
rect 10977 14660 11033 14716
rect 11033 14660 11037 14716
rect 10973 14656 11037 14660
rect 11053 14716 11117 14720
rect 11053 14660 11057 14716
rect 11057 14660 11113 14716
rect 11113 14660 11117 14716
rect 11053 14656 11117 14660
rect 9812 14512 9876 14516
rect 9812 14456 9826 14512
rect 9826 14456 9876 14512
rect 9812 14452 9876 14456
rect 11468 14588 11532 14652
rect 5580 14316 5644 14380
rect 9628 14180 9692 14244
rect 3417 14172 3481 14176
rect 3417 14116 3421 14172
rect 3421 14116 3477 14172
rect 3477 14116 3481 14172
rect 3417 14112 3481 14116
rect 3497 14172 3561 14176
rect 3497 14116 3501 14172
rect 3501 14116 3557 14172
rect 3557 14116 3561 14172
rect 3497 14112 3561 14116
rect 3577 14172 3641 14176
rect 3577 14116 3581 14172
rect 3581 14116 3637 14172
rect 3637 14116 3641 14172
rect 3577 14112 3641 14116
rect 3657 14172 3721 14176
rect 3657 14116 3661 14172
rect 3661 14116 3717 14172
rect 3717 14116 3721 14172
rect 3657 14112 3721 14116
rect 8348 14172 8412 14176
rect 8348 14116 8352 14172
rect 8352 14116 8408 14172
rect 8408 14116 8412 14172
rect 8348 14112 8412 14116
rect 8428 14172 8492 14176
rect 8428 14116 8432 14172
rect 8432 14116 8488 14172
rect 8488 14116 8492 14172
rect 8428 14112 8492 14116
rect 8508 14172 8572 14176
rect 8508 14116 8512 14172
rect 8512 14116 8568 14172
rect 8568 14116 8572 14172
rect 8508 14112 8572 14116
rect 8588 14172 8652 14176
rect 8588 14116 8592 14172
rect 8592 14116 8648 14172
rect 8648 14116 8652 14172
rect 8588 14112 8652 14116
rect 13278 14172 13342 14176
rect 13278 14116 13282 14172
rect 13282 14116 13338 14172
rect 13338 14116 13342 14172
rect 13278 14112 13342 14116
rect 13358 14172 13422 14176
rect 13358 14116 13362 14172
rect 13362 14116 13418 14172
rect 13418 14116 13422 14172
rect 13358 14112 13422 14116
rect 13438 14172 13502 14176
rect 13438 14116 13442 14172
rect 13442 14116 13498 14172
rect 13498 14116 13502 14172
rect 13438 14112 13502 14116
rect 13518 14172 13582 14176
rect 13518 14116 13522 14172
rect 13522 14116 13578 14172
rect 13578 14116 13582 14172
rect 13518 14112 13582 14116
rect 4476 14044 4540 14108
rect 9260 14104 9324 14108
rect 9260 14048 9310 14104
rect 9310 14048 9324 14104
rect 9260 14044 9324 14048
rect 10364 14044 10428 14108
rect 10548 14044 10612 14108
rect 6500 13636 6564 13700
rect 11836 13832 11900 13836
rect 11836 13776 11850 13832
rect 11850 13776 11900 13832
rect 11836 13772 11900 13776
rect 12388 13832 12452 13836
rect 12388 13776 12438 13832
rect 12438 13776 12452 13832
rect 12388 13772 12452 13776
rect 5882 13628 5946 13632
rect 5882 13572 5886 13628
rect 5886 13572 5942 13628
rect 5942 13572 5946 13628
rect 5882 13568 5946 13572
rect 5962 13628 6026 13632
rect 5962 13572 5966 13628
rect 5966 13572 6022 13628
rect 6022 13572 6026 13628
rect 5962 13568 6026 13572
rect 6042 13628 6106 13632
rect 6042 13572 6046 13628
rect 6046 13572 6102 13628
rect 6102 13572 6106 13628
rect 6042 13568 6106 13572
rect 6122 13628 6186 13632
rect 6122 13572 6126 13628
rect 6126 13572 6182 13628
rect 6182 13572 6186 13628
rect 6122 13568 6186 13572
rect 10813 13628 10877 13632
rect 10813 13572 10817 13628
rect 10817 13572 10873 13628
rect 10873 13572 10877 13628
rect 10813 13568 10877 13572
rect 10893 13628 10957 13632
rect 10893 13572 10897 13628
rect 10897 13572 10953 13628
rect 10953 13572 10957 13628
rect 10893 13568 10957 13572
rect 10973 13628 11037 13632
rect 10973 13572 10977 13628
rect 10977 13572 11033 13628
rect 11033 13572 11037 13628
rect 10973 13568 11037 13572
rect 11053 13628 11117 13632
rect 11053 13572 11057 13628
rect 11057 13572 11113 13628
rect 11113 13572 11117 13628
rect 11053 13568 11117 13572
rect 10548 13500 10612 13564
rect 12204 13500 12268 13564
rect 3417 13084 3481 13088
rect 3417 13028 3421 13084
rect 3421 13028 3477 13084
rect 3477 13028 3481 13084
rect 3417 13024 3481 13028
rect 3497 13084 3561 13088
rect 3497 13028 3501 13084
rect 3501 13028 3557 13084
rect 3557 13028 3561 13084
rect 3497 13024 3561 13028
rect 3577 13084 3641 13088
rect 3577 13028 3581 13084
rect 3581 13028 3637 13084
rect 3637 13028 3641 13084
rect 3577 13024 3641 13028
rect 3657 13084 3721 13088
rect 3657 13028 3661 13084
rect 3661 13028 3717 13084
rect 3717 13028 3721 13084
rect 3657 13024 3721 13028
rect 8348 13084 8412 13088
rect 8348 13028 8352 13084
rect 8352 13028 8408 13084
rect 8408 13028 8412 13084
rect 8348 13024 8412 13028
rect 8428 13084 8492 13088
rect 8428 13028 8432 13084
rect 8432 13028 8488 13084
rect 8488 13028 8492 13084
rect 8428 13024 8492 13028
rect 8508 13084 8572 13088
rect 8508 13028 8512 13084
rect 8512 13028 8568 13084
rect 8568 13028 8572 13084
rect 8508 13024 8572 13028
rect 8588 13084 8652 13088
rect 8588 13028 8592 13084
rect 8592 13028 8648 13084
rect 8648 13028 8652 13084
rect 8588 13024 8652 13028
rect 7236 12820 7300 12884
rect 9444 12956 9508 13020
rect 12020 13228 12084 13292
rect 13278 13084 13342 13088
rect 13278 13028 13282 13084
rect 13282 13028 13338 13084
rect 13338 13028 13342 13084
rect 13278 13024 13342 13028
rect 13358 13084 13422 13088
rect 13358 13028 13362 13084
rect 13362 13028 13418 13084
rect 13418 13028 13422 13084
rect 13358 13024 13422 13028
rect 13438 13084 13502 13088
rect 13438 13028 13442 13084
rect 13442 13028 13498 13084
rect 13498 13028 13502 13084
rect 13438 13024 13502 13028
rect 13518 13084 13582 13088
rect 13518 13028 13522 13084
rect 13522 13028 13578 13084
rect 13578 13028 13582 13084
rect 13518 13024 13582 13028
rect 13124 12880 13188 12884
rect 13124 12824 13174 12880
rect 13174 12824 13188 12880
rect 13124 12820 13188 12824
rect 4476 12608 4540 12612
rect 4476 12552 4490 12608
rect 4490 12552 4540 12608
rect 4476 12548 4540 12552
rect 8892 12548 8956 12612
rect 11652 12548 11716 12612
rect 12756 12548 12820 12612
rect 5882 12540 5946 12544
rect 5882 12484 5886 12540
rect 5886 12484 5942 12540
rect 5942 12484 5946 12540
rect 5882 12480 5946 12484
rect 5962 12540 6026 12544
rect 5962 12484 5966 12540
rect 5966 12484 6022 12540
rect 6022 12484 6026 12540
rect 5962 12480 6026 12484
rect 6042 12540 6106 12544
rect 6042 12484 6046 12540
rect 6046 12484 6102 12540
rect 6102 12484 6106 12540
rect 6042 12480 6106 12484
rect 6122 12540 6186 12544
rect 6122 12484 6126 12540
rect 6126 12484 6182 12540
rect 6182 12484 6186 12540
rect 6122 12480 6186 12484
rect 10813 12540 10877 12544
rect 10813 12484 10817 12540
rect 10817 12484 10873 12540
rect 10873 12484 10877 12540
rect 10813 12480 10877 12484
rect 10893 12540 10957 12544
rect 10893 12484 10897 12540
rect 10897 12484 10953 12540
rect 10953 12484 10957 12540
rect 10893 12480 10957 12484
rect 10973 12540 11037 12544
rect 10973 12484 10977 12540
rect 10977 12484 11033 12540
rect 11033 12484 11037 12540
rect 10973 12480 11037 12484
rect 11053 12540 11117 12544
rect 11053 12484 11057 12540
rect 11057 12484 11113 12540
rect 11113 12484 11117 12540
rect 11053 12480 11117 12484
rect 6684 12412 6748 12476
rect 9444 12472 9508 12476
rect 9444 12416 9458 12472
rect 9458 12416 9508 12472
rect 9444 12412 9508 12416
rect 5580 12004 5644 12068
rect 9260 12140 9324 12204
rect 9812 12140 9876 12204
rect 14412 12140 14476 12204
rect 11284 12004 11348 12068
rect 3417 11996 3481 12000
rect 3417 11940 3421 11996
rect 3421 11940 3477 11996
rect 3477 11940 3481 11996
rect 3417 11936 3481 11940
rect 3497 11996 3561 12000
rect 3497 11940 3501 11996
rect 3501 11940 3557 11996
rect 3557 11940 3561 11996
rect 3497 11936 3561 11940
rect 3577 11996 3641 12000
rect 3577 11940 3581 11996
rect 3581 11940 3637 11996
rect 3637 11940 3641 11996
rect 3577 11936 3641 11940
rect 3657 11996 3721 12000
rect 3657 11940 3661 11996
rect 3661 11940 3717 11996
rect 3717 11940 3721 11996
rect 3657 11936 3721 11940
rect 8348 11996 8412 12000
rect 8348 11940 8352 11996
rect 8352 11940 8408 11996
rect 8408 11940 8412 11996
rect 8348 11936 8412 11940
rect 8428 11996 8492 12000
rect 8428 11940 8432 11996
rect 8432 11940 8488 11996
rect 8488 11940 8492 11996
rect 8428 11936 8492 11940
rect 8508 11996 8572 12000
rect 8508 11940 8512 11996
rect 8512 11940 8568 11996
rect 8568 11940 8572 11996
rect 8508 11936 8572 11940
rect 8588 11996 8652 12000
rect 8588 11940 8592 11996
rect 8592 11940 8648 11996
rect 8648 11940 8652 11996
rect 8588 11936 8652 11940
rect 13278 11996 13342 12000
rect 13278 11940 13282 11996
rect 13282 11940 13338 11996
rect 13338 11940 13342 11996
rect 13278 11936 13342 11940
rect 13358 11996 13422 12000
rect 13358 11940 13362 11996
rect 13362 11940 13418 11996
rect 13418 11940 13422 11996
rect 13358 11936 13422 11940
rect 13438 11996 13502 12000
rect 13438 11940 13442 11996
rect 13442 11940 13498 11996
rect 13498 11940 13502 11996
rect 13438 11936 13502 11940
rect 13518 11996 13582 12000
rect 13518 11940 13522 11996
rect 13522 11940 13578 11996
rect 13578 11940 13582 11996
rect 13518 11936 13582 11940
rect 9076 11868 9140 11932
rect 9628 11868 9692 11932
rect 10364 11868 10428 11932
rect 9996 11732 10060 11796
rect 10364 11792 10428 11796
rect 10364 11736 10414 11792
rect 10414 11736 10428 11792
rect 10364 11732 10428 11736
rect 11652 11460 11716 11524
rect 5882 11452 5946 11456
rect 5882 11396 5886 11452
rect 5886 11396 5942 11452
rect 5942 11396 5946 11452
rect 5882 11392 5946 11396
rect 5962 11452 6026 11456
rect 5962 11396 5966 11452
rect 5966 11396 6022 11452
rect 6022 11396 6026 11452
rect 5962 11392 6026 11396
rect 6042 11452 6106 11456
rect 6042 11396 6046 11452
rect 6046 11396 6102 11452
rect 6102 11396 6106 11452
rect 6042 11392 6106 11396
rect 6122 11452 6186 11456
rect 6122 11396 6126 11452
rect 6126 11396 6182 11452
rect 6182 11396 6186 11452
rect 6122 11392 6186 11396
rect 10813 11452 10877 11456
rect 10813 11396 10817 11452
rect 10817 11396 10873 11452
rect 10873 11396 10877 11452
rect 10813 11392 10877 11396
rect 10893 11452 10957 11456
rect 10893 11396 10897 11452
rect 10897 11396 10953 11452
rect 10953 11396 10957 11452
rect 10893 11392 10957 11396
rect 10973 11452 11037 11456
rect 10973 11396 10977 11452
rect 10977 11396 11033 11452
rect 11033 11396 11037 11452
rect 10973 11392 11037 11396
rect 11053 11452 11117 11456
rect 11053 11396 11057 11452
rect 11057 11396 11113 11452
rect 11113 11396 11117 11452
rect 11053 11392 11117 11396
rect 7788 11324 7852 11388
rect 11652 11188 11716 11252
rect 14964 11188 15028 11252
rect 14044 11112 14108 11116
rect 14044 11056 14094 11112
rect 14094 11056 14108 11112
rect 14044 11052 14108 11056
rect 7420 10916 7484 10980
rect 9628 10916 9692 10980
rect 3417 10908 3481 10912
rect 3417 10852 3421 10908
rect 3421 10852 3477 10908
rect 3477 10852 3481 10908
rect 3417 10848 3481 10852
rect 3497 10908 3561 10912
rect 3497 10852 3501 10908
rect 3501 10852 3557 10908
rect 3557 10852 3561 10908
rect 3497 10848 3561 10852
rect 3577 10908 3641 10912
rect 3577 10852 3581 10908
rect 3581 10852 3637 10908
rect 3637 10852 3641 10908
rect 3577 10848 3641 10852
rect 3657 10908 3721 10912
rect 3657 10852 3661 10908
rect 3661 10852 3717 10908
rect 3717 10852 3721 10908
rect 3657 10848 3721 10852
rect 8348 10908 8412 10912
rect 8348 10852 8352 10908
rect 8352 10852 8408 10908
rect 8408 10852 8412 10908
rect 8348 10848 8412 10852
rect 8428 10908 8492 10912
rect 8428 10852 8432 10908
rect 8432 10852 8488 10908
rect 8488 10852 8492 10908
rect 8428 10848 8492 10852
rect 8508 10908 8572 10912
rect 8508 10852 8512 10908
rect 8512 10852 8568 10908
rect 8568 10852 8572 10908
rect 8508 10848 8572 10852
rect 8588 10908 8652 10912
rect 8588 10852 8592 10908
rect 8592 10852 8648 10908
rect 8648 10852 8652 10908
rect 8588 10848 8652 10852
rect 13278 10908 13342 10912
rect 13278 10852 13282 10908
rect 13282 10852 13338 10908
rect 13338 10852 13342 10908
rect 13278 10848 13342 10852
rect 13358 10908 13422 10912
rect 13358 10852 13362 10908
rect 13362 10852 13418 10908
rect 13418 10852 13422 10908
rect 13358 10848 13422 10852
rect 13438 10908 13502 10912
rect 13438 10852 13442 10908
rect 13442 10852 13498 10908
rect 13498 10852 13502 10908
rect 13438 10848 13502 10852
rect 13518 10908 13582 10912
rect 13518 10852 13522 10908
rect 13522 10852 13578 10908
rect 13578 10852 13582 10908
rect 13518 10848 13582 10852
rect 9996 10780 10060 10844
rect 12020 10780 12084 10844
rect 6500 10644 6564 10708
rect 3188 10372 3252 10436
rect 7236 10372 7300 10436
rect 10180 10372 10244 10436
rect 5882 10364 5946 10368
rect 5882 10308 5886 10364
rect 5886 10308 5942 10364
rect 5942 10308 5946 10364
rect 5882 10304 5946 10308
rect 5962 10364 6026 10368
rect 5962 10308 5966 10364
rect 5966 10308 6022 10364
rect 6022 10308 6026 10364
rect 5962 10304 6026 10308
rect 6042 10364 6106 10368
rect 6042 10308 6046 10364
rect 6046 10308 6102 10364
rect 6102 10308 6106 10364
rect 6042 10304 6106 10308
rect 6122 10364 6186 10368
rect 6122 10308 6126 10364
rect 6126 10308 6182 10364
rect 6182 10308 6186 10364
rect 6122 10304 6186 10308
rect 10813 10364 10877 10368
rect 10813 10308 10817 10364
rect 10817 10308 10873 10364
rect 10873 10308 10877 10364
rect 10813 10304 10877 10308
rect 10893 10364 10957 10368
rect 10893 10308 10897 10364
rect 10897 10308 10953 10364
rect 10953 10308 10957 10364
rect 10893 10304 10957 10308
rect 10973 10364 11037 10368
rect 10973 10308 10977 10364
rect 10977 10308 11033 10364
rect 11033 10308 11037 10364
rect 10973 10304 11037 10308
rect 11053 10364 11117 10368
rect 11053 10308 11057 10364
rect 11057 10308 11113 10364
rect 11113 10308 11117 10364
rect 11053 10304 11117 10308
rect 8892 10236 8956 10300
rect 6316 9964 6380 10028
rect 3417 9820 3481 9824
rect 3417 9764 3421 9820
rect 3421 9764 3477 9820
rect 3477 9764 3481 9820
rect 3417 9760 3481 9764
rect 3497 9820 3561 9824
rect 3497 9764 3501 9820
rect 3501 9764 3557 9820
rect 3557 9764 3561 9820
rect 3497 9760 3561 9764
rect 3577 9820 3641 9824
rect 3577 9764 3581 9820
rect 3581 9764 3637 9820
rect 3637 9764 3641 9820
rect 3577 9760 3641 9764
rect 3657 9820 3721 9824
rect 3657 9764 3661 9820
rect 3661 9764 3717 9820
rect 3717 9764 3721 9820
rect 3657 9760 3721 9764
rect 8348 9820 8412 9824
rect 8348 9764 8352 9820
rect 8352 9764 8408 9820
rect 8408 9764 8412 9820
rect 8348 9760 8412 9764
rect 8428 9820 8492 9824
rect 8428 9764 8432 9820
rect 8432 9764 8488 9820
rect 8488 9764 8492 9820
rect 8428 9760 8492 9764
rect 8508 9820 8572 9824
rect 8508 9764 8512 9820
rect 8512 9764 8568 9820
rect 8568 9764 8572 9820
rect 8508 9760 8572 9764
rect 8588 9820 8652 9824
rect 8588 9764 8592 9820
rect 8592 9764 8648 9820
rect 8648 9764 8652 9820
rect 8588 9760 8652 9764
rect 11652 9828 11716 9892
rect 11836 9828 11900 9892
rect 13278 9820 13342 9824
rect 13278 9764 13282 9820
rect 13282 9764 13338 9820
rect 13338 9764 13342 9820
rect 13278 9760 13342 9764
rect 13358 9820 13422 9824
rect 13358 9764 13362 9820
rect 13362 9764 13418 9820
rect 13418 9764 13422 9820
rect 13358 9760 13422 9764
rect 13438 9820 13502 9824
rect 13438 9764 13442 9820
rect 13442 9764 13498 9820
rect 13498 9764 13502 9820
rect 13438 9760 13502 9764
rect 13518 9820 13582 9824
rect 13518 9764 13522 9820
rect 13522 9764 13578 9820
rect 13578 9764 13582 9820
rect 13518 9760 13582 9764
rect 10364 9556 10428 9620
rect 14964 9616 15028 9620
rect 14964 9560 15014 9616
rect 15014 9560 15028 9616
rect 14964 9556 15028 9560
rect 9444 9284 9508 9348
rect 5882 9276 5946 9280
rect 5882 9220 5886 9276
rect 5886 9220 5942 9276
rect 5942 9220 5946 9276
rect 5882 9216 5946 9220
rect 5962 9276 6026 9280
rect 5962 9220 5966 9276
rect 5966 9220 6022 9276
rect 6022 9220 6026 9276
rect 5962 9216 6026 9220
rect 6042 9276 6106 9280
rect 6042 9220 6046 9276
rect 6046 9220 6102 9276
rect 6102 9220 6106 9276
rect 6042 9216 6106 9220
rect 6122 9276 6186 9280
rect 6122 9220 6126 9276
rect 6126 9220 6182 9276
rect 6182 9220 6186 9276
rect 6122 9216 6186 9220
rect 10813 9276 10877 9280
rect 10813 9220 10817 9276
rect 10817 9220 10873 9276
rect 10873 9220 10877 9276
rect 10813 9216 10877 9220
rect 10893 9276 10957 9280
rect 10893 9220 10897 9276
rect 10897 9220 10953 9276
rect 10953 9220 10957 9276
rect 10893 9216 10957 9220
rect 10973 9276 11037 9280
rect 10973 9220 10977 9276
rect 10977 9220 11033 9276
rect 11033 9220 11037 9276
rect 10973 9216 11037 9220
rect 11053 9276 11117 9280
rect 11053 9220 11057 9276
rect 11057 9220 11113 9276
rect 11113 9220 11117 9276
rect 11053 9216 11117 9220
rect 11652 9284 11716 9348
rect 12020 9012 12084 9076
rect 9812 8876 9876 8940
rect 11652 8740 11716 8804
rect 3417 8732 3481 8736
rect 3417 8676 3421 8732
rect 3421 8676 3477 8732
rect 3477 8676 3481 8732
rect 3417 8672 3481 8676
rect 3497 8732 3561 8736
rect 3497 8676 3501 8732
rect 3501 8676 3557 8732
rect 3557 8676 3561 8732
rect 3497 8672 3561 8676
rect 3577 8732 3641 8736
rect 3577 8676 3581 8732
rect 3581 8676 3637 8732
rect 3637 8676 3641 8732
rect 3577 8672 3641 8676
rect 3657 8732 3721 8736
rect 3657 8676 3661 8732
rect 3661 8676 3717 8732
rect 3717 8676 3721 8732
rect 3657 8672 3721 8676
rect 8348 8732 8412 8736
rect 8348 8676 8352 8732
rect 8352 8676 8408 8732
rect 8408 8676 8412 8732
rect 8348 8672 8412 8676
rect 8428 8732 8492 8736
rect 8428 8676 8432 8732
rect 8432 8676 8488 8732
rect 8488 8676 8492 8732
rect 8428 8672 8492 8676
rect 8508 8732 8572 8736
rect 8508 8676 8512 8732
rect 8512 8676 8568 8732
rect 8568 8676 8572 8732
rect 8508 8672 8572 8676
rect 8588 8732 8652 8736
rect 8588 8676 8592 8732
rect 8592 8676 8648 8732
rect 8648 8676 8652 8732
rect 8588 8672 8652 8676
rect 13278 8732 13342 8736
rect 13278 8676 13282 8732
rect 13282 8676 13338 8732
rect 13338 8676 13342 8732
rect 13278 8672 13342 8676
rect 13358 8732 13422 8736
rect 13358 8676 13362 8732
rect 13362 8676 13418 8732
rect 13418 8676 13422 8732
rect 13358 8672 13422 8676
rect 13438 8732 13502 8736
rect 13438 8676 13442 8732
rect 13442 8676 13498 8732
rect 13498 8676 13502 8732
rect 13438 8672 13502 8676
rect 13518 8732 13582 8736
rect 13518 8676 13522 8732
rect 13522 8676 13578 8732
rect 13578 8676 13582 8732
rect 13518 8672 13582 8676
rect 8156 8604 8220 8668
rect 13860 8332 13924 8396
rect 14228 8332 14292 8396
rect 7420 8196 7484 8260
rect 14964 8196 15028 8260
rect 5882 8188 5946 8192
rect 5882 8132 5886 8188
rect 5886 8132 5942 8188
rect 5942 8132 5946 8188
rect 5882 8128 5946 8132
rect 5962 8188 6026 8192
rect 5962 8132 5966 8188
rect 5966 8132 6022 8188
rect 6022 8132 6026 8188
rect 5962 8128 6026 8132
rect 6042 8188 6106 8192
rect 6042 8132 6046 8188
rect 6046 8132 6102 8188
rect 6102 8132 6106 8188
rect 6042 8128 6106 8132
rect 6122 8188 6186 8192
rect 6122 8132 6126 8188
rect 6126 8132 6182 8188
rect 6182 8132 6186 8188
rect 6122 8128 6186 8132
rect 10813 8188 10877 8192
rect 10813 8132 10817 8188
rect 10817 8132 10873 8188
rect 10873 8132 10877 8188
rect 10813 8128 10877 8132
rect 10893 8188 10957 8192
rect 10893 8132 10897 8188
rect 10897 8132 10953 8188
rect 10953 8132 10957 8188
rect 10893 8128 10957 8132
rect 10973 8188 11037 8192
rect 10973 8132 10977 8188
rect 10977 8132 11033 8188
rect 11033 8132 11037 8188
rect 10973 8128 11037 8132
rect 11053 8188 11117 8192
rect 11053 8132 11057 8188
rect 11057 8132 11113 8188
rect 11113 8132 11117 8188
rect 11053 8128 11117 8132
rect 10548 8060 10612 8124
rect 11284 8120 11348 8124
rect 11284 8064 11298 8120
rect 11298 8064 11348 8120
rect 11284 8060 11348 8064
rect 7052 7924 7116 7988
rect 13676 7924 13740 7988
rect 9076 7788 9140 7852
rect 3417 7644 3481 7648
rect 3417 7588 3421 7644
rect 3421 7588 3477 7644
rect 3477 7588 3481 7644
rect 3417 7584 3481 7588
rect 3497 7644 3561 7648
rect 3497 7588 3501 7644
rect 3501 7588 3557 7644
rect 3557 7588 3561 7644
rect 3497 7584 3561 7588
rect 3577 7644 3641 7648
rect 3577 7588 3581 7644
rect 3581 7588 3637 7644
rect 3637 7588 3641 7644
rect 3577 7584 3641 7588
rect 3657 7644 3721 7648
rect 3657 7588 3661 7644
rect 3661 7588 3717 7644
rect 3717 7588 3721 7644
rect 3657 7584 3721 7588
rect 8348 7644 8412 7648
rect 8348 7588 8352 7644
rect 8352 7588 8408 7644
rect 8408 7588 8412 7644
rect 8348 7584 8412 7588
rect 8428 7644 8492 7648
rect 8428 7588 8432 7644
rect 8432 7588 8488 7644
rect 8488 7588 8492 7644
rect 8428 7584 8492 7588
rect 8508 7644 8572 7648
rect 8508 7588 8512 7644
rect 8512 7588 8568 7644
rect 8568 7588 8572 7644
rect 8508 7584 8572 7588
rect 8588 7644 8652 7648
rect 8588 7588 8592 7644
rect 8592 7588 8648 7644
rect 8648 7588 8652 7644
rect 8588 7584 8652 7588
rect 8892 7576 8956 7580
rect 8892 7520 8942 7576
rect 8942 7520 8956 7576
rect 8892 7516 8956 7520
rect 11468 7652 11532 7716
rect 13278 7644 13342 7648
rect 13278 7588 13282 7644
rect 13282 7588 13338 7644
rect 13338 7588 13342 7644
rect 13278 7584 13342 7588
rect 13358 7644 13422 7648
rect 13358 7588 13362 7644
rect 13362 7588 13418 7644
rect 13418 7588 13422 7644
rect 13358 7584 13422 7588
rect 13438 7644 13502 7648
rect 13438 7588 13442 7644
rect 13442 7588 13498 7644
rect 13498 7588 13502 7644
rect 13438 7584 13502 7588
rect 13518 7644 13582 7648
rect 13518 7588 13522 7644
rect 13522 7588 13578 7644
rect 13578 7588 13582 7644
rect 13518 7584 13582 7588
rect 7604 7380 7668 7444
rect 11284 7380 11348 7444
rect 12940 7380 13004 7444
rect 12388 7244 12452 7308
rect 12940 7244 13004 7308
rect 10548 7108 10612 7172
rect 11468 7108 11532 7172
rect 12388 7108 12452 7172
rect 14780 7108 14844 7172
rect 5882 7100 5946 7104
rect 5882 7044 5886 7100
rect 5886 7044 5942 7100
rect 5942 7044 5946 7100
rect 5882 7040 5946 7044
rect 5962 7100 6026 7104
rect 5962 7044 5966 7100
rect 5966 7044 6022 7100
rect 6022 7044 6026 7100
rect 5962 7040 6026 7044
rect 6042 7100 6106 7104
rect 6042 7044 6046 7100
rect 6046 7044 6102 7100
rect 6102 7044 6106 7100
rect 6042 7040 6106 7044
rect 6122 7100 6186 7104
rect 6122 7044 6126 7100
rect 6126 7044 6182 7100
rect 6182 7044 6186 7100
rect 6122 7040 6186 7044
rect 10813 7100 10877 7104
rect 10813 7044 10817 7100
rect 10817 7044 10873 7100
rect 10873 7044 10877 7100
rect 10813 7040 10877 7044
rect 10893 7100 10957 7104
rect 10893 7044 10897 7100
rect 10897 7044 10953 7100
rect 10953 7044 10957 7100
rect 10893 7040 10957 7044
rect 10973 7100 11037 7104
rect 10973 7044 10977 7100
rect 10977 7044 11033 7100
rect 11033 7044 11037 7100
rect 10973 7040 11037 7044
rect 11053 7100 11117 7104
rect 11053 7044 11057 7100
rect 11057 7044 11113 7100
rect 11113 7044 11117 7100
rect 11053 7040 11117 7044
rect 5212 6972 5276 7036
rect 11836 6972 11900 7036
rect 14044 6700 14108 6764
rect 10180 6564 10244 6628
rect 11468 6564 11532 6628
rect 11836 6564 11900 6628
rect 3417 6556 3481 6560
rect 3417 6500 3421 6556
rect 3421 6500 3477 6556
rect 3477 6500 3481 6556
rect 3417 6496 3481 6500
rect 3497 6556 3561 6560
rect 3497 6500 3501 6556
rect 3501 6500 3557 6556
rect 3557 6500 3561 6556
rect 3497 6496 3561 6500
rect 3577 6556 3641 6560
rect 3577 6500 3581 6556
rect 3581 6500 3637 6556
rect 3637 6500 3641 6556
rect 3577 6496 3641 6500
rect 3657 6556 3721 6560
rect 3657 6500 3661 6556
rect 3661 6500 3717 6556
rect 3717 6500 3721 6556
rect 3657 6496 3721 6500
rect 8348 6556 8412 6560
rect 8348 6500 8352 6556
rect 8352 6500 8408 6556
rect 8408 6500 8412 6556
rect 8348 6496 8412 6500
rect 8428 6556 8492 6560
rect 8428 6500 8432 6556
rect 8432 6500 8488 6556
rect 8488 6500 8492 6556
rect 8428 6496 8492 6500
rect 8508 6556 8572 6560
rect 8508 6500 8512 6556
rect 8512 6500 8568 6556
rect 8568 6500 8572 6556
rect 8508 6496 8572 6500
rect 8588 6556 8652 6560
rect 8588 6500 8592 6556
rect 8592 6500 8648 6556
rect 8648 6500 8652 6556
rect 8588 6496 8652 6500
rect 13278 6556 13342 6560
rect 13278 6500 13282 6556
rect 13282 6500 13338 6556
rect 13338 6500 13342 6556
rect 13278 6496 13342 6500
rect 13358 6556 13422 6560
rect 13358 6500 13362 6556
rect 13362 6500 13418 6556
rect 13418 6500 13422 6556
rect 13358 6496 13422 6500
rect 13438 6556 13502 6560
rect 13438 6500 13442 6556
rect 13442 6500 13498 6556
rect 13498 6500 13502 6556
rect 13438 6496 13502 6500
rect 13518 6556 13582 6560
rect 13518 6500 13522 6556
rect 13522 6500 13578 6556
rect 13578 6500 13582 6556
rect 13518 6496 13582 6500
rect 9996 6428 10060 6492
rect 13676 6156 13740 6220
rect 11468 6080 11532 6084
rect 11468 6024 11518 6080
rect 11518 6024 11532 6080
rect 5882 6012 5946 6016
rect 5882 5956 5886 6012
rect 5886 5956 5942 6012
rect 5942 5956 5946 6012
rect 5882 5952 5946 5956
rect 5962 6012 6026 6016
rect 5962 5956 5966 6012
rect 5966 5956 6022 6012
rect 6022 5956 6026 6012
rect 5962 5952 6026 5956
rect 6042 6012 6106 6016
rect 6042 5956 6046 6012
rect 6046 5956 6102 6012
rect 6102 5956 6106 6012
rect 6042 5952 6106 5956
rect 6122 6012 6186 6016
rect 6122 5956 6126 6012
rect 6126 5956 6182 6012
rect 6182 5956 6186 6012
rect 6122 5952 6186 5956
rect 4476 5884 4540 5948
rect 7420 5884 7484 5948
rect 9260 5884 9324 5948
rect 4108 5748 4172 5812
rect 11468 6020 11532 6024
rect 12572 6080 12636 6084
rect 12572 6024 12586 6080
rect 12586 6024 12636 6080
rect 12572 6020 12636 6024
rect 10813 6012 10877 6016
rect 10813 5956 10817 6012
rect 10817 5956 10873 6012
rect 10873 5956 10877 6012
rect 10813 5952 10877 5956
rect 10893 6012 10957 6016
rect 10893 5956 10897 6012
rect 10897 5956 10953 6012
rect 10953 5956 10957 6012
rect 10893 5952 10957 5956
rect 10973 6012 11037 6016
rect 10973 5956 10977 6012
rect 10977 5956 11033 6012
rect 11033 5956 11037 6012
rect 10973 5952 11037 5956
rect 11053 6012 11117 6016
rect 11053 5956 11057 6012
rect 11057 5956 11113 6012
rect 11113 5956 11117 6012
rect 11053 5952 11117 5956
rect 7052 5672 7116 5676
rect 7052 5616 7066 5672
rect 7066 5616 7116 5672
rect 7052 5612 7116 5616
rect 6500 5476 6564 5540
rect 12388 5748 12452 5812
rect 13676 5748 13740 5812
rect 12020 5612 12084 5676
rect 12572 5612 12636 5676
rect 12204 5476 12268 5540
rect 3417 5468 3481 5472
rect 3417 5412 3421 5468
rect 3421 5412 3477 5468
rect 3477 5412 3481 5468
rect 3417 5408 3481 5412
rect 3497 5468 3561 5472
rect 3497 5412 3501 5468
rect 3501 5412 3557 5468
rect 3557 5412 3561 5468
rect 3497 5408 3561 5412
rect 3577 5468 3641 5472
rect 3577 5412 3581 5468
rect 3581 5412 3637 5468
rect 3637 5412 3641 5468
rect 3577 5408 3641 5412
rect 3657 5468 3721 5472
rect 3657 5412 3661 5468
rect 3661 5412 3717 5468
rect 3717 5412 3721 5468
rect 3657 5408 3721 5412
rect 8348 5468 8412 5472
rect 8348 5412 8352 5468
rect 8352 5412 8408 5468
rect 8408 5412 8412 5468
rect 8348 5408 8412 5412
rect 8428 5468 8492 5472
rect 8428 5412 8432 5468
rect 8432 5412 8488 5468
rect 8488 5412 8492 5468
rect 8428 5408 8492 5412
rect 8508 5468 8572 5472
rect 8508 5412 8512 5468
rect 8512 5412 8568 5468
rect 8568 5412 8572 5468
rect 8508 5408 8572 5412
rect 8588 5468 8652 5472
rect 8588 5412 8592 5468
rect 8592 5412 8648 5468
rect 8648 5412 8652 5468
rect 8588 5408 8652 5412
rect 13278 5468 13342 5472
rect 13278 5412 13282 5468
rect 13282 5412 13338 5468
rect 13338 5412 13342 5468
rect 13278 5408 13342 5412
rect 13358 5468 13422 5472
rect 13358 5412 13362 5468
rect 13362 5412 13418 5468
rect 13418 5412 13422 5468
rect 13358 5408 13422 5412
rect 13438 5468 13502 5472
rect 13438 5412 13442 5468
rect 13442 5412 13498 5468
rect 13498 5412 13502 5468
rect 13438 5408 13502 5412
rect 13518 5468 13582 5472
rect 13518 5412 13522 5468
rect 13522 5412 13578 5468
rect 13578 5412 13582 5468
rect 13518 5408 13582 5412
rect 8892 5340 8956 5404
rect 13860 5204 13924 5268
rect 6684 4932 6748 4996
rect 11836 4932 11900 4996
rect 5882 4924 5946 4928
rect 5882 4868 5886 4924
rect 5886 4868 5942 4924
rect 5942 4868 5946 4924
rect 5882 4864 5946 4868
rect 5962 4924 6026 4928
rect 5962 4868 5966 4924
rect 5966 4868 6022 4924
rect 6022 4868 6026 4924
rect 5962 4864 6026 4868
rect 6042 4924 6106 4928
rect 6042 4868 6046 4924
rect 6046 4868 6102 4924
rect 6102 4868 6106 4924
rect 6042 4864 6106 4868
rect 6122 4924 6186 4928
rect 6122 4868 6126 4924
rect 6126 4868 6182 4924
rect 6182 4868 6186 4924
rect 6122 4864 6186 4868
rect 10813 4924 10877 4928
rect 10813 4868 10817 4924
rect 10817 4868 10873 4924
rect 10873 4868 10877 4924
rect 10813 4864 10877 4868
rect 10893 4924 10957 4928
rect 10893 4868 10897 4924
rect 10897 4868 10953 4924
rect 10953 4868 10957 4924
rect 10893 4864 10957 4868
rect 10973 4924 11037 4928
rect 10973 4868 10977 4924
rect 10977 4868 11033 4924
rect 11033 4868 11037 4924
rect 10973 4864 11037 4868
rect 11053 4924 11117 4928
rect 11053 4868 11057 4924
rect 11057 4868 11113 4924
rect 11113 4868 11117 4924
rect 11053 4864 11117 4868
rect 5212 4796 5276 4860
rect 10364 4796 10428 4860
rect 11836 4796 11900 4860
rect 14780 4796 14844 4860
rect 3417 4380 3481 4384
rect 3417 4324 3421 4380
rect 3421 4324 3477 4380
rect 3477 4324 3481 4380
rect 3417 4320 3481 4324
rect 3497 4380 3561 4384
rect 3497 4324 3501 4380
rect 3501 4324 3557 4380
rect 3557 4324 3561 4380
rect 3497 4320 3561 4324
rect 3577 4380 3641 4384
rect 3577 4324 3581 4380
rect 3581 4324 3637 4380
rect 3637 4324 3641 4380
rect 3577 4320 3641 4324
rect 3657 4380 3721 4384
rect 3657 4324 3661 4380
rect 3661 4324 3717 4380
rect 3717 4324 3721 4380
rect 3657 4320 3721 4324
rect 9076 4388 9140 4452
rect 9628 4388 9692 4452
rect 9996 4388 10060 4452
rect 8348 4380 8412 4384
rect 8348 4324 8352 4380
rect 8352 4324 8408 4380
rect 8408 4324 8412 4380
rect 8348 4320 8412 4324
rect 8428 4380 8492 4384
rect 8428 4324 8432 4380
rect 8432 4324 8488 4380
rect 8488 4324 8492 4380
rect 8428 4320 8492 4324
rect 8508 4380 8572 4384
rect 8508 4324 8512 4380
rect 8512 4324 8568 4380
rect 8568 4324 8572 4380
rect 8508 4320 8572 4324
rect 8588 4380 8652 4384
rect 8588 4324 8592 4380
rect 8592 4324 8648 4380
rect 8648 4324 8652 4380
rect 8588 4320 8652 4324
rect 4476 4252 4540 4316
rect 9076 4312 9140 4316
rect 10548 4388 10612 4452
rect 13278 4380 13342 4384
rect 13278 4324 13282 4380
rect 13282 4324 13338 4380
rect 13338 4324 13342 4380
rect 13278 4320 13342 4324
rect 13358 4380 13422 4384
rect 13358 4324 13362 4380
rect 13362 4324 13418 4380
rect 13418 4324 13422 4380
rect 13358 4320 13422 4324
rect 13438 4380 13502 4384
rect 13438 4324 13442 4380
rect 13442 4324 13498 4380
rect 13498 4324 13502 4380
rect 13438 4320 13502 4324
rect 13518 4380 13582 4384
rect 13518 4324 13522 4380
rect 13522 4324 13578 4380
rect 13578 4324 13582 4380
rect 13518 4320 13582 4324
rect 9076 4256 9126 4312
rect 9126 4256 9140 4312
rect 9076 4252 9140 4256
rect 8892 4116 8956 4180
rect 9444 4176 9508 4180
rect 9444 4120 9494 4176
rect 9494 4120 9508 4176
rect 9444 4116 9508 4120
rect 9812 4176 9876 4180
rect 9812 4120 9826 4176
rect 9826 4120 9876 4176
rect 9812 4116 9876 4120
rect 12020 4252 12084 4316
rect 10364 3980 10428 4044
rect 5396 3904 5460 3908
rect 5396 3848 5446 3904
rect 5446 3848 5460 3904
rect 5396 3844 5460 3848
rect 6500 3844 6564 3908
rect 10548 3844 10612 3908
rect 14412 3980 14476 4044
rect 5882 3836 5946 3840
rect 5882 3780 5886 3836
rect 5886 3780 5942 3836
rect 5942 3780 5946 3836
rect 5882 3776 5946 3780
rect 5962 3836 6026 3840
rect 5962 3780 5966 3836
rect 5966 3780 6022 3836
rect 6022 3780 6026 3836
rect 5962 3776 6026 3780
rect 6042 3836 6106 3840
rect 6042 3780 6046 3836
rect 6046 3780 6102 3836
rect 6102 3780 6106 3836
rect 6042 3776 6106 3780
rect 6122 3836 6186 3840
rect 6122 3780 6126 3836
rect 6126 3780 6182 3836
rect 6182 3780 6186 3836
rect 6122 3776 6186 3780
rect 10813 3836 10877 3840
rect 10813 3780 10817 3836
rect 10817 3780 10873 3836
rect 10873 3780 10877 3836
rect 10813 3776 10877 3780
rect 10893 3836 10957 3840
rect 10893 3780 10897 3836
rect 10897 3780 10953 3836
rect 10953 3780 10957 3836
rect 10893 3776 10957 3780
rect 10973 3836 11037 3840
rect 10973 3780 10977 3836
rect 10977 3780 11033 3836
rect 11033 3780 11037 3836
rect 10973 3776 11037 3780
rect 11053 3836 11117 3840
rect 11053 3780 11057 3836
rect 11057 3780 11113 3836
rect 11113 3780 11117 3836
rect 11053 3776 11117 3780
rect 3188 3708 3252 3772
rect 8156 3708 8220 3772
rect 12020 3768 12084 3772
rect 12020 3712 12034 3768
rect 12034 3712 12084 3768
rect 12020 3708 12084 3712
rect 12388 3708 12452 3772
rect 12204 3360 12268 3364
rect 12204 3304 12254 3360
rect 12254 3304 12268 3360
rect 12204 3300 12268 3304
rect 12572 3300 12636 3364
rect 3417 3292 3481 3296
rect 3417 3236 3421 3292
rect 3421 3236 3477 3292
rect 3477 3236 3481 3292
rect 3417 3232 3481 3236
rect 3497 3292 3561 3296
rect 3497 3236 3501 3292
rect 3501 3236 3557 3292
rect 3557 3236 3561 3292
rect 3497 3232 3561 3236
rect 3577 3292 3641 3296
rect 3577 3236 3581 3292
rect 3581 3236 3637 3292
rect 3637 3236 3641 3292
rect 3577 3232 3641 3236
rect 3657 3292 3721 3296
rect 3657 3236 3661 3292
rect 3661 3236 3717 3292
rect 3717 3236 3721 3292
rect 3657 3232 3721 3236
rect 8348 3292 8412 3296
rect 8348 3236 8352 3292
rect 8352 3236 8408 3292
rect 8408 3236 8412 3292
rect 8348 3232 8412 3236
rect 8428 3292 8492 3296
rect 8428 3236 8432 3292
rect 8432 3236 8488 3292
rect 8488 3236 8492 3292
rect 8428 3232 8492 3236
rect 8508 3292 8572 3296
rect 8508 3236 8512 3292
rect 8512 3236 8568 3292
rect 8568 3236 8572 3292
rect 8508 3232 8572 3236
rect 8588 3292 8652 3296
rect 8588 3236 8592 3292
rect 8592 3236 8648 3292
rect 8648 3236 8652 3292
rect 8588 3232 8652 3236
rect 13278 3292 13342 3296
rect 13278 3236 13282 3292
rect 13282 3236 13338 3292
rect 13338 3236 13342 3292
rect 13278 3232 13342 3236
rect 13358 3292 13422 3296
rect 13358 3236 13362 3292
rect 13362 3236 13418 3292
rect 13418 3236 13422 3292
rect 13358 3232 13422 3236
rect 13438 3292 13502 3296
rect 13438 3236 13442 3292
rect 13442 3236 13498 3292
rect 13498 3236 13502 3292
rect 13438 3232 13502 3236
rect 13518 3292 13582 3296
rect 13518 3236 13522 3292
rect 13522 3236 13578 3292
rect 13578 3236 13582 3292
rect 13518 3232 13582 3236
rect 7604 3224 7668 3228
rect 7604 3168 7618 3224
rect 7618 3168 7668 3224
rect 7604 3164 7668 3168
rect 13124 3164 13188 3228
rect 11284 2892 11348 2956
rect 11652 3088 11716 3092
rect 11652 3032 11666 3088
rect 11666 3032 11716 3088
rect 11652 3028 11716 3032
rect 13676 3028 13740 3092
rect 14964 2892 15028 2956
rect 9444 2756 9508 2820
rect 5882 2748 5946 2752
rect 5882 2692 5886 2748
rect 5886 2692 5942 2748
rect 5942 2692 5946 2748
rect 5882 2688 5946 2692
rect 5962 2748 6026 2752
rect 5962 2692 5966 2748
rect 5966 2692 6022 2748
rect 6022 2692 6026 2748
rect 5962 2688 6026 2692
rect 6042 2748 6106 2752
rect 6042 2692 6046 2748
rect 6046 2692 6102 2748
rect 6102 2692 6106 2748
rect 6042 2688 6106 2692
rect 6122 2748 6186 2752
rect 6122 2692 6126 2748
rect 6126 2692 6182 2748
rect 6182 2692 6186 2748
rect 6122 2688 6186 2692
rect 10813 2748 10877 2752
rect 10813 2692 10817 2748
rect 10817 2692 10873 2748
rect 10873 2692 10877 2748
rect 10813 2688 10877 2692
rect 10893 2748 10957 2752
rect 10893 2692 10897 2748
rect 10897 2692 10953 2748
rect 10953 2692 10957 2748
rect 10893 2688 10957 2692
rect 10973 2748 11037 2752
rect 10973 2692 10977 2748
rect 10977 2692 11033 2748
rect 11033 2692 11037 2748
rect 10973 2688 11037 2692
rect 11053 2748 11117 2752
rect 11053 2692 11057 2748
rect 11057 2692 11113 2748
rect 11113 2692 11117 2748
rect 11053 2688 11117 2692
rect 5212 2680 5276 2684
rect 5212 2624 5226 2680
rect 5226 2624 5276 2680
rect 5212 2620 5276 2624
rect 5396 2680 5460 2684
rect 5396 2624 5446 2680
rect 5446 2624 5460 2680
rect 5396 2620 5460 2624
rect 7788 2620 7852 2684
rect 8892 2620 8956 2684
rect 12204 2620 12268 2684
rect 9260 2484 9324 2548
rect 12020 2484 12084 2548
rect 12940 2484 13004 2548
rect 6684 2348 6748 2412
rect 12756 2348 12820 2412
rect 3417 2204 3481 2208
rect 3417 2148 3421 2204
rect 3421 2148 3477 2204
rect 3477 2148 3481 2204
rect 3417 2144 3481 2148
rect 3497 2204 3561 2208
rect 3497 2148 3501 2204
rect 3501 2148 3557 2204
rect 3557 2148 3561 2204
rect 3497 2144 3561 2148
rect 3577 2204 3641 2208
rect 3577 2148 3581 2204
rect 3581 2148 3637 2204
rect 3637 2148 3641 2204
rect 3577 2144 3641 2148
rect 3657 2204 3721 2208
rect 3657 2148 3661 2204
rect 3661 2148 3717 2204
rect 3717 2148 3721 2204
rect 3657 2144 3721 2148
rect 8348 2204 8412 2208
rect 8348 2148 8352 2204
rect 8352 2148 8408 2204
rect 8408 2148 8412 2204
rect 8348 2144 8412 2148
rect 8428 2204 8492 2208
rect 8428 2148 8432 2204
rect 8432 2148 8488 2204
rect 8488 2148 8492 2204
rect 8428 2144 8492 2148
rect 8508 2204 8572 2208
rect 8508 2148 8512 2204
rect 8512 2148 8568 2204
rect 8568 2148 8572 2204
rect 8508 2144 8572 2148
rect 8588 2204 8652 2208
rect 8588 2148 8592 2204
rect 8592 2148 8648 2204
rect 8648 2148 8652 2204
rect 8588 2144 8652 2148
rect 13278 2204 13342 2208
rect 13278 2148 13282 2204
rect 13282 2148 13338 2204
rect 13338 2148 13342 2204
rect 13278 2144 13342 2148
rect 13358 2204 13422 2208
rect 13358 2148 13362 2204
rect 13362 2148 13418 2204
rect 13418 2148 13422 2204
rect 13358 2144 13422 2148
rect 13438 2204 13502 2208
rect 13438 2148 13442 2204
rect 13442 2148 13498 2204
rect 13498 2148 13502 2204
rect 13438 2144 13502 2148
rect 13518 2204 13582 2208
rect 13518 2148 13522 2204
rect 13522 2148 13578 2204
rect 13578 2148 13582 2204
rect 13518 2144 13582 2148
rect 11468 2076 11532 2140
rect 14228 1804 14292 1868
rect 11836 1532 11900 1596
rect 9076 1396 9140 1460
<< metal4 >>
rect 10179 16012 10245 16013
rect 10179 15948 10180 16012
rect 10244 15948 10245 16012
rect 10179 15947 10245 15948
rect 3409 15264 3729 15824
rect 3409 15200 3417 15264
rect 3481 15200 3497 15264
rect 3561 15200 3577 15264
rect 3641 15200 3657 15264
rect 3721 15200 3729 15264
rect 3187 14652 3253 14653
rect 3187 14588 3188 14652
rect 3252 14588 3253 14652
rect 3187 14587 3253 14588
rect 3190 10437 3250 14587
rect 3409 14176 3729 15200
rect 5874 15808 6195 15824
rect 5874 15744 5882 15808
rect 5946 15744 5962 15808
rect 6026 15744 6042 15808
rect 6106 15744 6122 15808
rect 6186 15744 6195 15808
rect 5874 14720 6195 15744
rect 7419 15332 7485 15333
rect 7419 15268 7420 15332
rect 7484 15268 7485 15332
rect 7419 15267 7485 15268
rect 6315 15060 6381 15061
rect 6315 14996 6316 15060
rect 6380 14996 6381 15060
rect 6315 14995 6381 14996
rect 5874 14656 5882 14720
rect 5946 14656 5962 14720
rect 6026 14656 6042 14720
rect 6106 14656 6122 14720
rect 6186 14656 6195 14720
rect 5579 14380 5645 14381
rect 5579 14316 5580 14380
rect 5644 14316 5645 14380
rect 5579 14315 5645 14316
rect 3409 14112 3417 14176
rect 3481 14112 3497 14176
rect 3561 14112 3577 14176
rect 3641 14112 3657 14176
rect 3721 14112 3729 14176
rect 3409 13088 3729 14112
rect 4475 14108 4541 14109
rect 4475 14044 4476 14108
rect 4540 14044 4541 14108
rect 4475 14043 4541 14044
rect 3409 13024 3417 13088
rect 3481 13024 3497 13088
rect 3561 13024 3577 13088
rect 3641 13024 3657 13088
rect 3721 13024 3729 13088
rect 3409 12000 3729 13024
rect 4478 12613 4538 14043
rect 4475 12612 4541 12613
rect 4475 12548 4476 12612
rect 4540 12548 4541 12612
rect 4475 12547 4541 12548
rect 5582 12069 5642 14315
rect 5874 13632 6195 14656
rect 5874 13568 5882 13632
rect 5946 13568 5962 13632
rect 6026 13568 6042 13632
rect 6106 13568 6122 13632
rect 6186 13568 6195 13632
rect 5874 12544 6195 13568
rect 5874 12480 5882 12544
rect 5946 12480 5962 12544
rect 6026 12480 6042 12544
rect 6106 12480 6122 12544
rect 6186 12480 6195 12544
rect 5579 12068 5645 12069
rect 5579 12004 5580 12068
rect 5644 12004 5645 12068
rect 5579 12003 5645 12004
rect 3409 11936 3417 12000
rect 3481 11936 3497 12000
rect 3561 11936 3577 12000
rect 3641 11936 3657 12000
rect 3721 11936 3729 12000
rect 3409 10912 3729 11936
rect 3409 10848 3417 10912
rect 3481 10848 3497 10912
rect 3561 10848 3577 10912
rect 3641 10848 3657 10912
rect 3721 10848 3729 10912
rect 3187 10436 3253 10437
rect 3187 10372 3188 10436
rect 3252 10372 3253 10436
rect 3187 10371 3253 10372
rect 3190 3773 3250 10371
rect 3409 9824 3729 10848
rect 3409 9760 3417 9824
rect 3481 9760 3497 9824
rect 3561 9760 3577 9824
rect 3641 9760 3657 9824
rect 3721 9760 3729 9824
rect 3409 8736 3729 9760
rect 3409 8672 3417 8736
rect 3481 8672 3497 8736
rect 3561 8672 3577 8736
rect 3641 8672 3657 8736
rect 3721 8672 3729 8736
rect 3409 7648 3729 8672
rect 3409 7584 3417 7648
rect 3481 7584 3497 7648
rect 3561 7584 3577 7648
rect 3641 7584 3657 7648
rect 3721 7584 3729 7648
rect 3409 6560 3729 7584
rect 5874 11456 6195 12480
rect 5874 11392 5882 11456
rect 5946 11392 5962 11456
rect 6026 11392 6042 11456
rect 6106 11392 6122 11456
rect 6186 11392 6195 11456
rect 5874 10368 6195 11392
rect 5874 10304 5882 10368
rect 5946 10304 5962 10368
rect 6026 10304 6042 10368
rect 6106 10304 6122 10368
rect 6186 10304 6195 10368
rect 5874 9280 6195 10304
rect 6318 10029 6378 14995
rect 6683 14652 6749 14653
rect 6683 14588 6684 14652
rect 6748 14588 6749 14652
rect 6683 14587 6749 14588
rect 6499 13700 6565 13701
rect 6499 13636 6500 13700
rect 6564 13636 6565 13700
rect 6499 13635 6565 13636
rect 6502 10709 6562 13635
rect 6686 12477 6746 14587
rect 7235 12884 7301 12885
rect 7235 12820 7236 12884
rect 7300 12820 7301 12884
rect 7235 12819 7301 12820
rect 6683 12476 6749 12477
rect 6683 12412 6684 12476
rect 6748 12412 6749 12476
rect 6683 12411 6749 12412
rect 6499 10708 6565 10709
rect 6499 10644 6500 10708
rect 6564 10644 6565 10708
rect 6499 10643 6565 10644
rect 7238 10437 7298 12819
rect 7422 10981 7482 15267
rect 8340 15264 8660 15824
rect 8340 15200 8348 15264
rect 8412 15200 8428 15264
rect 8492 15200 8508 15264
rect 8572 15200 8588 15264
rect 8652 15200 8660 15264
rect 8340 14176 8660 15200
rect 9075 14788 9141 14789
rect 9075 14724 9076 14788
rect 9140 14724 9141 14788
rect 9075 14723 9141 14724
rect 8340 14112 8348 14176
rect 8412 14112 8428 14176
rect 8492 14112 8508 14176
rect 8572 14112 8588 14176
rect 8652 14112 8660 14176
rect 8340 13088 8660 14112
rect 8340 13024 8348 13088
rect 8412 13024 8428 13088
rect 8492 13024 8508 13088
rect 8572 13024 8588 13088
rect 8652 13024 8660 13088
rect 8340 12000 8660 13024
rect 8891 12612 8957 12613
rect 8891 12548 8892 12612
rect 8956 12548 8957 12612
rect 8891 12547 8957 12548
rect 8340 11936 8348 12000
rect 8412 11936 8428 12000
rect 8492 11936 8508 12000
rect 8572 11936 8588 12000
rect 8652 11936 8660 12000
rect 7787 11388 7853 11389
rect 7787 11324 7788 11388
rect 7852 11324 7853 11388
rect 7787 11323 7853 11324
rect 7419 10980 7485 10981
rect 7419 10916 7420 10980
rect 7484 10916 7485 10980
rect 7419 10915 7485 10916
rect 7235 10436 7301 10437
rect 7235 10372 7236 10436
rect 7300 10372 7301 10436
rect 7235 10371 7301 10372
rect 6315 10028 6381 10029
rect 6315 9964 6316 10028
rect 6380 9964 6381 10028
rect 6315 9963 6381 9964
rect 5874 9216 5882 9280
rect 5946 9216 5962 9280
rect 6026 9216 6042 9280
rect 6106 9216 6122 9280
rect 6186 9216 6195 9280
rect 5874 8192 6195 9216
rect 7422 8261 7482 10915
rect 7419 8260 7485 8261
rect 7419 8196 7420 8260
rect 7484 8196 7485 8260
rect 7419 8195 7485 8196
rect 5874 8128 5882 8192
rect 5946 8128 5962 8192
rect 6026 8128 6042 8192
rect 6106 8128 6122 8192
rect 6186 8128 6195 8192
rect 5874 7104 6195 8128
rect 7051 7988 7117 7989
rect 7051 7924 7052 7988
rect 7116 7924 7117 7988
rect 7051 7923 7117 7924
rect 5874 7040 5882 7104
rect 5946 7040 5962 7104
rect 6026 7040 6042 7104
rect 6106 7040 6122 7104
rect 6186 7040 6195 7104
rect 5211 7036 5277 7037
rect 5211 6972 5212 7036
rect 5276 6972 5277 7036
rect 5211 6971 5277 6972
rect 3409 6496 3417 6560
rect 3481 6496 3497 6560
rect 3561 6496 3577 6560
rect 3641 6496 3657 6560
rect 3721 6496 3729 6560
rect 3409 5472 3729 6496
rect 4475 5948 4541 5949
rect 4475 5884 4476 5948
rect 4540 5884 4541 5948
rect 4475 5883 4541 5884
rect 3409 5408 3417 5472
rect 3481 5408 3497 5472
rect 3561 5408 3577 5472
rect 3641 5408 3657 5472
rect 3721 5408 3729 5472
rect 3409 4384 3729 5408
rect 3409 4320 3417 4384
rect 3481 4320 3497 4384
rect 3561 4320 3577 4384
rect 3641 4320 3657 4384
rect 3721 4320 3729 4384
rect 3187 3772 3253 3773
rect 3187 3708 3188 3772
rect 3252 3708 3253 3772
rect 3187 3707 3253 3708
rect 3409 3296 3729 4320
rect 4478 4317 4538 5883
rect 5214 4861 5274 6971
rect 5874 6016 6195 7040
rect 5874 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6122 6016
rect 6186 5952 6195 6016
rect 5874 4928 6195 5952
rect 7054 5677 7114 7923
rect 7422 5949 7482 8195
rect 7603 7444 7669 7445
rect 7603 7380 7604 7444
rect 7668 7380 7669 7444
rect 7603 7379 7669 7380
rect 7419 5948 7485 5949
rect 7419 5884 7420 5948
rect 7484 5884 7485 5948
rect 7419 5883 7485 5884
rect 7051 5676 7117 5677
rect 7051 5612 7052 5676
rect 7116 5612 7117 5676
rect 7051 5611 7117 5612
rect 6499 5540 6565 5541
rect 6499 5476 6500 5540
rect 6564 5476 6565 5540
rect 6499 5475 6565 5476
rect 5874 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6122 4928
rect 6186 4864 6195 4928
rect 5211 4860 5277 4861
rect 5211 4796 5212 4860
rect 5276 4796 5277 4860
rect 5211 4795 5277 4796
rect 4475 4316 4541 4317
rect 4475 4252 4476 4316
rect 4540 4252 4541 4316
rect 4475 4251 4541 4252
rect 3409 3232 3417 3296
rect 3481 3232 3497 3296
rect 3561 3232 3577 3296
rect 3641 3232 3657 3296
rect 3721 3232 3729 3296
rect 3409 2208 3729 3232
rect 5214 2685 5274 4795
rect 5395 3908 5461 3909
rect 5395 3844 5396 3908
rect 5460 3844 5461 3908
rect 5395 3843 5461 3844
rect 5398 2685 5458 3843
rect 5874 3840 6195 4864
rect 6502 3909 6562 5475
rect 6683 4996 6749 4997
rect 6683 4932 6684 4996
rect 6748 4932 6749 4996
rect 6683 4931 6749 4932
rect 6499 3908 6565 3909
rect 6499 3844 6500 3908
rect 6564 3844 6565 3908
rect 6499 3843 6565 3844
rect 5874 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6122 3840
rect 6186 3776 6195 3840
rect 5874 2752 6195 3776
rect 5874 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6122 2752
rect 6186 2688 6195 2752
rect 5211 2684 5277 2685
rect 5211 2620 5212 2684
rect 5276 2620 5277 2684
rect 5211 2619 5277 2620
rect 5395 2684 5461 2685
rect 5395 2620 5396 2684
rect 5460 2620 5461 2684
rect 5395 2619 5461 2620
rect 3409 2144 3417 2208
rect 3481 2144 3497 2208
rect 3561 2144 3577 2208
rect 3641 2144 3657 2208
rect 3721 2144 3729 2208
rect 3409 2128 3729 2144
rect 5874 2128 6195 2688
rect 6686 2413 6746 4931
rect 7606 3229 7666 7379
rect 7603 3228 7669 3229
rect 7603 3164 7604 3228
rect 7668 3164 7669 3228
rect 7603 3163 7669 3164
rect 7790 2685 7850 11323
rect 8340 10912 8660 11936
rect 8340 10848 8348 10912
rect 8412 10848 8428 10912
rect 8492 10848 8508 10912
rect 8572 10848 8588 10912
rect 8652 10848 8660 10912
rect 8340 9824 8660 10848
rect 8894 10301 8954 12547
rect 9078 11933 9138 14723
rect 9811 14516 9877 14517
rect 9811 14452 9812 14516
rect 9876 14452 9877 14516
rect 9811 14451 9877 14452
rect 9627 14244 9693 14245
rect 9627 14180 9628 14244
rect 9692 14180 9693 14244
rect 9627 14179 9693 14180
rect 9259 14108 9325 14109
rect 9259 14044 9260 14108
rect 9324 14044 9325 14108
rect 9259 14043 9325 14044
rect 9262 12205 9322 14043
rect 9443 13020 9509 13021
rect 9443 12956 9444 13020
rect 9508 12956 9509 13020
rect 9443 12955 9509 12956
rect 9446 12477 9506 12955
rect 9443 12476 9509 12477
rect 9443 12412 9444 12476
rect 9508 12412 9509 12476
rect 9443 12411 9509 12412
rect 9259 12204 9325 12205
rect 9259 12140 9260 12204
rect 9324 12140 9325 12204
rect 9259 12139 9325 12140
rect 9630 11933 9690 14179
rect 9814 12205 9874 14451
rect 9811 12204 9877 12205
rect 9811 12140 9812 12204
rect 9876 12140 9877 12204
rect 9811 12139 9877 12140
rect 9075 11932 9141 11933
rect 9075 11868 9076 11932
rect 9140 11868 9141 11932
rect 9075 11867 9141 11868
rect 9627 11932 9693 11933
rect 9627 11868 9628 11932
rect 9692 11868 9693 11932
rect 9627 11867 9693 11868
rect 9995 11796 10061 11797
rect 9995 11732 9996 11796
rect 10060 11732 10061 11796
rect 9995 11731 10061 11732
rect 9627 10980 9693 10981
rect 9627 10916 9628 10980
rect 9692 10916 9693 10980
rect 9627 10915 9693 10916
rect 8891 10300 8957 10301
rect 8891 10236 8892 10300
rect 8956 10236 8957 10300
rect 8891 10235 8957 10236
rect 8340 9760 8348 9824
rect 8412 9760 8428 9824
rect 8492 9760 8508 9824
rect 8572 9760 8588 9824
rect 8652 9760 8660 9824
rect 8340 8736 8660 9760
rect 9443 9348 9509 9349
rect 9443 9284 9444 9348
rect 9508 9284 9509 9348
rect 9443 9283 9509 9284
rect 8340 8672 8348 8736
rect 8412 8672 8428 8736
rect 8492 8672 8508 8736
rect 8572 8672 8588 8736
rect 8652 8672 8660 8736
rect 8155 8668 8221 8669
rect 8155 8604 8156 8668
rect 8220 8604 8221 8668
rect 8155 8603 8221 8604
rect 8158 3773 8218 8603
rect 8340 7648 8660 8672
rect 9075 7852 9141 7853
rect 9075 7788 9076 7852
rect 9140 7788 9141 7852
rect 9075 7787 9141 7788
rect 8340 7584 8348 7648
rect 8412 7584 8428 7648
rect 8492 7584 8508 7648
rect 8572 7584 8588 7648
rect 8652 7584 8660 7648
rect 8340 6560 8660 7584
rect 8891 7580 8957 7581
rect 8891 7516 8892 7580
rect 8956 7516 8957 7580
rect 8891 7515 8957 7516
rect 8340 6496 8348 6560
rect 8412 6496 8428 6560
rect 8492 6496 8508 6560
rect 8572 6496 8588 6560
rect 8652 6496 8660 6560
rect 8340 5472 8660 6496
rect 8894 5538 8954 7515
rect 8340 5408 8348 5472
rect 8412 5408 8428 5472
rect 8492 5408 8508 5472
rect 8572 5408 8588 5472
rect 8652 5408 8660 5472
rect 8340 4384 8660 5408
rect 8340 4320 8348 4384
rect 8412 4320 8428 4384
rect 8492 4320 8508 4384
rect 8572 4320 8588 4384
rect 8652 4320 8660 4384
rect 8155 3772 8221 3773
rect 8155 3708 8156 3772
rect 8220 3708 8221 3772
rect 8155 3707 8221 3708
rect 8340 3296 8660 4320
rect 8756 5478 8954 5538
rect 8756 4042 8816 5478
rect 8891 5404 8957 5405
rect 8891 5340 8892 5404
rect 8956 5340 8957 5404
rect 8891 5339 8957 5340
rect 8894 4181 8954 5339
rect 9078 4453 9138 7787
rect 9259 5948 9325 5949
rect 9259 5884 9260 5948
rect 9324 5884 9325 5948
rect 9259 5883 9325 5884
rect 9075 4452 9141 4453
rect 9075 4388 9076 4452
rect 9140 4388 9141 4452
rect 9075 4387 9141 4388
rect 9075 4316 9141 4317
rect 9075 4252 9076 4316
rect 9140 4252 9141 4316
rect 9075 4251 9141 4252
rect 8891 4180 8957 4181
rect 8891 4116 8892 4180
rect 8956 4116 8957 4180
rect 8891 4115 8957 4116
rect 8756 3982 8954 4042
rect 8340 3232 8348 3296
rect 8412 3232 8428 3296
rect 8492 3232 8508 3296
rect 8572 3232 8588 3296
rect 8652 3232 8660 3296
rect 7787 2684 7853 2685
rect 7787 2620 7788 2684
rect 7852 2620 7853 2684
rect 7787 2619 7853 2620
rect 6683 2412 6749 2413
rect 6683 2348 6684 2412
rect 6748 2348 6749 2412
rect 6683 2347 6749 2348
rect 8340 2208 8660 3232
rect 8894 2685 8954 3982
rect 8891 2684 8957 2685
rect 8891 2620 8892 2684
rect 8956 2620 8957 2684
rect 8891 2619 8957 2620
rect 8340 2144 8348 2208
rect 8412 2144 8428 2208
rect 8492 2144 8508 2208
rect 8572 2144 8588 2208
rect 8652 2144 8660 2208
rect 8340 2128 8660 2144
rect 9078 1461 9138 4251
rect 9262 2549 9322 5883
rect 9446 4314 9506 9283
rect 9630 4453 9690 10915
rect 9998 10845 10058 11731
rect 9995 10844 10061 10845
rect 9995 10780 9996 10844
rect 10060 10780 10061 10844
rect 9995 10779 10061 10780
rect 10182 10570 10242 15947
rect 10805 15808 11125 15824
rect 10805 15744 10813 15808
rect 10877 15744 10893 15808
rect 10957 15744 10973 15808
rect 11037 15744 11053 15808
rect 11117 15744 11125 15808
rect 10805 14720 11125 15744
rect 12571 15604 12637 15605
rect 12571 15540 12572 15604
rect 12636 15540 12637 15604
rect 12571 15539 12637 15540
rect 10805 14656 10813 14720
rect 10877 14656 10893 14720
rect 10957 14656 10973 14720
rect 11037 14656 11053 14720
rect 11117 14656 11125 14720
rect 10363 14108 10429 14109
rect 10363 14044 10364 14108
rect 10428 14044 10429 14108
rect 10363 14043 10429 14044
rect 10547 14108 10613 14109
rect 10547 14044 10548 14108
rect 10612 14044 10613 14108
rect 10547 14043 10613 14044
rect 10366 11933 10426 14043
rect 10550 13565 10610 14043
rect 10805 13632 11125 14656
rect 11467 14652 11533 14653
rect 11467 14588 11468 14652
rect 11532 14588 11533 14652
rect 11467 14587 11533 14588
rect 10805 13568 10813 13632
rect 10877 13568 10893 13632
rect 10957 13568 10973 13632
rect 11037 13568 11053 13632
rect 11117 13568 11125 13632
rect 10547 13564 10613 13565
rect 10547 13500 10548 13564
rect 10612 13500 10613 13564
rect 10547 13499 10613 13500
rect 10805 12544 11125 13568
rect 10805 12480 10813 12544
rect 10877 12480 10893 12544
rect 10957 12480 10973 12544
rect 11037 12480 11053 12544
rect 11117 12480 11125 12544
rect 10363 11932 10429 11933
rect 10363 11868 10364 11932
rect 10428 11868 10429 11932
rect 10363 11867 10429 11868
rect 10363 11796 10429 11797
rect 10363 11732 10364 11796
rect 10428 11732 10429 11796
rect 10363 11731 10429 11732
rect 9998 10510 10242 10570
rect 9811 8940 9877 8941
rect 9811 8876 9812 8940
rect 9876 8876 9877 8940
rect 9811 8875 9877 8876
rect 9814 6082 9874 8875
rect 9998 6493 10058 10510
rect 10179 10436 10245 10437
rect 10179 10372 10180 10436
rect 10244 10372 10245 10436
rect 10179 10371 10245 10372
rect 10182 6629 10242 10371
rect 10366 9621 10426 11731
rect 10805 11456 11125 12480
rect 11283 12068 11349 12069
rect 11283 12004 11284 12068
rect 11348 12004 11349 12068
rect 11283 12003 11349 12004
rect 10805 11392 10813 11456
rect 10877 11392 10893 11456
rect 10957 11392 10973 11456
rect 11037 11392 11053 11456
rect 11117 11392 11125 11456
rect 10805 10368 11125 11392
rect 10805 10304 10813 10368
rect 10877 10304 10893 10368
rect 10957 10304 10973 10368
rect 11037 10304 11053 10368
rect 11117 10304 11125 10368
rect 10363 9620 10429 9621
rect 10363 9556 10364 9620
rect 10428 9556 10429 9620
rect 10363 9555 10429 9556
rect 10179 6628 10245 6629
rect 10179 6564 10180 6628
rect 10244 6564 10245 6628
rect 10179 6563 10245 6564
rect 9995 6492 10061 6493
rect 9995 6428 9996 6492
rect 10060 6428 10061 6492
rect 9995 6427 10061 6428
rect 9768 6022 9874 6082
rect 9768 5538 9828 6022
rect 9998 5898 10058 6427
rect 9768 5478 9874 5538
rect 9627 4452 9693 4453
rect 9627 4388 9628 4452
rect 9692 4388 9693 4452
rect 9627 4387 9693 4388
rect 9446 4254 9690 4314
rect 9443 4180 9509 4181
rect 9443 4116 9444 4180
rect 9508 4116 9509 4180
rect 9443 4115 9509 4116
rect 9446 2821 9506 4115
rect 9630 4042 9690 4254
rect 9814 4181 9874 5478
rect 9998 4453 10058 5662
rect 10366 4861 10426 9555
rect 10805 9280 11125 10304
rect 10805 9216 10813 9280
rect 10877 9216 10893 9280
rect 10957 9216 10973 9280
rect 11037 9216 11053 9280
rect 11117 9216 11125 9280
rect 10805 8192 11125 9216
rect 10805 8128 10813 8192
rect 10877 8128 10893 8192
rect 10957 8128 10973 8192
rect 11037 8128 11053 8192
rect 11117 8128 11125 8192
rect 10547 8124 10613 8125
rect 10547 8060 10548 8124
rect 10612 8060 10613 8124
rect 10547 8059 10613 8060
rect 10550 7173 10610 8059
rect 10547 7172 10613 7173
rect 10547 7108 10548 7172
rect 10612 7108 10613 7172
rect 10547 7107 10613 7108
rect 10805 7104 11125 8128
rect 11286 8125 11346 12003
rect 11283 8124 11349 8125
rect 11283 8060 11284 8124
rect 11348 8060 11349 8124
rect 11283 8059 11349 8060
rect 11470 7717 11530 14587
rect 11835 13836 11901 13837
rect 11835 13772 11836 13836
rect 11900 13772 11901 13836
rect 11835 13771 11901 13772
rect 12387 13836 12453 13837
rect 12387 13772 12388 13836
rect 12452 13772 12453 13836
rect 12387 13771 12453 13772
rect 11651 12612 11717 12613
rect 11651 12548 11652 12612
rect 11716 12548 11717 12612
rect 11651 12547 11717 12548
rect 11654 11525 11714 12547
rect 11651 11524 11717 11525
rect 11651 11460 11652 11524
rect 11716 11460 11717 11524
rect 11651 11459 11717 11460
rect 11651 11252 11717 11253
rect 11651 11188 11652 11252
rect 11716 11188 11717 11252
rect 11651 11187 11717 11188
rect 11654 9893 11714 11187
rect 11838 9893 11898 13771
rect 12203 13564 12269 13565
rect 12203 13500 12204 13564
rect 12268 13500 12269 13564
rect 12203 13499 12269 13500
rect 12019 13292 12085 13293
rect 12019 13228 12020 13292
rect 12084 13228 12085 13292
rect 12019 13227 12085 13228
rect 12022 10845 12082 13227
rect 12019 10844 12085 10845
rect 12019 10780 12020 10844
rect 12084 10780 12085 10844
rect 12019 10779 12085 10780
rect 11651 9892 11717 9893
rect 11651 9828 11652 9892
rect 11716 9828 11717 9892
rect 11651 9827 11717 9828
rect 11835 9892 11901 9893
rect 11835 9828 11836 9892
rect 11900 9828 11901 9892
rect 11835 9827 11901 9828
rect 11654 9349 11714 9827
rect 11651 9348 11717 9349
rect 11651 9284 11652 9348
rect 11716 9284 11717 9348
rect 11651 9283 11717 9284
rect 12019 9076 12085 9077
rect 12019 9012 12020 9076
rect 12084 9012 12085 9076
rect 12019 9011 12085 9012
rect 11651 8804 11717 8805
rect 11651 8740 11652 8804
rect 11716 8740 11717 8804
rect 11651 8739 11717 8740
rect 11467 7716 11533 7717
rect 11467 7652 11468 7716
rect 11532 7652 11533 7716
rect 11467 7651 11533 7652
rect 11283 7444 11349 7445
rect 11283 7380 11284 7444
rect 11348 7380 11349 7444
rect 11283 7379 11349 7380
rect 10805 7040 10813 7104
rect 10877 7040 10893 7104
rect 10957 7040 10973 7104
rect 11037 7040 11053 7104
rect 11117 7040 11125 7104
rect 10805 6016 11125 7040
rect 10805 5952 10813 6016
rect 10877 5952 10893 6016
rect 10957 5952 10973 6016
rect 11037 5952 11053 6016
rect 11117 5952 11125 6016
rect 10805 4928 11125 5952
rect 10805 4864 10813 4928
rect 10877 4864 10893 4928
rect 10957 4864 10973 4928
rect 11037 4864 11053 4928
rect 11117 4864 11125 4928
rect 10363 4860 10429 4861
rect 10363 4796 10364 4860
rect 10428 4796 10429 4860
rect 10363 4795 10429 4796
rect 9995 4452 10061 4453
rect 9995 4388 9996 4452
rect 10060 4388 10061 4452
rect 9995 4387 10061 4388
rect 10547 4452 10613 4453
rect 10547 4388 10548 4452
rect 10612 4388 10613 4452
rect 10547 4387 10613 4388
rect 9811 4180 9877 4181
rect 9811 4116 9812 4180
rect 9876 4116 9877 4180
rect 9811 4115 9877 4116
rect 10363 4044 10429 4045
rect 10363 4042 10364 4044
rect 9630 3982 10364 4042
rect 10363 3980 10364 3982
rect 10428 3980 10429 4044
rect 10363 3979 10429 3980
rect 10550 3909 10610 4387
rect 10547 3908 10613 3909
rect 10547 3844 10548 3908
rect 10612 3844 10613 3908
rect 10547 3843 10613 3844
rect 10805 3840 11125 4864
rect 10805 3776 10813 3840
rect 10877 3776 10893 3840
rect 10957 3776 10973 3840
rect 11037 3776 11053 3840
rect 11117 3776 11125 3840
rect 9443 2820 9509 2821
rect 9443 2756 9444 2820
rect 9508 2756 9509 2820
rect 9443 2755 9509 2756
rect 10805 2752 11125 3776
rect 11286 2957 11346 7379
rect 11467 7172 11533 7173
rect 11467 7108 11468 7172
rect 11532 7108 11533 7172
rect 11467 7107 11533 7108
rect 11470 6629 11530 7107
rect 11654 7034 11714 8739
rect 11835 7036 11901 7037
rect 11835 7034 11836 7036
rect 11654 6974 11836 7034
rect 11467 6628 11533 6629
rect 11467 6564 11468 6628
rect 11532 6564 11533 6628
rect 11467 6563 11533 6564
rect 11467 6084 11533 6085
rect 11467 6020 11468 6084
rect 11532 6020 11533 6084
rect 11467 6019 11533 6020
rect 11283 2956 11349 2957
rect 11283 2892 11284 2956
rect 11348 2892 11349 2956
rect 11283 2891 11349 2892
rect 10805 2688 10813 2752
rect 10877 2688 10893 2752
rect 10957 2688 10973 2752
rect 11037 2688 11053 2752
rect 11117 2688 11125 2752
rect 9259 2548 9325 2549
rect 9259 2484 9260 2548
rect 9324 2484 9325 2548
rect 9259 2483 9325 2484
rect 10805 2128 11125 2688
rect 11470 2141 11530 6019
rect 11654 3093 11714 6974
rect 11835 6972 11836 6974
rect 11900 6972 11901 7036
rect 11835 6971 11901 6972
rect 11835 6628 11901 6629
rect 11835 6564 11836 6628
rect 11900 6564 11901 6628
rect 11835 6563 11901 6564
rect 11838 4997 11898 6563
rect 12022 5677 12082 9011
rect 12019 5676 12085 5677
rect 12019 5612 12020 5676
rect 12084 5612 12085 5676
rect 12019 5611 12085 5612
rect 11835 4996 11901 4997
rect 11835 4932 11836 4996
rect 11900 4932 11901 4996
rect 11835 4931 11901 4932
rect 11835 4860 11901 4861
rect 11835 4796 11836 4860
rect 11900 4796 11901 4860
rect 11835 4795 11901 4796
rect 11651 3092 11717 3093
rect 11651 3028 11652 3092
rect 11716 3028 11717 3092
rect 11651 3027 11717 3028
rect 11467 2140 11533 2141
rect 11467 2076 11468 2140
rect 11532 2076 11533 2140
rect 11467 2075 11533 2076
rect 11838 1597 11898 4795
rect 12022 4317 12082 5611
rect 12206 5541 12266 13499
rect 12390 7309 12450 13771
rect 12387 7308 12453 7309
rect 12387 7244 12388 7308
rect 12452 7244 12453 7308
rect 12387 7243 12453 7244
rect 12387 7172 12453 7173
rect 12387 7108 12388 7172
rect 12452 7108 12453 7172
rect 12387 7107 12453 7108
rect 12390 5813 12450 7107
rect 12574 6085 12634 15539
rect 12939 15468 13005 15469
rect 12939 15404 12940 15468
rect 13004 15404 13005 15468
rect 12939 15403 13005 15404
rect 12755 12612 12821 12613
rect 12755 12548 12756 12612
rect 12820 12548 12821 12612
rect 12755 12547 12821 12548
rect 12571 6084 12637 6085
rect 12571 6020 12572 6084
rect 12636 6020 12637 6084
rect 12571 6019 12637 6020
rect 12387 5812 12453 5813
rect 12387 5748 12388 5812
rect 12452 5748 12453 5812
rect 12387 5747 12453 5748
rect 12203 5540 12269 5541
rect 12203 5476 12204 5540
rect 12268 5476 12269 5540
rect 12203 5475 12269 5476
rect 12019 4316 12085 4317
rect 12019 4252 12020 4316
rect 12084 4252 12085 4316
rect 12019 4251 12085 4252
rect 12390 3773 12450 5747
rect 12571 5676 12637 5677
rect 12571 5612 12572 5676
rect 12636 5612 12637 5676
rect 12571 5611 12637 5612
rect 12019 3772 12085 3773
rect 12019 3708 12020 3772
rect 12084 3708 12085 3772
rect 12019 3707 12085 3708
rect 12387 3772 12453 3773
rect 12387 3708 12388 3772
rect 12452 3708 12453 3772
rect 12387 3707 12453 3708
rect 12022 2549 12082 3707
rect 12574 3365 12634 5611
rect 12203 3364 12269 3365
rect 12203 3300 12204 3364
rect 12268 3300 12269 3364
rect 12203 3299 12269 3300
rect 12571 3364 12637 3365
rect 12571 3300 12572 3364
rect 12636 3300 12637 3364
rect 12571 3299 12637 3300
rect 12206 2685 12266 3299
rect 12203 2684 12269 2685
rect 12203 2620 12204 2684
rect 12268 2620 12269 2684
rect 12203 2619 12269 2620
rect 12019 2548 12085 2549
rect 12019 2484 12020 2548
rect 12084 2484 12085 2548
rect 12019 2483 12085 2484
rect 12758 2413 12818 12547
rect 12942 7445 13002 15403
rect 13270 15264 13590 15824
rect 13270 15200 13278 15264
rect 13342 15200 13358 15264
rect 13422 15200 13438 15264
rect 13502 15200 13518 15264
rect 13582 15200 13590 15264
rect 13270 14176 13590 15200
rect 13270 14112 13278 14176
rect 13342 14112 13358 14176
rect 13422 14112 13438 14176
rect 13502 14112 13518 14176
rect 13582 14112 13590 14176
rect 13270 13088 13590 14112
rect 13270 13024 13278 13088
rect 13342 13024 13358 13088
rect 13422 13024 13438 13088
rect 13502 13024 13518 13088
rect 13582 13024 13590 13088
rect 13123 12884 13189 12885
rect 13123 12820 13124 12884
rect 13188 12820 13189 12884
rect 13123 12819 13189 12820
rect 12939 7444 13005 7445
rect 12939 7380 12940 7444
rect 13004 7380 13005 7444
rect 12939 7379 13005 7380
rect 12939 7308 13005 7309
rect 12939 7244 12940 7308
rect 13004 7244 13005 7308
rect 12939 7243 13005 7244
rect 12942 2549 13002 7243
rect 13126 3229 13186 12819
rect 13270 12000 13590 13024
rect 14411 12204 14477 12205
rect 14411 12140 14412 12204
rect 14476 12140 14477 12204
rect 14411 12139 14477 12140
rect 13270 11936 13278 12000
rect 13342 11936 13358 12000
rect 13422 11936 13438 12000
rect 13502 11936 13518 12000
rect 13582 11936 13590 12000
rect 13270 10912 13590 11936
rect 14043 11116 14109 11117
rect 14043 11052 14044 11116
rect 14108 11052 14109 11116
rect 14043 11051 14109 11052
rect 13270 10848 13278 10912
rect 13342 10848 13358 10912
rect 13422 10848 13438 10912
rect 13502 10848 13518 10912
rect 13582 10848 13590 10912
rect 13270 9824 13590 10848
rect 13270 9760 13278 9824
rect 13342 9760 13358 9824
rect 13422 9760 13438 9824
rect 13502 9760 13518 9824
rect 13582 9760 13590 9824
rect 13270 8736 13590 9760
rect 13270 8672 13278 8736
rect 13342 8672 13358 8736
rect 13422 8672 13438 8736
rect 13502 8672 13518 8736
rect 13582 8672 13590 8736
rect 13270 7648 13590 8672
rect 13859 8396 13925 8397
rect 13859 8332 13860 8396
rect 13924 8332 13925 8396
rect 13859 8331 13925 8332
rect 13675 7988 13741 7989
rect 13675 7924 13676 7988
rect 13740 7924 13741 7988
rect 13675 7923 13741 7924
rect 13270 7584 13278 7648
rect 13342 7584 13358 7648
rect 13422 7584 13438 7648
rect 13502 7584 13518 7648
rect 13582 7584 13590 7648
rect 13270 6560 13590 7584
rect 13270 6496 13278 6560
rect 13342 6496 13358 6560
rect 13422 6496 13438 6560
rect 13502 6496 13518 6560
rect 13582 6496 13590 6560
rect 13270 5472 13590 6496
rect 13678 6221 13738 7923
rect 13675 6220 13741 6221
rect 13675 6156 13676 6220
rect 13740 6156 13741 6220
rect 13675 6155 13741 6156
rect 13675 5812 13741 5813
rect 13675 5748 13676 5812
rect 13740 5748 13741 5812
rect 13675 5747 13741 5748
rect 13270 5408 13278 5472
rect 13342 5408 13358 5472
rect 13422 5408 13438 5472
rect 13502 5408 13518 5472
rect 13582 5408 13590 5472
rect 13270 4384 13590 5408
rect 13270 4320 13278 4384
rect 13342 4320 13358 4384
rect 13422 4320 13438 4384
rect 13502 4320 13518 4384
rect 13582 4320 13590 4384
rect 13270 3296 13590 4320
rect 13270 3232 13278 3296
rect 13342 3232 13358 3296
rect 13422 3232 13438 3296
rect 13502 3232 13518 3296
rect 13582 3232 13590 3296
rect 13123 3228 13189 3229
rect 13123 3164 13124 3228
rect 13188 3164 13189 3228
rect 13123 3163 13189 3164
rect 12939 2548 13005 2549
rect 12939 2484 12940 2548
rect 13004 2484 13005 2548
rect 12939 2483 13005 2484
rect 12755 2412 12821 2413
rect 12755 2348 12756 2412
rect 12820 2348 12821 2412
rect 12755 2347 12821 2348
rect 13270 2208 13590 3232
rect 13678 3093 13738 5747
rect 13862 5269 13922 8331
rect 14046 6765 14106 11051
rect 14227 8396 14293 8397
rect 14227 8332 14228 8396
rect 14292 8332 14293 8396
rect 14227 8331 14293 8332
rect 14043 6764 14109 6765
rect 14043 6700 14044 6764
rect 14108 6700 14109 6764
rect 14043 6699 14109 6700
rect 13859 5268 13925 5269
rect 13859 5204 13860 5268
rect 13924 5204 13925 5268
rect 13859 5203 13925 5204
rect 13675 3092 13741 3093
rect 13675 3028 13676 3092
rect 13740 3028 13741 3092
rect 13675 3027 13741 3028
rect 13270 2144 13278 2208
rect 13342 2144 13358 2208
rect 13422 2144 13438 2208
rect 13502 2144 13518 2208
rect 13582 2144 13590 2208
rect 13270 2128 13590 2144
rect 14230 1869 14290 8331
rect 14414 4045 14474 12139
rect 14963 11252 15029 11253
rect 14963 11188 14964 11252
rect 15028 11188 15029 11252
rect 14963 11187 15029 11188
rect 14966 9621 15026 11187
rect 14963 9620 15029 9621
rect 14963 9556 14964 9620
rect 15028 9556 15029 9620
rect 14963 9555 15029 9556
rect 14963 8260 15029 8261
rect 14963 8196 14964 8260
rect 15028 8196 15029 8260
rect 14963 8195 15029 8196
rect 14779 7172 14845 7173
rect 14779 7108 14780 7172
rect 14844 7108 14845 7172
rect 14779 7107 14845 7108
rect 14782 4861 14842 7107
rect 14779 4860 14845 4861
rect 14779 4796 14780 4860
rect 14844 4796 14845 4860
rect 14779 4795 14845 4796
rect 14411 4044 14477 4045
rect 14411 3980 14412 4044
rect 14476 3980 14477 4044
rect 14411 3979 14477 3980
rect 14966 2957 15026 8195
rect 14963 2956 15029 2957
rect 14963 2892 14964 2956
rect 15028 2892 15029 2956
rect 14963 2891 15029 2892
rect 14227 1868 14293 1869
rect 14227 1804 14228 1868
rect 14292 1804 14293 1868
rect 14227 1803 14293 1804
rect 11835 1596 11901 1597
rect 11835 1532 11836 1596
rect 11900 1532 11901 1596
rect 11835 1531 11901 1532
rect 9075 1460 9141 1461
rect 9075 1396 9076 1460
rect 9140 1396 9141 1460
rect 9075 1395 9141 1396
<< via4 >>
rect 4022 5812 4258 5898
rect 4022 5748 4108 5812
rect 4108 5748 4172 5812
rect 4172 5748 4258 5812
rect 4022 5662 4258 5748
rect 9910 5662 10146 5898
<< metal5 >>
rect 3980 5898 10188 5940
rect 3980 5662 4022 5898
rect 4258 5662 9910 5898
rect 10146 5662 10188 5898
rect 3980 5620 10188 5662
use sky130_fd_sc_hd__decap_3  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1380 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1605641404
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1605641404
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1472 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1656 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_15 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18
timestamp 1605641404
transform 1 0 2760 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10
timestamp 1605641404
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l1_in_0_
timestamp 1605641404
transform 1 0 2668 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2208 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_0_
timestamp 1605641404
transform 1 0 2944 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1605641404
transform 1 0 4692 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 4048 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_1_
timestamp 1605641404
transform 1 0 4784 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_0_
timestamp 1605641404
transform 1 0 3680 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1605641404
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38
timestamp 1605641404
transform 1 0 4600 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_26
timestamp 1605641404
transform 1 0 3496 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_37
timestamp 1605641404
transform 1 0 4508 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l1_in_0_
timestamp 1605641404
transform 1 0 5796 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_0_
timestamp 1605641404
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l4_in_0_
timestamp 1605641404
transform 1 0 5704 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1605641404
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1605641404
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49
timestamp 1605641404
transform 1 0 5612 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60
timestamp 1605641404
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_48
timestamp 1605641404
transform 1 0 5520 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1605641404
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_0_
timestamp 1605641404
transform 1 0 7084 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7820 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63
timestamp 1605641404
transform 1 0 6900 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74
timestamp 1605641404
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_71
timestamp 1605641404
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_82
timestamp 1605641404
transform 1 0 8648 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_93
timestamp 1605641404
transform 1 0 9660 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1605641404
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1605641404
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1605641404
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_1_
timestamp 1605641404
transform 1 0 8832 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _51_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 9108 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1605641404
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1605641404
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l3_in_0_
timestamp 1605641404
transform 1 0 9844 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_104
timestamp 1605641404
transform 1 0 10672 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114
timestamp 1605641404
transform 1 0 11592 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_1_
timestamp 1605641404
transform 1 0 10764 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1605641404
transform 1 0 10856 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1605641404
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_115
timestamp 1605641404
transform 1 0 11684 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 12144 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1605641404
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_1_
timestamp 1605641404
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1605641404
transform 1 0 11776 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _32_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 11868 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1605641404
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1605641404
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_129
timestamp 1605641404
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_132
timestamp 1605641404
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1605641404
transform 1 0 13432 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1605641404
transform 1 0 13156 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_138
timestamp 1605641404
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_135
timestamp 1605641404
transform 1 0 13524 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1605641404
transform 1 0 13708 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_144
timestamp 1605641404
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1605641404
transform 1 0 14076 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1605641404
transform 1 0 13984 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1605641404
transform 1 0 14260 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_150 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 14904 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1605641404
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1605641404
transform 1 0 14536 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1605641404
transform 1 0 14812 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_156
timestamp 1605641404
transform 1 0 15456 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156
timestamp 1605641404
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1605641404
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1605641404
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1605641404
transform -1 0 15824 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1605641404
transform -1 0 15824 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1605641404
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l4_in_0_
timestamp 1605641404
transform 1 0 1932 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_1_
timestamp 1605641404
transform 1 0 2944 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1605641404
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_7
timestamp 1605641404
transform 1 0 1748 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_18
timestamp 1605641404
transform 1 0 2760 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_0_
timestamp 1605641404
transform 1 0 4324 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1605641404
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1605641404
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_32
timestamp 1605641404
transform 1 0 4048 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l1_in_0_
timestamp 1605641404
transform 1 0 6716 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l4_in_0_
timestamp 1605641404
transform 1 0 5336 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6440 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_44
timestamp 1605641404
transform 1 0 5152 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_55
timestamp 1605641404
transform 1 0 6164 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1605641404
transform 1 0 8740 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_1_
timestamp 1605641404
transform 1 0 7728 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_70
timestamp 1605641404
transform 1 0 7544 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_81
timestamp 1605641404
transform 1 0 8556 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_2_
timestamp 1605641404
transform 1 0 10672 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_2_
timestamp 1605641404
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1605641404
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_87
timestamp 1605641404
transform 1 0 9108 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_91
timestamp 1605641404
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_102
timestamp 1605641404
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1605641404
transform 1 0 11684 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_113
timestamp 1605641404
transform 1 0 11500 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_124
timestamp 1605641404
transform 1 0 12512 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_1_
timestamp 1605641404
transform 1 0 13708 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_3_
timestamp 1605641404
transform 1 0 12696 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_135
timestamp 1605641404
transform 1 0 13524 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1605641404
transform -1 0 15824 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1605641404
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_146
timestamp 1605641404
transform 1 0 14536 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_152
timestamp 1605641404
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_154
timestamp 1605641404
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 2668 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_0_
timestamp 1605641404
transform 1 0 1656 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1605641404
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1605641404
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_15
timestamp 1605641404
transform 1 0 2484 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4692 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1605641404
transform 1 0 4416 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_33
timestamp 1605641404
transform 1 0 4140 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 6808 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_0_
timestamp 1605641404
transform 1 0 5704 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1605641404
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_48
timestamp 1605641404
transform 1 0 5520 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1605641404
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_2_
timestamp 1605641404
transform 1 0 8464 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_78
timestamp 1605641404
transform 1 0 8280 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_1_
timestamp 1605641404
transform 1 0 9476 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_1_
timestamp 1605641404
transform 1 0 10488 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_89
timestamp 1605641404
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_100
timestamp 1605641404
transform 1 0 10304 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1605641404
transform 1 0 11500 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1605641404
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1605641404
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_111
timestamp 1605641404
transform 1 0 11316 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_117
timestamp 1605641404
transform 1 0 11868 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_121
timestamp 1605641404
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_2_
timestamp 1605641404
transform 1 0 14444 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_2_
timestamp 1605641404
transform 1 0 13432 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_132
timestamp 1605641404
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_143
timestamp 1605641404
transform 1 0 14260 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1605641404
transform -1 0 15824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_154
timestamp 1605641404
transform 1 0 15272 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1605641404
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 2944 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1605641404
transform 1 0 1932 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1605641404
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_7
timestamp 1605641404
transform 1 0 1748 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_18
timestamp 1605641404
transform 1 0 2760 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1605641404
transform 1 0 4140 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_0_
timestamp 1605641404
transform 1 0 4692 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1605641404
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1605641404
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_32
timestamp 1605641404
transform 1 0 4048 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_37
timestamp 1605641404
transform 1 0 4508 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 6716 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_1_
timestamp 1605641404
transform 1 0 5704 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_48
timestamp 1605641404
transform 1 0 5520 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_59
timestamp 1605641404
transform 1 0 6532 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_1_
timestamp 1605641404
transform 1 0 8372 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_77
timestamp 1605641404
transform 1 0 8188 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_3_
timestamp 1605641404
transform 1 0 10672 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_2_
timestamp 1605641404
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1605641404
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_88
timestamp 1605641404
transform 1 0 9200 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_102
timestamp 1605641404
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 12512 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_0_
timestamp 1605641404
transform 1 0 11684 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_113
timestamp 1605641404
transform 1 0 11500 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_3_
timestamp 1605641404
transform 1 0 13708 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 13524 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_133
timestamp 1605641404
transform 1 0 13340 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1605641404
transform -1 0 15824 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1605641404
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_146
timestamp 1605641404
transform 1 0 14536 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1605641404
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_154
timestamp 1605641404
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1605641404
transform 1 0 1472 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1605641404
transform 1 0 1840 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1605641404
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1605641404
transform 1 0 2852 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp 1605641404
transform 1 0 1380 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_17
timestamp 1605641404
transform 1 0 2668 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_1_
timestamp 1605641404
transform 1 0 4048 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l4_in_0_
timestamp 1605641404
transform 1 0 3036 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_30
timestamp 1605641404
transform 1 0 3864 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_41
timestamp 1605641404
transform 1 0 4876 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 6808 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 5060 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1605641404
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1605641404
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 8464 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_78
timestamp 1605641404
transform 1 0 8280 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_3_
timestamp 1605641404
transform 1 0 10120 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_96
timestamp 1605641404
transform 1 0 9936 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_3_
timestamp 1605641404
transform 1 0 11132 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_1_
timestamp 1605641404
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1605641404
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_107
timestamp 1605641404
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_118
timestamp 1605641404
transform 1 0 11960 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_1_
timestamp 1605641404
transform 1 0 13432 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_2_
timestamp 1605641404
transform 1 0 14444 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_132
timestamp 1605641404
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_143
timestamp 1605641404
transform 1 0 14260 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1605641404
transform -1 0 15824 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_154
timestamp 1605641404
transform 1 0 15272 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_7
timestamp 1605641404
transform 1 0 1748 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1605641404
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1605641404
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l4_in_0_
timestamp 1605641404
transform 1 0 1932 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_0_
timestamp 1605641404
transform 1 0 1380 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1605641404
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_12
timestamp 1605641404
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_18
timestamp 1605641404
transform 1 0 2760 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_1_
timestamp 1605641404
transform 1 0 2392 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l4_in_0_
timestamp 1605641404
transform 1 0 2944 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1605641404
transform 1 0 4600 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 3404 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 4048 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1605641404
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1605641404
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_41
timestamp 1605641404
transform 1 0 4876 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_23
timestamp 1605641404
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_41
timestamp 1605641404
transform 1 0 4876 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6624 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 5060 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4968 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1605641404
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_58
timestamp 1605641404
transform 1 0 6440 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1605641404
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_62
timestamp 1605641404
transform 1 0 6808 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6900 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 8556 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8280 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_76
timestamp 1605641404
transform 1 0 8096 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_79
timestamp 1605641404
transform 1 0 8372 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 10212 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_3_
timestamp 1605641404
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_1_
timestamp 1605641404
transform 1 0 10672 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1605641404
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1605641404
transform 1 0 9292 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_87
timestamp 1605641404
transform 1 0 9108 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_102
timestamp 1605641404
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_97
timestamp 1605641404
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1605641404
transform 1 0 11868 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_0_
timestamp 1605641404
transform 1 0 11684 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_1_
timestamp 1605641404
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1605641404
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_113
timestamp 1605641404
transform 1 0 11500 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_124
timestamp 1605641404
transform 1 0 12512 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_115
timestamp 1605641404
transform 1 0 11684 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1605641404
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_2_
timestamp 1605641404
transform 1 0 14444 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1605641404
transform 1 0 13708 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_1_
timestamp 1605641404
transform 1 0 13432 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_2_
timestamp 1605641404
transform 1 0 12696 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_135
timestamp 1605641404
transform 1 0 13524 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_132
timestamp 1605641404
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_143
timestamp 1605641404
transform 1 0 14260 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1605641404
transform 1 0 14720 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1605641404
transform -1 0 15824 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1605641404
transform -1 0 15824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1605641404
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_146
timestamp 1605641404
transform 1 0 14536 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1605641404
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_154
timestamp 1605641404
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_154
timestamp 1605641404
transform 1 0 15272 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 2300 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1564 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1605641404
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1605641404
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_11
timestamp 1605641404
transform 1 0 2116 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1605641404
transform 1 0 4048 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l4_in_0_
timestamp 1605641404
transform 1 0 4508 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1605641404
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1605641404
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_35
timestamp 1605641404
transform 1 0 4324 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 5520 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_46
timestamp 1605641404
transform 1 0 5336 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7176 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8648 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_64
timestamp 1605641404
transform 1 0 6992 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9660 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1605641404
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1605641404
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_2_
timestamp 1605641404
transform 1 0 11316 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_1_
timestamp 1605641404
transform 1 0 12328 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_109
timestamp 1605641404
transform 1 0 11132 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_120
timestamp 1605641404
transform 1 0 12144 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1605641404
transform 1 0 14352 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_2_
timestamp 1605641404
transform 1 0 13340 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_131
timestamp 1605641404
transform 1 0 13156 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_142
timestamp 1605641404
transform 1 0 14168 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1605641404
transform -1 0 15824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1605641404
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1605641404
transform 1 0 14904 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_148
timestamp 1605641404
transform 1 0 14720 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_154
timestamp 1605641404
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_0_
timestamp 1605641404
transform 1 0 1380 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_0_
timestamp 1605641404
transform 1 0 2392 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1605641404
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_12
timestamp 1605641404
transform 1 0 2208 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 3404 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_23
timestamp 1605641404
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_41
timestamp 1605641404
transform 1 0 4876 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 5060 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 6808 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1605641404
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1605641404
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 8464 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_78
timestamp 1605641404
transform 1 0 8280 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 10120 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_96
timestamp 1605641404
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1605641404
transform 1 0 11776 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_2_
timestamp 1605641404
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1605641404
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_114
timestamp 1605641404
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1605641404
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_2_
timestamp 1605641404
transform 1 0 13432 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_1_
timestamp 1605641404
transform 1 0 14444 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_132
timestamp 1605641404
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_143
timestamp 1605641404
transform 1 0 14260 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1605641404
transform -1 0 15824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_154
timestamp 1605641404
transform 1 0 15272 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 2300 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1564 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1605641404
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1605641404
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_11
timestamp 1605641404
transform 1 0 2116 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4600 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 4048 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1605641404
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1605641404
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6072 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 7544 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 9660 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 9016 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1605641404
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 11316 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_109
timestamp 1605641404
transform 1 0 11132 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_0_
timestamp 1605641404
transform 1 0 13984 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_3_
timestamp 1605641404
transform 1 0 12972 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_127
timestamp 1605641404
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1605641404
transform 1 0 13800 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1605641404
transform -1 0 15824 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1605641404
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_149
timestamp 1605641404
transform 1 0 14812 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_154
timestamp 1605641404
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 1748 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1605641404
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1605641404
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 3404 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_23
timestamp 1605641404
transform 1 0 3220 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_41
timestamp 1605641404
transform 1 0 4876 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1605641404
transform 1 0 6808 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 5060 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1605641404
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1605641404
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7912 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1605641404
transform 1 0 7360 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_66
timestamp 1605641404
transform 1 0 7176 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_71
timestamp 1605641404
transform 1 0 7636 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9384 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1605641404
transform 1 0 11868 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 12420 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_0_
timestamp 1605641404
transform 1 0 10856 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1605641404
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_115
timestamp 1605641404
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1605641404
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_0_
timestamp 1605641404
transform 1 0 14076 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_139
timestamp 1605641404
transform 1 0 13892 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1605641404
transform 1 0 15088 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1605641404
transform -1 0 15824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_150
timestamp 1605641404
transform 1 0 14904 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_155
timestamp 1605641404
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 2300 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1564 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1605641404
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1605641404
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_11
timestamp 1605641404
transform 1 0 2116 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4232 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1605641404
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1605641404
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_32
timestamp 1605641404
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 5704 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 7360 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_12_66
timestamp 1605641404
transform 1 0 7176 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 9660 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1605641404
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_88
timestamp 1605641404
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 11316 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_109
timestamp 1605641404
transform 1 0 11132 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12972 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_127
timestamp 1605641404
transform 1 0 12788 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_145
timestamp 1605641404
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1605641404
transform 1 0 14628 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1605641404
transform -1 0 15824 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1605641404
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_150
timestamp 1605641404
transform 1 0 14904 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_154
timestamp 1605641404
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 2300 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 1748 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1564 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1605641404
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1605641404
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1605641404
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1605641404
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_11
timestamp 1605641404
transform 1 0 2116 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 3404 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4140 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1605641404
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_23
timestamp 1605641404
transform 1 0 3220 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_41
timestamp 1605641404
transform 1 0 4876 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1605641404
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_32
timestamp 1605641404
transform 1 0 4048 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 5796 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 5060 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1605641404
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1605641404
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_62
timestamp 1605641404
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_49
timestamp 1605641404
transform 1 0 5612 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1605641404
transform 1 0 7452 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 8280 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 7912 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_1_
timestamp 1605641404
transform 1 0 6992 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1605641404
transform 1 0 8004 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_73
timestamp 1605641404
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_67
timestamp 1605641404
transform 1 0 7268 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_72
timestamp 1605641404
transform 1 0 7728 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9936 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 9660 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1605641404
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_94
timestamp 1605641404
transform 1 0 9752 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1605641404
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1605641404
transform 1 0 11592 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 11316 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12420 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1605641404
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1605641404
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_112
timestamp 1605641404
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_117
timestamp 1605641404
transform 1 0 11868 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_109
timestamp 1605641404
transform 1 0 11132 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_2_
timestamp 1605641404
transform 1 0 12972 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_2_
timestamp 1605641404
transform 1 0 14076 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_2_
timestamp 1605641404
transform 1 0 13984 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_139
timestamp 1605641404
transform 1 0 13892 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_127
timestamp 1605641404
transform 1 0 12788 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1605641404
transform 1 0 13800 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1605641404
transform 1 0 15088 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1605641404
transform -1 0 15824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1605641404
transform -1 0 15824 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1605641404
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_150
timestamp 1605641404
transform 1 0 14904 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_155
timestamp 1605641404
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_149
timestamp 1605641404
transform 1 0 14812 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_154
timestamp 1605641404
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l4_in_0_
timestamp 1605641404
transform 1 0 1380 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_1_
timestamp 1605641404
transform 1 0 2392 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1605641404
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_12
timestamp 1605641404
transform 1 0 2208 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 3404 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_23
timestamp 1605641404
transform 1 0 3220 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_41
timestamp 1605641404
transform 1 0 4876 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 6808 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 5060 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1605641404
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1605641404
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8464 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_78
timestamp 1605641404
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 9476 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_89
timestamp 1605641404
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_3_
timestamp 1605641404
transform 1 0 11132 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_3_
timestamp 1605641404
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1605641404
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_107
timestamp 1605641404
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1605641404
transform 1 0 11960 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_2_
timestamp 1605641404
transform 1 0 14444 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_0_
timestamp 1605641404
transform 1 0 13432 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_132
timestamp 1605641404
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_143
timestamp 1605641404
transform 1 0 14260 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1605641404
transform -1 0 15824 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_154
timestamp 1605641404
transform 1 0 15272 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1605641404
transform 1 0 1472 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l4_in_0_
timestamp 1605641404
transform 1 0 2944 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_0_
timestamp 1605641404
transform 1 0 1932 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1605641404
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1605641404
transform 1 0 1748 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1605641404
transform 1 0 1380 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_18
timestamp 1605641404
transform 1 0 2760 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 4324 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1605641404
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1605641404
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_32
timestamp 1605641404
transform 1 0 4048 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 5980 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_51
timestamp 1605641404
transform 1 0 5796 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 7636 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_69
timestamp 1605641404
transform 1 0 7452 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 9660 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1605641404
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1605641404
transform 1 0 9292 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_87
timestamp 1605641404
transform 1 0 9108 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_1_
timestamp 1605641404
transform 1 0 11316 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l4_in_0_
timestamp 1605641404
transform 1 0 12328 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_109
timestamp 1605641404
transform 1 0 11132 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_120
timestamp 1605641404
transform 1 0 12144 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1605641404
transform 1 0 14352 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_3_
timestamp 1605641404
transform 1 0 13340 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_131
timestamp 1605641404
transform 1 0 13156 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_142
timestamp 1605641404
transform 1 0 14168 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1605641404
transform -1 0 15824 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1605641404
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1605641404
transform 1 0 14812 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_147
timestamp 1605641404
transform 1 0 14628 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1605641404
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_154
timestamp 1605641404
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_1_
timestamp 1605641404
transform 1 0 2024 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1605641404
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1605641404
transform 1 0 1748 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1605641404
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_19
timestamp 1605641404
transform 1 0 2852 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_1_
timestamp 1605641404
transform 1 0 4048 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_1_
timestamp 1605641404
transform 1 0 3036 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_30
timestamp 1605641404
transform 1 0 3864 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_41
timestamp 1605641404
transform 1 0 4876 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 5060 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 6808 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1605641404
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1605641404
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 8464 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_78
timestamp 1605641404
transform 1 0 8280 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 10120 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_96
timestamp 1605641404
transform 1 0 9936 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1605641404
transform 1 0 11776 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_0_
timestamp 1605641404
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1605641404
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_114
timestamp 1605641404
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_119
timestamp 1605641404
transform 1 0 12052 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_3_
timestamp 1605641404
transform 1 0 13432 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_3_
timestamp 1605641404
transform 1 0 14444 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_132
timestamp 1605641404
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_143
timestamp 1605641404
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1605641404
transform -1 0 15824 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_154
timestamp 1605641404
transform 1 0 15272 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_0_
timestamp 1605641404
transform 1 0 2944 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_1_
timestamp 1605641404
transform 1 0 1932 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1605641404
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1605641404
transform 1 0 1656 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1605641404
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_18
timestamp 1605641404
transform 1 0 2760 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l4_in_0_
timestamp 1605641404
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1605641404
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1605641404
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_41
timestamp 1605641404
transform 1 0 4876 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 5060 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 6716 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_59
timestamp 1605641404
transform 1 0 6532 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_2_
timestamp 1605641404
transform 1 0 8372 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_77
timestamp 1605641404
transform 1 0 8188 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_0_
timestamp 1605641404
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_0_
timestamp 1605641404
transform 1 0 10672 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1605641404
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_88
timestamp 1605641404
transform 1 0 9200 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_102
timestamp 1605641404
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_1_
timestamp 1605641404
transform 1 0 11684 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_113
timestamp 1605641404
transform 1 0 11500 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_124
timestamp 1605641404
transform 1 0 12512 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_2_
timestamp 1605641404
transform 1 0 12696 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_3_
timestamp 1605641404
transform 1 0 13708 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_135
timestamp 1605641404
transform 1 0 13524 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1605641404
transform 1 0 14720 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1605641404
transform -1 0 15824 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1605641404
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_146
timestamp 1605641404
transform 1 0 14536 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1605641404
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_154
timestamp 1605641404
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3
timestamp 1605641404
transform 1 0 1380 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp 1605641404
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1605641404
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1605641404
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l4_in_0_
timestamp 1605641404
transform 1 0 1656 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1472 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_18
timestamp 1605641404
transform 1 0 2760 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_10
timestamp 1605641404
transform 1 0 2024 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_15
timestamp 1605641404
transform 1 0 2484 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_0_
timestamp 1605641404
transform 1 0 2668 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2208 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_0_
timestamp 1605641404
transform 1 0 2944 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4692 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4232 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_0_
timestamp 1605641404
transform 1 0 3680 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1605641404
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_26
timestamp 1605641404
transform 1 0 3496 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_37
timestamp 1605641404
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1605641404
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_32
timestamp 1605641404
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 6256 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 6808 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_0_
timestamp 1605641404
transform 1 0 5704 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_0_
timestamp 1605641404
transform 1 0 5244 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1605641404
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_48
timestamp 1605641404
transform 1 0 5520 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1605641404
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_43
timestamp 1605641404
transform 1 0 5060 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_54
timestamp 1605641404
transform 1 0 6072 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7912 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_1_
timestamp 1605641404
transform 1 0 8464 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_78
timestamp 1605641404
transform 1 0 8280 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_72
timestamp 1605641404
transform 1 0 7728 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_83
timestamp 1605641404
transform 1 0 8740 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_89
timestamp 1605641404
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_89
timestamp 1605641404
transform 1 0 9292 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1605641404
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_2_
timestamp 1605641404
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_2_
timestamp 1605641404
transform 1 0 9476 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1605641404
transform 1 0 8924 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_102
timestamp 1605641404
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_100
timestamp 1605641404
transform 1 0 10304 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_3_
timestamp 1605641404
transform 1 0 10488 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_1_
timestamp 1605641404
transform 1 0 10672 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1605641404
transform 1 0 11500 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_0_
timestamp 1605641404
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_1_
timestamp 1605641404
transform 1 0 11684 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1605641404
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1605641404
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_111
timestamp 1605641404
transform 1 0 11316 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_117
timestamp 1605641404
transform 1 0 11868 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_113
timestamp 1605641404
transform 1 0 11500 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_124
timestamp 1605641404
transform 1 0 12512 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l3_in_1_
timestamp 1605641404
transform 1 0 13432 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l4_in_0_
timestamp 1605641404
transform 1 0 12696 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 13708 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_132
timestamp 1605641404
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_143 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 14260 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_135
timestamp 1605641404
transform 1 0 13524 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_143 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 14260 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1605641404
transform -1 0 15824 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1605641404
transform -1 0 15824 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1605641404
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_155
timestamp 1605641404
transform 1 0 15364 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1605641404
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_154
timestamp 1605641404
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1605641404
transform 1 0 1564 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2116 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2852 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1605641404
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1605641404
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_9
timestamp 1605641404
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_17
timestamp 1605641404
transform 1 0 2668 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l4_in_0_
timestamp 1605641404
transform 1 0 4692 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l4_in_0_
timestamp 1605641404
transform 1 0 3680 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_21_25
timestamp 1605641404
transform 1 0 3404 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_37
timestamp 1605641404
transform 1 0 4508 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l4_in_0_
timestamp 1605641404
transform 1 0 5704 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_0_
timestamp 1605641404
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1605641404
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_48
timestamp 1605641404
transform 1 0 5520 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1605641404
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_1_
timestamp 1605641404
transform 1 0 7820 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_71
timestamp 1605641404
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_82
timestamp 1605641404
transform 1 0 8648 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_3_
timestamp 1605641404
transform 1 0 9844 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_1_
timestamp 1605641404
transform 1 0 8832 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_93
timestamp 1605641404
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_104
timestamp 1605641404
transform 1 0 10672 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1605641404
transform 1 0 11868 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1605641404
transform 1 0 12420 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_2_
timestamp 1605641404
transform 1 0 10856 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1605641404
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_115
timestamp 1605641404
transform 1 0 11684 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_120
timestamp 1605641404
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_127
timestamp 1605641404
transform 1 0 12788 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_139
timestamp 1605641404
transform 1 0 13892 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1605641404
transform -1 0 15824 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_151
timestamp 1605641404
transform 1 0 14996 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1605641404
transform 1 0 1840 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1605641404
transform 1 0 2392 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2944 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1605641404
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1605641404
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_7
timestamp 1605641404
transform 1 0 1748 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_12
timestamp 1605641404
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_18
timestamp 1605641404
transform 1 0 2760 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4324 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1605641404
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_26
timestamp 1605641404
transform 1 0 3496 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_30
timestamp 1605641404
transform 1 0 3864 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_32
timestamp 1605641404
transform 1 0 4048 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_0_
timestamp 1605641404
transform 1 0 6348 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_0_
timestamp 1605641404
transform 1 0 5336 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_44
timestamp 1605641404
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_55
timestamp 1605641404
transform 1 0 6164 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_1_
timestamp 1605641404
transform 1 0 7360 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_1_
timestamp 1605641404
transform 1 0 8372 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_66
timestamp 1605641404
transform 1 0 7176 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_77
timestamp 1605641404
transform 1 0 8188 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_3_
timestamp 1605641404
transform 1 0 10672 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_1_
timestamp 1605641404
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1605641404
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_88
timestamp 1605641404
transform 1 0 9200 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_102
timestamp 1605641404
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1605641404
transform 1 0 11684 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1605641404
transform 1 0 12236 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_113
timestamp 1605641404
transform 1 0 11500 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_119
timestamp 1605641404
transform 1 0 12052 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_124
timestamp 1605641404
transform 1 0 12512 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_136
timestamp 1605641404
transform 1 0 13616 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1605641404
transform -1 0 15824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1605641404
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_148
timestamp 1605641404
transform 1 0 14720 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_152
timestamp 1605641404
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_154
timestamp 1605641404
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1605641404
transform 1 0 2208 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1605641404
transform 1 0 2760 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1605641404
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_3
timestamp 1605641404
transform 1 0 1380 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_11
timestamp 1605641404
transform 1 0 2116 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_16
timestamp 1605641404
transform 1 0 2576 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1605641404
transform 1 0 4600 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1605641404
transform 1 0 3312 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 3864 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_22
timestamp 1605641404
transform 1 0 3128 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_28
timestamp 1605641404
transform 1 0 3680 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_36
timestamp 1605641404
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1605641404
transform 1 0 6808 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1605641404
transform 1 0 5152 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_1_
timestamp 1605641404
transform 1 0 5704 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1605641404
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_42
timestamp 1605641404
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_48
timestamp 1605641404
transform 1 0 5520 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1605641404
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_1_
timestamp 1605641404
transform 1 0 7636 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_2_
timestamp 1605641404
transform 1 0 8648 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1605641404
transform 1 0 7360 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_66
timestamp 1605641404
transform 1 0 7176 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_80
timestamp 1605641404
transform 1 0 8464 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1605641404
transform 1 0 10672 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_2_
timestamp 1605641404
transform 1 0 9660 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_91
timestamp 1605641404
transform 1 0 9476 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_102
timestamp 1605641404
transform 1 0 10488 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1605641404
transform 1 0 11224 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1605641404
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_108
timestamp 1605641404
transform 1 0 11040 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_113
timestamp 1605641404
transform 1 0 11500 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1605641404
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1605641404
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1605641404
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1605641404
transform -1 0 15824 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_147
timestamp 1605641404
transform 1 0 14628 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_155
timestamp 1605641404
transform 1 0 15364 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1605641404
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1605641404
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_15
timestamp 1605641404
transform 1 0 2484 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1605641404
transform 1 0 4232 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1605641404
transform 1 0 4784 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1605641404
transform 1 0 3220 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1605641404
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1605641404
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_32
timestamp 1605641404
transform 1 0 4048 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_38
timestamp 1605641404
transform 1 0 4600 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 5796 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1605641404
transform 1 0 6808 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_44
timestamp 1605641404
transform 1 0 5152 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_50
timestamp 1605641404
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_60
timestamp 1605641404
transform 1 0 6624 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7084 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_1_
timestamp 1605641404
transform 1 0 8096 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_63
timestamp 1605641404
transform 1 0 6900 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_74
timestamp 1605641404
transform 1 0 7912 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1605641404
transform 1 0 9108 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1605641404
transform 1 0 9752 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1605641404
transform 1 0 10304 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1605641404
transform 1 0 9660 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1605641404
transform 1 0 8924 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_91
timestamp 1605641404
transform 1 0 9476 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_98
timestamp 1605641404
transform 1 0 10120 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_104
timestamp 1605641404
transform 1 0 10672 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1605641404
transform 1 0 12512 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_116
timestamp 1605641404
transform 1 0 11776 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_125
timestamp 1605641404
transform 1 0 12604 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_137
timestamp 1605641404
transform 1 0 13708 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1605641404
transform -1 0 15824 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1605641404
transform 1 0 15364 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_149
timestamp 1605641404
transform 1 0 14812 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_156
timestamp 1605641404
transform 1 0 15456 0 -1 15776
box -38 -48 130 592
<< labels >>
rlabel metal3 s 0 416 480 536 6 ccff_head
port 0 nsew default input
rlabel metal3 s 16520 8984 17000 9104 6 ccff_tail
port 1 nsew default tristate
rlabel metal2 s 8666 0 8722 480 6 chany_bottom_in[0]
port 2 nsew default input
rlabel metal2 s 12898 0 12954 480 6 chany_bottom_in[10]
port 3 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[11]
port 4 nsew default input
rlabel metal2 s 13818 0 13874 480 6 chany_bottom_in[12]
port 5 nsew default input
rlabel metal2 s 14186 0 14242 480 6 chany_bottom_in[13]
port 6 nsew default input
rlabel metal2 s 14646 0 14702 480 6 chany_bottom_in[14]
port 7 nsew default input
rlabel metal2 s 15014 0 15070 480 6 chany_bottom_in[15]
port 8 nsew default input
rlabel metal2 s 15474 0 15530 480 6 chany_bottom_in[16]
port 9 nsew default input
rlabel metal2 s 15934 0 15990 480 6 chany_bottom_in[17]
port 10 nsew default input
rlabel metal2 s 16302 0 16358 480 6 chany_bottom_in[18]
port 11 nsew default input
rlabel metal2 s 16762 0 16818 480 6 chany_bottom_in[19]
port 12 nsew default input
rlabel metal2 s 9126 0 9182 480 6 chany_bottom_in[1]
port 13 nsew default input
rlabel metal2 s 9494 0 9550 480 6 chany_bottom_in[2]
port 14 nsew default input
rlabel metal2 s 9954 0 10010 480 6 chany_bottom_in[3]
port 15 nsew default input
rlabel metal2 s 10414 0 10470 480 6 chany_bottom_in[4]
port 16 nsew default input
rlabel metal2 s 10782 0 10838 480 6 chany_bottom_in[5]
port 17 nsew default input
rlabel metal2 s 11242 0 11298 480 6 chany_bottom_in[6]
port 18 nsew default input
rlabel metal2 s 11610 0 11666 480 6 chany_bottom_in[7]
port 19 nsew default input
rlabel metal2 s 12070 0 12126 480 6 chany_bottom_in[8]
port 20 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[9]
port 21 nsew default input
rlabel metal2 s 202 0 258 480 6 chany_bottom_out[0]
port 22 nsew default tristate
rlabel metal2 s 4434 0 4490 480 6 chany_bottom_out[10]
port 23 nsew default tristate
rlabel metal2 s 4802 0 4858 480 6 chany_bottom_out[11]
port 24 nsew default tristate
rlabel metal2 s 5262 0 5318 480 6 chany_bottom_out[12]
port 25 nsew default tristate
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_out[13]
port 26 nsew default tristate
rlabel metal2 s 6090 0 6146 480 6 chany_bottom_out[14]
port 27 nsew default tristate
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_out[15]
port 28 nsew default tristate
rlabel metal2 s 7010 0 7066 480 6 chany_bottom_out[16]
port 29 nsew default tristate
rlabel metal2 s 7378 0 7434 480 6 chany_bottom_out[17]
port 30 nsew default tristate
rlabel metal2 s 7838 0 7894 480 6 chany_bottom_out[18]
port 31 nsew default tristate
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_out[19]
port 32 nsew default tristate
rlabel metal2 s 570 0 626 480 6 chany_bottom_out[1]
port 33 nsew default tristate
rlabel metal2 s 1030 0 1086 480 6 chany_bottom_out[2]
port 34 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_out[3]
port 35 nsew default tristate
rlabel metal2 s 1858 0 1914 480 6 chany_bottom_out[4]
port 36 nsew default tristate
rlabel metal2 s 2318 0 2374 480 6 chany_bottom_out[5]
port 37 nsew default tristate
rlabel metal2 s 2686 0 2742 480 6 chany_bottom_out[6]
port 38 nsew default tristate
rlabel metal2 s 3146 0 3202 480 6 chany_bottom_out[7]
port 39 nsew default tristate
rlabel metal2 s 3606 0 3662 480 6 chany_bottom_out[8]
port 40 nsew default tristate
rlabel metal2 s 3974 0 4030 480 6 chany_bottom_out[9]
port 41 nsew default tristate
rlabel metal2 s 8666 17520 8722 18000 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 12898 17520 12954 18000 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 13358 17520 13414 18000 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 13818 17520 13874 18000 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 14186 17520 14242 18000 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 14646 17520 14702 18000 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 15014 17520 15070 18000 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 15474 17520 15530 18000 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 15934 17520 15990 18000 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 16302 17520 16358 18000 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 16762 17520 16818 18000 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 9126 17520 9182 18000 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 9494 17520 9550 18000 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 9954 17520 10010 18000 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 10414 17520 10470 18000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 10782 17520 10838 18000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 11242 17520 11298 18000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 11610 17520 11666 18000 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 12070 17520 12126 18000 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 12530 17520 12586 18000 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 202 17520 258 18000 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 4434 17520 4490 18000 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 4802 17520 4858 18000 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 5262 17520 5318 18000 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 5722 17520 5778 18000 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 6090 17520 6146 18000 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 6550 17520 6606 18000 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 7010 17520 7066 18000 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 7378 17520 7434 18000 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 7838 17520 7894 18000 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 8206 17520 8262 18000 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 570 17520 626 18000 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 1030 17520 1086 18000 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 1398 17520 1454 18000 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 1858 17520 1914 18000 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 2318 17520 2374 18000 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 2686 17520 2742 18000 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 3146 17520 3202 18000 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 3606 17520 3662 18000 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 3974 17520 4030 18000 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 0 1368 480 1488 6 left_grid_pin_16_
port 82 nsew default tristate
rlabel metal3 s 0 2456 480 2576 6 left_grid_pin_17_
port 83 nsew default tristate
rlabel metal3 s 0 3544 480 3664 6 left_grid_pin_18_
port 84 nsew default tristate
rlabel metal3 s 0 4632 480 4752 6 left_grid_pin_19_
port 85 nsew default tristate
rlabel metal3 s 0 5584 480 5704 6 left_grid_pin_20_
port 86 nsew default tristate
rlabel metal3 s 0 6672 480 6792 6 left_grid_pin_21_
port 87 nsew default tristate
rlabel metal3 s 0 7760 480 7880 6 left_grid_pin_22_
port 88 nsew default tristate
rlabel metal3 s 0 8848 480 8968 6 left_grid_pin_23_
port 89 nsew default tristate
rlabel metal3 s 0 9800 480 9920 6 left_grid_pin_24_
port 90 nsew default tristate
rlabel metal3 s 0 10888 480 11008 6 left_grid_pin_25_
port 91 nsew default tristate
rlabel metal3 s 0 11976 480 12096 6 left_grid_pin_26_
port 92 nsew default tristate
rlabel metal3 s 0 13064 480 13184 6 left_grid_pin_27_
port 93 nsew default tristate
rlabel metal3 s 0 14016 480 14136 6 left_grid_pin_28_
port 94 nsew default tristate
rlabel metal3 s 0 15104 480 15224 6 left_grid_pin_29_
port 95 nsew default tristate
rlabel metal3 s 0 16192 480 16312 6 left_grid_pin_30_
port 96 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 left_grid_pin_31_
port 97 nsew default tristate
rlabel metal3 s 16520 3000 17000 3120 6 prog_clk
port 98 nsew default input
rlabel metal3 s 16520 14968 17000 15088 6 right_grid_pin_0_
port 99 nsew default tristate
rlabel metal4 s 3409 2128 3729 15824 6 VPWR
port 100 nsew default input
rlabel metal4 s 5875 2128 6195 15824 6 VGND
port 101 nsew default input
<< properties >>
string FIXED_BBOX 0 0 17000 18000
<< end >>
