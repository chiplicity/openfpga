* NGSPICE file created from cby_0__1_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor3_4 abstract view
.subckt scs8hd_nor3_4 A B C Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

.subckt cby_0__1_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] chany_bottom_in[0] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_out[0] chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3]
+ chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7]
+ chany_bottom_out[8] chany_top_in[0] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_out[0] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] data_in enable
+ left_grid_pin_0_ left_grid_pin_10_ left_grid_pin_12_ left_grid_pin_14_ left_grid_pin_2_
+ left_grid_pin_4_ left_grid_pin_6_ left_grid_pin_8_ right_grid_pin_3_ right_grid_pin_7_
+ vpwr vgnd
XFILLER_26_41 vgnd vpwr scs8hd_decap_3
XFILLER_9_115 vgnd vpwr scs8hd_decap_6
XANTENNA__113__B _112_/B vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_4.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[5] mux_right_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_6.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_39 vgnd vpwr scs8hd_decap_12
XFILLER_10_125 vgnd vpwr scs8hd_decap_12
XFILLER_37_62 vpwr vgnd scs8hd_fill_2
XANTENNA__108__B _109_/B vgnd vpwr scs8hd_diode_2
XANTENNA__124__A _088_/A vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_2_.latch/Q mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_ipin_6.LATCH_3_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_0.LATCH_1_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_062_ address[1] address[2] address[0] _062_/X vgnd vpwr scs8hd_or3_4
XFILLER_23_31 vgnd vpwr scs8hd_decap_4
X_131_ _131_/A _129_/B _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_75 vpwr vgnd scs8hd_fill_2
XFILLER_23_97 vpwr vgnd scs8hd_fill_2
XFILLER_48_83 vpwr vgnd scs8hd_fill_2
XANTENNA__110__C _118_/C vgnd vpwr scs8hd_diode_2
XFILLER_9_22 vgnd vpwr scs8hd_decap_3
XANTENNA__119__A _118_/X vgnd vpwr scs8hd_diode_2
XFILLER_50_3 vgnd vpwr scs8hd_decap_12
XFILLER_18_75 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_ipin_7.LATCH_0_.latch/Q mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_114_ _086_/A _112_/B _114_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__121__B _125_/B vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_2.LATCH_1_.latch data_in mem_right_ipin_2.LATCH_1_.latch/Q _097_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_32 vgnd vpwr scs8hd_decap_3
XFILLER_20_65 vpwr vgnd scs8hd_fill_2
XFILLER_29_96 vpwr vgnd scs8hd_fill_2
XFILLER_45_62 vgnd vpwr scs8hd_fill_1
XFILLER_45_51 vpwr vgnd scs8hd_fill_2
XFILLER_43_120 vpwr vgnd scs8hd_fill_2
XFILLER_35_109 vpwr vgnd scs8hd_fill_2
XANTENNA__116__B _112_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_89 vgnd vpwr scs8hd_decap_3
XANTENNA__132__A _166_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_3 vgnd vpwr scs8hd_decap_6
Xmem_right_ipin_4.LATCH_4_.latch data_in mem_right_ipin_4.LATCH_4_.latch/Q _113_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_109 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.INVTX1_5_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_4.LATCH_4_.latch_SLEEPB _113_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_145 vgnd vpwr scs8hd_fill_1
XFILLER_31_20 vgnd vpwr scs8hd_fill_1
XFILLER_31_53 vgnd vpwr scs8hd_decap_3
XFILLER_31_75 vgnd vpwr scs8hd_decap_4
XFILLER_56_83 vgnd vpwr scs8hd_decap_8
XFILLER_16_131 vgnd vpwr scs8hd_decap_12
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_101 vpwr vgnd scs8hd_fill_2
XFILLER_31_123 vgnd vpwr scs8hd_decap_12
XANTENNA__127__A address[5] vgnd vpwr scs8hd_diode_2
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_101 vgnd vpwr scs8hd_decap_4
XFILLER_13_112 vgnd vpwr scs8hd_decap_8
XFILLER_13_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_64 vgnd vpwr scs8hd_decap_4
XFILLER_26_86 vgnd vpwr scs8hd_fill_1
XFILLER_3_57 vpwr vgnd scs8hd_fill_2
XFILLER_10_137 vgnd vpwr scs8hd_decap_8
XFILLER_12_22 vgnd vpwr scs8hd_decap_8
XFILLER_12_66 vgnd vpwr scs8hd_decap_3
XFILLER_37_41 vgnd vpwr scs8hd_decap_3
XFILLER_37_96 vpwr vgnd scs8hd_fill_2
XFILLER_53_95 vpwr vgnd scs8hd_fill_2
XFILLER_53_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _175_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__124__B _125_/B vgnd vpwr scs8hd_diode_2
XANTENNA__140__A _166_/B vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_2.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[4] mux_right_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_130_ _159_/B _129_/B _130_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_10 vpwr vgnd scs8hd_fill_2
XFILLER_48_51 vgnd vpwr scs8hd_decap_4
XFILLER_64_94 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_2.LATCH_5_.latch_SLEEPB _093_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_58 vpwr vgnd scs8hd_fill_2
XFILLER_9_34 vpwr vgnd scs8hd_fill_2
XANTENNA__135__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_43_3 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_32 vgnd vpwr scs8hd_decap_4
XFILLER_18_43 vgnd vpwr scs8hd_decap_4
Xmux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _145_/A mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_ipin_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_113_ _085_/A _112_/B _113_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_50_41 vgnd vpwr scs8hd_decap_8
XFILLER_34_64 vpwr vgnd scs8hd_fill_2
XFILLER_59_72 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_46_140 vgnd vpwr scs8hd_decap_6
XFILLER_15_7 vgnd vpwr scs8hd_fill_1
Xmem_right_ipin_5.LATCH_0_.latch data_in mem_right_ipin_5.LATCH_0_.latch/Q _125_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_61_143 vgnd vpwr scs8hd_decap_3
XFILLER_61_121 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_29_75 vgnd vpwr scs8hd_fill_1
XFILLER_43_143 vgnd vpwr scs8hd_decap_3
XFILLER_61_51 vgnd vpwr scs8hd_decap_8
Xmem_right_ipin_7.LATCH_3_.latch data_in mem_right_ipin_7.LATCH_3_.latch/Q _139_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_4.INVTX1_3_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__132__B _129_/B vgnd vpwr scs8hd_diode_2
XFILLER_25_121 vgnd vpwr scs8hd_fill_1
XFILLER_31_32 vpwr vgnd scs8hd_fill_2
XFILLER_56_51 vpwr vgnd scs8hd_fill_2
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_143 vgnd vpwr scs8hd_decap_3
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_135 vgnd vpwr scs8hd_decap_8
XANTENNA__127__B _127_/B vgnd vpwr scs8hd_diode_2
XANTENNA__143__A _082_/C vgnd vpwr scs8hd_diode_2
XFILLER_22_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_5.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_26_10 vpwr vgnd scs8hd_fill_2
XFILLER_42_53 vgnd vpwr scs8hd_decap_8
XFILLER_13_135 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_ipin_6.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_36 vpwr vgnd scs8hd_fill_2
XFILLER_3_25 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__138__A _159_/B vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_ipin_6.LATCH_0_.latch/Q mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_78 vgnd vpwr scs8hd_decap_12
XFILLER_37_31 vpwr vgnd scs8hd_fill_2
XFILLER_37_53 vpwr vgnd scs8hd_fill_2
XFILLER_37_75 vpwr vgnd scs8hd_fill_2
XFILLER_53_74 vpwr vgnd scs8hd_fill_2
XFILLER_53_52 vpwr vgnd scs8hd_fill_2
XANTENNA__140__B _142_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_127 vpwr vgnd scs8hd_fill_2
XFILLER_59_105 vgnd vpwr scs8hd_decap_12
XFILLER_4_90 vpwr vgnd scs8hd_fill_2
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_145 vgnd vpwr scs8hd_fill_1
XFILLER_48_96 vpwr vgnd scs8hd_fill_2
XFILLER_0_15 vgnd vpwr scs8hd_decap_8
XFILLER_0_37 vpwr vgnd scs8hd_fill_2
X_189_ chany_bottom_in[8] chany_top_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_9_79 vpwr vgnd scs8hd_fill_2
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
XANTENNA__135__B _127_/B vgnd vpwr scs8hd_diode_2
XANTENNA__151__A _129_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_10 vpwr vgnd scs8hd_fill_2
XFILLER_34_32 vpwr vgnd scs8hd_fill_2
X_112_ _084_/A _112_/B _112_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_34_87 vgnd vpwr scs8hd_decap_4
XFILLER_59_95 vpwr vgnd scs8hd_fill_2
XFILLER_59_62 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_0.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[2] mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA__146__A _146_/A vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ right_grid_pin_7_ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_6.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_20_12 vpwr vgnd scs8hd_fill_2
XFILLER_20_23 vpwr vgnd scs8hd_fill_2
XFILLER_29_54 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_ipin_7.LATCH_5_.latch_SLEEPB _137_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_1.LATCH_0_.latch_SLEEPB _089_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_23 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_0.INVTX1_1_.scs8hd_inv_1 chany_top_in[0] mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_6.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__C _154_/C vgnd vpwr scs8hd_diode_2
XANTENNA__143__B _101_/X vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_7.INVTX1_3_.scs8hd_inv_1 chany_top_in[4] mux_right_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_87 vgnd vpwr scs8hd_decap_4
XFILLER_42_76 vpwr vgnd scs8hd_fill_2
XFILLER_42_32 vgnd vpwr scs8hd_decap_3
Xmem_right_ipin_0.LATCH_4_.latch data_in mem_right_ipin_0.LATCH_4_.latch/Q _072_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_15 vgnd vpwr scs8hd_decap_6
XANTENNA__138__B _142_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__154__A address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_left_ipin_0.LATCH_3_.latch/Q mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_12_46 vpwr vgnd scs8hd_fill_2
XANTENNA__064__A _156_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _176_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_143 vgnd vpwr scs8hd_decap_3
XFILLER_38_7 vgnd vpwr scs8hd_decap_12
XANTENNA__149__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_59_117 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_4.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_113 vgnd vpwr scs8hd_decap_12
XFILLER_2_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_27 vpwr vgnd scs8hd_fill_2
XFILLER_64_63 vgnd vpwr scs8hd_decap_12
X_188_ chany_top_in[0] chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA__135__C _099_/C vgnd vpwr scs8hd_diode_2
XFILLER_29_3 vgnd vpwr scs8hd_decap_4
XFILLER_18_12 vgnd vpwr scs8hd_decap_8
XFILLER_18_23 vpwr vgnd scs8hd_fill_2
XFILLER_18_56 vpwr vgnd scs8hd_fill_2
XFILLER_50_87 vgnd vpwr scs8hd_decap_4
XFILLER_50_76 vpwr vgnd scs8hd_fill_2
X_111_ _111_/A _112_/B vgnd vpwr scs8hd_buf_1
XFILLER_61_123 vgnd vpwr scs8hd_decap_12
XFILLER_61_101 vgnd vpwr scs8hd_decap_12
XANTENNA__162__A _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_109 vgnd vpwr scs8hd_decap_12
XFILLER_52_145 vgnd vpwr scs8hd_fill_1
XFILLER_1_70 vgnd vpwr scs8hd_decap_4
XFILLER_1_92 vpwr vgnd scs8hd_fill_2
XANTENNA__072__A _085_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_57 vgnd vpwr scs8hd_decap_6
XFILLER_29_33 vpwr vgnd scs8hd_fill_2
XFILLER_43_123 vgnd vpwr scs8hd_decap_12
XFILLER_43_112 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_61_86 vgnd vpwr scs8hd_decap_8
XFILLER_45_76 vpwr vgnd scs8hd_fill_2
XFILLER_61_97 vpwr vgnd scs8hd_fill_2
XFILLER_6_48 vgnd vpwr scs8hd_fill_1
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_7 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_ipin_5.LATCH_0_.latch/Q mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__157__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_1.LATCH_0_.latch data_in mem_right_ipin_1.LATCH_0_.latch/Q _089_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_25_123 vgnd vpwr scs8hd_decap_4
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
XFILLER_15_79 vpwr vgnd scs8hd_fill_2
XFILLER_25_145 vgnd vpwr scs8hd_fill_1
XANTENNA__067__A _066_/X vgnd vpwr scs8hd_diode_2
XFILLER_31_12 vpwr vgnd scs8hd_fill_2
XFILLER_56_64 vgnd vpwr scs8hd_fill_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__C _143_/C vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_1_.latch/Q mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_right_ipin_3.LATCH_3_.latch data_in mem_right_ipin_3.LATCH_3_.latch/Q _106_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_80 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_6.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_23 vpwr vgnd scs8hd_fill_2
XFILLER_26_89 vgnd vpwr scs8hd_decap_3
XFILLER_42_11 vgnd vpwr scs8hd_decap_3
XFILLER_59_3 vgnd vpwr scs8hd_decap_12
XANTENNA__154__B address[6] vgnd vpwr scs8hd_diode_2
XANTENNA__064__B _064_/B vgnd vpwr scs8hd_diode_2
XANTENNA__080__A _117_/A vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_5.INVTX1_3_.scs8hd_inv_1 chany_top_in[6] mux_right_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_53_21 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_ipin_6.LATCH_0_.latch_SLEEPB _134_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_111 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__149__B _147_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__165__A _164_/X vgnd vpwr scs8hd_diode_2
XANTENNA__075__A _166_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_79 vgnd vpwr scs8hd_decap_3
XFILLER_48_32 vpwr vgnd scs8hd_fill_2
XFILLER_2_125 vgnd vpwr scs8hd_decap_12
XFILLER_48_87 vgnd vpwr scs8hd_decap_4
XFILLER_64_75 vgnd vpwr scs8hd_decap_12
XFILLER_9_15 vgnd vpwr scs8hd_decap_4
X_187_ chany_top_in[1] chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_13_90 vpwr vgnd scs8hd_fill_2
XANTENNA__135__D _101_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_5.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_0.LATCH_4_.latch data_in mem_left_ipin_0.LATCH_4_.latch/Q _159_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_55_143 vgnd vpwr scs8hd_decap_3
XFILLER_55_121 vgnd vpwr scs8hd_fill_1
XFILLER_34_23 vpwr vgnd scs8hd_fill_2
X_110_ _118_/A address[3] _118_/C _111_/A vgnd vpwr scs8hd_or3_4
XFILLER_34_45 vpwr vgnd scs8hd_fill_2
XFILLER_50_55 vgnd vpwr scs8hd_decap_6
XFILLER_59_53 vpwr vgnd scs8hd_fill_2
XFILLER_61_135 vgnd vpwr scs8hd_decap_8
XFILLER_61_113 vgnd vpwr scs8hd_decap_8
XFILLER_46_110 vpwr vgnd scs8hd_fill_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_143 vgnd vpwr scs8hd_decap_3
XFILLER_52_113 vgnd vpwr scs8hd_decap_12
XFILLER_52_102 vpwr vgnd scs8hd_fill_2
XANTENNA__072__B _069_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_1.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_69 vgnd vpwr scs8hd_decap_6
XFILLER_29_12 vpwr vgnd scs8hd_fill_2
XFILLER_29_78 vgnd vpwr scs8hd_decap_3
XFILLER_45_55 vpwr vgnd scs8hd_fill_2
XFILLER_43_135 vgnd vpwr scs8hd_decap_8
XFILLER_61_65 vpwr vgnd scs8hd_fill_2
XFILLER_6_38 vpwr vgnd scs8hd_fill_2
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_ipin_4.LATCH_1_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_121 vgnd vpwr scs8hd_fill_1
XFILLER_19_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_5.INVTX1_5_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA__157__B _147_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_102 vgnd vpwr scs8hd_decap_12
XFILLER_25_102 vpwr vgnd scs8hd_fill_2
XFILLER_25_113 vpwr vgnd scs8hd_fill_2
XANTENNA__083__A _083_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
XFILLER_15_36 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_6.LATCH_2_.latch data_in mem_right_ipin_6.LATCH_2_.latch/Q _132_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_56_32 vgnd vpwr scs8hd_decap_6
XFILLER_56_98 vgnd vpwr scs8hd_decap_12
XFILLER_56_76 vgnd vpwr scs8hd_decap_4
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_102 vpwr vgnd scs8hd_fill_2
XFILLER_31_105 vgnd vpwr scs8hd_decap_12
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__168__A _167_/X vgnd vpwr scs8hd_diode_2
XANTENNA__078__A _088_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_46 vpwr vgnd scs8hd_fill_2
XFILLER_42_23 vpwr vgnd scs8hd_fill_2
XANTENNA__154__C _154_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_15 vgnd vpwr scs8hd_decap_4
XANTENNA__080__B _069_/X vgnd vpwr scs8hd_diode_2
XFILLER_53_66 vpwr vgnd scs8hd_fill_2
XFILLER_53_33 vpwr vgnd scs8hd_fill_2
XFILLER_5_123 vgnd vpwr scs8hd_decap_12
Xmem_left_ipin_1.LATCH_0_.latch data_in _146_/A _144_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _177_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_ipin_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__149__C _143_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_3.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__181__A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_2.LATCH_2_.latch_SLEEPB _096_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_82 vgnd vpwr scs8hd_decap_8
XFILLER_23_14 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_58 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__091__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_48_66 vpwr vgnd scs8hd_fill_2
XFILLER_2_137 vgnd vpwr scs8hd_decap_8
XFILLER_64_87 vgnd vpwr scs8hd_decap_6
XFILLER_64_32 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_ipin_4.LATCH_0_.latch/Q mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_38 vpwr vgnd scs8hd_fill_2
X_186_ chany_top_in[2] chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
Xmux_right_ipin_3.INVTX1_3_.scs8hd_inv_1 chany_top_in[4] mux_right_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_6 vpwr vgnd scs8hd_fill_2
XANTENNA__086__A _086_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_68 vpwr vgnd scs8hd_fill_2
XFILLER_1_3 vgnd vpwr scs8hd_decap_12
XFILLER_59_76 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_3.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
X_169_ _156_/B _169_/B _169_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_52_125 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_7.INVTX1_3_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_46 vpwr vgnd scs8hd_fill_2
XFILLER_29_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_89 vpwr vgnd scs8hd_fill_2
XFILLER_45_34 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_7.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_114 vgnd vpwr scs8hd_decap_12
XANTENNA__157__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_40_117 vgnd vpwr scs8hd_decap_12
XFILLER_31_36 vpwr vgnd scs8hd_fill_2
XFILLER_31_58 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_0.LATCH_3_.latch_SLEEPB _074_/Y vgnd vpwr scs8hd_diode_2
XFILLER_56_55 vgnd vpwr scs8hd_decap_3
XPHY_120 vgnd vpwr scs8hd_decap_3
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_117 vgnd vpwr scs8hd_decap_4
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_22_106 vgnd vpwr scs8hd_decap_12
XANTENNA__184__A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__078__B _069_/X vgnd vpwr scs8hd_diode_2
XANTENNA__094__A _085_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_29 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ _146_/A mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__089__A _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_35 vgnd vpwr scs8hd_decap_4
XFILLER_37_57 vpwr vgnd scs8hd_fill_2
XFILLER_37_79 vpwr vgnd scs8hd_fill_2
XFILLER_53_89 vgnd vpwr scs8hd_decap_4
XFILLER_53_56 vgnd vpwr scs8hd_decap_4
XFILLER_5_135 vgnd vpwr scs8hd_decap_8
XFILLER_64_3 vgnd vpwr scs8hd_decap_12
XFILLER_4_61 vpwr vgnd scs8hd_fill_2
XFILLER_23_37 vpwr vgnd scs8hd_fill_2
XANTENNA__091__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_48_23 vgnd vpwr scs8hd_decap_8
XFILLER_64_44 vgnd vpwr scs8hd_decap_12
X_185_ chany_top_in[3] chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_13_81 vpwr vgnd scs8hd_fill_2
XFILLER_64_145 vgnd vpwr scs8hd_fill_1
XANTENNA__192__A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_5.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_55_123 vgnd vpwr scs8hd_decap_12
XANTENNA__086__B _084_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_6.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_ipin_7.LATCH_3_.latch/Q mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
X_168_ _167_/X _169_/B vgnd vpwr scs8hd_buf_1
XFILLER_24_80 vgnd vpwr scs8hd_decap_3
XFILLER_27_3 vgnd vpwr scs8hd_decap_4
X_099_ _091_/A address[6] _099_/C _118_/C vgnd vpwr scs8hd_or3_4
XFILLER_52_137 vgnd vpwr scs8hd_decap_8
XANTENNA__187__A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_37_123 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_1.INVTX1_3_.scs8hd_inv_1 chany_top_in[3] mux_right_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_ipin_1.LATCH_0_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_7.LATCH_2_.latch_SLEEPB _140_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_16 vpwr vgnd scs8hd_fill_2
XFILLER_20_27 vgnd vpwr scs8hd_decap_4
XFILLER_20_38 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_2_ vgnd vpwr scs8hd_inv_1
XFILLER_28_145 vgnd vpwr scs8hd_fill_1
XANTENNA__097__A _088_/A vgnd vpwr scs8hd_diode_2
XFILLER_43_104 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_9 vgnd vpwr scs8hd_fill_1
XFILLER_19_123 vgnd vpwr scs8hd_decap_12
XFILLER_34_126 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_129 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_7.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_right_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_121 vgnd vpwr scs8hd_decap_3
XPHY_110 vgnd vpwr scs8hd_decap_3
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_92 vgnd vpwr scs8hd_fill_1
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_22_118 vgnd vpwr scs8hd_decap_12
XFILLER_7_72 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_ipin_3.LATCH_0_.latch/Q mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__094__B _093_/B vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_2.LATCH_2_.latch data_in mem_right_ipin_2.LATCH_2_.latch/Q _096_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_144 vpwr vgnd scs8hd_fill_2
XFILLER_32_80 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__195__A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__089__B _084_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_14 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_5.LATCH_3_.latch_SLEEPB _122_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_4.LATCH_5_.latch data_in mem_right_ipin_4.LATCH_5_.latch/Q _112_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _178_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_57_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_106 vgnd vpwr scs8hd_decap_4
XANTENNA__091__C _154_/C vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_ipin_7.LATCH_1_.latch/Q mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_64_56 vgnd vpwr scs8hd_decap_6
X_184_ chany_top_in[4] chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_3.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_27 vgnd vpwr scs8hd_decap_4
XFILLER_55_135 vgnd vpwr scs8hd_decap_8
XFILLER_59_89 vgnd vpwr scs8hd_decap_4
XFILLER_46_102 vgnd vpwr scs8hd_decap_8
X_098_ _117_/A _093_/B _098_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_40_91 vgnd vpwr scs8hd_fill_1
XFILLER_40_80 vgnd vpwr scs8hd_fill_1
X_167_ address[1] address[2] _143_/C _167_/X vgnd vpwr scs8hd_or3_4
XFILLER_1_74 vgnd vpwr scs8hd_fill_1
XFILLER_37_135 vgnd vpwr scs8hd_decap_8
XANTENNA__097__B _093_/B vgnd vpwr scs8hd_diode_2
XFILLER_28_102 vpwr vgnd scs8hd_fill_2
XFILLER_28_113 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_92 vgnd vpwr scs8hd_fill_1
XFILLER_19_135 vgnd vpwr scs8hd_decap_8
XFILLER_34_138 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_ipin_3.LATCH_4_.latch_SLEEPB _105_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_0_.latch/Q mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_16 vgnd vpwr scs8hd_decap_4
XFILLER_31_49 vpwr vgnd scs8hd_fill_2
XPHY_100 vgnd vpwr scs8hd_decap_3
XPHY_122 vgnd vpwr scs8hd_decap_3
XPHY_111 vgnd vpwr scs8hd_decap_3
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_71 vpwr vgnd scs8hd_fill_2
XFILLER_11_7 vpwr vgnd scs8hd_fill_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_30_130 vgnd vpwr scs8hd_decap_12
XFILLER_7_84 vgnd vpwr scs8hd_fill_1
XFILLER_7_62 vgnd vpwr scs8hd_fill_1
XFILLER_7_51 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_5.LATCH_1_.latch data_in mem_right_ipin_5.LATCH_1_.latch/Q _124_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
XFILLER_42_37 vgnd vpwr scs8hd_fill_1
XFILLER_13_108 vpwr vgnd scs8hd_fill_2
XFILLER_16_82 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_5.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[2] mux_right_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_5.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_7.LATCH_4_.latch data_in mem_right_ipin_7.LATCH_4_.latch/Q _138_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_ipin_6.LATCH_3_.latch/Q mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_43_91 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_6.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[8] mux_right_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_right_ipin_1.LATCH_5_.latch_SLEEPB _084_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_47 vpwr vgnd scs8hd_fill_2
XFILLER_48_36 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _171_/HI _145_/Y mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_19 vgnd vpwr scs8hd_fill_1
X_183_ chany_top_in[5] chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_49_111 vgnd vpwr scs8hd_decap_8
XFILLER_64_125 vgnd vpwr scs8hd_decap_12
XFILLER_18_39 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_34_27 vpwr vgnd scs8hd_fill_2
XFILLER_34_49 vgnd vpwr scs8hd_decap_6
XFILLER_50_15 vgnd vpwr scs8hd_decap_12
XFILLER_59_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_097_ _088_/A _093_/B _097_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_ipin_4.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
X_166_ _156_/B _166_/B _166_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_ipin_2.LATCH_0_.latch/Q mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_53 vpwr vgnd scs8hd_fill_2
XFILLER_34_6 vpwr vgnd scs8hd_fill_2
XFILLER_37_103 vpwr vgnd scs8hd_fill_2
XFILLER_52_106 vgnd vpwr scs8hd_decap_4
XFILLER_29_16 vpwr vgnd scs8hd_fill_2
XFILLER_45_59 vpwr vgnd scs8hd_fill_2
XFILLER_45_15 vgnd vpwr scs8hd_decap_8
XFILLER_28_125 vgnd vpwr scs8hd_decap_12
XFILLER_61_69 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_84 vgnd vpwr scs8hd_decap_3
XFILLER_19_71 vpwr vgnd scs8hd_fill_2
XFILLER_19_103 vgnd vpwr scs8hd_decap_12
X_149_ address[1] _147_/Y _143_/C _149_/X vgnd vpwr scs8hd_or3_4
XFILLER_25_117 vpwr vgnd scs8hd_fill_2
XPHY_123 vgnd vpwr scs8hd_decap_3
XPHY_112 vgnd vpwr scs8hd_decap_3
XPHY_101 vgnd vpwr scs8hd_decap_3
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_106 vgnd vpwr scs8hd_decap_4
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_30_142 vgnd vpwr scs8hd_decap_4
XFILLER_7_96 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_3.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_ipin_6.LATCH_1_.latch/Q mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_ipin_4.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_42_49 vpwr vgnd scs8hd_fill_2
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_42_16 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_ipin_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_8_102 vpwr vgnd scs8hd_fill_2
XFILLER_8_124 vgnd vpwr scs8hd_decap_12
XFILLER_8_113 vgnd vpwr scs8hd_decap_8
XFILLER_12_19 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_37 vpwr vgnd scs8hd_fill_2
XFILLER_53_15 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _179_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_3.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_right_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_40 vpwr vgnd scs8hd_fill_2
XFILLER_13_51 vpwr vgnd scs8hd_fill_2
X_182_ chany_top_in[6] chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_13_62 vpwr vgnd scs8hd_fill_2
XFILLER_13_73 vpwr vgnd scs8hd_fill_2
XFILLER_49_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_1_130 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_137 vgnd vpwr scs8hd_decap_8
XANTENNA__100__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_62_3 vgnd vpwr scs8hd_decap_12
Xmem_right_ipin_0.LATCH_5_.latch data_in mem_right_ipin_0.LATCH_5_.latch/Q _070_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_ipin_4.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[6] mux_right_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_6.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_50_49 vgnd vpwr scs8hd_decap_3
XFILLER_50_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_165_ _164_/X _166_/B vgnd vpwr scs8hd_buf_1
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
X_096_ _115_/A _093_/B _096_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_left_ipin_0.LATCH_3_.latch_SLEEPB _163_/Y vgnd vpwr scs8hd_diode_2
XFILLER_45_38 vpwr vgnd scs8hd_fill_2
XFILLER_28_137 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_ipin_6.LATCH_5_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
XFILLER_61_59 vpwr vgnd scs8hd_fill_2
XFILLER_61_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_115 vgnd vpwr scs8hd_decap_6
XFILLER_35_60 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_ipin_0.LATCH_0_.latch_SLEEPB _080_/Y vgnd vpwr scs8hd_diode_2
X_148_ address[0] _143_/C vgnd vpwr scs8hd_inv_8
X_079_ _064_/B _117_/A vgnd vpwr scs8hd_buf_1
Xmux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_ipin_5.LATCH_3_.latch/Q mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_15_19 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_129 vgnd vpwr scs8hd_decap_12
XFILLER_56_15 vgnd vpwr scs8hd_decap_12
XPHY_124 vgnd vpwr scs8hd_decap_3
XPHY_113 vgnd vpwr scs8hd_decap_3
XPHY_102 vgnd vpwr scs8hd_decap_3
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_95 vgnd vpwr scs8hd_fill_1
XFILLER_46_81 vpwr vgnd scs8hd_fill_2
XFILLER_62_80 vgnd vpwr scs8hd_decap_12
XPHY_4 vgnd vpwr scs8hd_decap_3
Xmux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_left_ipin_0.LATCH_4_.latch/Q mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_21_121 vgnd vpwr scs8hd_fill_1
XFILLER_21_143 vgnd vpwr scs8hd_decap_3
XFILLER_8_136 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__103__A _102_/X vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_1.LATCH_1_.latch data_in mem_right_ipin_1.LATCH_1_.latch/Q _088_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_ipin_1.LATCH_0_.latch/Q mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_83 vpwr vgnd scs8hd_fill_2
XFILLER_43_60 vgnd vpwr scs8hd_fill_1
XFILLER_4_65 vpwr vgnd scs8hd_fill_2
XFILLER_4_32 vgnd vpwr scs8hd_decap_3
XFILLER_58_102 vgnd vpwr scs8hd_decap_12
XFILLER_64_15 vgnd vpwr scs8hd_decap_12
Xmem_right_ipin_3.LATCH_4_.latch data_in mem_right_ipin_3.LATCH_4_.latch/Q _105_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_181_ chany_top_in[7] chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_1_142 vgnd vpwr scs8hd_decap_4
XFILLER_49_135 vgnd vpwr scs8hd_decap_8
XANTENNA__100__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_38_71 vpwr vgnd scs8hd_fill_2
XFILLER_54_81 vgnd vpwr scs8hd_decap_8
XFILLER_54_70 vpwr vgnd scs8hd_fill_2
XFILLER_55_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_6.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_105 vgnd vpwr scs8hd_decap_12
XFILLER_59_15 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_1.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[2] mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_46_116 vgnd vpwr scs8hd_decap_12
X_095_ _086_/A _093_/B _095_/Y vgnd vpwr scs8hd_nor2_4
X_164_ _161_/A address[2] address[0] _164_/X vgnd vpwr scs8hd_or3_4
Xmux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_8_ vgnd vpwr scs8hd_inv_1
XFILLER_40_83 vgnd vpwr scs8hd_decap_8
XFILLER_49_92 vgnd vpwr scs8hd_fill_1
XANTENNA__111__A _111_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_66 vpwr vgnd scs8hd_fill_2
XFILLER_1_88 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_ipin_5.LATCH_1_.latch/Q mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_108 vpwr vgnd scs8hd_fill_2
XFILLER_61_27 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_2.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[8] mux_right_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_95 vgnd vpwr scs8hd_fill_1
XFILLER_35_83 vpwr vgnd scs8hd_fill_2
XFILLER_35_94 vpwr vgnd scs8hd_fill_2
XFILLER_51_60 vgnd vpwr scs8hd_fill_1
X_078_ _088_/A _069_/X _078_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__106__A _086_/A vgnd vpwr scs8hd_diode_2
X_147_ address[2] _147_/Y vgnd vpwr scs8hd_inv_8
XFILLER_18_3 vgnd vpwr scs8hd_decap_3
Xmux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_2_.latch/Q mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_56_27 vgnd vpwr scs8hd_decap_4
XFILLER_16_119 vgnd vpwr scs8hd_decap_12
XPHY_125 vgnd vpwr scs8hd_decap_3
XPHY_114 vgnd vpwr scs8hd_decap_3
XPHY_103 vgnd vpwr scs8hd_decap_3
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_left_ipin_0.LATCH_5_.latch data_in mem_left_ipin_0.LATCH_5_.latch/Q _156_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_5.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_52 vgnd vpwr scs8hd_decap_3
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_7_76 vpwr vgnd scs8hd_fill_2
XFILLER_16_41 vgnd vpwr scs8hd_decap_3
XFILLER_16_63 vgnd vpwr scs8hd_fill_1
XFILLER_16_85 vgnd vpwr scs8hd_decap_4
XFILLER_32_84 vgnd vpwr scs8hd_decap_8
XFILLER_57_92 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_4.LATCH_0_.latch data_in mem_right_ipin_4.LATCH_0_.latch/Q _117_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_5.LATCH_0_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_ipin_7.LATCH_0_.latch/Q mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_40 vpwr vgnd scs8hd_fill_2
XFILLER_27_62 vgnd vpwr scs8hd_decap_4
XANTENNA__114__A _086_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_44 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_6.LATCH_3_.latch data_in mem_right_ipin_6.LATCH_3_.latch/Q _131_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_58_114 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_27 vgnd vpwr scs8hd_decap_4
X_180_ chany_top_in[8] chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_13_86 vpwr vgnd scs8hd_fill_2
XFILLER_13_97 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_right_ipin_4.LATCH_3_.latch/Q mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_1_121 vgnd vpwr scs8hd_fill_1
XFILLER_64_106 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__109__A _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_55_117 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_1.INVTX1_5_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_59_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_7.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_128 vgnd vpwr scs8hd_decap_12
XFILLER_24_52 vgnd vpwr scs8hd_decap_4
XFILLER_24_85 vpwr vgnd scs8hd_fill_2
X_094_ _085_/A _093_/B _094_/Y vgnd vpwr scs8hd_nor2_4
X_163_ _156_/B _131_/A _163_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_49_71 vpwr vgnd scs8hd_fill_2
XFILLER_1_34 vpwr vgnd scs8hd_fill_2
Xmem_left_ipin_1.LATCH_1_.latch data_in _145_/A _143_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_ipin_3.LATCH_1_.latch_SLEEPB _108_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_106 vgnd vpwr scs8hd_decap_4
XFILLER_61_39 vgnd vpwr scs8hd_decap_12
XFILLER_10_54 vpwr vgnd scs8hd_fill_2
XFILLER_10_65 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_52 vpwr vgnd scs8hd_fill_2
XFILLER_35_62 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__106__B _109_/B vgnd vpwr scs8hd_diode_2
X_077_ _169_/B _088_/A vgnd vpwr scs8hd_buf_1
X_146_ _146_/A _146_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__122__A _086_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_6 vpwr vgnd scs8hd_fill_2
XFILLER_25_109 vpwr vgnd scs8hd_fill_2
XFILLER_33_120 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_0_.latch/Q mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_126 vgnd vpwr scs8hd_decap_3
XPHY_115 vgnd vpwr scs8hd_decap_3
XPHY_104 vgnd vpwr scs8hd_decap_3
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_31 vpwr vgnd scs8hd_fill_2
XFILLER_21_75 vpwr vgnd scs8hd_fill_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_62_93 vgnd vpwr scs8hd_decap_12
XANTENNA__117__A _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_55 vgnd vpwr scs8hd_decap_4
XFILLER_7_33 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_0.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[6] mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_129_ _129_/A _129_/B _129_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_5.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_123 vgnd vpwr scs8hd_decap_12
XFILLER_12_145 vgnd vpwr scs8hd_fill_1
XFILLER_32_52 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_6.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_right_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_119 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_1.LATCH_2_.latch_SLEEPB _087_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_ipin_4.LATCH_1_.latch/Q mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_30 vgnd vpwr scs8hd_fill_1
XFILLER_43_73 vgnd vpwr scs8hd_fill_1
XFILLER_43_51 vgnd vpwr scs8hd_decap_3
Xmux_left_ipin_0.INVTX1_3_.scs8hd_inv_1 chany_top_in[4] mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_96 vpwr vgnd scs8hd_fill_2
XANTENNA__114__B _112_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_130 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_78 vpwr vgnd scs8hd_fill_2
XANTENNA__130__A _159_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_7.INVTX1_5_.scs8hd_inv_1 chany_top_in[8] mux_right_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_58_126 vgnd vpwr scs8hd_decap_12
XFILLER_8_3 vgnd vpwr scs8hd_decap_12
XFILLER_64_118 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_ipin_3.INVTX1_3_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_38_84 vpwr vgnd scs8hd_fill_2
XANTENNA__109__B _109_/B vgnd vpwr scs8hd_diode_2
XANTENNA__125__A _117_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_59_39 vgnd vpwr scs8hd_decap_8
X_162_ _162_/A _131_/A vgnd vpwr scs8hd_buf_1
XFILLER_24_64 vpwr vgnd scs8hd_fill_2
X_093_ _084_/A _093_/B _093_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_40_52 vpwr vgnd scs8hd_fill_2
XFILLER_27_9 vpwr vgnd scs8hd_fill_2
XFILLER_37_107 vgnd vpwr scs8hd_decap_12
XFILLER_60_121 vgnd vpwr scs8hd_decap_12
XFILLER_1_57 vpwr vgnd scs8hd_fill_2
XFILLER_60_3 vgnd vpwr scs8hd_decap_12
XFILLER_51_143 vgnd vpwr scs8hd_decap_3
XFILLER_51_110 vpwr vgnd scs8hd_fill_2
XFILLER_19_20 vpwr vgnd scs8hd_fill_2
XFILLER_19_31 vpwr vgnd scs8hd_fill_2
XFILLER_19_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_30 vgnd vpwr scs8hd_decap_3
XFILLER_35_52 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_5.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_51_95 vpwr vgnd scs8hd_fill_2
X_145_ _145_/A _145_/Y vgnd vpwr scs8hd_inv_8
X_076_ _115_/A _069_/X _076_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_right_ipin_6.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__122__B _125_/B vgnd vpwr scs8hd_diode_2
XFILLER_33_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_ipin_6.LATCH_0_.latch/Q mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_116 vgnd vpwr scs8hd_decap_3
XPHY_105 vgnd vpwr scs8hd_decap_3
XPHY_127 vgnd vpwr scs8hd_decap_3
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_143 vgnd vpwr scs8hd_decap_3
XFILLER_30_102 vpwr vgnd scs8hd_fill_2
XANTENNA__117__B _112_/B vgnd vpwr scs8hd_diode_2
XANTENNA__133__A _169_/B vgnd vpwr scs8hd_diode_2
X_128_ _127_/X _129_/B vgnd vpwr scs8hd_buf_1
XFILLER_21_135 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_ipin_3.LATCH_3_.latch/Q mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ _146_/Y mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_12_102 vgnd vpwr scs8hd_decap_8
XFILLER_12_113 vgnd vpwr scs8hd_decap_12
XFILLER_8_106 vgnd vpwr scs8hd_decap_4
XFILLER_32_64 vpwr vgnd scs8hd_fill_2
XANTENNA__128__A _127_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_4_142 vgnd vpwr scs8hd_decap_4
XANTENNA__130__B _129_/B vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ right_grid_pin_3_ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_19 vgnd vpwr scs8hd_fill_1
Xmem_right_ipin_0.LATCH_0_.latch data_in mem_right_ipin_0.LATCH_0_.latch/Q _080_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_5.INVTX1_1_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_58_138 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_4.INVTX1_1_.scs8hd_inv_1 chany_top_in[1] mux_right_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_44 vpwr vgnd scs8hd_fill_2
XFILLER_13_55 vgnd vpwr scs8hd_decap_4
XFILLER_13_77 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_ipin_7.LATCH_4_.latch/Q mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA__125__B _125_/B vgnd vpwr scs8hd_diode_2
XANTENNA__141__A _169_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_2.LATCH_3_.latch data_in mem_right_ipin_2.LATCH_3_.latch/Q _095_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_161_ _161_/A address[2] _143_/C _162_/A vgnd vpwr scs8hd_or3_4
XANTENNA_mem_left_ipin_0.LATCH_0_.latch_SLEEPB _064_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_32 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_5.INVTX1_5_.scs8hd_inv_1 chany_top_in[7] mux_right_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_092_ _091_/X _093_/B vgnd vpwr scs8hd_buf_1
XFILLER_40_64 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_6.LATCH_2_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
XFILLER_49_95 vpwr vgnd scs8hd_fill_2
XFILLER_37_119 vgnd vpwr scs8hd_decap_3
XFILLER_60_133 vgnd vpwr scs8hd_decap_12
XFILLER_53_3 vgnd vpwr scs8hd_decap_12
XANTENNA__136__A _135_/X vgnd vpwr scs8hd_diode_2
XFILLER_10_23 vpwr vgnd scs8hd_fill_2
XFILLER_10_89 vgnd vpwr scs8hd_decap_3
XFILLER_27_130 vgnd vpwr scs8hd_decap_4
XFILLER_51_74 vpwr vgnd scs8hd_fill_2
XFILLER_51_52 vpwr vgnd scs8hd_fill_2
X_075_ _166_/B _115_/A vgnd vpwr scs8hd_buf_1
X_144_ _082_/C _101_/X address[0] _144_/Y vgnd vpwr scs8hd_nor3_4
XANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_100 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_ipin_3.LATCH_1_.latch/Q mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_128 vgnd vpwr scs8hd_decap_3
XPHY_117 vgnd vpwr scs8hd_decap_3
XPHY_106 vgnd vpwr scs8hd_decap_3
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_3.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_11 vgnd vpwr scs8hd_decap_4
XFILLER_21_88 vgnd vpwr scs8hd_decap_4
XFILLER_21_99 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_85 vpwr vgnd scs8hd_fill_2
XFILLER_15_100 vpwr vgnd scs8hd_fill_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_7_46 vgnd vpwr scs8hd_decap_3
XANTENNA__133__B _129_/B vgnd vpwr scs8hd_diode_2
X_127_ address[5] _127_/B _154_/C _127_/X vgnd vpwr scs8hd_or3_4
XFILLER_21_103 vgnd vpwr scs8hd_decap_12
XFILLER_12_125 vgnd vpwr scs8hd_decap_12
XFILLER_16_66 vgnd vpwr scs8hd_fill_1
XFILLER_32_10 vpwr vgnd scs8hd_fill_2
XFILLER_32_32 vgnd vpwr scs8hd_decap_4
XFILLER_57_73 vpwr vgnd scs8hd_fill_2
XANTENNA__144__A _082_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_4.LATCH_3_.latch_SLEEPB _114_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_ipin_7.LATCH_2_.latch/Q mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__139__A _131_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_12 vpwr vgnd scs8hd_fill_2
XFILLER_13_23 vpwr vgnd scs8hd_fill_2
XFILLER_1_113 vgnd vpwr scs8hd_decap_8
Xmem_right_ipin_5.LATCH_2_.latch data_in mem_right_ipin_5.LATCH_2_.latch/Q _123_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_54_74 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_ipin_5.LATCH_0_.latch/Q mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__141__B _142_/B vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_14_ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_5.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_32 vgnd vpwr scs8hd_decap_3
Xmem_right_ipin_7.LATCH_5_.latch data_in mem_right_ipin_7.LATCH_5_.latch/Q _137_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_160_ address[1] _161_/A vgnd vpwr scs8hd_inv_8
X_091_ _091_/A address[6] _154_/C _091_/X vgnd vpwr scs8hd_or3_4
XFILLER_40_76 vgnd vpwr scs8hd_decap_4
XFILLER_1_15 vgnd vpwr scs8hd_decap_8
XFILLER_60_145 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_2.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_1_.latch/Q mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__152__A enable vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_right_ipin_2.LATCH_3_.latch/Q mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_46_3 vgnd vpwr scs8hd_decap_12
XFILLER_51_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_2.LATCH_4_.latch_SLEEPB _094_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_35 vpwr vgnd scs8hd_fill_2
XANTENNA__062__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_19_88 vgnd vpwr scs8hd_decap_4
XFILLER_19_99 vpwr vgnd scs8hd_fill_2
XFILLER_27_142 vgnd vpwr scs8hd_decap_4
XFILLER_42_145 vgnd vpwr scs8hd_fill_1
XFILLER_35_87 vgnd vpwr scs8hd_decap_4
XFILLER_35_98 vpwr vgnd scs8hd_fill_2
XFILLER_51_31 vpwr vgnd scs8hd_fill_2
X_074_ _086_/A _069_/X _074_/Y vgnd vpwr scs8hd_nor2_4
X_143_ _082_/C _101_/X _143_/C _143_/Y vgnd vpwr scs8hd_nor3_4
Xmem_left_ipin_0.LATCH_0_.latch data_in mem_left_ipin_0.LATCH_0_.latch/Q _064_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_3.INVTX1_5_.scs8hd_inv_1 chany_top_in[5] mux_right_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_33_123 vgnd vpwr scs8hd_decap_12
XANTENNA__147__A address[2] vgnd vpwr scs8hd_diode_2
XPHY_129 vgnd vpwr scs8hd_decap_3
XPHY_118 vgnd vpwr scs8hd_decap_3
XPHY_107 vgnd vpwr scs8hd_decap_3
XFILLER_46_53 vgnd vpwr scs8hd_decap_4
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_112 vpwr vgnd scs8hd_fill_2
XFILLER_15_123 vgnd vpwr scs8hd_decap_12
X_126_ address[6] _127_/B vgnd vpwr scs8hd_inv_8
XFILLER_30_6 vpwr vgnd scs8hd_fill_2
XFILLER_21_115 vgnd vpwr scs8hd_decap_6
Xmux_right_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_ipin_6.LATCH_4_.latch/Q mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_16_23 vgnd vpwr scs8hd_decap_4
XFILLER_12_137 vgnd vpwr scs8hd_decap_8
XFILLER_16_78 vgnd vpwr scs8hd_decap_4
XFILLER_16_89 vgnd vpwr scs8hd_fill_1
XFILLER_57_96 vpwr vgnd scs8hd_fill_2
XANTENNA__144__B _101_/X vgnd vpwr scs8hd_diode_2
X_109_ _117_/A _109_/B _109_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__160__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_7.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__070__A _084_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_22 vpwr vgnd scs8hd_fill_2
XFILLER_43_87 vpwr vgnd scs8hd_fill_2
XFILLER_43_65 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_0.LATCH_5_.latch_SLEEPB _070_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_48 vgnd vpwr scs8hd_decap_4
XFILLER_4_15 vgnd vpwr scs8hd_decap_12
XANTENNA__139__B _142_/B vgnd vpwr scs8hd_diode_2
XANTENNA__155__A _154_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _171_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__065__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_38_32 vgnd vpwr scs8hd_decap_3
XFILLER_54_53 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.INVTX1_5_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_48_7 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_ipin_2.LATCH_1_.latch/Q mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_143 vgnd vpwr scs8hd_decap_3
XFILLER_63_110 vgnd vpwr scs8hd_decap_12
XFILLER_24_23 vpwr vgnd scs8hd_fill_2
XFILLER_40_44 vpwr vgnd scs8hd_fill_2
XFILLER_24_89 vgnd vpwr scs8hd_decap_3
X_090_ address[5] _091_/A vgnd vpwr scs8hd_inv_8
XFILLER_49_75 vpwr vgnd scs8hd_fill_2
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
XFILLER_45_143 vgnd vpwr scs8hd_decap_3
XFILLER_45_110 vpwr vgnd scs8hd_fill_2
XFILLER_1_38 vpwr vgnd scs8hd_fill_2
XFILLER_51_135 vgnd vpwr scs8hd_decap_8
XFILLER_10_58 vpwr vgnd scs8hd_fill_2
XFILLER_10_69 vgnd vpwr scs8hd_decap_4
XANTENNA__062__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_42_102 vpwr vgnd scs8hd_fill_2
XFILLER_19_56 vgnd vpwr scs8hd_decap_3
XFILLER_27_121 vgnd vpwr scs8hd_fill_1
XFILLER_42_113 vgnd vpwr scs8hd_decap_12
X_142_ _064_/B _142_/B _142_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_51_65 vpwr vgnd scs8hd_fill_2
X_073_ _131_/A _086_/A vgnd vpwr scs8hd_buf_1
XFILLER_18_8 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_135 vgnd vpwr scs8hd_decap_8
XANTENNA__163__A _156_/B vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_ipin_6.LATCH_2_.latch/Q mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_ipin_0.INVTX1_1_.scs8hd_inv_1 chany_top_in[1] mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_102 vgnd vpwr scs8hd_decap_8
XPHY_119 vgnd vpwr scs8hd_decap_3
XPHY_108 vgnd vpwr scs8hd_decap_3
XFILLER_24_113 vgnd vpwr scs8hd_decap_8
XFILLER_24_124 vgnd vpwr scs8hd_decap_12
XANTENNA__073__A _131_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_35 vpwr vgnd scs8hd_fill_2
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
XFILLER_46_76 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_32 vpwr vgnd scs8hd_fill_2
XFILLER_15_135 vgnd vpwr scs8hd_decap_8
X_125_ _117_/A _125_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__158__A _157_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_1.INVTX1_5_.scs8hd_inv_1 chany_top_in[7] mux_right_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_right_ipin_7.LATCH_4_.latch_SLEEPB _138_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_46 vpwr vgnd scs8hd_fill_2
XANTENNA__068__A _118_/A vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_ipin_4.LATCH_0_.latch/Q mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_ipin_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_32_23 vpwr vgnd scs8hd_fill_2
XFILLER_57_53 vpwr vgnd scs8hd_fill_2
X_108_ _088_/A _109_/B _108_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__144__C address[0] vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__070__B _069_/X vgnd vpwr scs8hd_diode_2
XFILLER_43_22 vgnd vpwr scs8hd_decap_3
XFILLER_43_11 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_7.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[4] mux_right_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_right_ipin_1.LATCH_3_.latch/Q mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_2.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_6.INVTX1_3_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_49_119 vgnd vpwr scs8hd_decap_3
XFILLER_1_126 vpwr vgnd scs8hd_fill_2
XANTENNA__081__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_54_32 vgnd vpwr scs8hd_decap_8
XFILLER_38_88 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_6.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__166__A _156_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_7.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_92 vgnd vpwr scs8hd_fill_1
XANTENNA__076__A _115_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_68 vgnd vpwr scs8hd_fill_1
XFILLER_40_12 vgnd vpwr scs8hd_decap_8
XFILLER_40_23 vpwr vgnd scs8hd_fill_2
XFILLER_49_54 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_ipin_5.LATCH_5_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_1.LATCH_2_.latch data_in mem_right_ipin_1.LATCH_2_.latch/Q _087_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_ipin_5.LATCH_4_.latch/Q mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_51_114 vgnd vpwr scs8hd_decap_8
XFILLER_10_15 vgnd vpwr scs8hd_decap_4
XANTENNA__062__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_19_13 vpwr vgnd scs8hd_fill_2
XFILLER_19_24 vpwr vgnd scs8hd_fill_2
XFILLER_19_35 vpwr vgnd scs8hd_fill_2
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
XFILLER_27_100 vpwr vgnd scs8hd_fill_2
XFILLER_35_56 vpwr vgnd scs8hd_fill_2
X_141_ _169_/B _142_/B _141_/Y vgnd vpwr scs8hd_nor2_4
X_072_ _085_/A _069_/X _072_/Y vgnd vpwr scs8hd_nor2_4
Xmem_right_ipin_3.LATCH_5_.latch data_in mem_right_ipin_3.LATCH_5_.latch/Q _104_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__163__B _131_/A vgnd vpwr scs8hd_diode_2
XFILLER_51_3 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _170_/HI mem_left_ipin_0.LATCH_5_.latch/Q
+ mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XPHY_109 vgnd vpwr scs8hd_decap_3
XFILLER_24_136 vgnd vpwr scs8hd_decap_8
XFILLER_62_32 vgnd vpwr scs8hd_decap_12
XFILLER_30_106 vgnd vpwr scs8hd_decap_12
XFILLER_7_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
X_124_ _088_/A _125_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_16_6 vgnd vpwr scs8hd_decap_6
XANTENNA__068__B address[3] vgnd vpwr scs8hd_diode_2
XANTENNA__084__A _084_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_68 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_ipin_1.LATCH_1_.latch/Q mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_107_ _115_/A _109_/B _107_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_3 vpwr vgnd scs8hd_fill_2
XANTENNA__169__A _156_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_8_70 vgnd vpwr scs8hd_fill_1
XANTENNA__079__A _064_/B vgnd vpwr scs8hd_diode_2
XFILLER_27_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_56 vpwr vgnd scs8hd_fill_2
XFILLER_43_34 vpwr vgnd scs8hd_fill_2
XFILLER_27_79 vpwr vgnd scs8hd_fill_2
XFILLER_4_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_5.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_0_ vgnd vpwr scs8hd_inv_1
XFILLER_57_120 vpwr vgnd scs8hd_fill_2
XFILLER_1_105 vpwr vgnd scs8hd_fill_2
XFILLER_38_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_67 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_ipin_5.LATCH_2_.latch/Q mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_ipin_5.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[6] mux_right_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_63_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__166__B _166_/B vgnd vpwr scs8hd_diode_2
XANTENNA__182__A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_5_71 vpwr vgnd scs8hd_fill_2
XFILLER_54_145 vgnd vpwr scs8hd_fill_1
Xmem_right_ipin_4.LATCH_1_.latch data_in mem_right_ipin_4.LATCH_1_.latch/Q _116_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_142 vgnd vpwr scs8hd_decap_4
XFILLER_39_131 vgnd vpwr scs8hd_decap_3
XANTENNA__076__B _069_/X vgnd vpwr scs8hd_diode_2
XANTENNA__092__A _091_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_99 vgnd vpwr scs8hd_decap_12
XFILLER_49_88 vgnd vpwr scs8hd_decap_4
XFILLER_49_44 vgnd vpwr scs8hd_decap_8
XFILLER_45_123 vgnd vpwr scs8hd_decap_12
XFILLER_36_145 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_ipin_3.LATCH_0_.latch/Q mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_27 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_6.LATCH_4_.latch data_in mem_right_ipin_6.LATCH_4_.latch/Q _130_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_42_137 vgnd vpwr scs8hd_decap_8
XANTENNA__087__A _115_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_13 vpwr vgnd scs8hd_fill_2
XFILLER_35_35 vgnd vpwr scs8hd_decap_4
XFILLER_35_68 vpwr vgnd scs8hd_fill_2
XFILLER_51_89 vgnd vpwr scs8hd_decap_4
XFILLER_51_56 vgnd vpwr scs8hd_decap_4
X_140_ _166_/B _142_/B _140_/Y vgnd vpwr scs8hd_nor2_4
X_071_ _159_/B _085_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_145 vgnd vpwr scs8hd_fill_1
XPHY_90 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_104 vpwr vgnd scs8hd_fill_2
XFILLER_44_3 vgnd vpwr scs8hd_decap_6
XFILLER_21_15 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_ipin_0.LATCH_3_.latch/Q mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_21_48 vpwr vgnd scs8hd_fill_2
XFILLER_46_23 vpwr vgnd scs8hd_fill_2
XFILLER_62_44 vgnd vpwr scs8hd_decap_12
XFILLER_46_89 vgnd vpwr scs8hd_decap_3
XFILLER_15_104 vgnd vpwr scs8hd_decap_6
XFILLER_30_118 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_123_ _115_/A _125_/B _123_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_7.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__190__A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_4.LATCH_0_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_59 vgnd vpwr scs8hd_decap_4
XANTENNA__068__C _082_/C vgnd vpwr scs8hd_diode_2
XANTENNA__084__B _084_/B vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_ipin_7.LATCH_1_.latch/Q mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_57_77 vpwr vgnd scs8hd_fill_2
XFILLER_7_111 vgnd vpwr scs8hd_decap_8
XFILLER_7_100 vpwr vgnd scs8hd_fill_2
X_106_ _086_/A _109_/B _106_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__169__B _169_/B vgnd vpwr scs8hd_diode_2
XANTENNA__185__A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _146_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_36 vpwr vgnd scs8hd_fill_2
XANTENNA__095__A _086_/A vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_right_ipin_4.LATCH_4_.latch/Q mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_13_16 vpwr vgnd scs8hd_fill_2
XFILLER_13_27 vpwr vgnd scs8hd_fill_2
XFILLER_57_143 vgnd vpwr scs8hd_decap_3
XFILLER_54_89 vgnd vpwr scs8hd_decap_3
XFILLER_54_78 vgnd vpwr scs8hd_fill_1
Xmem_right_ipin_7.LATCH_0_.latch data_in mem_right_ipin_7.LATCH_0_.latch/Q _142_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_5.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_135 vgnd vpwr scs8hd_decap_8
XFILLER_39_121 vgnd vpwr scs8hd_fill_1
XFILLER_54_113 vgnd vpwr scs8hd_decap_12
XFILLER_54_102 vpwr vgnd scs8hd_fill_2
XFILLER_24_48 vpwr vgnd scs8hd_fill_2
XFILLER_24_59 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_2.LATCH_1_.latch_SLEEPB _097_/Y vgnd vpwr scs8hd_diode_2
XFILLER_45_135 vgnd vpwr scs8hd_decap_8
XFILLER_30_91 vgnd vpwr scs8hd_fill_1
XFILLER_39_6 vgnd vpwr scs8hd_decap_3
XFILLER_36_102 vgnd vpwr scs8hd_decap_8
XFILLER_36_113 vgnd vpwr scs8hd_decap_12
XANTENNA__193__A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_39 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_1_.latch/Q mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_ipin_3.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[4] mux_right_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_48 vpwr vgnd scs8hd_fill_2
XFILLER_27_113 vpwr vgnd scs8hd_fill_2
XANTENNA__087__B _084_/B vgnd vpwr scs8hd_diode_2
XFILLER_51_35 vpwr vgnd scs8hd_fill_2
X_070_ _084_/A _069_/X _070_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
XFILLER_18_102 vgnd vpwr scs8hd_decap_8
XFILLER_18_113 vgnd vpwr scs8hd_decap_12
XPHY_91 vgnd vpwr scs8hd_decap_3
XPHY_80 vgnd vpwr scs8hd_decap_3
XFILLER_2_84 vpwr vgnd scs8hd_fill_2
XANTENNA__188__A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_37_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_4.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_68 vgnd vpwr scs8hd_decap_6
XANTENNA__098__A _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_116 vgnd vpwr scs8hd_decap_6
XFILLER_62_56 vgnd vpwr scs8hd_decap_12
XFILLER_11_71 vpwr vgnd scs8hd_fill_2
X_122_ _086_/A _125_/B _122_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_32_48 vpwr vgnd scs8hd_fill_2
XFILLER_32_59 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_ipin_0.LATCH_5_.latch_SLEEPB _156_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_ipin_4.LATCH_2_.latch/Q mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_7.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_145 vgnd vpwr scs8hd_fill_1
XFILLER_7_123 vpwr vgnd scs8hd_fill_2
X_105_ _085_/A _109_/B _105_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_right_ipin_0.LATCH_2_.latch_SLEEPB _076_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_26 vgnd vpwr scs8hd_decap_4
XANTENNA__095__B _093_/B vgnd vpwr scs8hd_diode_2
XFILLER_43_69 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_3.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_92 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_ipin_2.LATCH_0_.latch/Q mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__196__A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.INVTX1_5_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_57_100 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_100 vgnd vpwr scs8hd_decap_12
XFILLER_48_144 vpwr vgnd scs8hd_fill_2
XFILLER_5_95 vpwr vgnd scs8hd_fill_2
XFILLER_54_125 vgnd vpwr scs8hd_decap_12
XFILLER_24_27 vpwr vgnd scs8hd_fill_2
XFILLER_40_59 vgnd vpwr scs8hd_decap_3
XFILLER_40_48 vpwr vgnd scs8hd_fill_2
XFILLER_45_114 vgnd vpwr scs8hd_decap_8
XFILLER_39_90 vgnd vpwr scs8hd_decap_8
XFILLER_51_106 vpwr vgnd scs8hd_fill_2
XFILLER_36_125 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_ipin_6.LATCH_1_.latch/Q mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_106 vgnd vpwr scs8hd_decap_4
XFILLER_51_69 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_3.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_0.LATCH_1_.latch data_in mem_right_ipin_0.LATCH_1_.latch/Q _078_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_ipin_4.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_125 vgnd vpwr scs8hd_decap_12
XPHY_92 vgnd vpwr scs8hd_decap_3
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_63 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_ipin_3.LATCH_4_.latch/Q mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmem_right_ipin_2.LATCH_4_.latch data_in mem_right_ipin_2.LATCH_4_.latch/Q _094_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_46_36 vpwr vgnd scs8hd_fill_2
XANTENNA__098__B _093_/B vgnd vpwr scs8hd_diode_2
XFILLER_62_68 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_1.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[3] mux_right_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_121_ _085_/A _125_/B _121_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_7.LATCH_1_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_27 vpwr vgnd scs8hd_fill_2
XFILLER_32_38 vgnd vpwr scs8hd_fill_1
XFILLER_57_57 vpwr vgnd scs8hd_fill_2
XFILLER_57_35 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
X_104_ _084_/A _109_/B _104_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_21_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_5.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_8_84 vpwr vgnd scs8hd_fill_2
XFILLER_8_62 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _179_/HI mem_right_ipin_7.LATCH_5_.latch/Q
+ mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_left_ipin_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[1] mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_92 vgnd vpwr scs8hd_fill_1
XFILLER_12_3 vgnd vpwr scs8hd_decap_12
XFILLER_57_123 vgnd vpwr scs8hd_decap_12
XFILLER_57_112 vgnd vpwr scs8hd_decap_8
XFILLER_38_37 vpwr vgnd scs8hd_fill_2
XFILLER_38_48 vgnd vpwr scs8hd_decap_8
XFILLER_48_112 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_5.LATCH_2_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
XFILLER_39_123 vgnd vpwr scs8hd_decap_8
XFILLER_39_101 vpwr vgnd scs8hd_fill_2
XFILLER_54_137 vgnd vpwr scs8hd_decap_8
XFILLER_40_27 vpwr vgnd scs8hd_fill_2
XFILLER_49_58 vgnd vpwr scs8hd_fill_1
XFILLER_49_25 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_3.LATCH_0_.latch data_in mem_right_ipin_3.LATCH_0_.latch/Q _109_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_36_137 vgnd vpwr scs8hd_decap_8
XFILLER_10_19 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_ipin_3.LATCH_2_.latch/Q mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_126 vpwr vgnd scs8hd_fill_2
XFILLER_51_48 vpwr vgnd scs8hd_fill_2
XFILLER_51_15 vgnd vpwr scs8hd_decap_12
XPHY_82 vgnd vpwr scs8hd_decap_3
XFILLER_18_137 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XPHY_60 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_93 vgnd vpwr scs8hd_decap_3
X_197_ chany_bottom_in[0] chany_top_out[0] vgnd vpwr scs8hd_buf_2
Xmem_right_ipin_5.LATCH_3_.latch data_in mem_right_ipin_5.LATCH_3_.latch/Q _122_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_15 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_ipin_1.LATCH_0_.latch/Q mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
X_120_ _129_/A _125_/B _120_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_40 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_5.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_8
XFILLER_16_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_3.LATCH_3_.latch_SLEEPB _106_/Y vgnd vpwr scs8hd_diode_2
XFILLER_57_47 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_7.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_11_121 vgnd vpwr scs8hd_fill_1
X_103_ _102_/X _109_/B vgnd vpwr scs8hd_buf_1
XFILLER_11_143 vgnd vpwr scs8hd_decap_3
XFILLER_22_72 vgnd vpwr scs8hd_decap_8
XFILLER_22_83 vpwr vgnd scs8hd_fill_2
XFILLER_47_91 vpwr vgnd scs8hd_fill_2
XFILLER_14_7 vgnd vpwr scs8hd_decap_4
Xmem_left_ipin_0.LATCH_1_.latch data_in mem_left_ipin_0.LATCH_1_.latch/Q _169_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_43_38 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_106 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_6_ vgnd vpwr scs8hd_inv_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_ipin_5.LATCH_1_.latch/Q mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_109 vpwr vgnd scs8hd_fill_2
XFILLER_38_27 vpwr vgnd scs8hd_fill_2
XFILLER_57_135 vgnd vpwr scs8hd_decap_8
XFILLER_54_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_124 vgnd vpwr scs8hd_decap_12
XFILLER_28_82 vgnd vpwr scs8hd_fill_1
XFILLER_60_91 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_right_ipin_2.LATCH_4_.latch/Q mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_2_.latch/Q mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_75 vpwr vgnd scs8hd_fill_2
XFILLER_5_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_6.INVTX1_3_.scs8hd_inv_1 chany_top_in[7] mux_right_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_49_15 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_ipin_1.LATCH_4_.latch_SLEEPB _085_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_7.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_72 vgnd vpwr scs8hd_decap_4
XFILLER_30_83 vgnd vpwr scs8hd_decap_8
Xmux_left_ipin_0.INVTX1_5_.scs8hd_inv_1 chany_top_in[8] mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__101__A _100_/X vgnd vpwr scs8hd_diode_2
XFILLER_27_138 vpwr vgnd scs8hd_fill_2
XFILLER_35_17 vpwr vgnd scs8hd_fill_2
XFILLER_51_27 vpwr vgnd scs8hd_fill_2
XFILLER_50_130 vgnd vpwr scs8hd_decap_12
XPHY_94 vgnd vpwr scs8hd_decap_3
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_50 vgnd vpwr scs8hd_decap_3
XFILLER_25_83 vpwr vgnd scs8hd_fill_2
XPHY_61 vgnd vpwr scs8hd_decap_3
XFILLER_33_108 vgnd vpwr scs8hd_decap_12
XPHY_72 vgnd vpwr scs8hd_decap_3
X_196_ chany_bottom_in[1] chany_top_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_2_32 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _145_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _178_/HI mem_right_ipin_6.LATCH_5_.latch/Q
+ mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_46_49 vpwr vgnd scs8hd_fill_2
XFILLER_46_27 vgnd vpwr scs8hd_decap_4
XFILLER_62_15 vgnd vpwr scs8hd_decap_12
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XFILLER_11_96 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_71 vpwr vgnd scs8hd_fill_2
X_179_ _179_/HI _179_/LO vgnd vpwr scs8hd_conb_1
XFILLER_35_3 vgnd vpwr scs8hd_fill_1
XFILLER_20_100 vgnd vpwr scs8hd_decap_12
XFILLER_20_144 vpwr vgnd scs8hd_fill_2
XFILLER_57_15 vgnd vpwr scs8hd_decap_12
XFILLER_11_100 vpwr vgnd scs8hd_fill_2
XFILLER_11_111 vpwr vgnd scs8hd_fill_2
X_102_ _118_/C _101_/X _102_/X vgnd vpwr scs8hd_or2_4
XANTENNA_mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_43_17 vgnd vpwr scs8hd_decap_3
XFILLER_4_118 vgnd vpwr scs8hd_decap_12
XFILLER_17_62 vpwr vgnd scs8hd_fill_2
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_ipin_2.LATCH_2_.latch/Q mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__104__A _084_/A vgnd vpwr scs8hd_diode_2
XFILLER_58_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_110 vpwr vgnd scs8hd_fill_2
XFILLER_48_136 vgnd vpwr scs8hd_decap_8
XFILLER_0_132 vgnd vpwr scs8hd_decap_12
XFILLER_54_106 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_4.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_0_.latch/Q mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_45_106 vpwr vgnd scs8hd_fill_2
XFILLER_60_109 vgnd vpwr scs8hd_decap_12
XFILLER_14_41 vgnd vpwr scs8hd_decap_3
XFILLER_14_96 vgnd vpwr scs8hd_decap_12
XFILLER_30_51 vpwr vgnd scs8hd_fill_2
XFILLER_27_117 vgnd vpwr scs8hd_decap_4
XFILLER_50_142 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_4.INVTX1_3_.scs8hd_inv_1 chany_top_in[5] mux_right_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_95 vgnd vpwr scs8hd_decap_3
XPHY_84 vgnd vpwr scs8hd_decap_3
XFILLER_41_120 vpwr vgnd scs8hd_fill_2
XPHY_40 vgnd vpwr scs8hd_decap_3
XFILLER_25_62 vgnd vpwr scs8hd_decap_4
XPHY_51 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
X_195_ chany_bottom_in[2] chany_top_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA__112__A _084_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_44 vpwr vgnd scs8hd_fill_2
XFILLER_37_7 vgnd vpwr scs8hd_decap_4
XFILLER_2_88 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_27 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_ipin_4.LATCH_1_.latch/Q mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_53 vpwr vgnd scs8hd_fill_2
XFILLER_11_75 vpwr vgnd scs8hd_fill_2
XFILLER_14_120 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_6.LATCH_4_.latch_SLEEPB _130_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_0.LATCH_2_.latch_SLEEPB _166_/Y vgnd vpwr scs8hd_diode_2
XFILLER_36_50 vgnd vpwr scs8hd_decap_6
XANTENNA__107__A _115_/A vgnd vpwr scs8hd_diode_2
X_178_ _178_/HI _178_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mem_right_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_3 vpwr vgnd scs8hd_fill_2
XFILLER_20_112 vgnd vpwr scs8hd_decap_12
Xmem_right_ipin_1.LATCH_3_.latch data_in mem_right_ipin_1.LATCH_3_.latch/Q _086_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_57_27 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_ipin_1.LATCH_4_.latch/Q mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_7_127 vgnd vpwr scs8hd_decap_12
XFILLER_11_123 vgnd vpwr scs8hd_decap_12
XFILLER_22_41 vgnd vpwr scs8hd_decap_3
X_101_ _100_/X _101_/X vgnd vpwr scs8hd_buf_1
XANTENNA_mux_right_ipin_2.INVTX1_3_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_8_32 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_6.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_96 vpwr vgnd scs8hd_fill_2
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_73 vpwr vgnd scs8hd_fill_2
XFILLER_33_95 vgnd vpwr scs8hd_fill_1
XANTENNA__104__B _109_/B vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _129_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_122 vpwr vgnd scs8hd_fill_2
XFILLER_0_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_4.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_44_50 vgnd vpwr scs8hd_decap_4
XANTENNA__115__A _115_/A vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _177_/HI mem_right_ipin_5.LATCH_5_.latch/Q
+ mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
XFILLER_5_99 vgnd vpwr scs8hd_decap_12
XFILLER_5_88 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_5.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_4.LATCH_5_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_86 vgnd vpwr scs8hd_fill_1
XFILLER_55_71 vpwr vgnd scs8hd_fill_2
XFILLER_58_3 vgnd vpwr scs8hd_decap_12
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_143 vgnd vpwr scs8hd_decap_3
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_74 vgnd vpwr scs8hd_decap_3
XFILLER_41_95 vpwr vgnd scs8hd_fill_2
XFILLER_41_84 vpwr vgnd scs8hd_fill_2
XFILLER_41_73 vpwr vgnd scs8hd_fill_2
XFILLER_41_62 vpwr vgnd scs8hd_fill_2
X_194_ chany_bottom_in[3] chany_top_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA__112__B _112_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_110 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_ipin_1.LATCH_2_.latch/Q mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_4.LATCH_2_.latch data_in mem_right_ipin_4.LATCH_2_.latch/Q _115_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_132 vgnd vpwr scs8hd_decap_12
XFILLER_36_84 vpwr vgnd scs8hd_fill_2
XFILLER_52_72 vgnd vpwr scs8hd_fill_1
XANTENNA__107__B _109_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_177_ _177_/HI _177_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__123__A _115_/A vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_2.INVTX1_3_.scs8hd_inv_1 chany_top_in[4] mux_right_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_4.INVTX1_1_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_20_124 vgnd vpwr scs8hd_decap_12
XFILLER_7_139 vgnd vpwr scs8hd_decap_6
XFILLER_11_135 vgnd vpwr scs8hd_decap_8
X_100_ address[4] _118_/B _100_/X vgnd vpwr scs8hd_or2_4
Xmem_right_ipin_6.LATCH_5_.latch data_in mem_right_ipin_6.LATCH_5_.latch/Q _129_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_47_50 vgnd vpwr scs8hd_decap_4
XANTENNA__118__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_88 vpwr vgnd scs8hd_fill_2
XFILLER_8_66 vgnd vpwr scs8hd_decap_4
XFILLER_40_3 vpwr vgnd scs8hd_fill_2
XFILLER_17_31 vpwr vgnd scs8hd_fill_2
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_53 vpwr vgnd scs8hd_fill_2
XFILLER_17_75 vpwr vgnd scs8hd_fill_2
XFILLER_33_30 vpwr vgnd scs8hd_fill_2
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_58_60 vgnd vpwr scs8hd_decap_3
XANTENNA__120__B _125_/B vgnd vpwr scs8hd_diode_2
XFILLER_38_19 vgnd vpwr scs8hd_fill_1
XFILLER_54_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_7.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_30 vgnd vpwr scs8hd_fill_1
XFILLER_28_63 vpwr vgnd scs8hd_fill_2
XFILLER_28_85 vgnd vpwr scs8hd_decap_4
XFILLER_44_84 vpwr vgnd scs8hd_fill_2
XFILLER_60_83 vgnd vpwr scs8hd_decap_8
XFILLER_60_72 vgnd vpwr scs8hd_decap_4
XANTENNA__115__B _112_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_138 vpwr vgnd scs8hd_fill_2
XFILLER_39_105 vgnd vpwr scs8hd_decap_12
XANTENNA__131__A _131_/A vgnd vpwr scs8hd_diode_2
XFILLER_62_141 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_ipin_3.LATCH_1_.latch/Q mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_49_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _146_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_39_73 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__126__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_ipin_0.LATCH_4_.latch/Q mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_25_31 vpwr vgnd scs8hd_fill_2
XFILLER_25_53 vpwr vgnd scs8hd_fill_2
XFILLER_26_130 vgnd vpwr scs8hd_decap_12
XPHY_53 vgnd vpwr scs8hd_decap_3
XPHY_64 vgnd vpwr scs8hd_decap_3
X_193_ chany_bottom_in[4] chany_top_out[4] vgnd vpwr scs8hd_buf_2
XPHY_97 vgnd vpwr scs8hd_decap_3
XPHY_86 vgnd vpwr scs8hd_decap_3
XFILLER_41_52 vgnd vpwr scs8hd_decap_3
XPHY_75 vgnd vpwr scs8hd_decap_3
Xmem_right_ipin_7.LATCH_1_.latch data_in mem_right_ipin_7.LATCH_1_.latch/Q _141_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_5.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_ipin_7.LATCH_2_.latch/Q mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_11 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_ipin_3.LATCH_0_.latch_SLEEPB _109_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_144 vpwr vgnd scs8hd_fill_2
X_176_ _176_/HI _176_/LO vgnd vpwr scs8hd_conb_1
XFILLER_52_84 vgnd vpwr scs8hd_decap_8
XANTENNA__123__B _125_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_136 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _176_/HI mem_right_ipin_4.LATCH_5_.latch/Q
+ mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_7_107 vpwr vgnd scs8hd_fill_2
XFILLER_22_10 vpwr vgnd scs8hd_fill_2
XFILLER_22_32 vgnd vpwr scs8hd_fill_1
XFILLER_22_87 vgnd vpwr scs8hd_decap_3
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_73 vgnd vpwr scs8hd_fill_1
XFILLER_8_45 vpwr vgnd scs8hd_fill_2
XFILLER_8_23 vpwr vgnd scs8hd_fill_2
XANTENNA__118__B _118_/B vgnd vpwr scs8hd_diode_2
XANTENNA__134__A _064_/B vgnd vpwr scs8hd_diode_2
X_159_ _156_/B _159_/B _159_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_3 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_12_ vgnd vpwr scs8hd_inv_1
Xmux_right_ipin_0.INVTX1_3_.scs8hd_inv_1 chany_top_in[2] mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_53 vpwr vgnd scs8hd_fill_2
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_143 vgnd vpwr scs8hd_decap_3
XFILLER_3_121 vgnd vpwr scs8hd_fill_1
XFILLER_58_83 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_4.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__129__A _129_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_102 vgnd vpwr scs8hd_decap_4
XFILLER_28_42 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_6.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[3] mux_right_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_63 vpwr vgnd scs8hd_fill_2
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
XFILLER_5_35 vgnd vpwr scs8hd_fill_1
XANTENNA__131__B _129_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_117 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_ipin_1.LATCH_1_.latch_SLEEPB _088_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_2_.latch/Q mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_7.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[4] mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_11 vgnd vpwr scs8hd_fill_1
XFILLER_30_10 vpwr vgnd scs8hd_fill_2
XFILLER_30_32 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_7.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[8] mux_right_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__142__A _064_/B vgnd vpwr scs8hd_diode_2
XPHY_98 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_87 vgnd vpwr scs8hd_decap_3
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XFILLER_41_112 vgnd vpwr scs8hd_decap_8
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_26_142 vgnd vpwr scs8hd_decap_4
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_76 vgnd vpwr scs8hd_decap_3
X_192_ chany_bottom_in[5] chany_top_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_25_98 vpwr vgnd scs8hd_fill_2
XFILLER_2_69 vpwr vgnd scs8hd_fill_2
XANTENNA__137__A _129_/A vgnd vpwr scs8hd_diode_2
XFILLER_63_3 vgnd vpwr scs8hd_decap_12
XFILLER_23_123 vpwr vgnd scs8hd_fill_2
XFILLER_23_145 vgnd vpwr scs8hd_fill_1
XFILLER_36_42 vpwr vgnd scs8hd_fill_2
XFILLER_52_30 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_6.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_175_ _175_/HI _175_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_115 vgnd vpwr scs8hd_decap_6
XFILLER_7_119 vgnd vpwr scs8hd_decap_3
XFILLER_22_55 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_3.INVTX1_5_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_63_51 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_ipin_2.LATCH_1_.latch/Q mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_63_62 vgnd vpwr scs8hd_decap_12
XANTENNA__118__C _118_/C vgnd vpwr scs8hd_diode_2
X_089_ _117_/A _084_/B _089_/Y vgnd vpwr scs8hd_nor2_4
Xmem_right_ipin_0.LATCH_2_.latch data_in mem_right_ipin_0.LATCH_2_.latch/Q _076_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_158_ _157_/X _159_/B vgnd vpwr scs8hd_buf_1
XANTENNA__134__B _129_/B vgnd vpwr scs8hd_diode_2
XANTENNA__150__A _149_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_11 vpwr vgnd scs8hd_fill_2
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_43 vpwr vgnd scs8hd_fill_2
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_right_ipin_2.LATCH_5_.latch data_in mem_right_ipin_2.LATCH_5_.latch/Q _093_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__129__B _129_/B vgnd vpwr scs8hd_diode_2
XANTENNA__145__A _145_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_4.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_114 vgnd vpwr scs8hd_decap_8
XFILLER_28_32 vgnd vpwr scs8hd_fill_1
XFILLER_28_76 vgnd vpwr scs8hd_decap_6
Xmux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_ipin_6.LATCH_2_.latch/Q mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_53_143 vgnd vpwr scs8hd_decap_3
XFILLER_53_110 vpwr vgnd scs8hd_fill_2
XFILLER_14_23 vgnd vpwr scs8hd_decap_4
XFILLER_14_78 vgnd vpwr scs8hd_decap_8
XFILLER_14_89 vgnd vpwr scs8hd_decap_3
XFILLER_30_55 vpwr vgnd scs8hd_fill_2
XFILLER_39_53 vgnd vpwr scs8hd_decap_3
XANTENNA__142__B _142_/B vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_4.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[1] mux_right_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_50_102 vpwr vgnd scs8hd_fill_2
XFILLER_35_121 vgnd vpwr scs8hd_fill_1
XFILLER_35_143 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _175_/HI mem_right_ipin_3.LATCH_5_.latch/Q
+ mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_ipin_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_99 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_decap_3
XFILLER_41_135 vgnd vpwr scs8hd_decap_8
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_77 vgnd vpwr scs8hd_decap_3
X_191_ chany_bottom_in[6] chany_top_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_right_ipin_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_48 vpwr vgnd scs8hd_fill_2
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_17_121 vgnd vpwr scs8hd_fill_1
XFILLER_17_143 vgnd vpwr scs8hd_decap_3
XFILLER_32_102 vgnd vpwr scs8hd_decap_12
XANTENNA__137__B _142_/B vgnd vpwr scs8hd_diode_2
XFILLER_56_3 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_5.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[7] mux_right_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__153__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_6.LATCH_1_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_57 vpwr vgnd scs8hd_fill_2
XANTENNA__063__A _062_/X vgnd vpwr scs8hd_diode_2
XFILLER_11_79 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_ipin_1.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_36_10 vpwr vgnd scs8hd_fill_2
XFILLER_36_32 vgnd vpwr scs8hd_fill_1
X_174_ _174_/HI _174_/LO vgnd vpwr scs8hd_conb_1
XFILLER_28_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_5.INVTX1_3_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__148__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _170_/HI vgnd vpwr
+ scs8hd_diode_2
Xmem_right_ipin_3.LATCH_1_.latch data_in mem_right_ipin_3.LATCH_1_.latch/Q _108_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_23 vpwr vgnd scs8hd_fill_2
XFILLER_63_74 vgnd vpwr scs8hd_decap_12
X_157_ address[1] _147_/Y address[0] _157_/X vgnd vpwr scs8hd_or3_4
X_088_ _088_/A _084_/B _088_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_19_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_6.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_5.LATCH_4_.latch data_in mem_right_ipin_5.LATCH_4_.latch/Q _121_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_right_ipin_7.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_88 vgnd vpwr scs8hd_decap_4
XFILLER_3_123 vgnd vpwr scs8hd_decap_12
XANTENNA__161__A _161_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_4.LATCH_2_.latch_SLEEPB _115_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__071__A _159_/B vgnd vpwr scs8hd_diode_2
XFILLER_28_11 vpwr vgnd scs8hd_fill_2
XFILLER_28_22 vpwr vgnd scs8hd_fill_2
XFILLER_44_32 vgnd vpwr scs8hd_decap_3
XFILLER_60_97 vgnd vpwr scs8hd_decap_12
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__156__A _084_/A vgnd vpwr scs8hd_diode_2
XANTENNA__066__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_14_46 vpwr vgnd scs8hd_fill_2
Xmem_left_ipin_0.LATCH_2_.latch data_in mem_left_ipin_0.LATCH_2_.latch/Q _166_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_30_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_39_21 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_75 vpwr vgnd scs8hd_fill_2
XFILLER_55_53 vpwr vgnd scs8hd_fill_2
XFILLER_55_42 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_ipin_1.LATCH_1_.latch/Q mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_25_12 vpwr vgnd scs8hd_fill_2
XPHY_89 vgnd vpwr scs8hd_decap_3
XFILLER_41_103 vgnd vpwr scs8hd_decap_6
X_190_ chany_bottom_in[7] chany_top_out[7] vgnd vpwr scs8hd_buf_2
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_78 vgnd vpwr scs8hd_decap_3
XFILLER_41_99 vpwr vgnd scs8hd_fill_2
XFILLER_41_88 vpwr vgnd scs8hd_fill_2
XFILLER_41_77 vpwr vgnd scs8hd_fill_2
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XFILLER_32_114 vgnd vpwr scs8hd_decap_12
XANTENNA__153__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_49_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_3.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_23_114 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_2.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[3] mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_25 vpwr vgnd scs8hd_fill_2
XFILLER_11_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_7.INVTX1_1_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_36_88 vgnd vpwr scs8hd_decap_4
X_173_ _173_/HI _173_/LO vgnd vpwr scs8hd_conb_1
XFILLER_52_32 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_2.LATCH_3_.latch_SLEEPB _095_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_6.LATCH_0_.latch data_in mem_right_ipin_6.LATCH_0_.latch/Q _134_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__164__A _161_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_92 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_7.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__074__A _086_/A vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_3.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[5] mux_right_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_47_87 vpwr vgnd scs8hd_fill_2
XFILLER_47_65 vpwr vgnd scs8hd_fill_2
XFILLER_47_54 vgnd vpwr scs8hd_fill_1
XFILLER_63_86 vgnd vpwr scs8hd_decap_12
XFILLER_8_15 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_ipin_5.LATCH_2_.latch/Q mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_087_ _115_/A _084_/B _087_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_12_90 vpwr vgnd scs8hd_fill_2
X_156_ _084_/A _156_/B _156_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_40_7 vpwr vgnd scs8hd_fill_2
XANTENNA__159__A _156_/B vgnd vpwr scs8hd_diode_2
XANTENNA__069__A _068_/X vgnd vpwr scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_35 vpwr vgnd scs8hd_fill_2
XFILLER_17_57 vpwr vgnd scs8hd_fill_2
XFILLER_17_79 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _145_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_135 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _174_/HI mem_right_ipin_2.LATCH_5_.latch/Q
+ mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_139_ _131_/A _142_/B _139_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__161__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_28_89 vgnd vpwr scs8hd_fill_1
XFILLER_44_88 vpwr vgnd scs8hd_fill_2
XFILLER_60_76 vgnd vpwr scs8hd_fill_1
XFILLER_60_32 vgnd vpwr scs8hd_decap_12
XFILLER_5_38 vpwr vgnd scs8hd_fill_2
XFILLER_5_27 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_145 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_ipin_0.LATCH_4_.latch_SLEEPB _072_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__156__B _156_/B vgnd vpwr scs8hd_diode_2
XFILLER_53_123 vgnd vpwr scs8hd_decap_12
XANTENNA__066__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_30_68 vpwr vgnd scs8hd_fill_2
XFILLER_30_79 vpwr vgnd scs8hd_fill_2
XANTENNA__082__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_77 vpwr vgnd scs8hd_fill_2
XFILLER_39_11 vgnd vpwr scs8hd_decap_8
XFILLER_44_145 vgnd vpwr scs8hd_fill_1
XANTENNA__167__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_35_123 vgnd vpwr scs8hd_decap_12
XFILLER_6_81 vgnd vpwr scs8hd_decap_6
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XANTENNA__077__A _169_/B vgnd vpwr scs8hd_diode_2
XPHY_46 vgnd vpwr scs8hd_decap_3
XFILLER_25_35 vpwr vgnd scs8hd_fill_2
XFILLER_41_23 vpwr vgnd scs8hd_fill_2
XPHY_79 vgnd vpwr scs8hd_decap_3
XFILLER_25_57 vpwr vgnd scs8hd_fill_2
XFILLER_25_79 vpwr vgnd scs8hd_fill_2
XPHY_57 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XFILLER_9_3 vgnd vpwr scs8hd_decap_12
XFILLER_17_123 vgnd vpwr scs8hd_decap_12
XFILLER_32_126 vgnd vpwr scs8hd_decap_12
XANTENNA__153__C _099_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_23 vpwr vgnd scs8hd_fill_2
XFILLER_36_67 vpwr vgnd scs8hd_fill_2
XFILLER_52_44 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_4.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_172_ _172_/HI _172_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__164__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_61_3 vgnd vpwr scs8hd_decap_12
XANTENNA__180__A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_3_71 vgnd vpwr scs8hd_decap_4
XANTENNA__074__B _069_/X vgnd vpwr scs8hd_diode_2
XFILLER_11_107 vpwr vgnd scs8hd_fill_2
XFILLER_22_36 vgnd vpwr scs8hd_decap_3
XANTENNA__090__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_47_33 vpwr vgnd scs8hd_fill_2
XFILLER_47_22 vpwr vgnd scs8hd_fill_2
XFILLER_63_98 vgnd vpwr scs8hd_decap_12
XFILLER_8_49 vpwr vgnd scs8hd_fill_2
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_0.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[1] mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_086_ _086_/A _084_/B _086_/Y vgnd vpwr scs8hd_nor2_4
X_155_ _154_/X _156_/B vgnd vpwr scs8hd_buf_1
XFILLER_26_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__159__B _159_/B vgnd vpwr scs8hd_diode_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__085__A _085_/A vgnd vpwr scs8hd_diode_2
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_13 vpwr vgnd scs8hd_fill_2
XFILLER_33_57 vpwr vgnd scs8hd_fill_2
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_58_65 vgnd vpwr scs8hd_decap_3
XFILLER_58_43 vgnd vpwr scs8hd_decap_8
XFILLER_58_32 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_1.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[7] mux_right_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_ipin_1.LATCH_1_.latch_SLEEPB _143_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_7.LATCH_3_.latch_SLEEPB _139_/Y vgnd vpwr scs8hd_diode_2
X_069_ _068_/X _069_/X vgnd vpwr scs8hd_buf_1
XANTENNA__161__C _143_/C vgnd vpwr scs8hd_diode_2
X_138_ _159_/B _142_/B _138_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_3 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_1_.latch/Q mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_128 vpwr vgnd scs8hd_fill_2
XFILLER_56_110 vgnd vpwr scs8hd_decap_12
XFILLER_44_23 vpwr vgnd scs8hd_fill_2
XFILLER_44_12 vgnd vpwr scs8hd_decap_8
XFILLER_28_46 vpwr vgnd scs8hd_fill_2
XFILLER_60_55 vpwr vgnd scs8hd_fill_2
XFILLER_60_44 vgnd vpwr scs8hd_decap_8
Xmem_right_ipin_1.LATCH_4_.latch data_in mem_right_ipin_1.LATCH_4_.latch/Q _085_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_44_67 vgnd vpwr scs8hd_decap_6
XFILLER_47_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_7.INVTX1_1_.scs8hd_inv_1 chany_top_in[0] mux_right_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_53_135 vgnd vpwr scs8hd_decap_8
XFILLER_14_59 vgnd vpwr scs8hd_decap_6
XANTENNA__066__C _099_/C vgnd vpwr scs8hd_diode_2
XFILLER_30_36 vgnd vpwr scs8hd_fill_1
XANTENNA__082__B _118_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_34 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_6.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_121 vgnd vpwr scs8hd_fill_1
XFILLER_29_143 vgnd vpwr scs8hd_decap_3
XFILLER_55_88 vgnd vpwr scs8hd_decap_6
XFILLER_44_113 vgnd vpwr scs8hd_decap_12
XFILLER_44_102 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_113 vgnd vpwr scs8hd_decap_8
XFILLER_35_135 vgnd vpwr scs8hd_decap_8
XANTENNA__167__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__183__A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_6_60 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_ipin_4.LATCH_2_.latch/Q mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XFILLER_26_102 vpwr vgnd scs8hd_fill_2
XPHY_58 vgnd vpwr scs8hd_decap_3
XPHY_69 vgnd vpwr scs8hd_decap_3
XANTENNA__093__A _084_/A vgnd vpwr scs8hd_diode_2
XFILLER_41_57 vpwr vgnd scs8hd_fill_2
XFILLER_41_35 vpwr vgnd scs8hd_fill_2
XFILLER_17_113 vgnd vpwr scs8hd_decap_8
XFILLER_17_135 vgnd vpwr scs8hd_decap_8
XFILLER_32_138 vgnd vpwr scs8hd_decap_8
XFILLER_31_90 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_127 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_5.LATCH_4_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__088__A _088_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_46 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _173_/HI mem_right_ipin_1.LATCH_5_.latch/Q
+ mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_52_56 vgnd vpwr scs8hd_decap_12
XFILLER_52_23 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_2.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
X_171_ _171_/HI _171_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__164__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_54_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_6.INVTX1_5_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
X_085_ _085_/A _084_/B _085_/Y vgnd vpwr scs8hd_nor2_4
X_154_ address[5] address[6] _154_/C _154_/X vgnd vpwr scs8hd_or3_4
XANTENNA__191__A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_2.LATCH_0_.latch data_in mem_right_ipin_2.LATCH_0_.latch/Q _098_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_15 vgnd vpwr scs8hd_decap_4
XANTENNA__085__B _084_/B vgnd vpwr scs8hd_diode_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_47 vgnd vpwr scs8hd_decap_4
XFILLER_33_69 vpwr vgnd scs8hd_fill_2
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_137_ _129_/A _142_/B _137_/Y vgnd vpwr scs8hd_nor2_4
X_068_ _118_/A address[3] _082_/C _068_/X vgnd vpwr scs8hd_or3_4
Xmem_right_ipin_4.LATCH_3_.latch data_in mem_right_ipin_4.LATCH_3_.latch/Q _114_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__186__A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_56_122 vgnd vpwr scs8hd_decap_12
XFILLER_44_46 vpwr vgnd scs8hd_fill_2
XANTENNA__096__A _115_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_3.LATCH_5_.latch_SLEEPB _104_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_3.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_ipin_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_53_114 vgnd vpwr scs8hd_decap_8
XANTENNA__082__C _082_/C vgnd vpwr scs8hd_diode_2
XFILLER_55_23 vpwr vgnd scs8hd_fill_2
XFILLER_44_125 vgnd vpwr scs8hd_decap_12
XFILLER_50_106 vgnd vpwr scs8hd_decap_12
XANTENNA__167__C _143_/C vgnd vpwr scs8hd_diode_2
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XFILLER_25_48 vgnd vpwr scs8hd_decap_3
XPHY_59 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_5.INVTX1_1_.scs8hd_inv_1 chany_top_in[2] mux_right_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__093__B _093_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__194__A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_23_139 vgnd vpwr scs8hd_decap_6
XANTENNA__088__B _084_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_6.INVTX1_5_.scs8hd_inv_1 chany_top_in[8] mux_right_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_52_68 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_ipin_7.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_170_ _170_/HI _170_/LO vgnd vpwr scs8hd_conb_1
XFILLER_9_143 vgnd vpwr scs8hd_decap_3
XFILLER_9_121 vgnd vpwr scs8hd_fill_1
XFILLER_47_3 vpwr vgnd scs8hd_fill_2
XFILLER_3_40 vpwr vgnd scs8hd_fill_2
XANTENNA__189__A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_3_95 vgnd vpwr scs8hd_fill_1
XFILLER_22_27 vgnd vpwr scs8hd_decap_4
XANTENNA__099__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_47_57 vpwr vgnd scs8hd_fill_2
XFILLER_6_102 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _172_/HI vgnd vpwr
+ scs8hd_diode_2
X_153_ address[4] address[3] _099_/C _154_/C vgnd vpwr scs8hd_or3_4
X_084_ _084_/A _084_/B _084_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_9 vpwr vgnd scs8hd_fill_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_26 vpwr vgnd scs8hd_fill_2
XFILLER_3_105 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_7.LATCH_2_.latch data_in mem_right_ipin_7.LATCH_2_.latch/Q _140_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_59_131 vgnd vpwr scs8hd_decap_12
X_136_ _135_/X _142_/B vgnd vpwr scs8hd_buf_1
X_067_ _066_/X _082_/C vgnd vpwr scs8hd_buf_1
XFILLER_0_41 vpwr vgnd scs8hd_fill_2
XFILLER_0_74 vpwr vgnd scs8hd_fill_2
XFILLER_0_85 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_ipin_3.LATCH_2_.latch/Q mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_94 vpwr vgnd scs8hd_fill_2
XFILLER_56_134 vgnd vpwr scs8hd_decap_12
XFILLER_28_26 vgnd vpwr scs8hd_decap_4
XFILLER_28_59 vpwr vgnd scs8hd_fill_2
XANTENNA__096__B _093_/B vgnd vpwr scs8hd_diode_2
XFILLER_60_79 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_123 vgnd vpwr scs8hd_decap_12
XFILLER_18_81 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_91 vgnd vpwr scs8hd_fill_1
X_119_ _118_/X _125_/B vgnd vpwr scs8hd_buf_1
Xmux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _172_/HI mem_right_ipin_0.LATCH_5_.latch/Q
+ mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__197__A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_30_27 vpwr vgnd scs8hd_fill_2
XFILLER_55_57 vpwr vgnd scs8hd_fill_2
XFILLER_44_137 vgnd vpwr scs8hd_decap_8
XFILLER_39_58 vgnd vpwr scs8hd_decap_3
XFILLER_29_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_50_118 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_4.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_decap_3
XFILLER_25_16 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_6.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_2.LATCH_0_.latch_SLEEPB _098_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_29 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_4_ vgnd vpwr scs8hd_inv_1
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_3.INVTX1_1_.scs8hd_inv_1 chany_top_in[0] mux_right_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_7.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_70 vgnd vpwr scs8hd_fill_1
XFILLER_42_91 vgnd vpwr scs8hd_fill_1
XFILLER_9_111 vpwr vgnd scs8hd_fill_2
XFILLER_47_69 vgnd vpwr scs8hd_decap_4
XANTENNA__099__B address[6] vgnd vpwr scs8hd_diode_2
X_083_ _083_/A _084_/B vgnd vpwr scs8hd_buf_1
XFILLER_6_114 vgnd vpwr scs8hd_decap_12
XFILLER_12_50 vpwr vgnd scs8hd_fill_2
XFILLER_12_61 vgnd vpwr scs8hd_decap_3
X_152_ enable _099_/C vgnd vpwr scs8hd_inv_8
Xmux_right_ipin_4.INVTX1_5_.scs8hd_inv_1 chany_top_in[6] mux_right_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_39 vgnd vpwr scs8hd_decap_3
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_59_121 vgnd vpwr scs8hd_fill_1
XFILLER_59_143 vgnd vpwr scs8hd_decap_3
XFILLER_58_79 vpwr vgnd scs8hd_fill_2
XFILLER_23_71 vpwr vgnd scs8hd_fill_2
XFILLER_23_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_ipin_0.LATCH_4_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
X_066_ address[5] address[6] _099_/C _066_/X vgnd vpwr scs8hd_or3_4
X_135_ address[5] _127_/B _099_/C _101_/X _135_/X vgnd vpwr scs8hd_or4_4
XFILLER_9_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_6.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_0.LATCH_1_.latch_SLEEPB _078_/Y vgnd vpwr scs8hd_diode_2
XFILLER_62_105 vgnd vpwr scs8hd_decap_12
XFILLER_47_135 vgnd vpwr scs8hd_decap_8
XFILLER_18_60 vpwr vgnd scs8hd_fill_2
XFILLER_50_91 vgnd vpwr scs8hd_fill_1
X_118_ _118_/A _118_/B _118_/C _118_/X vgnd vpwr scs8hd_or3_4
XFILLER_38_102 vgnd vpwr scs8hd_decap_12
XFILLER_14_29 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_0.LATCH_3_.latch data_in mem_right_ipin_0.LATCH_3_.latch/Q _074_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_39 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_36 vgnd vpwr scs8hd_decap_4
XFILLER_29_135 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_92 vpwr vgnd scs8hd_fill_2
XFILLER_35_105 vpwr vgnd scs8hd_fill_2
XFILLER_6_52 vgnd vpwr scs8hd_decap_8
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_41_27 vpwr vgnd scs8hd_fill_2
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_40_141 vgnd vpwr scs8hd_decap_4
XFILLER_15_83 vpwr vgnd scs8hd_fill_2
XFILLER_31_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_4.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_19 vgnd vpwr scs8hd_decap_3
XFILLER_52_15 vgnd vpwr scs8hd_decap_8
XFILLER_14_108 vgnd vpwr scs8hd_decap_12
XFILLER_36_27 vpwr vgnd scs8hd_fill_2
XFILLER_52_26 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_130 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_ipin_2.LATCH_2_.latch/Q mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_123 vgnd vpwr scs8hd_decap_12
XFILLER_26_60 vpwr vgnd scs8hd_fill_2
XFILLER_26_82 vgnd vpwr scs8hd_decap_4
XFILLER_3_53 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_0_.latch/Q mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_47_37 vpwr vgnd scs8hd_fill_2
XFILLER_47_26 vpwr vgnd scs8hd_fill_2
XANTENNA__099__C _099_/C vgnd vpwr scs8hd_diode_2
XFILLER_6_126 vgnd vpwr scs8hd_decap_12
X_151_ _129_/A _084_/A vgnd vpwr scs8hd_buf_1
X_082_ _118_/A _118_/B _082_/C _083_/A vgnd vpwr scs8hd_or3_4
XANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _173_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_9 vpwr vgnd scs8hd_fill_2
XFILLER_37_92 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[2] mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_52_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_7.LATCH_0_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_134_ _064_/B _129_/B _134_/Y vgnd vpwr scs8hd_nor2_4
X_065_ address[4] _118_/A vgnd vpwr scs8hd_inv_8
XFILLER_48_91 vgnd vpwr scs8hd_fill_1
XFILLER_24_7 vgnd vpwr scs8hd_decap_3
XFILLER_0_32 vgnd vpwr scs8hd_fill_1
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
XFILLER_0_98 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_2.INVTX1_5_.scs8hd_inv_1 chany_top_in[8] mux_right_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_60_15 vgnd vpwr scs8hd_decap_12
XFILLER_44_27 vgnd vpwr scs8hd_decap_4
XFILLER_60_59 vpwr vgnd scs8hd_fill_2
XFILLER_62_117 vgnd vpwr scs8hd_decap_12
Xmem_right_ipin_3.LATCH_2_.latch data_in mem_right_ipin_3.LATCH_2_.latch/Q _107_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_117_ _117_/A _112_/B _117_/Y vgnd vpwr scs8hd_nor2_4
Xmux_left_ipin_1.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[1] mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_6.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_106 vpwr vgnd scs8hd_fill_2
XFILLER_15_3 vgnd vpwr scs8hd_decap_4
XFILLER_38_114 vgnd vpwr scs8hd_decap_12
XFILLER_39_38 vgnd vpwr scs8hd_decap_4
XFILLER_55_15 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_84 vgnd vpwr scs8hd_decap_8
Xmem_right_ipin_5.LATCH_5_.latch data_in mem_right_ipin_5.LATCH_5_.latch/Q _120_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_71 vgnd vpwr scs8hd_decap_4
XFILLER_6_42 vgnd vpwr scs8hd_decap_6
XFILLER_41_109 vgnd vpwr scs8hd_fill_1
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_26_106 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_39 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_1.INVTX1_3_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_5.LATCH_1_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_40 vpwr vgnd scs8hd_fill_2
XFILLER_15_62 vgnd vpwr scs8hd_decap_4
XANTENNA__102__A _118_/C vgnd vpwr scs8hd_diode_2
XFILLER_56_91 vgnd vpwr scs8hd_fill_1
XFILLER_56_80 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_5.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_52_38 vgnd vpwr scs8hd_decap_4
XFILLER_22_142 vgnd vpwr scs8hd_decap_4
XFILLER_26_50 vgnd vpwr scs8hd_fill_1
XFILLER_9_135 vgnd vpwr scs8hd_decap_8
XFILLER_13_120 vpwr vgnd scs8hd_fill_2
Xmem_left_ipin_0.LATCH_3_.latch data_in mem_left_ipin_0.LATCH_3_.latch/Q _163_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_65 vgnd vpwr scs8hd_decap_4
XFILLER_3_21 vgnd vpwr scs8hd_fill_1
XFILLER_63_15 vgnd vpwr scs8hd_decap_12
XFILLER_63_59 vpwr vgnd scs8hd_fill_2
X_150_ _149_/X _129_/A vgnd vpwr scs8hd_buf_1
XFILLER_6_138 vgnd vpwr scs8hd_decap_8
XFILLER_10_145 vgnd vpwr scs8hd_fill_1
XFILLER_12_30 vgnd vpwr scs8hd_fill_1
XFILLER_12_41 vgnd vpwr scs8hd_decap_3
X_081_ address[3] _118_/B vgnd vpwr scs8hd_inv_8
XFILLER_53_70 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_4.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_45_3 vgnd vpwr scs8hd_decap_12
XFILLER_17_19 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_ipin_5.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_59_101 vpwr vgnd scs8hd_fill_2
XFILLER_58_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_133_ _169_/B _129_/B _133_/Y vgnd vpwr scs8hd_nor2_4
X_064_ _156_/B _064_/B _064_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_48_70 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_3.LATCH_2_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_7 vpwr vgnd scs8hd_fill_2
XANTENNA__110__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_53 vpwr vgnd scs8hd_fill_2
XFILLER_9_75 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_6.LATCH_1_.latch data_in mem_right_ipin_6.LATCH_1_.latch/Q _133_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_60_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_47_104 vgnd vpwr scs8hd_decap_12
XFILLER_62_129 vgnd vpwr scs8hd_decap_12
X_116_ _088_/A _112_/B _116_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__105__A _085_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_83 vpwr vgnd scs8hd_fill_2
XFILLER_38_126 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_ipin_1.LATCH_2_.latch/Q mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_ipin_0.INVTX1_5_.scs8hd_inv_1 chany_top_in[6] mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_96 vpwr vgnd scs8hd_fill_2
XFILLER_29_50 vgnd vpwr scs8hd_decap_4
XFILLER_45_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_3.INVTX1_1_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_6_76 vgnd vpwr scs8hd_decap_3
XFILLER_6_65 vpwr vgnd scs8hd_fill_2
XFILLER_6_32 vgnd vpwr scs8hd_decap_4
XPHY_19 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_7.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_15_96 vpwr vgnd scs8hd_fill_2
XFILLER_31_95 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_6.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[7] mux_right_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__102__B _101_/X vgnd vpwr scs8hd_diode_2
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_121 vgnd vpwr scs8hd_fill_1
XFILLER_31_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_1.LATCH_3_.latch_SLEEPB _086_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[8] mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_83 vpwr vgnd scs8hd_fill_2
XFILLER_42_72 vpwr vgnd scs8hd_fill_2
XFILLER_13_143 vgnd vpwr scs8hd_decap_3
XANTENNA__113__A _085_/A vgnd vpwr scs8hd_diode_2
XFILLER_47_7 vgnd vpwr scs8hd_decap_12
XFILLER_3_88 vgnd vpwr scs8hd_decap_4
XFILLER_63_27 vgnd vpwr scs8hd_decap_12
X_080_ _117_/A _069_/X _080_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_102 vgnd vpwr scs8hd_decap_8
XFILLER_10_113 vgnd vpwr scs8hd_decap_12
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _174_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_53_60 vgnd vpwr scs8hd_fill_1
XANTENNA__108__A _088_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_109 vgnd vpwr scs8hd_decap_12
XFILLER_58_27 vgnd vpwr scs8hd_decap_4
X_063_ _062_/X _064_/B vgnd vpwr scs8hd_buf_1
XFILLER_23_52 vgnd vpwr scs8hd_decap_4
X_132_ _166_/B _129_/B _132_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_0_23 vpwr vgnd scs8hd_fill_2
XFILLER_0_78 vpwr vgnd scs8hd_fill_2
XANTENNA__110__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_0_89 vgnd vpwr scs8hd_decap_4
XFILLER_9_98 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_4.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_116 vgnd vpwr scs8hd_decap_6
XFILLER_18_85 vgnd vpwr scs8hd_decap_6
XFILLER_50_83 vpwr vgnd scs8hd_fill_2
XFILLER_50_72 vpwr vgnd scs8hd_fill_2
X_115_ _115_/A _112_/B _115_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__105__B _109_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_6 vpwr vgnd scs8hd_fill_2
XANTENNA__121__A _085_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_138 vgnd vpwr scs8hd_decap_8
XFILLER_20_42 vpwr vgnd scs8hd_fill_2
XFILLER_45_72 vpwr vgnd scs8hd_fill_2
XANTENNA__116__A _088_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_3 vpwr vgnd scs8hd_fill_2
XFILLER_26_119 vgnd vpwr scs8hd_decap_8
XFILLER_41_19 vgnd vpwr scs8hd_fill_1
XFILLER_25_141 vgnd vpwr scs8hd_decap_4
XFILLER_15_53 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_1.LATCH_5_.latch data_in mem_right_ipin_1.LATCH_5_.latch/Q _084_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_56_93 vgnd vpwr scs8hd_decap_3
XFILLER_56_60 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_10_ vgnd vpwr scs8hd_inv_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
.ends

