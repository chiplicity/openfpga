magic
tech EFS8A
magscale 1 2
timestamp 1602095458
<< locali >>
rect 7423 19873 7550 19907
rect 11063 17833 11069 17867
rect 11063 17765 11097 17833
rect 6043 16609 6078 16643
rect 15335 16609 15370 16643
rect 14467 15895 14501 15963
rect 14467 15861 14473 15895
rect 10419 15657 10425 15691
rect 10419 15589 10453 15657
rect 8251 15521 8286 15555
rect 2047 14569 2053 14603
rect 2047 14501 2081 14569
rect 8677 13787 8711 14025
rect 6739 13481 6745 13515
rect 6739 13413 6773 13481
rect 8159 13345 8194 13379
rect 15243 13345 15370 13379
rect 12811 12631 12845 12699
rect 12811 12597 12817 12631
rect 10419 12393 10425 12427
rect 10419 12325 10453 12393
rect 2139 11305 2145 11339
rect 4439 11305 4445 11339
rect 2139 11237 2173 11305
rect 4439 11237 4473 11305
rect 16859 10217 16865 10251
rect 16859 10149 16893 10217
rect 14007 9367 14041 9435
rect 14007 9333 14013 9367
rect 15663 9129 15669 9163
rect 15663 9061 15697 9129
rect 3801 8347 3835 8449
rect 9137 8279 9171 8517
rect 13823 8041 13829 8075
rect 13823 7973 13857 8041
rect 16899 7905 16934 7939
rect 3801 7191 3835 7497
rect 5089 7327 5123 7497
rect 15853 7259 15887 7497
rect 18003 6205 18130 6239
rect 15163 6069 15301 6103
rect 7751 4777 7757 4811
rect 7751 4709 7785 4777
rect 18423 3927 18457 3995
rect 18423 3893 18429 3927
rect 3007 3553 3042 3587
rect 2697 2839 2731 2941
<< viali >>
rect 10517 21097 10551 21131
rect 10333 20961 10367 20995
rect 13804 20961 13838 20995
rect 8677 20757 8711 20791
rect 13875 20757 13909 20791
rect 3801 20553 3835 20587
rect 8125 20553 8159 20587
rect 10333 20553 10367 20587
rect 14105 20553 14139 20587
rect 14473 20553 14507 20587
rect 15669 20553 15703 20587
rect 18889 20553 18923 20587
rect 21465 20553 21499 20587
rect 8677 20417 8711 20451
rect 1476 20349 1510 20383
rect 1869 20349 1903 20383
rect 2548 20349 2582 20383
rect 2973 20349 3007 20383
rect 3617 20349 3651 20383
rect 7640 20349 7674 20383
rect 10149 20349 10183 20383
rect 10701 20349 10735 20383
rect 13620 20349 13654 20383
rect 15184 20349 15218 20383
rect 18404 20349 18438 20383
rect 20980 20349 21014 20383
rect 8493 20281 8527 20315
rect 8769 20281 8803 20315
rect 9321 20281 9355 20315
rect 1547 20213 1581 20247
rect 2651 20213 2685 20247
rect 4261 20213 4295 20247
rect 7711 20213 7745 20247
rect 11069 20213 11103 20247
rect 13691 20213 13725 20247
rect 15255 20213 15289 20247
rect 18475 20213 18509 20247
rect 21051 20213 21085 20247
rect 1593 20009 1627 20043
rect 7619 20009 7653 20043
rect 10057 19941 10091 19975
rect 13730 19941 13764 19975
rect 15485 19941 15519 19975
rect 2120 19873 2154 19907
rect 7389 19873 7423 19907
rect 8528 19873 8562 19907
rect 12608 19873 12642 19907
rect 16932 19873 16966 19907
rect 20980 19873 21014 19907
rect 9965 19805 9999 19839
rect 10241 19805 10275 19839
rect 11437 19805 11471 19839
rect 13461 19805 13495 19839
rect 13645 19805 13679 19839
rect 14289 19805 14323 19839
rect 15393 19805 15427 19839
rect 15669 19805 15703 19839
rect 2191 19669 2225 19703
rect 6837 19669 6871 19703
rect 8631 19669 8665 19703
rect 8953 19669 8987 19703
rect 12679 19669 12713 19703
rect 17003 19669 17037 19703
rect 21051 19669 21085 19703
rect 2145 19465 2179 19499
rect 7849 19465 7883 19499
rect 8493 19465 8527 19499
rect 9781 19465 9815 19499
rect 16405 19465 16439 19499
rect 16957 19465 16991 19499
rect 19257 19465 19291 19499
rect 21097 19465 21131 19499
rect 21465 19465 21499 19499
rect 22109 19465 22143 19499
rect 6653 19397 6687 19431
rect 16037 19397 16071 19431
rect 7205 19329 7239 19363
rect 8861 19329 8895 19363
rect 9505 19329 9539 19363
rect 10241 19329 10275 19363
rect 10425 19329 10459 19363
rect 10701 19329 10735 19363
rect 14381 19329 14415 19363
rect 1444 19261 1478 19295
rect 12608 19261 12642 19295
rect 13001 19261 13035 19295
rect 13369 19261 13403 19295
rect 15612 19261 15646 19295
rect 18772 19261 18806 19295
rect 20612 19261 20646 19295
rect 21624 19261 21658 19295
rect 1547 19193 1581 19227
rect 6929 19193 6963 19227
rect 7021 19193 7055 19227
rect 8953 19193 8987 19227
rect 10517 19193 10551 19227
rect 14105 19193 14139 19227
rect 14197 19193 14231 19227
rect 15301 19193 15335 19227
rect 12679 19125 12713 19159
rect 13737 19125 13771 19159
rect 15715 19125 15749 19159
rect 18843 19125 18877 19159
rect 20683 19125 20717 19159
rect 21695 19125 21729 19159
rect 1593 18921 1627 18955
rect 14473 18921 14507 18955
rect 16313 18921 16347 18955
rect 18153 18921 18187 18955
rect 5273 18853 5307 18887
rect 5365 18853 5399 18887
rect 6929 18853 6963 18887
rect 10977 18853 11011 18887
rect 13001 18853 13035 18887
rect 13093 18853 13127 18887
rect 13645 18853 13679 18887
rect 15485 18853 15519 18887
rect 16957 18853 16991 18887
rect 17049 18853 17083 18887
rect 1409 18785 1443 18819
rect 8344 18785 8378 18819
rect 9965 18785 9999 18819
rect 2513 18717 2547 18751
rect 6837 18717 6871 18751
rect 7113 18717 7147 18751
rect 10885 18717 10919 18751
rect 11161 18717 11195 18751
rect 15393 18717 15427 18751
rect 16037 18717 16071 18751
rect 17233 18717 17267 18751
rect 5825 18649 5859 18683
rect 8447 18581 8481 18615
rect 8861 18581 8895 18615
rect 10425 18581 10459 18615
rect 14105 18581 14139 18615
rect 1961 18377 1995 18411
rect 2651 18377 2685 18411
rect 5549 18377 5583 18411
rect 6653 18377 6687 18411
rect 8309 18377 8343 18411
rect 17325 18377 17359 18411
rect 5273 18309 5307 18343
rect 9321 18309 9355 18343
rect 9965 18309 9999 18343
rect 15025 18309 15059 18343
rect 17049 18309 17083 18343
rect 6929 18241 6963 18275
rect 8769 18241 8803 18275
rect 10333 18241 10367 18275
rect 12541 18241 12575 18275
rect 12817 18241 12851 18275
rect 13921 18241 13955 18275
rect 14473 18241 14507 18275
rect 16037 18241 16071 18275
rect 16681 18241 16715 18275
rect 18153 18241 18187 18275
rect 18429 18241 18463 18275
rect 1409 18173 1443 18207
rect 2580 18173 2614 18207
rect 2973 18173 3007 18207
rect 7021 18105 7055 18139
rect 7573 18105 7607 18139
rect 8033 18105 8067 18139
rect 8861 18105 8895 18139
rect 10885 18105 10919 18139
rect 10977 18105 11011 18139
rect 11529 18105 11563 18139
rect 12633 18105 12667 18139
rect 14289 18105 14323 18139
rect 14565 18105 14599 18139
rect 16129 18105 16163 18139
rect 18245 18105 18279 18139
rect 1593 18037 1627 18071
rect 2421 18037 2455 18071
rect 4537 18037 4571 18071
rect 6285 18037 6319 18071
rect 10609 18037 10643 18071
rect 11805 18037 11839 18071
rect 12173 18037 12207 18071
rect 13461 18037 13495 18071
rect 15485 18037 15519 18071
rect 15853 18037 15887 18071
rect 17785 18037 17819 18071
rect 6561 17833 6595 17867
rect 7573 17833 7607 17867
rect 9045 17833 9079 17867
rect 11069 17833 11103 17867
rect 11621 17833 11655 17867
rect 12541 17833 12575 17867
rect 12909 17833 12943 17867
rect 15485 17833 15519 17867
rect 5962 17765 5996 17799
rect 7205 17765 7239 17799
rect 15853 17765 15887 17799
rect 17417 17765 17451 17799
rect 2237 17697 2271 17731
rect 3893 17697 3927 17731
rect 4169 17697 4203 17731
rect 4537 17697 4571 17731
rect 8033 17697 8067 17731
rect 8493 17697 8527 17731
rect 13093 17697 13127 17731
rect 13553 17697 13587 17731
rect 4629 17629 4663 17663
rect 5641 17629 5675 17663
rect 8585 17629 8619 17663
rect 10701 17629 10735 17663
rect 13829 17629 13863 17663
rect 14105 17629 14139 17663
rect 15761 17629 15795 17663
rect 17325 17629 17359 17663
rect 18797 17629 18831 17663
rect 16313 17561 16347 17595
rect 17877 17561 17911 17595
rect 1961 17493 1995 17527
rect 6929 17493 6963 17527
rect 10517 17493 10551 17527
rect 18337 17493 18371 17527
rect 2605 17289 2639 17323
rect 5181 17289 5215 17323
rect 8125 17289 8159 17323
rect 9505 17289 9539 17323
rect 11345 17289 11379 17323
rect 13185 17289 13219 17323
rect 14841 17289 14875 17323
rect 15577 17289 15611 17323
rect 17325 17289 17359 17323
rect 21097 17289 21131 17323
rect 12725 17221 12759 17255
rect 1685 17153 1719 17187
rect 2329 17153 2363 17187
rect 8585 17153 8619 17187
rect 11621 17153 11655 17187
rect 13921 17153 13955 17187
rect 18245 17153 18279 17187
rect 18705 17153 18739 17187
rect 3192 17085 3226 17119
rect 3617 17085 3651 17119
rect 4261 17085 4295 17119
rect 6561 17085 6595 17119
rect 7113 17085 7147 17119
rect 7297 17085 7331 17119
rect 10425 17085 10459 17119
rect 20913 17085 20947 17119
rect 21465 17085 21499 17119
rect 1777 17017 1811 17051
rect 4582 17017 4616 17051
rect 5641 17017 5675 17051
rect 6101 17017 6135 17051
rect 8906 17017 8940 17051
rect 10787 17017 10821 17051
rect 14242 17017 14276 17051
rect 16129 17017 16163 17051
rect 16221 17017 16255 17051
rect 16773 17017 16807 17051
rect 18337 17017 18371 17051
rect 2973 16949 3007 16983
rect 3295 16949 3329 16983
rect 4169 16949 4203 16983
rect 6929 16949 6963 16983
rect 8401 16949 8435 16983
rect 9965 16949 9999 16983
rect 10333 16949 10367 16983
rect 13737 16949 13771 16983
rect 15209 16949 15243 16983
rect 15853 16949 15887 16983
rect 17601 16949 17635 16983
rect 1685 16745 1719 16779
rect 4353 16745 4387 16779
rect 5089 16745 5123 16779
rect 7941 16745 7975 16779
rect 8585 16745 8619 16779
rect 11713 16745 11747 16779
rect 15439 16745 15473 16779
rect 16129 16745 16163 16779
rect 18245 16745 18279 16779
rect 2145 16677 2179 16711
rect 6837 16677 6871 16711
rect 7383 16677 7417 16711
rect 10793 16677 10827 16711
rect 16451 16677 16485 16711
rect 17646 16677 17680 16711
rect 4169 16609 4203 16643
rect 4629 16609 4663 16643
rect 6009 16609 6043 16643
rect 10333 16609 10367 16643
rect 10517 16609 10551 16643
rect 11069 16609 11103 16643
rect 11621 16609 11655 16643
rect 12081 16609 12115 16643
rect 13277 16609 13311 16643
rect 13829 16609 13863 16643
rect 15301 16609 15335 16643
rect 16348 16609 16382 16643
rect 18521 16609 18555 16643
rect 2053 16541 2087 16575
rect 2329 16541 2363 16575
rect 7021 16541 7055 16575
rect 14013 16541 14047 16575
rect 17325 16541 17359 16575
rect 2973 16473 3007 16507
rect 8217 16473 8251 16507
rect 3893 16405 3927 16439
rect 6147 16405 6181 16439
rect 9045 16405 9079 16439
rect 5365 16201 5399 16235
rect 8861 16201 8895 16235
rect 15025 16201 15059 16235
rect 16129 16201 16163 16235
rect 20131 16201 20165 16235
rect 3893 16133 3927 16167
rect 10057 16133 10091 16167
rect 18705 16133 18739 16167
rect 2053 16065 2087 16099
rect 2421 16065 2455 16099
rect 3617 16065 3651 16099
rect 4445 16065 4479 16099
rect 5641 16065 5675 16099
rect 9045 16065 9079 16099
rect 12265 16065 12299 16099
rect 14105 16065 14139 16099
rect 17049 16065 17083 16099
rect 17693 16065 17727 16099
rect 18153 16065 18187 16099
rect 19073 16065 19107 16099
rect 6653 15997 6687 16031
rect 7113 15997 7147 16031
rect 7297 15997 7331 16031
rect 7849 15997 7883 16031
rect 10793 15997 10827 16031
rect 10977 15997 11011 16031
rect 12633 15997 12667 16031
rect 12909 15997 12943 16031
rect 15393 15997 15427 16031
rect 16313 15997 16347 16031
rect 16773 15997 16807 16031
rect 20028 15997 20062 16031
rect 20453 15997 20487 16031
rect 2145 15929 2179 15963
rect 4807 15929 4841 15963
rect 7573 15929 7607 15963
rect 9137 15929 9171 15963
rect 9689 15929 9723 15963
rect 11897 15929 11931 15963
rect 18245 15929 18279 15963
rect 1869 15861 1903 15895
rect 2973 15861 3007 15895
rect 4353 15861 4387 15895
rect 6101 15861 6135 15895
rect 10609 15861 10643 15895
rect 12541 15861 12575 15895
rect 13461 15861 13495 15895
rect 14013 15861 14047 15895
rect 14473 15861 14507 15895
rect 15761 15861 15795 15895
rect 17325 15861 17359 15895
rect 1961 15657 1995 15691
rect 2697 15657 2731 15691
rect 5273 15657 5307 15691
rect 7665 15657 7699 15691
rect 10425 15657 10459 15691
rect 11621 15657 11655 15691
rect 11989 15657 12023 15691
rect 14105 15657 14139 15691
rect 16589 15657 16623 15691
rect 18061 15657 18095 15691
rect 18337 15657 18371 15691
rect 21097 15657 21131 15691
rect 4353 15589 4387 15623
rect 6745 15589 6779 15623
rect 6837 15589 6871 15623
rect 9965 15589 9999 15623
rect 12811 15589 12845 15623
rect 17462 15589 17496 15623
rect 2329 15521 2363 15555
rect 8217 15521 8251 15555
rect 10057 15521 10091 15555
rect 12449 15521 12483 15555
rect 15577 15521 15611 15555
rect 16037 15521 16071 15555
rect 20913 15521 20947 15555
rect 4261 15453 4295 15487
rect 7389 15453 7423 15487
rect 11345 15453 11379 15487
rect 16313 15453 16347 15487
rect 17141 15453 17175 15487
rect 4813 15385 4847 15419
rect 8355 15317 8389 15351
rect 8769 15317 8803 15351
rect 10977 15317 11011 15351
rect 13369 15317 13403 15351
rect 13737 15317 13771 15351
rect 4261 15113 4295 15147
rect 4629 15113 4663 15147
rect 6285 15113 6319 15147
rect 6653 15113 6687 15147
rect 11437 15113 11471 15147
rect 13461 15113 13495 15147
rect 15117 15113 15151 15147
rect 17509 15113 17543 15147
rect 21097 15113 21131 15147
rect 2421 15045 2455 15079
rect 7757 15045 7791 15079
rect 15393 15045 15427 15079
rect 20729 15045 20763 15079
rect 1869 14977 1903 15011
rect 3157 14977 3191 15011
rect 3479 14977 3513 15011
rect 4905 14977 4939 15011
rect 5181 14977 5215 15011
rect 7205 14977 7239 15011
rect 10425 14977 10459 15011
rect 11713 14977 11747 15011
rect 3392 14909 3426 14943
rect 8953 14909 8987 14943
rect 9229 14909 9263 14943
rect 12516 14909 12550 14943
rect 13553 14909 13587 14943
rect 15577 14909 15611 14943
rect 16037 14909 16071 14943
rect 20913 14909 20947 14943
rect 1961 14841 1995 14875
rect 4997 14841 5031 14875
rect 7297 14841 7331 14875
rect 8309 14841 8343 14875
rect 9781 14841 9815 14875
rect 10517 14841 10551 14875
rect 11069 14841 11103 14875
rect 13874 14841 13908 14875
rect 16313 14841 16347 14875
rect 21465 14841 21499 14875
rect 1685 14773 1719 14807
rect 2789 14773 2823 14807
rect 3801 14773 3835 14807
rect 8769 14773 8803 14807
rect 10149 14773 10183 14807
rect 12173 14773 12207 14807
rect 12587 14773 12621 14807
rect 12909 14773 12943 14807
rect 14473 14773 14507 14807
rect 17141 14773 17175 14807
rect 2053 14569 2087 14603
rect 2605 14569 2639 14603
rect 4629 14569 4663 14603
rect 7481 14569 7515 14603
rect 7941 14569 7975 14603
rect 11391 14569 11425 14603
rect 12541 14569 12575 14603
rect 15945 14569 15979 14603
rect 4997 14501 5031 14535
rect 5089 14501 5123 14535
rect 6653 14501 6687 14535
rect 8217 14501 8251 14535
rect 9137 14501 9171 14535
rect 9873 14501 9907 14535
rect 10793 14501 10827 14535
rect 12817 14501 12851 14535
rect 15669 14501 15703 14535
rect 16583 14501 16617 14535
rect 5641 14433 5675 14467
rect 11320 14433 11354 14467
rect 14232 14433 14266 14467
rect 1685 14365 1719 14399
rect 6561 14365 6595 14399
rect 6837 14365 6871 14399
rect 8125 14365 8159 14399
rect 8401 14365 8435 14399
rect 9781 14365 9815 14399
rect 10057 14365 10091 14399
rect 12725 14365 12759 14399
rect 13369 14365 13403 14399
rect 16221 14365 16255 14399
rect 4261 14229 4295 14263
rect 6285 14229 6319 14263
rect 13645 14229 13679 14263
rect 14335 14229 14369 14263
rect 14657 14229 14691 14263
rect 17141 14229 17175 14263
rect 2513 14025 2547 14059
rect 5181 14025 5215 14059
rect 5457 14025 5491 14059
rect 6561 14025 6595 14059
rect 8033 14025 8067 14059
rect 8401 14025 8435 14059
rect 8677 14025 8711 14059
rect 8769 14025 8803 14059
rect 9873 14025 9907 14059
rect 10149 14025 10183 14059
rect 11805 14025 11839 14059
rect 12265 14025 12299 14059
rect 4261 13889 4295 13923
rect 7021 13889 7055 13923
rect 7665 13889 7699 13923
rect 1593 13821 1627 13855
rect 4077 13821 4111 13855
rect 16313 13957 16347 13991
rect 8953 13889 8987 13923
rect 13461 13889 13495 13923
rect 14657 13889 14691 13923
rect 14933 13889 14967 13923
rect 15945 13889 15979 13923
rect 10885 13821 10919 13855
rect 11253 13821 11287 13855
rect 12725 13821 12759 13855
rect 13185 13821 13219 13855
rect 17141 13821 17175 13855
rect 1934 13753 1968 13787
rect 2789 13753 2823 13787
rect 3249 13753 3283 13787
rect 4582 13753 4616 13787
rect 6193 13753 6227 13787
rect 7113 13753 7147 13787
rect 8677 13753 8711 13787
rect 9274 13753 9308 13787
rect 10701 13753 10735 13787
rect 11529 13753 11563 13787
rect 13829 13753 13863 13787
rect 14197 13753 14231 13787
rect 14749 13753 14783 13787
rect 16497 13753 16531 13787
rect 16589 13753 16623 13787
rect 17509 13685 17543 13719
rect 1593 13481 1627 13515
rect 2651 13481 2685 13515
rect 4261 13481 4295 13515
rect 5641 13481 5675 13515
rect 6745 13481 6779 13515
rect 7297 13481 7331 13515
rect 7573 13481 7607 13515
rect 8263 13481 8297 13515
rect 8953 13481 8987 13515
rect 12173 13481 12207 13515
rect 12449 13481 12483 13515
rect 14657 13481 14691 13515
rect 16497 13481 16531 13515
rect 17601 13481 17635 13515
rect 21097 13481 21131 13515
rect 10701 13413 10735 13447
rect 11253 13413 11287 13447
rect 12995 13413 13029 13447
rect 17002 13413 17036 13447
rect 18613 13413 18647 13447
rect 1409 13345 1443 13379
rect 2580 13345 2614 13379
rect 4169 13345 4203 13379
rect 4721 13345 4755 13379
rect 8125 13345 8159 13379
rect 12633 13345 12667 13379
rect 15209 13345 15243 13379
rect 20913 13345 20947 13379
rect 6377 13277 6411 13311
rect 10609 13277 10643 13311
rect 16681 13277 16715 13311
rect 18521 13277 18555 13311
rect 18797 13277 18831 13311
rect 16129 13209 16163 13243
rect 1961 13141 1995 13175
rect 2329 13141 2363 13175
rect 5273 13141 5307 13175
rect 9873 13141 9907 13175
rect 13553 13141 13587 13175
rect 14289 13141 14323 13175
rect 15439 13141 15473 13175
rect 15853 13141 15887 13175
rect 4307 12937 4341 12971
rect 8723 12937 8757 12971
rect 10977 12937 11011 12971
rect 11299 12937 11333 12971
rect 13645 12937 13679 12971
rect 14013 12937 14047 12971
rect 18199 12937 18233 12971
rect 18889 12937 18923 12971
rect 6377 12869 6411 12903
rect 19257 12869 19291 12903
rect 20683 12869 20717 12903
rect 21373 12869 21407 12903
rect 12449 12801 12483 12835
rect 14565 12801 14599 12835
rect 16497 12801 16531 12835
rect 17141 12801 17175 12835
rect 1961 12733 1995 12767
rect 2145 12733 2179 12767
rect 4204 12733 4238 12767
rect 4629 12733 4663 12767
rect 5365 12733 5399 12767
rect 5733 12733 5767 12767
rect 5917 12733 5951 12767
rect 6929 12733 6963 12767
rect 8217 12733 8251 12767
rect 8652 12733 8686 12767
rect 9137 12733 9171 12767
rect 9597 12733 9631 12767
rect 10149 12733 10183 12767
rect 11196 12733 11230 12767
rect 11621 12733 11655 12767
rect 15761 12733 15795 12767
rect 16221 12733 16255 12767
rect 18096 12733 18130 12767
rect 19568 12733 19602 12767
rect 19993 12733 20027 12767
rect 20612 12733 20646 12767
rect 21005 12733 21039 12767
rect 4077 12665 4111 12699
rect 5089 12665 5123 12699
rect 6837 12665 6871 12699
rect 9505 12665 9539 12699
rect 14289 12665 14323 12699
rect 14381 12665 14415 12699
rect 18521 12665 18555 12699
rect 2513 12597 2547 12631
rect 3157 12597 3191 12631
rect 3709 12597 3743 12631
rect 9873 12597 9907 12631
rect 10701 12597 10735 12631
rect 12265 12597 12299 12631
rect 12817 12597 12851 12631
rect 13369 12597 13403 12631
rect 15301 12597 15335 12631
rect 16865 12597 16899 12631
rect 19671 12597 19705 12631
rect 6377 12393 6411 12427
rect 8769 12393 8803 12427
rect 9873 12393 9907 12427
rect 10425 12393 10459 12427
rect 10977 12393 11011 12427
rect 12541 12393 12575 12427
rect 14749 12393 14783 12427
rect 2513 12325 2547 12359
rect 4997 12325 5031 12359
rect 13461 12325 13495 12359
rect 14013 12325 14047 12359
rect 15485 12325 15519 12359
rect 8033 12257 8067 12291
rect 10057 12257 10091 12291
rect 20913 12257 20947 12291
rect 2421 12189 2455 12223
rect 4905 12189 4939 12223
rect 7757 12189 7791 12223
rect 13369 12189 13403 12223
rect 15393 12189 15427 12223
rect 16865 12189 16899 12223
rect 2973 12121 3007 12155
rect 4261 12121 4295 12155
rect 5457 12121 5491 12155
rect 15945 12121 15979 12155
rect 1685 12053 1719 12087
rect 2145 12053 2179 12087
rect 6837 12053 6871 12087
rect 7205 12053 7239 12087
rect 12817 12053 12851 12087
rect 21097 12053 21131 12087
rect 1547 11849 1581 11883
rect 2329 11849 2363 11883
rect 5641 11849 5675 11883
rect 6653 11849 6687 11883
rect 9965 11849 9999 11883
rect 11069 11849 11103 11883
rect 12265 11849 12299 11883
rect 13461 11849 13495 11883
rect 14565 11849 14599 11883
rect 15669 11849 15703 11883
rect 20913 11849 20947 11883
rect 3065 11781 3099 11815
rect 4353 11713 4387 11747
rect 4997 11713 5031 11747
rect 7113 11713 7147 11747
rect 7389 11713 7423 11747
rect 8677 11713 8711 11747
rect 8953 11713 8987 11747
rect 13001 11713 13035 11747
rect 13921 11713 13955 11747
rect 15025 11713 15059 11747
rect 1476 11645 1510 11679
rect 10216 11645 10250 11679
rect 12449 11645 12483 11679
rect 12909 11645 12943 11679
rect 16129 11645 16163 11679
rect 16221 11645 16255 11679
rect 16681 11645 16715 11679
rect 2513 11577 2547 11611
rect 2605 11577 2639 11611
rect 3433 11577 3467 11611
rect 4169 11577 4203 11611
rect 4445 11577 4479 11611
rect 7205 11577 7239 11611
rect 8769 11577 8803 11611
rect 11805 11577 11839 11611
rect 14749 11577 14783 11611
rect 14841 11577 14875 11611
rect 1961 11509 1995 11543
rect 5365 11509 5399 11543
rect 8033 11509 8067 11543
rect 8401 11509 8435 11543
rect 10287 11509 10321 11543
rect 10701 11509 10735 11543
rect 16497 11509 16531 11543
rect 2145 11305 2179 11339
rect 2973 11305 3007 11339
rect 4445 11305 4479 11339
rect 4997 11305 5031 11339
rect 5825 11305 5859 11339
rect 12449 11305 12483 11339
rect 7113 11237 7147 11271
rect 10701 11237 10735 11271
rect 11891 11237 11925 11271
rect 13461 11237 13495 11271
rect 14013 11237 14047 11271
rect 14749 11237 14783 11271
rect 15117 11237 15151 11271
rect 15485 11237 15519 11271
rect 18705 11237 18739 11271
rect 2697 11169 2731 11203
rect 9965 11169 9999 11203
rect 10241 11169 10275 11203
rect 20980 11169 21014 11203
rect 1777 11101 1811 11135
rect 4077 11101 4111 11135
rect 7021 11101 7055 11135
rect 7389 11101 7423 11135
rect 8033 11101 8067 11135
rect 8493 11101 8527 11135
rect 11529 11101 11563 11135
rect 13369 11101 13403 11135
rect 15393 11101 15427 11135
rect 15669 11101 15703 11135
rect 18613 11101 18647 11135
rect 10057 11033 10091 11067
rect 19165 11033 19199 11067
rect 16497 10965 16531 10999
rect 21051 10965 21085 10999
rect 1593 10761 1627 10795
rect 2329 10761 2363 10795
rect 2651 10761 2685 10795
rect 6285 10761 6319 10795
rect 7757 10761 7791 10795
rect 11161 10761 11195 10795
rect 11621 10761 11655 10795
rect 13369 10761 13403 10795
rect 14841 10761 14875 10795
rect 15301 10761 15335 10795
rect 16221 10761 16255 10795
rect 20913 10761 20947 10795
rect 4169 10693 4203 10727
rect 6975 10693 7009 10727
rect 13001 10693 13035 10727
rect 5089 10625 5123 10659
rect 7941 10625 7975 10659
rect 8401 10625 8435 10659
rect 9505 10625 9539 10659
rect 9781 10625 9815 10659
rect 17877 10625 17911 10659
rect 1409 10557 1443 10591
rect 2548 10557 2582 10591
rect 2973 10557 3007 10591
rect 3801 10557 3835 10591
rect 4813 10557 4847 10591
rect 6904 10557 6938 10591
rect 12516 10557 12550 10591
rect 13921 10557 13955 10591
rect 16405 10557 16439 10591
rect 16957 10557 16991 10591
rect 7297 10489 7331 10523
rect 8033 10489 8067 10523
rect 9597 10489 9631 10523
rect 13829 10489 13863 10523
rect 14283 10489 14317 10523
rect 17141 10489 17175 10523
rect 18613 10489 18647 10523
rect 18705 10489 18739 10523
rect 19257 10489 19291 10523
rect 2053 10421 2087 10455
rect 3341 10421 3375 10455
rect 5457 10421 5491 10455
rect 6653 10421 6687 10455
rect 9229 10421 9263 10455
rect 10425 10421 10459 10455
rect 10793 10421 10827 10455
rect 11897 10421 11931 10455
rect 12587 10421 12621 10455
rect 15761 10421 15795 10455
rect 18337 10421 18371 10455
rect 19533 10421 19567 10455
rect 19901 10421 19935 10455
rect 2651 10217 2685 10251
rect 3801 10217 3835 10251
rect 4261 10217 4295 10251
rect 7941 10217 7975 10251
rect 9505 10217 9539 10251
rect 12541 10217 12575 10251
rect 16865 10217 16899 10251
rect 19165 10217 19199 10251
rect 7342 10149 7376 10183
rect 11621 10149 11655 10183
rect 18566 10149 18600 10183
rect 1409 10081 1443 10115
rect 2580 10081 2614 10115
rect 4813 10081 4847 10115
rect 5181 10081 5215 10115
rect 5549 10081 5583 10115
rect 6101 10081 6135 10115
rect 10977 10081 11011 10115
rect 11437 10081 11471 10115
rect 13185 10081 13219 10115
rect 13369 10081 13403 10115
rect 13645 10081 13679 10115
rect 13921 10081 13955 10115
rect 15368 10081 15402 10115
rect 16497 10081 16531 10115
rect 20913 10081 20947 10115
rect 2053 10013 2087 10047
rect 6193 10013 6227 10047
rect 7021 10013 7055 10047
rect 14289 10013 14323 10047
rect 18245 10013 18279 10047
rect 1593 9945 1627 9979
rect 3341 9945 3375 9979
rect 10333 9945 10367 9979
rect 21097 9945 21131 9979
rect 2329 9877 2363 9911
rect 3065 9877 3099 9911
rect 8217 9877 8251 9911
rect 10609 9877 10643 9911
rect 15439 9877 15473 9911
rect 15853 9877 15887 9911
rect 17417 9877 17451 9911
rect 6285 9673 6319 9707
rect 7113 9673 7147 9707
rect 7389 9673 7423 9707
rect 10406 9673 10440 9707
rect 10885 9673 10919 9707
rect 11345 9673 11379 9707
rect 13553 9673 13587 9707
rect 17049 9673 17083 9707
rect 17785 9673 17819 9707
rect 5549 9605 5583 9639
rect 10517 9605 10551 9639
rect 16313 9605 16347 9639
rect 3617 9537 3651 9571
rect 8769 9537 8803 9571
rect 10609 9537 10643 9571
rect 19165 9537 19199 9571
rect 2145 9469 2179 9503
rect 2421 9469 2455 9503
rect 2697 9469 2731 9503
rect 3157 9469 3191 9503
rect 4169 9469 4203 9503
rect 4629 9469 4663 9503
rect 5181 9469 5215 9503
rect 5549 9469 5583 9503
rect 12700 9469 12734 9503
rect 13645 9469 13679 9503
rect 15209 9469 15243 9503
rect 8125 9401 8159 9435
rect 8217 9401 8251 9435
rect 10241 9401 10275 9435
rect 15761 9401 15795 9435
rect 15853 9401 15887 9435
rect 18889 9401 18923 9435
rect 19257 9401 19291 9435
rect 19809 9401 19843 9435
rect 1777 9333 1811 9367
rect 2145 9333 2179 9367
rect 4077 9333 4111 9367
rect 6009 9333 6043 9367
rect 7941 9333 7975 9367
rect 9689 9333 9723 9367
rect 10149 9333 10183 9367
rect 11621 9333 11655 9367
rect 12265 9333 12299 9367
rect 12771 9333 12805 9367
rect 13185 9333 13219 9367
rect 14013 9333 14047 9367
rect 14565 9333 14599 9367
rect 15577 9333 15611 9367
rect 16773 9333 16807 9367
rect 18337 9333 18371 9367
rect 20913 9333 20947 9367
rect 3525 9129 3559 9163
rect 4353 9129 4387 9163
rect 8401 9129 8435 9163
rect 10333 9129 10367 9163
rect 12909 9129 12943 9163
rect 14841 9129 14875 9163
rect 15669 9129 15703 9163
rect 16221 9129 16255 9163
rect 19165 9129 19199 9163
rect 21051 9129 21085 9163
rect 3157 9061 3191 9095
rect 4813 9061 4847 9095
rect 7802 9061 7836 9095
rect 9137 9061 9171 9095
rect 18061 9061 18095 9095
rect 1961 8993 1995 9027
rect 2329 8993 2363 9027
rect 2513 8993 2547 9027
rect 2973 8993 3007 9027
rect 5457 8993 5491 9027
rect 5641 8993 5675 9027
rect 6009 8993 6043 9027
rect 6377 8993 6411 9027
rect 9689 8993 9723 9027
rect 9836 8993 9870 9027
rect 11253 8993 11287 9027
rect 11529 8993 11563 9027
rect 11989 8993 12023 9027
rect 13921 8993 13955 9027
rect 14197 8993 14231 9027
rect 20980 8993 21014 9027
rect 3801 8925 3835 8959
rect 6653 8925 6687 8959
rect 7481 8925 7515 8959
rect 10057 8925 10091 8959
rect 14381 8925 14415 8959
rect 15301 8925 15335 8959
rect 17969 8925 18003 8959
rect 18613 8925 18647 8959
rect 11345 8857 11379 8891
rect 9505 8789 9539 8823
rect 9965 8789 9999 8823
rect 3985 8585 4019 8619
rect 4445 8585 4479 8619
rect 5549 8585 5583 8619
rect 6469 8585 6503 8619
rect 14657 8585 14691 8619
rect 17417 8585 17451 8619
rect 4813 8517 4847 8551
rect 9137 8517 9171 8551
rect 9505 8517 9539 8551
rect 10793 8517 10827 8551
rect 11115 8517 11149 8551
rect 19257 8517 19291 8551
rect 1777 8449 1811 8483
rect 3341 8449 3375 8483
rect 3801 8449 3835 8483
rect 5181 8449 5215 8483
rect 7113 8449 7147 8483
rect 8861 8449 8895 8483
rect 1961 8381 1995 8415
rect 2329 8381 2363 8415
rect 2697 8381 2731 8415
rect 3249 8381 3283 8415
rect 5457 8381 5491 8415
rect 7573 8381 7607 8415
rect 8217 8381 8251 8415
rect 3617 8313 3651 8347
rect 3801 8313 3835 8347
rect 5273 8313 5307 8347
rect 6193 8313 6227 8347
rect 9873 8449 9907 8483
rect 12725 8449 12759 8483
rect 13553 8449 13587 8483
rect 14933 8449 14967 8483
rect 15945 8449 15979 8483
rect 20177 8449 20211 8483
rect 9413 8381 9447 8415
rect 9689 8381 9723 8415
rect 11012 8381 11046 8415
rect 11805 8381 11839 8415
rect 13001 8381 13035 8415
rect 13369 8381 13403 8415
rect 16405 8381 16439 8415
rect 16865 8381 16899 8415
rect 17141 8381 17175 8415
rect 18061 8381 18095 8415
rect 9229 8313 9263 8347
rect 15025 8313 15059 8347
rect 15577 8313 15611 8347
rect 18382 8313 18416 8347
rect 19901 8313 19935 8347
rect 19993 8313 20027 8347
rect 7481 8245 7515 8279
rect 9137 8245 9171 8279
rect 10425 8245 10459 8279
rect 11437 8245 11471 8279
rect 13921 8245 13955 8279
rect 14289 8245 14323 8279
rect 16221 8245 16255 8279
rect 17785 8245 17819 8279
rect 18981 8245 19015 8279
rect 19625 8245 19659 8279
rect 21005 8245 21039 8279
rect 2329 8041 2363 8075
rect 3065 8041 3099 8075
rect 3525 8041 3559 8075
rect 7481 8041 7515 8075
rect 9413 8041 9447 8075
rect 9873 8041 9907 8075
rect 11621 8041 11655 8075
rect 13829 8041 13863 8075
rect 15025 8041 15059 8075
rect 15393 8041 15427 8075
rect 16497 8041 16531 8075
rect 18061 8041 18095 8075
rect 5365 7973 5399 8007
rect 5549 7973 5583 8007
rect 8585 7973 8619 8007
rect 18613 7973 18647 8007
rect 19165 7973 19199 8007
rect 2145 7905 2179 7939
rect 8493 7905 8527 7939
rect 10241 7905 10275 7939
rect 10388 7905 10422 7939
rect 11253 7905 11287 7939
rect 11805 7905 11839 7939
rect 12265 7905 12299 7939
rect 12909 7905 12943 7939
rect 15577 7905 15611 7939
rect 15853 7905 15887 7939
rect 16865 7905 16899 7939
rect 5917 7837 5951 7871
rect 10609 7837 10643 7871
rect 12449 7837 12483 7871
rect 13461 7837 13495 7871
rect 18521 7837 18555 7871
rect 20913 7837 20947 7871
rect 5825 7769 5859 7803
rect 10517 7769 10551 7803
rect 10885 7769 10919 7803
rect 1961 7701 1995 7735
rect 5687 7701 5721 7735
rect 6193 7701 6227 7735
rect 14381 7701 14415 7735
rect 17003 7701 17037 7735
rect 19441 7701 19475 7735
rect 19809 7701 19843 7735
rect 1593 7497 1627 7531
rect 2513 7497 2547 7531
rect 3617 7497 3651 7531
rect 3801 7497 3835 7531
rect 1409 7293 1443 7327
rect 5089 7497 5123 7531
rect 5273 7497 5307 7531
rect 6653 7497 6687 7531
rect 7481 7497 7515 7531
rect 8585 7497 8619 7531
rect 9413 7497 9447 7531
rect 11161 7497 11195 7531
rect 11897 7497 11931 7531
rect 14105 7497 14139 7531
rect 15669 7497 15703 7531
rect 15853 7497 15887 7531
rect 17877 7497 17911 7531
rect 18475 7497 18509 7531
rect 4261 7361 4295 7395
rect 4905 7361 4939 7395
rect 6285 7429 6319 7463
rect 13737 7429 13771 7463
rect 14381 7429 14415 7463
rect 15209 7429 15243 7463
rect 7941 7361 7975 7395
rect 9229 7361 9263 7395
rect 12449 7361 12483 7395
rect 5089 7293 5123 7327
rect 5549 7293 5583 7327
rect 5784 7293 5818 7327
rect 9597 7293 9631 7327
rect 9965 7293 9999 7327
rect 10057 7293 10091 7327
rect 16773 7429 16807 7463
rect 19165 7429 19199 7463
rect 15945 7361 15979 7395
rect 16221 7361 16255 7395
rect 18889 7361 18923 7395
rect 19901 7361 19935 7395
rect 18404 7293 18438 7327
rect 4353 7225 4387 7259
rect 5871 7225 5905 7259
rect 7021 7225 7055 7259
rect 7665 7225 7699 7259
rect 7757 7225 7791 7259
rect 12265 7225 12299 7259
rect 12811 7225 12845 7259
rect 14657 7225 14691 7259
rect 14749 7225 14783 7259
rect 15853 7225 15887 7259
rect 16313 7225 16347 7259
rect 19441 7225 19475 7259
rect 19533 7225 19567 7259
rect 2145 7157 2179 7191
rect 3801 7157 3835 7191
rect 4077 7157 4111 7191
rect 10793 7157 10827 7191
rect 11345 7157 11379 7191
rect 13369 7157 13403 7191
rect 17141 7157 17175 7191
rect 20913 7157 20947 7191
rect 1593 6953 1627 6987
rect 4997 6953 5031 6987
rect 5641 6953 5675 6987
rect 9965 6953 9999 6987
rect 11161 6953 11195 6987
rect 11805 6953 11839 6987
rect 12449 6953 12483 6987
rect 15577 6953 15611 6987
rect 21097 6953 21131 6987
rect 4439 6885 4473 6919
rect 6831 6885 6865 6919
rect 8769 6885 8803 6919
rect 10885 6885 10919 6919
rect 13001 6885 13035 6919
rect 16589 6885 16623 6919
rect 18613 6885 18647 6919
rect 2421 6817 2455 6851
rect 2881 6817 2915 6851
rect 8217 6817 8251 6851
rect 8401 6817 8435 6851
rect 10149 6817 10183 6851
rect 10425 6817 10459 6851
rect 15736 6817 15770 6851
rect 16748 6817 16782 6851
rect 20913 6817 20947 6851
rect 3157 6749 3191 6783
rect 4077 6749 4111 6783
rect 6469 6749 6503 6783
rect 12909 6749 12943 6783
rect 13553 6749 13587 6783
rect 18521 6749 18555 6783
rect 18797 6749 18831 6783
rect 10241 6681 10275 6715
rect 13921 6681 13955 6715
rect 18337 6681 18371 6715
rect 3433 6613 3467 6647
rect 7389 6613 7423 6647
rect 9321 6613 9355 6647
rect 14565 6613 14599 6647
rect 15807 6613 15841 6647
rect 16221 6613 16255 6647
rect 16819 6613 16853 6647
rect 19441 6613 19475 6647
rect 4629 6409 4663 6443
rect 5733 6409 5767 6443
rect 6561 6409 6595 6443
rect 7389 6409 7423 6443
rect 8585 6409 8619 6443
rect 10425 6409 10459 6443
rect 12173 6409 12207 6443
rect 14473 6409 14507 6443
rect 17141 6409 17175 6443
rect 18889 6409 18923 6443
rect 21465 6409 21499 6443
rect 9229 6341 9263 6375
rect 12587 6341 12621 6375
rect 1547 6273 1581 6307
rect 2973 6273 3007 6307
rect 3617 6273 3651 6307
rect 7573 6273 7607 6307
rect 8953 6273 8987 6307
rect 9413 6273 9447 6307
rect 13001 6273 13035 6307
rect 19441 6273 19475 6307
rect 1460 6205 1494 6239
rect 1869 6205 1903 6239
rect 9505 6205 9539 6239
rect 11012 6205 11046 6239
rect 11437 6205 11471 6239
rect 12516 6205 12550 6239
rect 13277 6205 13311 6239
rect 13461 6205 13495 6239
rect 13921 6205 13955 6239
rect 15060 6205 15094 6239
rect 15485 6205 15519 6239
rect 16129 6205 16163 6239
rect 16589 6205 16623 6239
rect 17969 6205 18003 6239
rect 18521 6205 18555 6239
rect 20672 6205 20706 6239
rect 3065 6137 3099 6171
rect 4813 6137 4847 6171
rect 4905 6137 4939 6171
rect 5457 6137 5491 6171
rect 7665 6137 7699 6171
rect 8217 6137 8251 6171
rect 10885 6137 10919 6171
rect 14197 6137 14231 6171
rect 16865 6137 16899 6171
rect 19165 6137 19199 6171
rect 19257 6137 19291 6171
rect 21097 6137 21131 6171
rect 2513 6069 2547 6103
rect 4077 6069 4111 6103
rect 6101 6069 6135 6103
rect 11115 6069 11149 6103
rect 15301 6069 15335 6103
rect 15945 6069 15979 6103
rect 18199 6069 18233 6103
rect 20177 6069 20211 6103
rect 20775 6069 20809 6103
rect 3433 5865 3467 5899
rect 4169 5865 4203 5899
rect 5549 5865 5583 5899
rect 6101 5865 6135 5899
rect 7665 5865 7699 5899
rect 10793 5865 10827 5899
rect 14197 5865 14231 5899
rect 16681 5865 16715 5899
rect 18521 5865 18555 5899
rect 21051 5865 21085 5899
rect 5273 5797 5307 5831
rect 8217 5797 8251 5831
rect 13093 5797 13127 5831
rect 15485 5797 15519 5831
rect 17227 5797 17261 5831
rect 18889 5797 18923 5831
rect 3008 5729 3042 5763
rect 3111 5729 3145 5763
rect 4353 5729 4387 5763
rect 4629 5729 4663 5763
rect 6101 5729 6135 5763
rect 6285 5729 6319 5763
rect 10057 5729 10091 5763
rect 10333 5729 10367 5763
rect 11345 5729 11379 5763
rect 11897 5729 11931 5763
rect 16865 5729 16899 5763
rect 20980 5729 21014 5763
rect 8125 5661 8159 5695
rect 8401 5661 8435 5695
rect 10425 5661 10459 5695
rect 12081 5661 12115 5695
rect 13001 5661 13035 5695
rect 13277 5661 13311 5695
rect 15393 5661 15427 5695
rect 16037 5661 16071 5695
rect 18797 5661 18831 5695
rect 16313 5593 16347 5627
rect 19349 5593 19383 5627
rect 2513 5525 2547 5559
rect 7297 5525 7331 5559
rect 11161 5525 11195 5559
rect 17785 5525 17819 5559
rect 3525 5321 3559 5355
rect 4261 5321 4295 5355
rect 6193 5321 6227 5355
rect 7113 5321 7147 5355
rect 8493 5321 8527 5355
rect 9873 5321 9907 5355
rect 11713 5321 11747 5355
rect 12265 5321 12299 5355
rect 13369 5321 13403 5355
rect 13645 5321 13679 5355
rect 18521 5321 18555 5355
rect 19625 5321 19659 5355
rect 3801 5253 3835 5287
rect 14013 5253 14047 5287
rect 19257 5253 19291 5287
rect 2145 5185 2179 5219
rect 2605 5185 2639 5219
rect 5917 5185 5951 5219
rect 7297 5185 7331 5219
rect 10425 5185 10459 5219
rect 12449 5185 12483 5219
rect 14197 5185 14231 5219
rect 16313 5185 16347 5219
rect 16589 5185 16623 5219
rect 18705 5185 18739 5219
rect 19993 5185 20027 5219
rect 20637 5185 20671 5219
rect 5089 5117 5123 5151
rect 5457 5117 5491 5151
rect 5733 5117 5767 5151
rect 8217 5117 8251 5151
rect 20228 5117 20262 5151
rect 21224 5117 21258 5151
rect 21649 5117 21683 5151
rect 2926 5049 2960 5083
rect 7659 5049 7693 5083
rect 9045 5049 9079 5083
rect 10333 5049 10367 5083
rect 10787 5049 10821 5083
rect 12770 5049 12804 5083
rect 14518 5049 14552 5083
rect 16129 5049 16163 5083
rect 16405 5049 16439 5083
rect 17877 5049 17911 5083
rect 18797 5049 18831 5083
rect 20315 5049 20349 5083
rect 21327 5049 21361 5083
rect 2421 4981 2455 5015
rect 4537 4981 4571 5015
rect 6653 4981 6687 5015
rect 8861 4981 8895 5015
rect 11345 4981 11379 5015
rect 15117 4981 15151 5015
rect 15485 4981 15519 5015
rect 17325 4981 17359 5015
rect 21097 4981 21131 5015
rect 3433 4777 3467 4811
rect 7757 4777 7791 4811
rect 8309 4777 8343 4811
rect 8585 4777 8619 4811
rect 10701 4777 10735 4811
rect 12449 4777 12483 4811
rect 12909 4777 12943 4811
rect 13231 4777 13265 4811
rect 15117 4777 15151 4811
rect 15393 4777 15427 4811
rect 16773 4777 16807 4811
rect 3157 4709 3191 4743
rect 11437 4709 11471 4743
rect 18797 4709 18831 4743
rect 19349 4709 19383 4743
rect 2421 4641 2455 4675
rect 2697 4641 2731 4675
rect 4353 4641 4387 4675
rect 6101 4641 6135 4675
rect 6285 4641 6319 4675
rect 9781 4641 9815 4675
rect 10149 4641 10183 4675
rect 13160 4641 13194 4675
rect 14105 4641 14139 4675
rect 15485 4641 15519 4675
rect 15853 4641 15887 4675
rect 17049 4641 17083 4675
rect 17325 4641 17359 4675
rect 20948 4641 20982 4675
rect 4261 4573 4295 4607
rect 6561 4573 6595 4607
rect 7389 4573 7423 4607
rect 10241 4573 10275 4607
rect 11345 4573 11379 4607
rect 11989 4573 12023 4607
rect 17601 4573 17635 4607
rect 18521 4573 18555 4607
rect 18705 4573 18739 4607
rect 21051 4573 21085 4607
rect 2513 4505 2547 4539
rect 14289 4505 14323 4539
rect 1685 4437 1719 4471
rect 5273 4437 5307 4471
rect 7297 4437 7331 4471
rect 9045 4437 9079 4471
rect 14657 4437 14691 4471
rect 16313 4437 16347 4471
rect 1593 4233 1627 4267
rect 6561 4233 6595 4267
rect 11253 4233 11287 4267
rect 13461 4233 13495 4267
rect 14105 4233 14139 4267
rect 15577 4233 15611 4267
rect 17141 4233 17175 4267
rect 19257 4233 19291 4267
rect 21511 4233 21545 4267
rect 5825 4165 5859 4199
rect 7481 4165 7515 4199
rect 7757 4165 7791 4199
rect 9229 4165 9263 4199
rect 10885 4165 10919 4199
rect 17417 4165 17451 4199
rect 20913 4165 20947 4199
rect 2145 4097 2179 4131
rect 3341 4097 3375 4131
rect 3985 4097 4019 4131
rect 8953 4097 8987 4131
rect 9689 4097 9723 4131
rect 16773 4097 16807 4131
rect 18061 4097 18095 4131
rect 20177 4097 20211 4131
rect 1409 4029 1443 4063
rect 3249 4029 3283 4063
rect 3525 4029 3559 4063
rect 4813 4029 4847 4063
rect 4905 4029 4939 4063
rect 5089 4029 5123 4063
rect 6837 4029 6871 4063
rect 9965 4029 9999 4063
rect 10241 4029 10275 4063
rect 11380 4029 11414 4063
rect 11805 4029 11839 4063
rect 12173 4029 12207 4063
rect 12449 4029 12483 4063
rect 12909 4029 12943 4063
rect 21408 4029 21442 4063
rect 3157 3961 3191 3995
rect 4721 3961 4755 3995
rect 5549 3961 5583 3995
rect 8309 3961 8343 3995
rect 8401 3961 8435 3995
rect 14565 3961 14599 3995
rect 14657 3961 14691 3995
rect 15209 3961 15243 3995
rect 16129 3961 16163 3995
rect 16221 3961 16255 3995
rect 19901 3961 19935 3995
rect 19993 3961 20027 3995
rect 2421 3893 2455 3927
rect 4353 3893 4387 3927
rect 6285 3893 6319 3927
rect 7021 3893 7055 3927
rect 9873 3893 9907 3927
rect 11483 3893 11517 3927
rect 12541 3893 12575 3927
rect 15853 3893 15887 3927
rect 17877 3893 17911 3927
rect 18429 3893 18463 3927
rect 18981 3893 19015 3927
rect 19625 3893 19659 3927
rect 21833 3893 21867 3927
rect 2513 3689 2547 3723
rect 3433 3689 3467 3723
rect 5273 3689 5307 3723
rect 6469 3689 6503 3723
rect 7757 3689 7791 3723
rect 9321 3689 9355 3723
rect 11253 3689 11287 3723
rect 12449 3689 12483 3723
rect 14565 3689 14599 3723
rect 16221 3689 16255 3723
rect 18061 3689 18095 3723
rect 19901 3689 19935 3723
rect 8677 3621 8711 3655
rect 10333 3621 10367 3655
rect 13093 3621 13127 3655
rect 15663 3621 15697 3655
rect 16497 3621 16531 3655
rect 18705 3621 18739 3655
rect 1409 3553 1443 3587
rect 2973 3553 3007 3587
rect 4905 3553 4939 3587
rect 6561 3553 6595 3587
rect 6837 3553 6871 3587
rect 7941 3553 7975 3587
rect 8217 3553 8251 3587
rect 9873 3553 9907 3587
rect 11805 3553 11839 3587
rect 15301 3553 15335 3587
rect 17049 3553 17083 3587
rect 17601 3553 17635 3587
rect 20980 3553 21014 3587
rect 3111 3485 3145 3519
rect 10241 3485 10275 3519
rect 13001 3485 13035 3519
rect 13921 3485 13955 3519
rect 18613 3485 18647 3519
rect 18981 3485 19015 3519
rect 8033 3417 8067 3451
rect 10793 3417 10827 3451
rect 13553 3417 13587 3451
rect 1593 3349 1627 3383
rect 4721 3349 4755 3383
rect 11713 3349 11747 3383
rect 11989 3349 12023 3383
rect 17233 3349 17267 3383
rect 21051 3349 21085 3383
rect 1685 3145 1719 3179
rect 3249 3145 3283 3179
rect 6377 3145 6411 3179
rect 10057 3145 10091 3179
rect 13369 3145 13403 3179
rect 15117 3145 15151 3179
rect 15761 3145 15795 3179
rect 18429 3145 18463 3179
rect 19901 3145 19935 3179
rect 4721 3077 4755 3111
rect 8677 3077 8711 3111
rect 10517 3077 10551 3111
rect 19533 3077 19567 3111
rect 5365 3009 5399 3043
rect 7113 3009 7147 3043
rect 7757 3009 7791 3043
rect 8401 3009 8435 3043
rect 10609 3009 10643 3043
rect 11897 3009 11931 3043
rect 12449 3009 12483 3043
rect 14013 3009 14047 3043
rect 18889 3009 18923 3043
rect 2697 2941 2731 2975
rect 3065 2941 3099 2975
rect 4445 2941 4479 2975
rect 4629 2941 4663 2975
rect 4905 2941 4939 2975
rect 9229 2941 9263 2975
rect 12173 2941 12207 2975
rect 14197 2941 14231 2975
rect 16221 2941 16255 2975
rect 16405 2941 16439 2975
rect 20085 2941 20119 2975
rect 20545 2941 20579 2975
rect 2513 2873 2547 2907
rect 7849 2873 7883 2907
rect 9045 2873 9079 2907
rect 10930 2873 10964 2907
rect 12770 2873 12804 2907
rect 13737 2873 13771 2907
rect 14518 2873 14552 2907
rect 15485 2873 15519 2907
rect 16957 2873 16991 2907
rect 17509 2873 17543 2907
rect 18613 2873 18647 2907
rect 18705 2873 18739 2907
rect 2697 2805 2731 2839
rect 2789 2805 2823 2839
rect 4169 2805 4203 2839
rect 5733 2805 5767 2839
rect 7573 2805 7607 2839
rect 9413 2805 9447 2839
rect 11529 2805 11563 2839
rect 16037 2805 16071 2839
rect 17877 2805 17911 2839
rect 20177 2805 20211 2839
rect 21189 2805 21223 2839
rect 3525 2601 3559 2635
rect 4353 2601 4387 2635
rect 6377 2601 6411 2635
rect 7941 2601 7975 2635
rect 10701 2601 10735 2635
rect 10977 2601 11011 2635
rect 11345 2601 11379 2635
rect 11667 2601 11701 2635
rect 12357 2601 12391 2635
rect 13645 2601 13679 2635
rect 15301 2601 15335 2635
rect 17417 2601 17451 2635
rect 5825 2533 5859 2567
rect 6653 2533 6687 2567
rect 7342 2533 7376 2567
rect 9505 2533 9539 2567
rect 10143 2533 10177 2567
rect 12817 2533 12851 2567
rect 15623 2533 15657 2567
rect 16405 2533 16439 2567
rect 16859 2533 16893 2567
rect 17785 2533 17819 2567
rect 18153 2533 18187 2567
rect 19073 2533 19107 2567
rect 19165 2533 19199 2567
rect 20085 2533 20119 2567
rect 1409 2465 1443 2499
rect 2881 2465 2915 2499
rect 4445 2465 4479 2499
rect 4721 2465 4755 2499
rect 5181 2465 5215 2499
rect 7021 2465 7055 2499
rect 9229 2465 9263 2499
rect 9781 2465 9815 2499
rect 11564 2465 11598 2499
rect 11989 2465 12023 2499
rect 14197 2465 14231 2499
rect 15520 2465 15554 2499
rect 15945 2465 15979 2499
rect 16497 2465 16531 2499
rect 21189 2465 21223 2499
rect 21741 2465 21775 2499
rect 2053 2397 2087 2431
rect 3893 2397 3927 2431
rect 5457 2397 5491 2431
rect 12725 2397 12759 2431
rect 14013 2397 14047 2431
rect 18797 2397 18831 2431
rect 19349 2397 19383 2431
rect 3065 2329 3099 2363
rect 4537 2329 4571 2363
rect 13277 2329 13311 2363
rect 14381 2329 14415 2363
rect 14841 2329 14875 2363
rect 21373 2329 21407 2363
rect 1593 2261 1627 2295
rect 8309 2261 8343 2295
<< metal1 >>
rect 22094 23536 22100 23588
rect 22152 23576 22158 23588
rect 23290 23576 23296 23588
rect 22152 23548 23296 23576
rect 22152 23536 22158 23548
rect 23290 23536 23296 23548
rect 23348 23536 23354 23588
rect 1104 21786 22816 21808
rect 1104 21734 4982 21786
rect 5034 21734 5046 21786
rect 5098 21734 5110 21786
rect 5162 21734 5174 21786
rect 5226 21734 12982 21786
rect 13034 21734 13046 21786
rect 13098 21734 13110 21786
rect 13162 21734 13174 21786
rect 13226 21734 20982 21786
rect 21034 21734 21046 21786
rect 21098 21734 21110 21786
rect 21162 21734 21174 21786
rect 21226 21734 22816 21786
rect 1104 21712 22816 21734
rect 1104 21242 22816 21264
rect 1104 21190 8982 21242
rect 9034 21190 9046 21242
rect 9098 21190 9110 21242
rect 9162 21190 9174 21242
rect 9226 21190 16982 21242
rect 17034 21190 17046 21242
rect 17098 21190 17110 21242
rect 17162 21190 17174 21242
rect 17226 21190 22816 21242
rect 1104 21168 22816 21190
rect 566 21088 572 21140
rect 624 21128 630 21140
rect 6454 21128 6460 21140
rect 624 21100 6460 21128
rect 624 21088 630 21100
rect 6454 21088 6460 21100
rect 6512 21088 6518 21140
rect 10505 21131 10563 21137
rect 10505 21097 10517 21131
rect 10551 21128 10563 21131
rect 11422 21128 11428 21140
rect 10551 21100 11428 21128
rect 10551 21097 10563 21100
rect 10505 21091 10563 21097
rect 11422 21088 11428 21100
rect 11480 21088 11486 21140
rect 10321 20995 10379 21001
rect 10321 20961 10333 20995
rect 10367 20992 10379 20995
rect 11054 20992 11060 21004
rect 10367 20964 11060 20992
rect 10367 20961 10379 20964
rect 10321 20955 10379 20961
rect 11054 20952 11060 20964
rect 11112 20952 11118 21004
rect 13792 20995 13850 21001
rect 13792 20961 13804 20995
rect 13838 20992 13850 20995
rect 15010 20992 15016 21004
rect 13838 20964 15016 20992
rect 13838 20961 13850 20964
rect 13792 20955 13850 20961
rect 15010 20952 15016 20964
rect 15068 20952 15074 21004
rect 8662 20788 8668 20800
rect 8623 20760 8668 20788
rect 8662 20748 8668 20760
rect 8720 20748 8726 20800
rect 13722 20748 13728 20800
rect 13780 20788 13786 20800
rect 13863 20791 13921 20797
rect 13863 20788 13875 20791
rect 13780 20760 13875 20788
rect 13780 20748 13786 20760
rect 13863 20757 13875 20760
rect 13909 20757 13921 20791
rect 13863 20751 13921 20757
rect 1104 20698 22816 20720
rect 1104 20646 4982 20698
rect 5034 20646 5046 20698
rect 5098 20646 5110 20698
rect 5162 20646 5174 20698
rect 5226 20646 12982 20698
rect 13034 20646 13046 20698
rect 13098 20646 13110 20698
rect 13162 20646 13174 20698
rect 13226 20646 20982 20698
rect 21034 20646 21046 20698
rect 21098 20646 21110 20698
rect 21162 20646 21174 20698
rect 21226 20646 22816 20698
rect 1104 20624 22816 20646
rect 3789 20587 3847 20593
rect 3789 20553 3801 20587
rect 3835 20584 3847 20587
rect 4338 20584 4344 20596
rect 3835 20556 4344 20584
rect 3835 20553 3847 20556
rect 3789 20547 3847 20553
rect 4338 20544 4344 20556
rect 4396 20544 4402 20596
rect 8113 20587 8171 20593
rect 8113 20553 8125 20587
rect 8159 20584 8171 20587
rect 8386 20584 8392 20596
rect 8159 20556 8392 20584
rect 8159 20553 8171 20556
rect 8113 20547 8171 20553
rect 1464 20383 1522 20389
rect 1464 20349 1476 20383
rect 1510 20380 1522 20383
rect 1854 20380 1860 20392
rect 1510 20352 1860 20380
rect 1510 20349 1522 20352
rect 1464 20343 1522 20349
rect 1854 20340 1860 20352
rect 1912 20340 1918 20392
rect 2222 20340 2228 20392
rect 2280 20380 2286 20392
rect 2536 20383 2594 20389
rect 2536 20380 2548 20383
rect 2280 20352 2548 20380
rect 2280 20340 2286 20352
rect 2536 20349 2548 20352
rect 2582 20380 2594 20383
rect 2961 20383 3019 20389
rect 2961 20380 2973 20383
rect 2582 20352 2973 20380
rect 2582 20349 2594 20352
rect 2536 20343 2594 20349
rect 2961 20349 2973 20352
rect 3007 20349 3019 20383
rect 2961 20343 3019 20349
rect 3605 20383 3663 20389
rect 3605 20349 3617 20383
rect 3651 20380 3663 20383
rect 3694 20380 3700 20392
rect 3651 20352 3700 20380
rect 3651 20349 3663 20352
rect 3605 20343 3663 20349
rect 3694 20340 3700 20352
rect 3752 20340 3758 20392
rect 7628 20383 7686 20389
rect 7628 20349 7640 20383
rect 7674 20380 7686 20383
rect 8128 20380 8156 20547
rect 8386 20544 8392 20556
rect 8444 20544 8450 20596
rect 10134 20544 10140 20596
rect 10192 20584 10198 20596
rect 10321 20587 10379 20593
rect 10321 20584 10333 20587
rect 10192 20556 10333 20584
rect 10192 20544 10198 20556
rect 10321 20553 10333 20556
rect 10367 20553 10379 20587
rect 14090 20584 14096 20596
rect 14051 20556 14096 20584
rect 10321 20547 10379 20553
rect 14090 20544 14096 20556
rect 14148 20544 14154 20596
rect 14461 20587 14519 20593
rect 14461 20553 14473 20587
rect 14507 20584 14519 20587
rect 15010 20584 15016 20596
rect 14507 20556 15016 20584
rect 14507 20553 14519 20556
rect 14461 20547 14519 20553
rect 15010 20544 15016 20556
rect 15068 20544 15074 20596
rect 15657 20587 15715 20593
rect 15657 20553 15669 20587
rect 15703 20584 15715 20587
rect 16390 20584 16396 20596
rect 15703 20556 16396 20584
rect 15703 20553 15715 20556
rect 15657 20547 15715 20553
rect 8662 20448 8668 20460
rect 8623 20420 8668 20448
rect 8662 20408 8668 20420
rect 8720 20408 8726 20460
rect 10137 20383 10195 20389
rect 10137 20380 10149 20383
rect 7674 20352 8156 20380
rect 9416 20352 10149 20380
rect 7674 20349 7686 20352
rect 7628 20343 7686 20349
rect 6454 20272 6460 20324
rect 6512 20312 6518 20324
rect 8481 20315 8539 20321
rect 6512 20284 8386 20312
rect 6512 20272 6518 20284
rect 1535 20247 1593 20253
rect 1535 20213 1547 20247
rect 1581 20244 1593 20247
rect 2498 20244 2504 20256
rect 1581 20216 2504 20244
rect 1581 20213 1593 20216
rect 1535 20207 1593 20213
rect 2498 20204 2504 20216
rect 2556 20204 2562 20256
rect 2639 20247 2697 20253
rect 2639 20213 2651 20247
rect 2685 20244 2697 20247
rect 2774 20244 2780 20256
rect 2685 20216 2780 20244
rect 2685 20213 2697 20216
rect 2639 20207 2697 20213
rect 2774 20204 2780 20216
rect 2832 20204 2838 20256
rect 3694 20204 3700 20256
rect 3752 20244 3758 20256
rect 4249 20247 4307 20253
rect 4249 20244 4261 20247
rect 3752 20216 4261 20244
rect 3752 20204 3758 20216
rect 4249 20213 4261 20216
rect 4295 20244 4307 20247
rect 7374 20244 7380 20256
rect 4295 20216 7380 20244
rect 4295 20213 4307 20216
rect 4249 20207 4307 20213
rect 7374 20204 7380 20216
rect 7432 20204 7438 20256
rect 7699 20247 7757 20253
rect 7699 20213 7711 20247
rect 7745 20244 7757 20247
rect 7834 20244 7840 20256
rect 7745 20216 7840 20244
rect 7745 20213 7757 20216
rect 7699 20207 7757 20213
rect 7834 20204 7840 20216
rect 7892 20204 7898 20256
rect 8358 20244 8386 20284
rect 8481 20281 8493 20315
rect 8527 20312 8539 20315
rect 8754 20312 8760 20324
rect 8527 20284 8760 20312
rect 8527 20281 8539 20284
rect 8481 20275 8539 20281
rect 8754 20272 8760 20284
rect 8812 20272 8818 20324
rect 9306 20312 9312 20324
rect 9267 20284 9312 20312
rect 9306 20272 9312 20284
rect 9364 20272 9370 20324
rect 9416 20244 9444 20352
rect 10137 20349 10149 20352
rect 10183 20380 10195 20383
rect 10689 20383 10747 20389
rect 10689 20380 10701 20383
rect 10183 20352 10701 20380
rect 10183 20349 10195 20352
rect 10137 20343 10195 20349
rect 10689 20349 10701 20352
rect 10735 20349 10747 20383
rect 10689 20343 10747 20349
rect 13608 20383 13666 20389
rect 13608 20349 13620 20383
rect 13654 20380 13666 20383
rect 14090 20380 14096 20392
rect 13654 20352 14096 20380
rect 13654 20349 13666 20352
rect 13608 20343 13666 20349
rect 14090 20340 14096 20352
rect 14148 20340 14154 20392
rect 15172 20383 15230 20389
rect 15172 20349 15184 20383
rect 15218 20380 15230 20383
rect 15672 20380 15700 20547
rect 16390 20544 16396 20556
rect 16448 20544 16454 20596
rect 18877 20587 18935 20593
rect 18877 20553 18889 20587
rect 18923 20584 18935 20587
rect 19058 20584 19064 20596
rect 18923 20556 19064 20584
rect 18923 20553 18935 20556
rect 18877 20547 18935 20553
rect 15218 20352 15700 20380
rect 18392 20383 18450 20389
rect 15218 20349 15230 20352
rect 15172 20343 15230 20349
rect 18392 20349 18404 20383
rect 18438 20380 18450 20383
rect 18892 20380 18920 20547
rect 19058 20544 19064 20556
rect 19116 20544 19122 20596
rect 21450 20584 21456 20596
rect 21411 20556 21456 20584
rect 21450 20544 21456 20556
rect 21508 20544 21514 20596
rect 18438 20352 18920 20380
rect 20968 20383 21026 20389
rect 18438 20349 18450 20352
rect 18392 20343 18450 20349
rect 20968 20349 20980 20383
rect 21014 20380 21026 20383
rect 21450 20380 21456 20392
rect 21014 20352 21456 20380
rect 21014 20349 21026 20352
rect 20968 20343 21026 20349
rect 21450 20340 21456 20352
rect 21508 20340 21514 20392
rect 11054 20244 11060 20256
rect 8358 20216 9444 20244
rect 11015 20216 11060 20244
rect 11054 20204 11060 20216
rect 11112 20204 11118 20256
rect 13679 20247 13737 20253
rect 13679 20213 13691 20247
rect 13725 20244 13737 20247
rect 13814 20244 13820 20256
rect 13725 20216 13820 20244
rect 13725 20213 13737 20216
rect 13679 20207 13737 20213
rect 13814 20204 13820 20216
rect 13872 20204 13878 20256
rect 15243 20247 15301 20253
rect 15243 20213 15255 20247
rect 15289 20244 15301 20247
rect 15378 20244 15384 20256
rect 15289 20216 15384 20244
rect 15289 20213 15301 20216
rect 15243 20207 15301 20213
rect 15378 20204 15384 20216
rect 15436 20204 15442 20256
rect 18463 20247 18521 20253
rect 18463 20213 18475 20247
rect 18509 20244 18521 20247
rect 18598 20244 18604 20256
rect 18509 20216 18604 20244
rect 18509 20213 18521 20216
rect 18463 20207 18521 20213
rect 18598 20204 18604 20216
rect 18656 20204 18662 20256
rect 18690 20204 18696 20256
rect 18748 20244 18754 20256
rect 21039 20247 21097 20253
rect 21039 20244 21051 20247
rect 18748 20216 21051 20244
rect 18748 20204 18754 20216
rect 21039 20213 21051 20216
rect 21085 20213 21097 20247
rect 21039 20207 21097 20213
rect 1104 20154 22816 20176
rect 1104 20102 8982 20154
rect 9034 20102 9046 20154
rect 9098 20102 9110 20154
rect 9162 20102 9174 20154
rect 9226 20102 16982 20154
rect 17034 20102 17046 20154
rect 17098 20102 17110 20154
rect 17162 20102 17174 20154
rect 17226 20102 22816 20154
rect 1104 20080 22816 20102
rect 1578 20040 1584 20052
rect 1539 20012 1584 20040
rect 1578 20000 1584 20012
rect 1636 20000 1642 20052
rect 7607 20043 7665 20049
rect 7607 20009 7619 20043
rect 7653 20040 7665 20043
rect 8662 20040 8668 20052
rect 7653 20012 8668 20040
rect 7653 20009 7665 20012
rect 7607 20003 7665 20009
rect 8662 20000 8668 20012
rect 8720 20000 8726 20052
rect 13538 20000 13544 20052
rect 13596 20000 13602 20052
rect 106 19932 112 19984
rect 164 19972 170 19984
rect 164 19944 8559 19972
rect 164 19932 170 19944
rect 8531 19916 8559 19944
rect 8754 19932 8760 19984
rect 8812 19972 8818 19984
rect 9766 19972 9772 19984
rect 8812 19944 9772 19972
rect 8812 19932 8818 19944
rect 9766 19932 9772 19944
rect 9824 19972 9830 19984
rect 10045 19975 10103 19981
rect 10045 19972 10057 19975
rect 9824 19944 10057 19972
rect 9824 19932 9830 19944
rect 10045 19941 10057 19944
rect 10091 19941 10103 19975
rect 13556 19972 13584 20000
rect 13718 19975 13776 19981
rect 13718 19972 13730 19975
rect 13556 19944 13730 19972
rect 10045 19935 10103 19941
rect 13718 19941 13730 19944
rect 13764 19941 13776 19975
rect 15470 19972 15476 19984
rect 15431 19944 15476 19972
rect 13718 19935 13776 19941
rect 15470 19932 15476 19944
rect 15528 19932 15534 19984
rect 2130 19913 2136 19916
rect 2108 19907 2136 19913
rect 2108 19904 2120 19907
rect 2043 19876 2120 19904
rect 2108 19873 2120 19876
rect 2188 19904 2194 19916
rect 3050 19904 3056 19916
rect 2188 19876 3056 19904
rect 2108 19867 2136 19873
rect 2130 19864 2136 19867
rect 2188 19864 2194 19876
rect 3050 19864 3056 19876
rect 3108 19864 3114 19916
rect 7374 19904 7380 19916
rect 7335 19876 7380 19904
rect 7374 19864 7380 19876
rect 7432 19864 7438 19916
rect 8478 19904 8484 19916
rect 8536 19913 8559 19916
rect 8536 19907 8574 19913
rect 8426 19876 8484 19904
rect 8478 19864 8484 19876
rect 8562 19873 8574 19907
rect 8536 19867 8574 19873
rect 12596 19907 12654 19913
rect 12596 19873 12608 19907
rect 12642 19904 12654 19907
rect 12710 19904 12716 19916
rect 12642 19876 12716 19904
rect 12642 19873 12654 19876
rect 12596 19867 12654 19873
rect 8536 19864 8542 19867
rect 12710 19864 12716 19876
rect 12768 19864 12774 19916
rect 16942 19913 16948 19916
rect 16920 19907 16948 19913
rect 16920 19904 16932 19907
rect 16855 19876 16932 19904
rect 16920 19873 16932 19876
rect 17000 19904 17006 19916
rect 17678 19904 17684 19916
rect 17000 19876 17684 19904
rect 16920 19867 16948 19873
rect 16942 19864 16948 19867
rect 17000 19864 17006 19876
rect 17678 19864 17684 19876
rect 17736 19864 17742 19916
rect 20968 19907 21026 19913
rect 20968 19873 20980 19907
rect 21014 19904 21026 19907
rect 21174 19904 21180 19916
rect 21014 19876 21180 19904
rect 21014 19873 21026 19876
rect 20968 19867 21026 19873
rect 21174 19864 21180 19876
rect 21232 19864 21238 19916
rect 9950 19836 9956 19848
rect 9911 19808 9956 19836
rect 9950 19796 9956 19808
rect 10008 19796 10014 19848
rect 10134 19796 10140 19848
rect 10192 19836 10198 19848
rect 10229 19839 10287 19845
rect 10229 19836 10241 19839
rect 10192 19808 10241 19836
rect 10192 19796 10198 19808
rect 10229 19805 10241 19808
rect 10275 19805 10287 19839
rect 10229 19799 10287 19805
rect 10410 19796 10416 19848
rect 10468 19836 10474 19848
rect 11425 19839 11483 19845
rect 11425 19836 11437 19839
rect 10468 19808 11437 19836
rect 10468 19796 10474 19808
rect 11425 19805 11437 19808
rect 11471 19805 11483 19839
rect 11425 19799 11483 19805
rect 13449 19839 13507 19845
rect 13449 19805 13461 19839
rect 13495 19836 13507 19839
rect 13633 19839 13691 19845
rect 13633 19836 13645 19839
rect 13495 19808 13645 19836
rect 13495 19805 13507 19808
rect 13449 19799 13507 19805
rect 13633 19805 13645 19808
rect 13679 19836 13691 19839
rect 13722 19836 13728 19848
rect 13679 19808 13728 19836
rect 13679 19805 13691 19808
rect 13633 19799 13691 19805
rect 13722 19796 13728 19808
rect 13780 19796 13786 19848
rect 14274 19836 14280 19848
rect 14235 19808 14280 19836
rect 14274 19796 14280 19808
rect 14332 19796 14338 19848
rect 15378 19836 15384 19848
rect 15339 19808 15384 19836
rect 15378 19796 15384 19808
rect 15436 19796 15442 19848
rect 15657 19839 15715 19845
rect 15657 19805 15669 19839
rect 15703 19805 15715 19839
rect 15657 19799 15715 19805
rect 14292 19768 14320 19796
rect 15672 19768 15700 19799
rect 14292 19740 15700 19768
rect 2038 19660 2044 19712
rect 2096 19700 2102 19712
rect 2179 19703 2237 19709
rect 2179 19700 2191 19703
rect 2096 19672 2191 19700
rect 2096 19660 2102 19672
rect 2179 19669 2191 19672
rect 2225 19669 2237 19703
rect 6822 19700 6828 19712
rect 6783 19672 6828 19700
rect 2179 19663 2237 19669
rect 6822 19660 6828 19672
rect 6880 19660 6886 19712
rect 8619 19703 8677 19709
rect 8619 19669 8631 19703
rect 8665 19700 8677 19703
rect 8846 19700 8852 19712
rect 8665 19672 8852 19700
rect 8665 19669 8677 19672
rect 8619 19663 8677 19669
rect 8846 19660 8852 19672
rect 8904 19700 8910 19712
rect 8941 19703 8999 19709
rect 8941 19700 8953 19703
rect 8904 19672 8953 19700
rect 8904 19660 8910 19672
rect 8941 19669 8953 19672
rect 8987 19669 8999 19703
rect 8941 19663 8999 19669
rect 12667 19703 12725 19709
rect 12667 19669 12679 19703
rect 12713 19700 12725 19703
rect 13354 19700 13360 19712
rect 12713 19672 13360 19700
rect 12713 19669 12725 19672
rect 12667 19663 12725 19669
rect 13354 19660 13360 19672
rect 13412 19660 13418 19712
rect 16850 19660 16856 19712
rect 16908 19700 16914 19712
rect 16991 19703 17049 19709
rect 16991 19700 17003 19703
rect 16908 19672 17003 19700
rect 16908 19660 16914 19672
rect 16991 19669 17003 19672
rect 17037 19669 17049 19703
rect 16991 19663 17049 19669
rect 17402 19660 17408 19712
rect 17460 19700 17466 19712
rect 21039 19703 21097 19709
rect 21039 19700 21051 19703
rect 17460 19672 21051 19700
rect 17460 19660 17466 19672
rect 21039 19669 21051 19672
rect 21085 19669 21097 19703
rect 21039 19663 21097 19669
rect 1104 19610 22816 19632
rect 1104 19558 4982 19610
rect 5034 19558 5046 19610
rect 5098 19558 5110 19610
rect 5162 19558 5174 19610
rect 5226 19558 12982 19610
rect 13034 19558 13046 19610
rect 13098 19558 13110 19610
rect 13162 19558 13174 19610
rect 13226 19558 20982 19610
rect 21034 19558 21046 19610
rect 21098 19558 21110 19610
rect 21162 19558 21174 19610
rect 21226 19558 22816 19610
rect 1104 19536 22816 19558
rect 2130 19496 2136 19508
rect 2091 19468 2136 19496
rect 2130 19456 2136 19468
rect 2188 19456 2194 19508
rect 7374 19456 7380 19508
rect 7432 19496 7438 19508
rect 7837 19499 7895 19505
rect 7837 19496 7849 19499
rect 7432 19468 7849 19496
rect 7432 19456 7438 19468
rect 7837 19465 7849 19468
rect 7883 19465 7895 19499
rect 8478 19496 8484 19508
rect 8439 19468 8484 19496
rect 7837 19459 7895 19465
rect 8478 19456 8484 19468
rect 8536 19456 8542 19508
rect 9766 19496 9772 19508
rect 9727 19468 9772 19496
rect 9766 19456 9772 19468
rect 9824 19456 9830 19508
rect 15378 19456 15384 19508
rect 15436 19496 15442 19508
rect 16393 19499 16451 19505
rect 16393 19496 16405 19499
rect 15436 19468 16405 19496
rect 15436 19456 15442 19468
rect 16393 19465 16405 19468
rect 16439 19465 16451 19499
rect 16942 19496 16948 19508
rect 16903 19468 16948 19496
rect 16393 19459 16451 19465
rect 16942 19456 16948 19468
rect 17000 19456 17006 19508
rect 19245 19499 19303 19505
rect 19245 19465 19257 19499
rect 19291 19496 19303 19499
rect 20714 19496 20720 19508
rect 19291 19468 20720 19496
rect 19291 19465 19303 19468
rect 19245 19459 19303 19465
rect 6641 19431 6699 19437
rect 6641 19397 6653 19431
rect 6687 19428 6699 19431
rect 7006 19428 7012 19440
rect 6687 19400 7012 19428
rect 6687 19397 6699 19400
rect 6641 19391 6699 19397
rect 7006 19388 7012 19400
rect 7064 19388 7070 19440
rect 10152 19400 10732 19428
rect 10152 19372 10180 19400
rect 1578 19360 1584 19372
rect 1447 19332 1584 19360
rect 1447 19301 1475 19332
rect 1578 19320 1584 19332
rect 1636 19320 1642 19372
rect 6914 19320 6920 19372
rect 6972 19360 6978 19372
rect 7193 19363 7251 19369
rect 7193 19360 7205 19363
rect 6972 19332 7205 19360
rect 6972 19320 6978 19332
rect 7193 19329 7205 19332
rect 7239 19329 7251 19363
rect 8846 19360 8852 19372
rect 8807 19332 8852 19360
rect 7193 19323 7251 19329
rect 8846 19320 8852 19332
rect 8904 19320 8910 19372
rect 9493 19363 9551 19369
rect 9493 19329 9505 19363
rect 9539 19360 9551 19363
rect 10134 19360 10140 19372
rect 9539 19332 10140 19360
rect 9539 19329 9551 19332
rect 9493 19323 9551 19329
rect 10134 19320 10140 19332
rect 10192 19320 10198 19372
rect 10229 19363 10287 19369
rect 10229 19329 10241 19363
rect 10275 19360 10287 19363
rect 10410 19360 10416 19372
rect 10275 19332 10416 19360
rect 10275 19329 10287 19332
rect 10229 19323 10287 19329
rect 10410 19320 10416 19332
rect 10468 19320 10474 19372
rect 10704 19369 10732 19400
rect 14090 19388 14096 19440
rect 14148 19428 14154 19440
rect 16025 19431 16083 19437
rect 16025 19428 16037 19431
rect 14148 19400 16037 19428
rect 14148 19388 14154 19400
rect 10689 19363 10747 19369
rect 10689 19329 10701 19363
rect 10735 19360 10747 19363
rect 12066 19360 12072 19372
rect 10735 19332 12072 19360
rect 10735 19329 10747 19332
rect 10689 19323 10747 19329
rect 12066 19320 12072 19332
rect 12124 19320 12130 19372
rect 14366 19360 14372 19372
rect 14327 19332 14372 19360
rect 14366 19320 14372 19332
rect 14424 19320 14430 19372
rect 1432 19295 1490 19301
rect 1432 19261 1444 19295
rect 1478 19261 1490 19295
rect 1432 19255 1490 19261
rect 12596 19295 12654 19301
rect 12596 19261 12608 19295
rect 12642 19292 12654 19295
rect 12710 19292 12716 19304
rect 12642 19264 12716 19292
rect 12642 19261 12654 19264
rect 12596 19255 12654 19261
rect 12710 19252 12716 19264
rect 12768 19292 12774 19304
rect 12989 19295 13047 19301
rect 12989 19292 13001 19295
rect 12768 19264 13001 19292
rect 12768 19252 12774 19264
rect 12989 19261 13001 19264
rect 13035 19292 13047 19295
rect 13357 19295 13415 19301
rect 13357 19292 13369 19295
rect 13035 19264 13369 19292
rect 13035 19261 13047 19264
rect 12989 19255 13047 19261
rect 13357 19261 13369 19264
rect 13403 19261 13415 19295
rect 13357 19255 13415 19261
rect 13722 19252 13728 19304
rect 13780 19252 13786 19304
rect 15615 19301 15643 19400
rect 16025 19397 16037 19400
rect 16071 19397 16083 19431
rect 16025 19391 16083 19397
rect 15600 19295 15658 19301
rect 15600 19261 15612 19295
rect 15646 19261 15658 19295
rect 15600 19255 15658 19261
rect 18760 19295 18818 19301
rect 18760 19261 18772 19295
rect 18806 19292 18818 19295
rect 19260 19292 19288 19459
rect 20714 19456 20720 19468
rect 20772 19456 20778 19508
rect 21085 19499 21143 19505
rect 21085 19465 21097 19499
rect 21131 19496 21143 19499
rect 21266 19496 21272 19508
rect 21131 19468 21272 19496
rect 21131 19465 21143 19468
rect 21085 19459 21143 19465
rect 21266 19456 21272 19468
rect 21324 19456 21330 19508
rect 21453 19499 21511 19505
rect 21453 19465 21465 19499
rect 21499 19496 21511 19499
rect 21726 19496 21732 19508
rect 21499 19468 21732 19496
rect 21499 19465 21511 19468
rect 21453 19459 21511 19465
rect 18806 19264 19288 19292
rect 20600 19295 20658 19301
rect 18806 19261 18818 19264
rect 18760 19255 18818 19261
rect 20600 19261 20612 19295
rect 20646 19292 20658 19295
rect 21468 19292 21496 19459
rect 21726 19456 21732 19468
rect 21784 19456 21790 19508
rect 22097 19499 22155 19505
rect 22097 19465 22109 19499
rect 22143 19496 22155 19499
rect 22462 19496 22468 19508
rect 22143 19468 22468 19496
rect 22143 19465 22155 19468
rect 22097 19459 22155 19465
rect 20646 19264 21496 19292
rect 21612 19295 21670 19301
rect 20646 19261 20658 19264
rect 20600 19255 20658 19261
rect 21612 19261 21624 19295
rect 21658 19292 21670 19295
rect 22112 19292 22140 19459
rect 22462 19456 22468 19468
rect 22520 19456 22526 19508
rect 21658 19264 22140 19292
rect 21658 19261 21670 19264
rect 21612 19255 21670 19261
rect 1535 19227 1593 19233
rect 1535 19193 1547 19227
rect 1581 19224 1593 19227
rect 5258 19224 5264 19236
rect 1581 19196 5264 19224
rect 1581 19193 1593 19196
rect 1535 19187 1593 19193
rect 5258 19184 5264 19196
rect 5316 19184 5322 19236
rect 6917 19227 6975 19233
rect 6917 19193 6929 19227
rect 6963 19193 6975 19227
rect 6917 19187 6975 19193
rect 6822 19116 6828 19168
rect 6880 19156 6886 19168
rect 6932 19156 6960 19187
rect 7006 19184 7012 19236
rect 7064 19224 7070 19236
rect 7064 19196 7109 19224
rect 7064 19184 7070 19196
rect 8846 19184 8852 19236
rect 8904 19224 8910 19236
rect 8941 19227 8999 19233
rect 8941 19224 8953 19227
rect 8904 19196 8953 19224
rect 8904 19184 8910 19196
rect 8941 19193 8953 19196
rect 8987 19193 8999 19227
rect 10502 19224 10508 19236
rect 10463 19196 10508 19224
rect 8941 19187 8999 19193
rect 10502 19184 10508 19196
rect 10560 19184 10566 19236
rect 13740 19224 13768 19252
rect 14090 19224 14096 19236
rect 13740 19196 14096 19224
rect 14090 19184 14096 19196
rect 14148 19184 14154 19236
rect 14182 19184 14188 19236
rect 14240 19224 14246 19236
rect 15289 19227 15347 19233
rect 15289 19224 15301 19227
rect 14240 19196 15301 19224
rect 14240 19184 14246 19196
rect 15289 19193 15301 19196
rect 15335 19224 15347 19227
rect 15470 19224 15476 19236
rect 15335 19196 15476 19224
rect 15335 19193 15347 19196
rect 15289 19187 15347 19193
rect 15470 19184 15476 19196
rect 15528 19184 15534 19236
rect 7374 19156 7380 19168
rect 6880 19128 7380 19156
rect 6880 19116 6886 19128
rect 7374 19116 7380 19128
rect 7432 19116 7438 19168
rect 12667 19159 12725 19165
rect 12667 19125 12679 19159
rect 12713 19156 12725 19159
rect 12802 19156 12808 19168
rect 12713 19128 12808 19156
rect 12713 19125 12725 19128
rect 12667 19119 12725 19125
rect 12802 19116 12808 19128
rect 12860 19116 12866 19168
rect 13446 19116 13452 19168
rect 13504 19156 13510 19168
rect 13630 19156 13636 19168
rect 13504 19128 13636 19156
rect 13504 19116 13510 19128
rect 13630 19116 13636 19128
rect 13688 19156 13694 19168
rect 13725 19159 13783 19165
rect 13725 19156 13737 19159
rect 13688 19128 13737 19156
rect 13688 19116 13694 19128
rect 13725 19125 13737 19128
rect 13771 19125 13783 19159
rect 13725 19119 13783 19125
rect 15378 19116 15384 19168
rect 15436 19156 15442 19168
rect 15703 19159 15761 19165
rect 15703 19156 15715 19159
rect 15436 19128 15715 19156
rect 15436 19116 15442 19128
rect 15703 19125 15715 19128
rect 15749 19125 15761 19159
rect 15703 19119 15761 19125
rect 18138 19116 18144 19168
rect 18196 19156 18202 19168
rect 18831 19159 18889 19165
rect 18831 19156 18843 19159
rect 18196 19128 18843 19156
rect 18196 19116 18202 19128
rect 18831 19125 18843 19128
rect 18877 19125 18889 19159
rect 18831 19119 18889 19125
rect 18966 19116 18972 19168
rect 19024 19156 19030 19168
rect 20671 19159 20729 19165
rect 20671 19156 20683 19159
rect 19024 19128 20683 19156
rect 19024 19116 19030 19128
rect 20671 19125 20683 19128
rect 20717 19125 20729 19159
rect 20671 19119 20729 19125
rect 20806 19116 20812 19168
rect 20864 19156 20870 19168
rect 21683 19159 21741 19165
rect 21683 19156 21695 19159
rect 20864 19128 21695 19156
rect 20864 19116 20870 19128
rect 21683 19125 21695 19128
rect 21729 19125 21741 19159
rect 21683 19119 21741 19125
rect 1104 19066 22816 19088
rect 1104 19014 8982 19066
rect 9034 19014 9046 19066
rect 9098 19014 9110 19066
rect 9162 19014 9174 19066
rect 9226 19014 16982 19066
rect 17034 19014 17046 19066
rect 17098 19014 17110 19066
rect 17162 19014 17174 19066
rect 17226 19014 22816 19066
rect 1104 18992 22816 19014
rect 198 18912 204 18964
rect 256 18952 262 18964
rect 1581 18955 1639 18961
rect 1581 18952 1593 18955
rect 256 18924 1593 18952
rect 256 18912 262 18924
rect 1581 18921 1593 18924
rect 1627 18921 1639 18955
rect 1581 18915 1639 18921
rect 14090 18912 14096 18964
rect 14148 18952 14154 18964
rect 14461 18955 14519 18961
rect 14461 18952 14473 18955
rect 14148 18924 14473 18952
rect 14148 18912 14154 18924
rect 14461 18921 14473 18924
rect 14507 18921 14519 18955
rect 16298 18952 16304 18964
rect 16259 18924 16304 18952
rect 14461 18915 14519 18921
rect 16298 18912 16304 18924
rect 16356 18912 16362 18964
rect 16850 18912 16856 18964
rect 16908 18952 16914 18964
rect 18138 18952 18144 18964
rect 16908 18924 16988 18952
rect 18099 18924 18144 18952
rect 16908 18912 16914 18924
rect 5258 18884 5264 18896
rect 5219 18856 5264 18884
rect 5258 18844 5264 18856
rect 5316 18844 5322 18896
rect 5353 18887 5411 18893
rect 5353 18853 5365 18887
rect 5399 18884 5411 18887
rect 5442 18884 5448 18896
rect 5399 18856 5448 18884
rect 5399 18853 5411 18856
rect 5353 18847 5411 18853
rect 5442 18844 5448 18856
rect 5500 18844 5506 18896
rect 6638 18844 6644 18896
rect 6696 18884 6702 18896
rect 6917 18887 6975 18893
rect 6917 18884 6929 18887
rect 6696 18856 6929 18884
rect 6696 18844 6702 18856
rect 6917 18853 6929 18856
rect 6963 18853 6975 18887
rect 6917 18847 6975 18853
rect 10502 18844 10508 18896
rect 10560 18884 10566 18896
rect 10965 18887 11023 18893
rect 10965 18884 10977 18887
rect 10560 18856 10977 18884
rect 10560 18844 10566 18856
rect 10965 18853 10977 18856
rect 11011 18853 11023 18887
rect 10965 18847 11023 18853
rect 12802 18844 12808 18896
rect 12860 18884 12866 18896
rect 12989 18887 13047 18893
rect 12989 18884 13001 18887
rect 12860 18856 13001 18884
rect 12860 18844 12866 18856
rect 12989 18853 13001 18856
rect 13035 18853 13047 18887
rect 12989 18847 13047 18853
rect 13081 18887 13139 18893
rect 13081 18853 13093 18887
rect 13127 18884 13139 18887
rect 13446 18884 13452 18896
rect 13127 18856 13452 18884
rect 13127 18853 13139 18856
rect 13081 18847 13139 18853
rect 13446 18844 13452 18856
rect 13504 18844 13510 18896
rect 13633 18887 13691 18893
rect 13633 18853 13645 18887
rect 13679 18884 13691 18887
rect 13722 18884 13728 18896
rect 13679 18856 13728 18884
rect 13679 18853 13691 18856
rect 13633 18847 13691 18853
rect 13722 18844 13728 18856
rect 13780 18884 13786 18896
rect 14366 18884 14372 18896
rect 13780 18856 14372 18884
rect 13780 18844 13786 18856
rect 14366 18844 14372 18856
rect 14424 18844 14430 18896
rect 15473 18887 15531 18893
rect 15473 18853 15485 18887
rect 15519 18884 15531 18887
rect 15838 18884 15844 18896
rect 15519 18856 15844 18884
rect 15519 18853 15531 18856
rect 15473 18847 15531 18853
rect 15838 18844 15844 18856
rect 15896 18844 15902 18896
rect 16960 18893 16988 18924
rect 18138 18912 18144 18924
rect 18196 18912 18202 18964
rect 16945 18887 17003 18893
rect 16945 18853 16957 18887
rect 16991 18853 17003 18887
rect 16945 18847 17003 18853
rect 17034 18844 17040 18896
rect 17092 18884 17098 18896
rect 17092 18856 17137 18884
rect 17092 18844 17098 18856
rect 1397 18819 1455 18825
rect 1397 18785 1409 18819
rect 1443 18816 1455 18819
rect 1946 18816 1952 18828
rect 1443 18788 1952 18816
rect 1443 18785 1455 18788
rect 1397 18779 1455 18785
rect 1946 18776 1952 18788
rect 2004 18776 2010 18828
rect 7558 18776 7564 18828
rect 7616 18816 7622 18828
rect 8294 18816 8300 18828
rect 8352 18825 8358 18828
rect 8352 18819 8390 18825
rect 7616 18788 8300 18816
rect 7616 18776 7622 18788
rect 8294 18776 8300 18788
rect 8378 18785 8390 18819
rect 9950 18816 9956 18828
rect 9911 18788 9956 18816
rect 8352 18779 8390 18785
rect 8352 18776 8358 18779
rect 9950 18776 9956 18788
rect 10008 18776 10014 18828
rect 2498 18748 2504 18760
rect 2459 18720 2504 18748
rect 2498 18708 2504 18720
rect 2556 18708 2562 18760
rect 6822 18748 6828 18760
rect 6783 18720 6828 18748
rect 6822 18708 6828 18720
rect 6880 18708 6886 18760
rect 7101 18751 7159 18757
rect 7101 18717 7113 18751
rect 7147 18717 7159 18751
rect 10870 18748 10876 18760
rect 10831 18720 10876 18748
rect 7101 18711 7159 18717
rect 5813 18683 5871 18689
rect 5813 18649 5825 18683
rect 5859 18680 5871 18683
rect 6914 18680 6920 18692
rect 5859 18652 6920 18680
rect 5859 18649 5871 18652
rect 5813 18643 5871 18649
rect 6914 18640 6920 18652
rect 6972 18680 6978 18692
rect 7116 18680 7144 18711
rect 10870 18708 10876 18720
rect 10928 18708 10934 18760
rect 11149 18751 11207 18757
rect 11149 18717 11161 18751
rect 11195 18717 11207 18751
rect 11149 18711 11207 18717
rect 6972 18652 7144 18680
rect 6972 18640 6978 18652
rect 10686 18640 10692 18692
rect 10744 18680 10750 18692
rect 11164 18680 11192 18711
rect 13354 18708 13360 18760
rect 13412 18748 13418 18760
rect 15381 18751 15439 18757
rect 15381 18748 15393 18751
rect 13412 18720 15393 18748
rect 13412 18708 13418 18720
rect 15381 18717 15393 18720
rect 15427 18748 15439 18751
rect 15470 18748 15476 18760
rect 15427 18720 15476 18748
rect 15427 18717 15439 18720
rect 15381 18711 15439 18717
rect 15470 18708 15476 18720
rect 15528 18708 15534 18760
rect 15562 18708 15568 18760
rect 15620 18748 15626 18760
rect 16025 18751 16083 18757
rect 16025 18748 16037 18751
rect 15620 18720 16037 18748
rect 15620 18708 15626 18720
rect 16025 18717 16037 18720
rect 16071 18748 16083 18751
rect 16666 18748 16672 18760
rect 16071 18720 16672 18748
rect 16071 18717 16083 18720
rect 16025 18711 16083 18717
rect 16666 18708 16672 18720
rect 16724 18708 16730 18760
rect 17218 18748 17224 18760
rect 17179 18720 17224 18748
rect 17218 18708 17224 18720
rect 17276 18708 17282 18760
rect 10744 18652 11192 18680
rect 10744 18640 10750 18652
rect 8435 18615 8493 18621
rect 8435 18581 8447 18615
rect 8481 18612 8493 18615
rect 8570 18612 8576 18624
rect 8481 18584 8576 18612
rect 8481 18581 8493 18584
rect 8435 18575 8493 18581
rect 8570 18572 8576 18584
rect 8628 18572 8634 18624
rect 8846 18612 8852 18624
rect 8807 18584 8852 18612
rect 8846 18572 8852 18584
rect 8904 18572 8910 18624
rect 10413 18615 10471 18621
rect 10413 18581 10425 18615
rect 10459 18612 10471 18615
rect 10502 18612 10508 18624
rect 10459 18584 10508 18612
rect 10459 18581 10471 18584
rect 10413 18575 10471 18581
rect 10502 18572 10508 18584
rect 10560 18572 10566 18624
rect 14093 18615 14151 18621
rect 14093 18581 14105 18615
rect 14139 18612 14151 18615
rect 14182 18612 14188 18624
rect 14139 18584 14188 18612
rect 14139 18581 14151 18584
rect 14093 18575 14151 18581
rect 14182 18572 14188 18584
rect 14240 18612 14246 18624
rect 14734 18612 14740 18624
rect 14240 18584 14740 18612
rect 14240 18572 14246 18584
rect 14734 18572 14740 18584
rect 14792 18572 14798 18624
rect 1104 18522 22816 18544
rect 1104 18470 4982 18522
rect 5034 18470 5046 18522
rect 5098 18470 5110 18522
rect 5162 18470 5174 18522
rect 5226 18470 12982 18522
rect 13034 18470 13046 18522
rect 13098 18470 13110 18522
rect 13162 18470 13174 18522
rect 13226 18470 20982 18522
rect 21034 18470 21046 18522
rect 21098 18470 21110 18522
rect 21162 18470 21174 18522
rect 21226 18470 22816 18522
rect 1104 18448 22816 18470
rect 1946 18408 1952 18420
rect 1907 18380 1952 18408
rect 1946 18368 1952 18380
rect 2004 18408 2010 18420
rect 2639 18411 2697 18417
rect 2639 18408 2651 18411
rect 2004 18380 2651 18408
rect 2004 18368 2010 18380
rect 2639 18377 2651 18380
rect 2685 18377 2697 18411
rect 2639 18371 2697 18377
rect 5350 18368 5356 18420
rect 5408 18408 5414 18420
rect 5537 18411 5595 18417
rect 5537 18408 5549 18411
rect 5408 18380 5549 18408
rect 5408 18368 5414 18380
rect 5537 18377 5549 18380
rect 5583 18377 5595 18411
rect 6638 18408 6644 18420
rect 6599 18380 6644 18408
rect 5537 18371 5595 18377
rect 6638 18368 6644 18380
rect 6696 18368 6702 18420
rect 8294 18408 8300 18420
rect 8255 18380 8300 18408
rect 8294 18368 8300 18380
rect 8352 18368 8358 18420
rect 16850 18368 16856 18420
rect 16908 18408 16914 18420
rect 17313 18411 17371 18417
rect 17313 18408 17325 18411
rect 16908 18380 17325 18408
rect 16908 18368 16914 18380
rect 17313 18377 17325 18380
rect 17359 18377 17371 18411
rect 17313 18371 17371 18377
rect 5261 18343 5319 18349
rect 5261 18309 5273 18343
rect 5307 18340 5319 18343
rect 5442 18340 5448 18352
rect 5307 18312 5448 18340
rect 5307 18309 5319 18312
rect 5261 18303 5319 18309
rect 5442 18300 5448 18312
rect 5500 18300 5506 18352
rect 9306 18340 9312 18352
rect 9267 18312 9312 18340
rect 9306 18300 9312 18312
rect 9364 18300 9370 18352
rect 9953 18343 10011 18349
rect 9953 18309 9965 18343
rect 9999 18340 10011 18343
rect 10870 18340 10876 18352
rect 9999 18312 10876 18340
rect 9999 18309 10011 18312
rect 9953 18303 10011 18309
rect 10870 18300 10876 18312
rect 10928 18300 10934 18352
rect 15013 18343 15071 18349
rect 11992 18312 12848 18340
rect 6914 18272 6920 18284
rect 6875 18244 6920 18272
rect 6914 18232 6920 18244
rect 6972 18232 6978 18284
rect 8570 18232 8576 18284
rect 8628 18272 8634 18284
rect 8757 18275 8815 18281
rect 8757 18272 8769 18275
rect 8628 18244 8769 18272
rect 8628 18232 8634 18244
rect 8757 18241 8769 18244
rect 8803 18241 8815 18275
rect 9324 18272 9352 18300
rect 10321 18275 10379 18281
rect 9324 18244 9674 18272
rect 8757 18235 8815 18241
rect 1397 18207 1455 18213
rect 1397 18173 1409 18207
rect 1443 18173 1455 18207
rect 1397 18167 1455 18173
rect 1412 18136 1440 18167
rect 2314 18164 2320 18216
rect 2372 18204 2378 18216
rect 2568 18207 2626 18213
rect 2568 18204 2580 18207
rect 2372 18176 2580 18204
rect 2372 18164 2378 18176
rect 2568 18173 2580 18176
rect 2614 18204 2626 18207
rect 2961 18207 3019 18213
rect 2961 18204 2973 18207
rect 2614 18176 2973 18204
rect 2614 18173 2626 18176
rect 2568 18167 2626 18173
rect 2961 18173 2973 18176
rect 3007 18173 3019 18207
rect 9646 18204 9674 18244
rect 10321 18241 10333 18275
rect 10367 18272 10379 18275
rect 10962 18272 10968 18284
rect 10367 18244 10968 18272
rect 10367 18241 10379 18244
rect 10321 18235 10379 18241
rect 10962 18232 10968 18244
rect 11020 18232 11026 18284
rect 10686 18204 10692 18216
rect 9646 18176 10692 18204
rect 2961 18167 3019 18173
rect 10686 18164 10692 18176
rect 10744 18164 10750 18216
rect 11992 18204 12020 18312
rect 12066 18232 12072 18284
rect 12124 18272 12130 18284
rect 12526 18272 12532 18284
rect 12124 18244 12532 18272
rect 12124 18232 12130 18244
rect 12526 18232 12532 18244
rect 12584 18232 12590 18284
rect 12820 18281 12848 18312
rect 15013 18309 15025 18343
rect 15059 18340 15071 18343
rect 15562 18340 15568 18352
rect 15059 18312 15568 18340
rect 15059 18309 15071 18312
rect 15013 18303 15071 18309
rect 15562 18300 15568 18312
rect 15620 18300 15626 18352
rect 15930 18300 15936 18352
rect 15988 18340 15994 18352
rect 17034 18340 17040 18352
rect 15988 18312 17040 18340
rect 15988 18300 15994 18312
rect 17034 18300 17040 18312
rect 17092 18300 17098 18352
rect 18230 18340 18236 18352
rect 17236 18312 18236 18340
rect 17236 18284 17264 18312
rect 18230 18300 18236 18312
rect 18288 18340 18294 18352
rect 18288 18312 18460 18340
rect 18288 18300 18294 18312
rect 12805 18275 12863 18281
rect 12805 18241 12817 18275
rect 12851 18241 12863 18275
rect 12805 18235 12863 18241
rect 13909 18275 13967 18281
rect 13909 18241 13921 18275
rect 13955 18272 13967 18275
rect 14461 18275 14519 18281
rect 14461 18272 14473 18275
rect 13955 18244 14473 18272
rect 13955 18241 13967 18244
rect 13909 18235 13967 18241
rect 14461 18241 14473 18244
rect 14507 18272 14519 18275
rect 15378 18272 15384 18284
rect 14507 18244 15384 18272
rect 14507 18241 14519 18244
rect 14461 18235 14519 18241
rect 15378 18232 15384 18244
rect 15436 18232 15442 18284
rect 16025 18275 16083 18281
rect 16025 18241 16037 18275
rect 16071 18272 16083 18275
rect 16298 18272 16304 18284
rect 16071 18244 16304 18272
rect 16071 18241 16083 18244
rect 16025 18235 16083 18241
rect 16298 18232 16304 18244
rect 16356 18232 16362 18284
rect 16669 18275 16727 18281
rect 16669 18241 16681 18275
rect 16715 18272 16727 18275
rect 17218 18272 17224 18284
rect 16715 18244 17224 18272
rect 16715 18241 16727 18244
rect 16669 18235 16727 18241
rect 17218 18232 17224 18244
rect 17276 18232 17282 18284
rect 18138 18272 18144 18284
rect 18099 18244 18144 18272
rect 18138 18232 18144 18244
rect 18196 18232 18202 18284
rect 18432 18281 18460 18312
rect 18417 18275 18475 18281
rect 18417 18241 18429 18275
rect 18463 18241 18475 18275
rect 18417 18235 18475 18241
rect 11532 18176 12020 18204
rect 7009 18139 7067 18145
rect 1412 18108 2452 18136
rect 106 18028 112 18080
rect 164 18068 170 18080
rect 2424 18077 2452 18108
rect 6288 18108 6868 18136
rect 6288 18080 6316 18108
rect 1581 18071 1639 18077
rect 1581 18068 1593 18071
rect 164 18040 1593 18068
rect 164 18028 170 18040
rect 1581 18037 1593 18040
rect 1627 18037 1639 18071
rect 1581 18031 1639 18037
rect 2409 18071 2467 18077
rect 2409 18037 2421 18071
rect 2455 18068 2467 18071
rect 2774 18068 2780 18080
rect 2455 18040 2780 18068
rect 2455 18037 2467 18040
rect 2409 18031 2467 18037
rect 2774 18028 2780 18040
rect 2832 18028 2838 18080
rect 4522 18068 4528 18080
rect 4483 18040 4528 18068
rect 4522 18028 4528 18040
rect 4580 18028 4586 18080
rect 6270 18068 6276 18080
rect 6231 18040 6276 18068
rect 6270 18028 6276 18040
rect 6328 18028 6334 18080
rect 6840 18068 6868 18108
rect 7009 18105 7021 18139
rect 7055 18105 7067 18139
rect 7009 18099 7067 18105
rect 7561 18139 7619 18145
rect 7561 18105 7573 18139
rect 7607 18136 7619 18139
rect 7650 18136 7656 18148
rect 7607 18108 7656 18136
rect 7607 18105 7619 18108
rect 7561 18099 7619 18105
rect 7024 18068 7052 18099
rect 7650 18096 7656 18108
rect 7708 18096 7714 18148
rect 8021 18139 8079 18145
rect 8021 18105 8033 18139
rect 8067 18136 8079 18139
rect 8846 18136 8852 18148
rect 8067 18108 8852 18136
rect 8067 18105 8079 18108
rect 8021 18099 8079 18105
rect 8846 18096 8852 18108
rect 8904 18136 8910 18148
rect 9858 18136 9864 18148
rect 8904 18108 9864 18136
rect 8904 18096 8910 18108
rect 9858 18096 9864 18108
rect 9916 18096 9922 18148
rect 10873 18139 10931 18145
rect 10873 18105 10885 18139
rect 10919 18105 10931 18139
rect 10873 18099 10931 18105
rect 6840 18040 7052 18068
rect 10502 18028 10508 18080
rect 10560 18068 10566 18080
rect 10597 18071 10655 18077
rect 10597 18068 10609 18071
rect 10560 18040 10609 18068
rect 10560 18028 10566 18040
rect 10597 18037 10609 18040
rect 10643 18037 10655 18071
rect 10597 18031 10655 18037
rect 10778 18028 10784 18080
rect 10836 18068 10842 18080
rect 10888 18068 10916 18099
rect 10962 18096 10968 18148
rect 11020 18136 11026 18148
rect 11146 18136 11152 18148
rect 11020 18108 11152 18136
rect 11020 18096 11026 18108
rect 11146 18096 11152 18108
rect 11204 18096 11210 18148
rect 11238 18096 11244 18148
rect 11296 18136 11302 18148
rect 11532 18145 11560 18176
rect 11517 18139 11575 18145
rect 11517 18136 11529 18139
rect 11296 18108 11529 18136
rect 11296 18096 11302 18108
rect 11517 18105 11529 18108
rect 11563 18105 11575 18139
rect 11517 18099 11575 18105
rect 12621 18139 12679 18145
rect 12621 18105 12633 18139
rect 12667 18105 12679 18139
rect 12621 18099 12679 18105
rect 14277 18139 14335 18145
rect 14277 18105 14289 18139
rect 14323 18136 14335 18139
rect 14550 18136 14556 18148
rect 14323 18108 14556 18136
rect 14323 18105 14335 18108
rect 14277 18099 14335 18105
rect 11793 18071 11851 18077
rect 11793 18068 11805 18071
rect 10836 18040 11805 18068
rect 10836 18028 10842 18040
rect 11793 18037 11805 18040
rect 11839 18037 11851 18071
rect 12158 18068 12164 18080
rect 12119 18040 12164 18068
rect 11793 18031 11851 18037
rect 12158 18028 12164 18040
rect 12216 18068 12222 18080
rect 12636 18068 12664 18099
rect 14550 18096 14556 18108
rect 14608 18096 14614 18148
rect 16117 18139 16175 18145
rect 16117 18105 16129 18139
rect 16163 18105 16175 18139
rect 18233 18139 18291 18145
rect 18233 18136 18245 18139
rect 16117 18099 16175 18105
rect 17788 18108 18245 18136
rect 13446 18068 13452 18080
rect 12216 18040 12664 18068
rect 13407 18040 13452 18068
rect 12216 18028 12222 18040
rect 13446 18028 13452 18040
rect 13504 18028 13510 18080
rect 15473 18071 15531 18077
rect 15473 18037 15485 18071
rect 15519 18068 15531 18071
rect 15838 18068 15844 18080
rect 15519 18040 15844 18068
rect 15519 18037 15531 18040
rect 15473 18031 15531 18037
rect 15838 18028 15844 18040
rect 15896 18068 15902 18080
rect 16132 18068 16160 18099
rect 15896 18040 16160 18068
rect 15896 18028 15902 18040
rect 17586 18028 17592 18080
rect 17644 18068 17650 18080
rect 17788 18077 17816 18108
rect 18233 18105 18245 18108
rect 18279 18105 18291 18139
rect 18233 18099 18291 18105
rect 17773 18071 17831 18077
rect 17773 18068 17785 18071
rect 17644 18040 17785 18068
rect 17644 18028 17650 18040
rect 17773 18037 17785 18040
rect 17819 18037 17831 18071
rect 17773 18031 17831 18037
rect 1104 17978 22816 18000
rect 1104 17926 8982 17978
rect 9034 17926 9046 17978
rect 9098 17926 9110 17978
rect 9162 17926 9174 17978
rect 9226 17926 16982 17978
rect 17034 17926 17046 17978
rect 17098 17926 17110 17978
rect 17162 17926 17174 17978
rect 17226 17926 22816 17978
rect 1104 17904 22816 17926
rect 6270 17824 6276 17876
rect 6328 17864 6334 17876
rect 6549 17867 6607 17873
rect 6549 17864 6561 17867
rect 6328 17836 6561 17864
rect 6328 17824 6334 17836
rect 6549 17833 6561 17836
rect 6595 17833 6607 17867
rect 6549 17827 6607 17833
rect 6914 17824 6920 17876
rect 6972 17864 6978 17876
rect 7561 17867 7619 17873
rect 7561 17864 7573 17867
rect 6972 17836 7573 17864
rect 6972 17824 6978 17836
rect 7561 17833 7573 17836
rect 7607 17833 7619 17867
rect 7561 17827 7619 17833
rect 8570 17824 8576 17876
rect 8628 17864 8634 17876
rect 9033 17867 9091 17873
rect 9033 17864 9045 17867
rect 8628 17836 9045 17864
rect 8628 17824 8634 17836
rect 9033 17833 9045 17836
rect 9079 17833 9091 17867
rect 9033 17827 9091 17833
rect 10962 17824 10968 17876
rect 11020 17864 11026 17876
rect 11057 17867 11115 17873
rect 11057 17864 11069 17867
rect 11020 17836 11069 17864
rect 11020 17824 11026 17836
rect 11057 17833 11069 17836
rect 11103 17833 11115 17867
rect 11057 17827 11115 17833
rect 11146 17824 11152 17876
rect 11204 17864 11210 17876
rect 11609 17867 11667 17873
rect 11609 17864 11621 17867
rect 11204 17836 11621 17864
rect 11204 17824 11210 17836
rect 11609 17833 11621 17836
rect 11655 17833 11667 17867
rect 12526 17864 12532 17876
rect 12487 17836 12532 17864
rect 11609 17827 11667 17833
rect 12526 17824 12532 17836
rect 12584 17824 12590 17876
rect 12802 17824 12808 17876
rect 12860 17864 12866 17876
rect 12897 17867 12955 17873
rect 12897 17864 12909 17867
rect 12860 17836 12909 17864
rect 12860 17824 12866 17836
rect 12897 17833 12909 17836
rect 12943 17833 12955 17867
rect 15470 17864 15476 17876
rect 15431 17836 15476 17864
rect 12897 17827 12955 17833
rect 15470 17824 15476 17836
rect 15528 17824 15534 17876
rect 5626 17756 5632 17808
rect 5684 17796 5690 17808
rect 5950 17799 6008 17805
rect 5950 17796 5962 17799
rect 5684 17768 5962 17796
rect 5684 17756 5690 17768
rect 5950 17765 5962 17768
rect 5996 17765 6008 17799
rect 5950 17759 6008 17765
rect 6822 17756 6828 17808
rect 6880 17796 6886 17808
rect 7193 17799 7251 17805
rect 7193 17796 7205 17799
rect 6880 17768 7205 17796
rect 6880 17756 6886 17768
rect 7193 17765 7205 17768
rect 7239 17765 7251 17799
rect 7193 17759 7251 17765
rect 15841 17799 15899 17805
rect 15841 17765 15853 17799
rect 15887 17796 15899 17799
rect 15930 17796 15936 17808
rect 15887 17768 15936 17796
rect 15887 17765 15899 17768
rect 15841 17759 15899 17765
rect 15930 17756 15936 17768
rect 15988 17756 15994 17808
rect 17405 17799 17463 17805
rect 17405 17765 17417 17799
rect 17451 17796 17463 17799
rect 17586 17796 17592 17808
rect 17451 17768 17592 17796
rect 17451 17765 17463 17768
rect 17405 17759 17463 17765
rect 17586 17756 17592 17768
rect 17644 17756 17650 17808
rect 2222 17728 2228 17740
rect 2183 17700 2228 17728
rect 2222 17688 2228 17700
rect 2280 17688 2286 17740
rect 3881 17731 3939 17737
rect 3881 17697 3893 17731
rect 3927 17728 3939 17731
rect 4157 17731 4215 17737
rect 4157 17728 4169 17731
rect 3927 17700 4169 17728
rect 3927 17697 3939 17700
rect 3881 17691 3939 17697
rect 4157 17697 4169 17700
rect 4203 17697 4215 17731
rect 4157 17691 4215 17697
rect 4525 17731 4583 17737
rect 4525 17697 4537 17731
rect 4571 17728 4583 17731
rect 4706 17728 4712 17740
rect 4571 17700 4712 17728
rect 4571 17697 4583 17700
rect 4525 17691 4583 17697
rect 4172 17592 4200 17691
rect 4706 17688 4712 17700
rect 4764 17688 4770 17740
rect 8018 17728 8024 17740
rect 7979 17700 8024 17728
rect 8018 17688 8024 17700
rect 8076 17688 8082 17740
rect 8478 17728 8484 17740
rect 8439 17700 8484 17728
rect 8478 17688 8484 17700
rect 8536 17688 8542 17740
rect 12710 17688 12716 17740
rect 12768 17728 12774 17740
rect 13081 17731 13139 17737
rect 13081 17728 13093 17731
rect 12768 17700 13093 17728
rect 12768 17688 12774 17700
rect 13081 17697 13093 17700
rect 13127 17697 13139 17731
rect 13538 17728 13544 17740
rect 13499 17700 13544 17728
rect 13081 17691 13139 17697
rect 13538 17688 13544 17700
rect 13596 17688 13602 17740
rect 4614 17660 4620 17672
rect 4575 17632 4620 17660
rect 4614 17620 4620 17632
rect 4672 17620 4678 17672
rect 5629 17663 5687 17669
rect 5629 17629 5641 17663
rect 5675 17660 5687 17663
rect 6086 17660 6092 17672
rect 5675 17632 6092 17660
rect 5675 17629 5687 17632
rect 5629 17623 5687 17629
rect 6086 17620 6092 17632
rect 6144 17620 6150 17672
rect 8570 17660 8576 17672
rect 8531 17632 8576 17660
rect 8570 17620 8576 17632
rect 8628 17620 8634 17672
rect 10686 17660 10692 17672
rect 10647 17632 10692 17660
rect 10686 17620 10692 17632
rect 10744 17620 10750 17672
rect 13817 17663 13875 17669
rect 13817 17629 13829 17663
rect 13863 17660 13875 17663
rect 13906 17660 13912 17672
rect 13863 17632 13912 17660
rect 13863 17629 13875 17632
rect 13817 17623 13875 17629
rect 13906 17620 13912 17632
rect 13964 17660 13970 17672
rect 14093 17663 14151 17669
rect 14093 17660 14105 17663
rect 13964 17632 14105 17660
rect 13964 17620 13970 17632
rect 14093 17629 14105 17632
rect 14139 17629 14151 17663
rect 14093 17623 14151 17629
rect 15194 17620 15200 17672
rect 15252 17660 15258 17672
rect 15749 17663 15807 17669
rect 15749 17660 15761 17663
rect 15252 17632 15761 17660
rect 15252 17620 15258 17632
rect 15749 17629 15761 17632
rect 15795 17629 15807 17663
rect 17310 17660 17316 17672
rect 17223 17632 17316 17660
rect 15749 17623 15807 17629
rect 17310 17620 17316 17632
rect 17368 17660 17374 17672
rect 18785 17663 18843 17669
rect 18785 17660 18797 17663
rect 17368 17632 18797 17660
rect 17368 17620 17374 17632
rect 18785 17629 18797 17632
rect 18831 17629 18843 17663
rect 18785 17623 18843 17629
rect 11606 17592 11612 17604
rect 4172 17564 11612 17592
rect 11606 17552 11612 17564
rect 11664 17552 11670 17604
rect 16301 17595 16359 17601
rect 16301 17561 16313 17595
rect 16347 17592 16359 17595
rect 17862 17592 17868 17604
rect 16347 17564 17868 17592
rect 16347 17561 16359 17564
rect 16301 17555 16359 17561
rect 17862 17552 17868 17564
rect 17920 17552 17926 17604
rect 1946 17524 1952 17536
rect 1907 17496 1952 17524
rect 1946 17484 1952 17496
rect 2004 17484 2010 17536
rect 6917 17527 6975 17533
rect 6917 17493 6929 17527
rect 6963 17524 6975 17527
rect 7098 17524 7104 17536
rect 6963 17496 7104 17524
rect 6963 17493 6975 17496
rect 6917 17487 6975 17493
rect 7098 17484 7104 17496
rect 7156 17484 7162 17536
rect 10505 17527 10563 17533
rect 10505 17493 10517 17527
rect 10551 17524 10563 17527
rect 10594 17524 10600 17536
rect 10551 17496 10600 17524
rect 10551 17493 10563 17496
rect 10505 17487 10563 17493
rect 10594 17484 10600 17496
rect 10652 17484 10658 17536
rect 18322 17524 18328 17536
rect 18283 17496 18328 17524
rect 18322 17484 18328 17496
rect 18380 17484 18386 17536
rect 1104 17434 22816 17456
rect 1104 17382 4982 17434
rect 5034 17382 5046 17434
rect 5098 17382 5110 17434
rect 5162 17382 5174 17434
rect 5226 17382 12982 17434
rect 13034 17382 13046 17434
rect 13098 17382 13110 17434
rect 13162 17382 13174 17434
rect 13226 17382 20982 17434
rect 21034 17382 21046 17434
rect 21098 17382 21110 17434
rect 21162 17382 21174 17434
rect 21226 17382 22816 17434
rect 1104 17360 22816 17382
rect 2498 17280 2504 17332
rect 2556 17320 2562 17332
rect 2593 17323 2651 17329
rect 2593 17320 2605 17323
rect 2556 17292 2605 17320
rect 2556 17280 2562 17292
rect 2593 17289 2605 17292
rect 2639 17289 2651 17323
rect 2593 17283 2651 17289
rect 5169 17323 5227 17329
rect 5169 17289 5181 17323
rect 5215 17320 5227 17323
rect 7006 17320 7012 17332
rect 5215 17292 7012 17320
rect 5215 17289 5227 17292
rect 5169 17283 5227 17289
rect 7006 17280 7012 17292
rect 7064 17280 7070 17332
rect 8113 17323 8171 17329
rect 8113 17289 8125 17323
rect 8159 17320 8171 17323
rect 8478 17320 8484 17332
rect 8159 17292 8484 17320
rect 8159 17289 8171 17292
rect 8113 17283 8171 17289
rect 8478 17280 8484 17292
rect 8536 17280 8542 17332
rect 9493 17323 9551 17329
rect 9493 17289 9505 17323
rect 9539 17320 9551 17323
rect 9766 17320 9772 17332
rect 9539 17292 9772 17320
rect 9539 17289 9551 17292
rect 9493 17283 9551 17289
rect 9766 17280 9772 17292
rect 9824 17280 9830 17332
rect 11333 17323 11391 17329
rect 11333 17289 11345 17323
rect 11379 17320 11391 17323
rect 12158 17320 12164 17332
rect 11379 17292 12164 17320
rect 11379 17289 11391 17292
rect 11333 17283 11391 17289
rect 12158 17280 12164 17292
rect 12216 17280 12222 17332
rect 13173 17323 13231 17329
rect 13173 17289 13185 17323
rect 13219 17320 13231 17323
rect 13538 17320 13544 17332
rect 13219 17292 13544 17320
rect 13219 17289 13231 17292
rect 13173 17283 13231 17289
rect 13538 17280 13544 17292
rect 13596 17280 13602 17332
rect 14550 17280 14556 17332
rect 14608 17320 14614 17332
rect 14829 17323 14887 17329
rect 14829 17320 14841 17323
rect 14608 17292 14841 17320
rect 14608 17280 14614 17292
rect 14829 17289 14841 17292
rect 14875 17320 14887 17323
rect 15565 17323 15623 17329
rect 15565 17320 15577 17323
rect 14875 17292 15577 17320
rect 14875 17289 14887 17292
rect 14829 17283 14887 17289
rect 15565 17289 15577 17292
rect 15611 17320 15623 17323
rect 15930 17320 15936 17332
rect 15611 17292 15936 17320
rect 15611 17289 15623 17292
rect 15565 17283 15623 17289
rect 15930 17280 15936 17292
rect 15988 17280 15994 17332
rect 17310 17320 17316 17332
rect 17271 17292 17316 17320
rect 17310 17280 17316 17292
rect 17368 17280 17374 17332
rect 21085 17323 21143 17329
rect 21085 17289 21097 17323
rect 21131 17320 21143 17323
rect 21266 17320 21272 17332
rect 21131 17292 21272 17320
rect 21131 17289 21143 17292
rect 21085 17283 21143 17289
rect 21266 17280 21272 17292
rect 21324 17280 21330 17332
rect 2516 17252 2544 17280
rect 1688 17224 2544 17252
rect 1688 17193 1716 17224
rect 8018 17212 8024 17264
rect 8076 17252 8082 17264
rect 12710 17252 12716 17264
rect 8076 17224 12716 17252
rect 8076 17212 8082 17224
rect 12710 17212 12716 17224
rect 12768 17212 12774 17264
rect 1673 17187 1731 17193
rect 1673 17153 1685 17187
rect 1719 17153 1731 17187
rect 2314 17184 2320 17196
rect 2275 17156 2320 17184
rect 1673 17147 1731 17153
rect 2314 17144 2320 17156
rect 2372 17144 2378 17196
rect 8570 17184 8576 17196
rect 8531 17156 8576 17184
rect 8570 17144 8576 17156
rect 8628 17144 8634 17196
rect 10686 17144 10692 17196
rect 10744 17184 10750 17196
rect 11609 17187 11667 17193
rect 11609 17184 11621 17187
rect 10744 17156 11621 17184
rect 10744 17144 10750 17156
rect 11609 17153 11621 17156
rect 11655 17153 11667 17187
rect 13906 17184 13912 17196
rect 13867 17156 13912 17184
rect 11609 17147 11667 17153
rect 13906 17144 13912 17156
rect 13964 17144 13970 17196
rect 18230 17184 18236 17196
rect 18191 17156 18236 17184
rect 18230 17144 18236 17156
rect 18288 17144 18294 17196
rect 18690 17184 18696 17196
rect 18651 17156 18696 17184
rect 18690 17144 18696 17156
rect 18748 17144 18754 17196
rect 2866 17076 2872 17128
rect 2924 17116 2930 17128
rect 3180 17119 3238 17125
rect 3180 17116 3192 17119
rect 2924 17088 3192 17116
rect 2924 17076 2930 17088
rect 3180 17085 3192 17088
rect 3226 17116 3238 17119
rect 3605 17119 3663 17125
rect 3605 17116 3617 17119
rect 3226 17088 3617 17116
rect 3226 17085 3238 17088
rect 3180 17079 3238 17085
rect 3605 17085 3617 17088
rect 3651 17085 3663 17119
rect 4246 17116 4252 17128
rect 4207 17088 4252 17116
rect 3605 17079 3663 17085
rect 4246 17076 4252 17088
rect 4304 17076 4310 17128
rect 4706 17076 4712 17128
rect 4764 17116 4770 17128
rect 6546 17116 6552 17128
rect 4764 17088 6552 17116
rect 4764 17076 4770 17088
rect 6546 17076 6552 17088
rect 6604 17076 6610 17128
rect 7098 17116 7104 17128
rect 7059 17088 7104 17116
rect 7098 17076 7104 17088
rect 7156 17076 7162 17128
rect 7190 17076 7196 17128
rect 7248 17116 7254 17128
rect 7285 17119 7343 17125
rect 7285 17116 7297 17119
rect 7248 17088 7297 17116
rect 7248 17076 7254 17088
rect 7285 17085 7297 17088
rect 7331 17085 7343 17119
rect 7285 17079 7343 17085
rect 10413 17119 10471 17125
rect 10413 17085 10425 17119
rect 10459 17116 10471 17119
rect 10594 17116 10600 17128
rect 10459 17088 10600 17116
rect 10459 17085 10471 17088
rect 10413 17079 10471 17085
rect 10594 17076 10600 17088
rect 10652 17076 10658 17128
rect 20806 17076 20812 17128
rect 20864 17116 20870 17128
rect 20901 17119 20959 17125
rect 20901 17116 20913 17119
rect 20864 17088 20913 17116
rect 20864 17076 20870 17088
rect 20901 17085 20913 17088
rect 20947 17116 20959 17119
rect 21453 17119 21511 17125
rect 21453 17116 21465 17119
rect 20947 17088 21465 17116
rect 20947 17085 20959 17088
rect 20901 17079 20959 17085
rect 21453 17085 21465 17088
rect 21499 17085 21511 17119
rect 21453 17079 21511 17085
rect 1765 17051 1823 17057
rect 1765 17017 1777 17051
rect 1811 17048 1823 17051
rect 1946 17048 1952 17060
rect 1811 17020 1952 17048
rect 1811 17017 1823 17020
rect 1765 17011 1823 17017
rect 1946 17008 1952 17020
rect 2004 17008 2010 17060
rect 4570 17051 4628 17057
rect 4570 17048 4582 17051
rect 4356 17020 4582 17048
rect 4356 16992 4384 17020
rect 4570 17017 4582 17020
rect 4616 17048 4628 17051
rect 5626 17048 5632 17060
rect 4616 17020 5632 17048
rect 4616 17017 4628 17020
rect 4570 17011 4628 17017
rect 5626 17008 5632 17020
rect 5684 17008 5690 17060
rect 6086 17048 6092 17060
rect 5999 17020 6092 17048
rect 6086 17008 6092 17020
rect 6144 17048 6150 17060
rect 8894 17051 8952 17057
rect 8894 17048 8906 17051
rect 6144 17020 6770 17048
rect 6144 17008 6150 17020
rect 2958 16980 2964 16992
rect 2919 16952 2964 16980
rect 2958 16940 2964 16952
rect 3016 16940 3022 16992
rect 3283 16983 3341 16989
rect 3283 16949 3295 16983
rect 3329 16980 3341 16983
rect 3510 16980 3516 16992
rect 3329 16952 3516 16980
rect 3329 16949 3341 16952
rect 3283 16943 3341 16949
rect 3510 16940 3516 16952
rect 3568 16940 3574 16992
rect 4157 16983 4215 16989
rect 4157 16949 4169 16983
rect 4203 16980 4215 16983
rect 4338 16980 4344 16992
rect 4203 16952 4344 16980
rect 4203 16949 4215 16952
rect 4157 16943 4215 16949
rect 4338 16940 4344 16952
rect 4396 16940 4402 16992
rect 6742 16980 6770 17020
rect 8404 17020 8906 17048
rect 8404 16992 8432 17020
rect 8894 17017 8906 17020
rect 8940 17048 8952 17051
rect 10775 17051 10833 17057
rect 8940 17020 9674 17048
rect 8940 17017 8952 17020
rect 8894 17011 8952 17017
rect 6917 16983 6975 16989
rect 6917 16980 6929 16983
rect 6742 16952 6929 16980
rect 6917 16949 6929 16952
rect 6963 16949 6975 16983
rect 8386 16980 8392 16992
rect 8347 16952 8392 16980
rect 6917 16943 6975 16949
rect 8386 16940 8392 16952
rect 8444 16940 8450 16992
rect 9646 16980 9674 17020
rect 10775 17017 10787 17051
rect 10821 17017 10833 17051
rect 10775 17011 10833 17017
rect 9953 16983 10011 16989
rect 9953 16980 9965 16983
rect 9646 16952 9965 16980
rect 9953 16949 9965 16952
rect 9999 16980 10011 16983
rect 10321 16983 10379 16989
rect 10321 16980 10333 16983
rect 9999 16952 10333 16980
rect 9999 16949 10011 16952
rect 9953 16943 10011 16949
rect 10321 16949 10333 16952
rect 10367 16980 10379 16983
rect 10790 16980 10818 17011
rect 13538 17008 13544 17060
rect 13596 17048 13602 17060
rect 13814 17048 13820 17060
rect 13596 17020 13820 17048
rect 13596 17008 13602 17020
rect 13814 17008 13820 17020
rect 13872 17008 13878 17060
rect 14230 17051 14288 17057
rect 14230 17048 14242 17051
rect 13924 17020 14242 17048
rect 13924 16992 13952 17020
rect 14230 17017 14242 17020
rect 14276 17017 14288 17051
rect 16114 17048 16120 17060
rect 16075 17020 16120 17048
rect 14230 17011 14288 17017
rect 16114 17008 16120 17020
rect 16172 17008 16178 17060
rect 16209 17051 16267 17057
rect 16209 17017 16221 17051
rect 16255 17017 16267 17051
rect 16209 17011 16267 17017
rect 16761 17051 16819 17057
rect 16761 17017 16773 17051
rect 16807 17048 16819 17051
rect 17862 17048 17868 17060
rect 16807 17020 17868 17048
rect 16807 17017 16819 17020
rect 16761 17011 16819 17017
rect 10962 16980 10968 16992
rect 10367 16952 10968 16980
rect 10367 16949 10379 16952
rect 10321 16943 10379 16949
rect 10962 16940 10968 16952
rect 11020 16980 11026 16992
rect 13725 16983 13783 16989
rect 13725 16980 13737 16983
rect 11020 16952 13737 16980
rect 11020 16940 11026 16952
rect 13725 16949 13737 16952
rect 13771 16980 13783 16983
rect 13906 16980 13912 16992
rect 13771 16952 13912 16980
rect 13771 16949 13783 16952
rect 13725 16943 13783 16949
rect 13906 16940 13912 16952
rect 13964 16940 13970 16992
rect 15194 16980 15200 16992
rect 15155 16952 15200 16980
rect 15194 16940 15200 16952
rect 15252 16940 15258 16992
rect 15838 16980 15844 16992
rect 15799 16952 15844 16980
rect 15838 16940 15844 16952
rect 15896 16980 15902 16992
rect 16224 16980 16252 17011
rect 17862 17008 17868 17020
rect 17920 17008 17926 17060
rect 18322 17008 18328 17060
rect 18380 17048 18386 17060
rect 18380 17020 18425 17048
rect 18380 17008 18386 17020
rect 17586 16980 17592 16992
rect 15896 16952 16252 16980
rect 17547 16952 17592 16980
rect 15896 16940 15902 16952
rect 17586 16940 17592 16952
rect 17644 16940 17650 16992
rect 1104 16890 22816 16912
rect 1104 16838 8982 16890
rect 9034 16838 9046 16890
rect 9098 16838 9110 16890
rect 9162 16838 9174 16890
rect 9226 16838 16982 16890
rect 17034 16838 17046 16890
rect 17098 16838 17110 16890
rect 17162 16838 17174 16890
rect 17226 16838 22816 16890
rect 1104 16816 22816 16838
rect 1673 16779 1731 16785
rect 1673 16745 1685 16779
rect 1719 16776 1731 16779
rect 1946 16776 1952 16788
rect 1719 16748 1952 16776
rect 1719 16745 1731 16748
rect 1673 16739 1731 16745
rect 1946 16736 1952 16748
rect 2004 16736 2010 16788
rect 4246 16736 4252 16788
rect 4304 16776 4310 16788
rect 4341 16779 4399 16785
rect 4341 16776 4353 16779
rect 4304 16748 4353 16776
rect 4304 16736 4310 16748
rect 4341 16745 4353 16748
rect 4387 16776 4399 16779
rect 5077 16779 5135 16785
rect 5077 16776 5089 16779
rect 4387 16748 5089 16776
rect 4387 16745 4399 16748
rect 4341 16739 4399 16745
rect 5077 16745 5089 16748
rect 5123 16745 5135 16779
rect 5077 16739 5135 16745
rect 5442 16736 5448 16788
rect 5500 16776 5506 16788
rect 6730 16776 6736 16788
rect 5500 16748 6736 16776
rect 5500 16736 5506 16748
rect 6730 16736 6736 16748
rect 6788 16776 6794 16788
rect 7929 16779 7987 16785
rect 7929 16776 7941 16779
rect 6788 16748 7941 16776
rect 6788 16736 6794 16748
rect 7929 16745 7941 16748
rect 7975 16745 7987 16779
rect 8570 16776 8576 16788
rect 8531 16748 8576 16776
rect 7929 16739 7987 16745
rect 8570 16736 8576 16748
rect 8628 16736 8634 16788
rect 11698 16776 11704 16788
rect 11659 16748 11704 16776
rect 11698 16736 11704 16748
rect 11756 16736 11762 16788
rect 15427 16779 15485 16785
rect 15427 16745 15439 16779
rect 15473 16776 15485 16779
rect 16114 16776 16120 16788
rect 15473 16748 16120 16776
rect 15473 16745 15485 16748
rect 15427 16739 15485 16745
rect 16114 16736 16120 16748
rect 16172 16736 16178 16788
rect 18233 16779 18291 16785
rect 18233 16745 18245 16779
rect 18279 16776 18291 16779
rect 18322 16776 18328 16788
rect 18279 16748 18328 16776
rect 18279 16745 18291 16748
rect 18233 16739 18291 16745
rect 18322 16736 18328 16748
rect 18380 16736 18386 16788
rect 2133 16711 2191 16717
rect 2133 16677 2145 16711
rect 2179 16708 2191 16711
rect 2222 16708 2228 16720
rect 2179 16680 2228 16708
rect 2179 16677 2191 16680
rect 2133 16671 2191 16677
rect 2222 16668 2228 16680
rect 2280 16708 2286 16720
rect 2958 16708 2964 16720
rect 2280 16680 2964 16708
rect 2280 16668 2286 16680
rect 2958 16668 2964 16680
rect 3016 16668 3022 16720
rect 6546 16668 6552 16720
rect 6604 16708 6610 16720
rect 6825 16711 6883 16717
rect 6825 16708 6837 16711
rect 6604 16680 6837 16708
rect 6604 16668 6610 16680
rect 6825 16677 6837 16680
rect 6871 16708 6883 16711
rect 7190 16708 7196 16720
rect 6871 16680 7196 16708
rect 6871 16677 6883 16680
rect 6825 16671 6883 16677
rect 7190 16668 7196 16680
rect 7248 16668 7254 16720
rect 7371 16711 7429 16717
rect 7371 16677 7383 16711
rect 7417 16708 7429 16711
rect 8386 16708 8392 16720
rect 7417 16680 8392 16708
rect 7417 16677 7429 16680
rect 7371 16671 7429 16677
rect 8386 16668 8392 16680
rect 8444 16668 8450 16720
rect 10686 16668 10692 16720
rect 10744 16708 10750 16720
rect 10781 16711 10839 16717
rect 10781 16708 10793 16711
rect 10744 16680 10793 16708
rect 10744 16668 10750 16680
rect 10781 16677 10793 16680
rect 10827 16677 10839 16711
rect 10781 16671 10839 16677
rect 11072 16680 12112 16708
rect 4154 16600 4160 16652
rect 4212 16640 4218 16652
rect 4617 16643 4675 16649
rect 4212 16612 4257 16640
rect 4212 16600 4218 16612
rect 4617 16609 4629 16643
rect 4663 16640 4675 16643
rect 4706 16640 4712 16652
rect 4663 16612 4712 16640
rect 4663 16609 4675 16612
rect 4617 16603 4675 16609
rect 4706 16600 4712 16612
rect 4764 16600 4770 16652
rect 5997 16643 6055 16649
rect 5997 16609 6009 16643
rect 6043 16640 6055 16643
rect 6086 16640 6092 16652
rect 6043 16612 6092 16640
rect 6043 16609 6055 16612
rect 5997 16603 6055 16609
rect 6086 16600 6092 16612
rect 6144 16600 6150 16652
rect 7098 16600 7104 16652
rect 7156 16640 7162 16652
rect 10318 16640 10324 16652
rect 7156 16612 10324 16640
rect 7156 16600 7162 16612
rect 10318 16600 10324 16612
rect 10376 16600 10382 16652
rect 10410 16600 10416 16652
rect 10468 16640 10474 16652
rect 11072 16649 11100 16680
rect 10505 16643 10563 16649
rect 10505 16640 10517 16643
rect 10468 16612 10517 16640
rect 10468 16600 10474 16612
rect 10505 16609 10517 16612
rect 10551 16640 10563 16643
rect 11057 16643 11115 16649
rect 11057 16640 11069 16643
rect 10551 16612 11069 16640
rect 10551 16609 10563 16612
rect 10505 16603 10563 16609
rect 11057 16609 11069 16612
rect 11103 16609 11115 16643
rect 11606 16640 11612 16652
rect 11567 16612 11612 16640
rect 11057 16603 11115 16609
rect 11606 16600 11612 16612
rect 11664 16640 11670 16652
rect 11974 16640 11980 16652
rect 11664 16612 11980 16640
rect 11664 16600 11670 16612
rect 11974 16600 11980 16612
rect 12032 16600 12038 16652
rect 12084 16649 12112 16680
rect 15194 16668 15200 16720
rect 15252 16708 15258 16720
rect 16439 16711 16497 16717
rect 16439 16708 16451 16711
rect 15252 16680 16451 16708
rect 15252 16668 15258 16680
rect 16439 16677 16451 16680
rect 16485 16677 16497 16711
rect 16439 16671 16497 16677
rect 17402 16668 17408 16720
rect 17460 16708 17466 16720
rect 17634 16711 17692 16717
rect 17634 16708 17646 16711
rect 17460 16680 17646 16708
rect 17460 16668 17466 16680
rect 17634 16677 17646 16680
rect 17680 16677 17692 16711
rect 17634 16671 17692 16677
rect 12069 16643 12127 16649
rect 12069 16609 12081 16643
rect 12115 16609 12127 16643
rect 13262 16640 13268 16652
rect 13223 16612 13268 16640
rect 12069 16603 12127 16609
rect 13262 16600 13268 16612
rect 13320 16600 13326 16652
rect 13814 16600 13820 16652
rect 13872 16640 13878 16652
rect 15289 16643 15347 16649
rect 13872 16612 13917 16640
rect 13872 16600 13878 16612
rect 15289 16609 15301 16643
rect 15335 16640 15347 16643
rect 15378 16640 15384 16652
rect 15335 16612 15384 16640
rect 15335 16609 15347 16612
rect 15289 16603 15347 16609
rect 15378 16600 15384 16612
rect 15436 16600 15442 16652
rect 16336 16643 16394 16649
rect 16336 16640 16348 16643
rect 16132 16612 16348 16640
rect 2041 16575 2099 16581
rect 2041 16541 2053 16575
rect 2087 16541 2099 16575
rect 2314 16572 2320 16584
rect 2275 16544 2320 16572
rect 2041 16535 2099 16541
rect 2056 16504 2084 16535
rect 2314 16532 2320 16544
rect 2372 16532 2378 16584
rect 7009 16575 7067 16581
rect 7009 16541 7021 16575
rect 7055 16572 7067 16575
rect 7558 16572 7564 16584
rect 7055 16544 7564 16572
rect 7055 16541 7067 16544
rect 7009 16535 7067 16541
rect 7558 16532 7564 16544
rect 7616 16532 7622 16584
rect 13998 16572 14004 16584
rect 13959 16544 14004 16572
rect 13998 16532 14004 16544
rect 14056 16532 14062 16584
rect 16132 16516 16160 16612
rect 16336 16609 16348 16612
rect 16382 16609 16394 16643
rect 16336 16603 16394 16609
rect 18230 16600 18236 16652
rect 18288 16640 18294 16652
rect 18509 16643 18567 16649
rect 18509 16640 18521 16643
rect 18288 16612 18521 16640
rect 18288 16600 18294 16612
rect 18509 16609 18521 16612
rect 18555 16609 18567 16643
rect 18509 16603 18567 16609
rect 17310 16572 17316 16584
rect 17271 16544 17316 16572
rect 17310 16532 17316 16544
rect 17368 16532 17374 16584
rect 2406 16504 2412 16516
rect 2056 16476 2412 16504
rect 2406 16464 2412 16476
rect 2464 16504 2470 16516
rect 2961 16507 3019 16513
rect 2961 16504 2973 16507
rect 2464 16476 2973 16504
rect 2464 16464 2470 16476
rect 2961 16473 2973 16476
rect 3007 16473 3019 16507
rect 2961 16467 3019 16473
rect 4154 16464 4160 16516
rect 4212 16504 4218 16516
rect 8018 16504 8024 16516
rect 4212 16476 8024 16504
rect 4212 16464 4218 16476
rect 8018 16464 8024 16476
rect 8076 16504 8082 16516
rect 8205 16507 8263 16513
rect 8205 16504 8217 16507
rect 8076 16476 8217 16504
rect 8076 16464 8082 16476
rect 8205 16473 8217 16476
rect 8251 16473 8263 16507
rect 8205 16467 8263 16473
rect 10870 16464 10876 16516
rect 10928 16504 10934 16516
rect 11054 16504 11060 16516
rect 10928 16476 11060 16504
rect 10928 16464 10934 16476
rect 11054 16464 11060 16476
rect 11112 16504 11118 16516
rect 16114 16504 16120 16516
rect 11112 16476 16120 16504
rect 11112 16464 11118 16476
rect 16114 16464 16120 16476
rect 16172 16464 16178 16516
rect 3878 16436 3884 16448
rect 3839 16408 3884 16436
rect 3878 16396 3884 16408
rect 3936 16396 3942 16448
rect 6135 16439 6193 16445
rect 6135 16405 6147 16439
rect 6181 16436 6193 16439
rect 6270 16436 6276 16448
rect 6181 16408 6276 16436
rect 6181 16405 6193 16408
rect 6135 16399 6193 16405
rect 6270 16396 6276 16408
rect 6328 16396 6334 16448
rect 9033 16439 9091 16445
rect 9033 16405 9045 16439
rect 9079 16436 9091 16439
rect 9306 16436 9312 16448
rect 9079 16408 9312 16436
rect 9079 16405 9091 16408
rect 9033 16399 9091 16405
rect 9306 16396 9312 16408
rect 9364 16396 9370 16448
rect 1104 16346 22816 16368
rect 1104 16294 4982 16346
rect 5034 16294 5046 16346
rect 5098 16294 5110 16346
rect 5162 16294 5174 16346
rect 5226 16294 12982 16346
rect 13034 16294 13046 16346
rect 13098 16294 13110 16346
rect 13162 16294 13174 16346
rect 13226 16294 20982 16346
rect 21034 16294 21046 16346
rect 21098 16294 21110 16346
rect 21162 16294 21174 16346
rect 21226 16294 22816 16346
rect 1104 16272 22816 16294
rect 106 16192 112 16244
rect 164 16232 170 16244
rect 5350 16232 5356 16244
rect 164 16204 4154 16232
rect 5263 16204 5356 16232
rect 164 16192 170 16204
rect 3878 16164 3884 16176
rect 3839 16136 3884 16164
rect 3878 16124 3884 16136
rect 3936 16124 3942 16176
rect 4126 16164 4154 16204
rect 5350 16192 5356 16204
rect 5408 16232 5414 16244
rect 6638 16232 6644 16244
rect 5408 16204 6644 16232
rect 5408 16192 5414 16204
rect 6638 16192 6644 16204
rect 6696 16192 6702 16244
rect 8849 16235 8907 16241
rect 8849 16201 8861 16235
rect 8895 16232 8907 16235
rect 9122 16232 9128 16244
rect 8895 16204 9128 16232
rect 8895 16201 8907 16204
rect 8849 16195 8907 16201
rect 9122 16192 9128 16204
rect 9180 16232 9186 16244
rect 9766 16232 9772 16244
rect 9180 16204 9772 16232
rect 9180 16192 9186 16204
rect 9766 16192 9772 16204
rect 9824 16192 9830 16244
rect 10318 16192 10324 16244
rect 10376 16232 10382 16244
rect 15013 16235 15071 16241
rect 10376 16204 13814 16232
rect 10376 16192 10382 16204
rect 6086 16164 6092 16176
rect 4126 16136 6092 16164
rect 6086 16124 6092 16136
rect 6144 16124 6150 16176
rect 8478 16124 8484 16176
rect 8536 16164 8542 16176
rect 9398 16164 9404 16176
rect 8536 16136 9404 16164
rect 8536 16124 8542 16136
rect 9398 16124 9404 16136
rect 9456 16164 9462 16176
rect 10045 16167 10103 16173
rect 10045 16164 10057 16167
rect 9456 16136 10057 16164
rect 9456 16124 9462 16136
rect 10045 16133 10057 16136
rect 10091 16164 10103 16167
rect 10410 16164 10416 16176
rect 10091 16136 10416 16164
rect 10091 16133 10103 16136
rect 10045 16127 10103 16133
rect 10410 16124 10416 16136
rect 10468 16124 10474 16176
rect 13786 16164 13814 16204
rect 15013 16201 15025 16235
rect 15059 16232 15071 16235
rect 15838 16232 15844 16244
rect 15059 16204 15844 16232
rect 15059 16201 15071 16204
rect 15013 16195 15071 16201
rect 15838 16192 15844 16204
rect 15896 16192 15902 16244
rect 16114 16232 16120 16244
rect 16075 16204 16120 16232
rect 16114 16192 16120 16204
rect 16172 16192 16178 16244
rect 20119 16235 20177 16241
rect 20119 16201 20131 16235
rect 20165 16232 20177 16235
rect 20806 16232 20812 16244
rect 20165 16204 20812 16232
rect 20165 16201 20177 16204
rect 20119 16195 20177 16201
rect 20806 16192 20812 16204
rect 20864 16192 20870 16244
rect 18690 16164 18696 16176
rect 13786 16136 16344 16164
rect 18651 16136 18696 16164
rect 2038 16096 2044 16108
rect 1999 16068 2044 16096
rect 2038 16056 2044 16068
rect 2096 16056 2102 16108
rect 2406 16096 2412 16108
rect 2367 16068 2412 16096
rect 2406 16056 2412 16068
rect 2464 16056 2470 16108
rect 3605 16099 3663 16105
rect 3605 16065 3617 16099
rect 3651 16096 3663 16099
rect 4154 16096 4160 16108
rect 3651 16068 4160 16096
rect 3651 16065 3663 16068
rect 3605 16059 3663 16065
rect 4154 16056 4160 16068
rect 4212 16056 4218 16108
rect 4433 16099 4491 16105
rect 4433 16065 4445 16099
rect 4479 16096 4491 16099
rect 4614 16096 4620 16108
rect 4479 16068 4620 16096
rect 4479 16065 4491 16068
rect 4433 16059 4491 16065
rect 4614 16056 4620 16068
rect 4672 16096 4678 16108
rect 5629 16099 5687 16105
rect 5629 16096 5641 16099
rect 4672 16068 5641 16096
rect 4672 16056 4678 16068
rect 5629 16065 5641 16068
rect 5675 16065 5687 16099
rect 8754 16096 8760 16108
rect 5629 16059 5687 16065
rect 7116 16068 8760 16096
rect 4338 15988 4344 16040
rect 4396 16028 4402 16040
rect 7116 16037 7144 16068
rect 8754 16056 8760 16068
rect 8812 16056 8818 16108
rect 9033 16099 9091 16105
rect 9033 16065 9045 16099
rect 9079 16096 9091 16099
rect 9306 16096 9312 16108
rect 9079 16068 9312 16096
rect 9079 16065 9091 16068
rect 9033 16059 9091 16065
rect 9306 16056 9312 16068
rect 9364 16056 9370 16108
rect 10428 16096 10456 16124
rect 12253 16099 12311 16105
rect 10428 16068 11008 16096
rect 6641 16031 6699 16037
rect 4396 16000 4844 16028
rect 4396 15988 4402 16000
rect 2133 15963 2191 15969
rect 2133 15929 2145 15963
rect 2179 15929 2191 15963
rect 2133 15923 2191 15929
rect 1854 15892 1860 15904
rect 1815 15864 1860 15892
rect 1854 15852 1860 15864
rect 1912 15892 1918 15904
rect 2148 15892 2176 15923
rect 3878 15920 3884 15972
rect 3936 15960 3942 15972
rect 4614 15960 4620 15972
rect 3936 15932 4620 15960
rect 3936 15920 3942 15932
rect 4614 15920 4620 15932
rect 4672 15920 4678 15972
rect 4816 15969 4844 16000
rect 6641 15997 6653 16031
rect 6687 16028 6699 16031
rect 7101 16031 7159 16037
rect 7101 16028 7113 16031
rect 6687 16000 7113 16028
rect 6687 15997 6699 16000
rect 6641 15991 6699 15997
rect 7101 15997 7113 16000
rect 7147 15997 7159 16031
rect 7101 15991 7159 15997
rect 7190 15988 7196 16040
rect 7248 16028 7254 16040
rect 7285 16031 7343 16037
rect 7285 16028 7297 16031
rect 7248 16000 7297 16028
rect 7248 15988 7254 16000
rect 7285 15997 7297 16000
rect 7331 15997 7343 16031
rect 7837 16031 7895 16037
rect 7837 16028 7849 16031
rect 7285 15991 7343 15997
rect 7392 16000 7849 16028
rect 4795 15963 4853 15969
rect 4795 15929 4807 15963
rect 4841 15960 4853 15963
rect 7392 15960 7420 16000
rect 7837 15997 7849 16000
rect 7883 16028 7895 16031
rect 8386 16028 8392 16040
rect 7883 16000 8392 16028
rect 7883 15997 7895 16000
rect 7837 15991 7895 15997
rect 8386 15988 8392 16000
rect 8444 15988 8450 16040
rect 10778 16028 10784 16040
rect 10739 16000 10784 16028
rect 10778 15988 10784 16000
rect 10836 15988 10842 16040
rect 10980 16037 11008 16068
rect 12253 16065 12265 16099
rect 12299 16096 12311 16099
rect 13262 16096 13268 16108
rect 12299 16068 13268 16096
rect 12299 16065 12311 16068
rect 12253 16059 12311 16065
rect 10965 16031 11023 16037
rect 10965 15997 10977 16031
rect 11011 16028 11023 16031
rect 11606 16028 11612 16040
rect 11011 16000 11612 16028
rect 11011 15997 11023 16000
rect 10965 15991 11023 15997
rect 11606 15988 11612 16000
rect 11664 15988 11670 16040
rect 12636 16037 12664 16068
rect 13262 16056 13268 16068
rect 13320 16056 13326 16108
rect 13998 16056 14004 16108
rect 14056 16096 14062 16108
rect 14093 16099 14151 16105
rect 14093 16096 14105 16099
rect 14056 16068 14105 16096
rect 14056 16056 14062 16068
rect 14093 16065 14105 16068
rect 14139 16065 14151 16099
rect 14093 16059 14151 16065
rect 12621 16031 12679 16037
rect 12621 15997 12633 16031
rect 12667 15997 12679 16031
rect 12897 16031 12955 16037
rect 12897 16028 12909 16031
rect 12621 15991 12679 15997
rect 12774 16000 12909 16028
rect 7558 15960 7564 15972
rect 4841 15932 7420 15960
rect 7519 15932 7564 15960
rect 4841 15929 4853 15932
rect 4795 15923 4853 15929
rect 7558 15920 7564 15932
rect 7616 15920 7622 15972
rect 9122 15960 9128 15972
rect 9083 15932 9128 15960
rect 9122 15920 9128 15932
rect 9180 15920 9186 15972
rect 9677 15963 9735 15969
rect 9677 15929 9689 15963
rect 9723 15960 9735 15963
rect 9950 15960 9956 15972
rect 9723 15932 9956 15960
rect 9723 15929 9735 15932
rect 9677 15923 9735 15929
rect 9950 15920 9956 15932
rect 10008 15920 10014 15972
rect 11885 15963 11943 15969
rect 11885 15929 11897 15963
rect 11931 15960 11943 15963
rect 12250 15960 12256 15972
rect 11931 15932 12256 15960
rect 11931 15929 11943 15932
rect 11885 15923 11943 15929
rect 12250 15920 12256 15932
rect 12308 15960 12314 15972
rect 12774 15960 12802 16000
rect 12897 15997 12909 16000
rect 12943 15997 12955 16031
rect 15378 16028 15384 16040
rect 15291 16000 15384 16028
rect 12897 15991 12955 15997
rect 15378 15988 15384 16000
rect 15436 16028 15442 16040
rect 16114 16028 16120 16040
rect 15436 16000 16120 16028
rect 15436 15988 15442 16000
rect 16114 15988 16120 16000
rect 16172 15988 16178 16040
rect 16316 16037 16344 16136
rect 18690 16124 18696 16136
rect 18748 16124 18754 16176
rect 17037 16099 17095 16105
rect 17037 16065 17049 16099
rect 17083 16096 17095 16099
rect 17310 16096 17316 16108
rect 17083 16068 17316 16096
rect 17083 16065 17095 16068
rect 17037 16059 17095 16065
rect 17310 16056 17316 16068
rect 17368 16096 17374 16108
rect 17681 16099 17739 16105
rect 17681 16096 17693 16099
rect 17368 16068 17693 16096
rect 17368 16056 17374 16068
rect 17681 16065 17693 16068
rect 17727 16065 17739 16099
rect 17681 16059 17739 16065
rect 17862 16056 17868 16108
rect 17920 16096 17926 16108
rect 18141 16099 18199 16105
rect 18141 16096 18153 16099
rect 17920 16068 18153 16096
rect 17920 16056 17926 16068
rect 18141 16065 18153 16068
rect 18187 16096 18199 16099
rect 19061 16099 19119 16105
rect 19061 16096 19073 16099
rect 18187 16068 19073 16096
rect 18187 16065 18199 16068
rect 18141 16059 18199 16065
rect 19061 16065 19073 16068
rect 19107 16065 19119 16099
rect 19061 16059 19119 16065
rect 16301 16031 16359 16037
rect 16301 15997 16313 16031
rect 16347 16028 16359 16031
rect 16574 16028 16580 16040
rect 16347 16000 16580 16028
rect 16347 15997 16359 16000
rect 16301 15991 16359 15997
rect 16574 15988 16580 16000
rect 16632 15988 16638 16040
rect 16761 16031 16819 16037
rect 16761 15997 16773 16031
rect 16807 15997 16819 16031
rect 20016 16031 20074 16037
rect 20016 16028 20028 16031
rect 16761 15991 16819 15997
rect 18984 16000 20028 16028
rect 16776 15960 16804 15991
rect 12308 15932 12802 15960
rect 15764 15932 16804 15960
rect 12308 15920 12314 15932
rect 15764 15904 15792 15932
rect 18230 15920 18236 15972
rect 18288 15960 18294 15972
rect 18288 15932 18333 15960
rect 18288 15920 18294 15932
rect 1912 15864 2176 15892
rect 1912 15852 1918 15864
rect 2590 15852 2596 15904
rect 2648 15892 2654 15904
rect 2958 15892 2964 15904
rect 2648 15864 2964 15892
rect 2648 15852 2654 15864
rect 2958 15852 2964 15864
rect 3016 15852 3022 15904
rect 4341 15895 4399 15901
rect 4341 15861 4353 15895
rect 4387 15892 4399 15895
rect 4430 15892 4436 15904
rect 4387 15864 4436 15892
rect 4387 15861 4399 15864
rect 4341 15855 4399 15861
rect 4430 15852 4436 15864
rect 4488 15852 4494 15904
rect 6086 15892 6092 15904
rect 6047 15864 6092 15892
rect 6086 15852 6092 15864
rect 6144 15852 6150 15904
rect 10594 15892 10600 15904
rect 10555 15864 10600 15892
rect 10594 15852 10600 15864
rect 10652 15852 10658 15904
rect 12526 15892 12532 15904
rect 12487 15864 12532 15892
rect 12526 15852 12532 15864
rect 12584 15852 12590 15904
rect 13262 15852 13268 15904
rect 13320 15892 13326 15904
rect 13449 15895 13507 15901
rect 13449 15892 13461 15895
rect 13320 15864 13461 15892
rect 13320 15852 13326 15864
rect 13449 15861 13461 15864
rect 13495 15861 13507 15895
rect 13449 15855 13507 15861
rect 13906 15852 13912 15904
rect 13964 15892 13970 15904
rect 14001 15895 14059 15901
rect 14001 15892 14013 15895
rect 13964 15864 14013 15892
rect 13964 15852 13970 15864
rect 14001 15861 14013 15864
rect 14047 15892 14059 15895
rect 14458 15892 14464 15904
rect 14047 15864 14464 15892
rect 14047 15861 14059 15864
rect 14001 15855 14059 15861
rect 14458 15852 14464 15864
rect 14516 15852 14522 15904
rect 15746 15892 15752 15904
rect 15707 15864 15752 15892
rect 15746 15852 15752 15864
rect 15804 15852 15810 15904
rect 17310 15892 17316 15904
rect 17271 15864 17316 15892
rect 17310 15852 17316 15864
rect 17368 15852 17374 15904
rect 17954 15852 17960 15904
rect 18012 15892 18018 15904
rect 18984 15892 19012 16000
rect 20016 15997 20028 16000
rect 20062 16028 20074 16031
rect 20441 16031 20499 16037
rect 20441 16028 20453 16031
rect 20062 16000 20453 16028
rect 20062 15997 20074 16000
rect 20016 15991 20074 15997
rect 20441 15997 20453 16000
rect 20487 15997 20499 16031
rect 20441 15991 20499 15997
rect 18012 15864 19012 15892
rect 18012 15852 18018 15864
rect 1104 15802 22816 15824
rect 1104 15750 8982 15802
rect 9034 15750 9046 15802
rect 9098 15750 9110 15802
rect 9162 15750 9174 15802
rect 9226 15750 16982 15802
rect 17034 15750 17046 15802
rect 17098 15750 17110 15802
rect 17162 15750 17174 15802
rect 17226 15750 22816 15802
rect 1104 15728 22816 15750
rect 1854 15648 1860 15700
rect 1912 15688 1918 15700
rect 1949 15691 2007 15697
rect 1949 15688 1961 15691
rect 1912 15660 1961 15688
rect 1912 15648 1918 15660
rect 1949 15657 1961 15660
rect 1995 15657 2007 15691
rect 1949 15651 2007 15657
rect 2038 15648 2044 15700
rect 2096 15688 2102 15700
rect 2685 15691 2743 15697
rect 2685 15688 2697 15691
rect 2096 15660 2697 15688
rect 2096 15648 2102 15660
rect 2685 15657 2697 15660
rect 2731 15657 2743 15691
rect 2685 15651 2743 15657
rect 5261 15691 5319 15697
rect 5261 15657 5273 15691
rect 5307 15688 5319 15691
rect 5350 15688 5356 15700
rect 5307 15660 5356 15688
rect 5307 15657 5319 15660
rect 5261 15651 5319 15657
rect 5350 15648 5356 15660
rect 5408 15648 5414 15700
rect 5828 15660 6868 15688
rect 3510 15580 3516 15632
rect 3568 15620 3574 15632
rect 4246 15620 4252 15632
rect 3568 15592 4252 15620
rect 3568 15580 3574 15592
rect 4246 15580 4252 15592
rect 4304 15580 4310 15632
rect 4338 15580 4344 15632
rect 4396 15620 4402 15632
rect 5828 15620 5856 15660
rect 4396 15592 5856 15620
rect 4396 15580 4402 15592
rect 6270 15580 6276 15632
rect 6328 15620 6334 15632
rect 6840 15629 6868 15660
rect 7558 15648 7564 15700
rect 7616 15688 7622 15700
rect 7653 15691 7711 15697
rect 7653 15688 7665 15691
rect 7616 15660 7665 15688
rect 7616 15648 7622 15660
rect 7653 15657 7665 15660
rect 7699 15657 7711 15691
rect 10410 15688 10416 15700
rect 10371 15660 10416 15688
rect 7653 15651 7711 15657
rect 10410 15648 10416 15660
rect 10468 15648 10474 15700
rect 11606 15688 11612 15700
rect 11567 15660 11612 15688
rect 11606 15648 11612 15660
rect 11664 15648 11670 15700
rect 11974 15688 11980 15700
rect 11935 15660 11980 15688
rect 11974 15648 11980 15660
rect 12032 15648 12038 15700
rect 13998 15648 14004 15700
rect 14056 15688 14062 15700
rect 14093 15691 14151 15697
rect 14093 15688 14105 15691
rect 14056 15660 14105 15688
rect 14056 15648 14062 15660
rect 14093 15657 14105 15660
rect 14139 15657 14151 15691
rect 16574 15688 16580 15700
rect 16535 15660 16580 15688
rect 14093 15651 14151 15657
rect 16574 15648 16580 15660
rect 16632 15648 16638 15700
rect 18049 15691 18107 15697
rect 18049 15657 18061 15691
rect 18095 15688 18107 15691
rect 18230 15688 18236 15700
rect 18095 15660 18236 15688
rect 18095 15657 18107 15660
rect 18049 15651 18107 15657
rect 18230 15648 18236 15660
rect 18288 15688 18294 15700
rect 18325 15691 18383 15697
rect 18325 15688 18337 15691
rect 18288 15660 18337 15688
rect 18288 15648 18294 15660
rect 18325 15657 18337 15660
rect 18371 15657 18383 15691
rect 18325 15651 18383 15657
rect 21085 15691 21143 15697
rect 21085 15657 21097 15691
rect 21131 15688 21143 15691
rect 21450 15688 21456 15700
rect 21131 15660 21456 15688
rect 21131 15657 21143 15660
rect 21085 15651 21143 15657
rect 21450 15648 21456 15660
rect 21508 15648 21514 15700
rect 6733 15623 6791 15629
rect 6733 15620 6745 15623
rect 6328 15592 6745 15620
rect 6328 15580 6334 15592
rect 6733 15589 6745 15592
rect 6779 15589 6791 15623
rect 6733 15583 6791 15589
rect 6825 15623 6883 15629
rect 6825 15589 6837 15623
rect 6871 15620 6883 15623
rect 7006 15620 7012 15632
rect 6871 15592 7012 15620
rect 6871 15589 6883 15592
rect 6825 15583 6883 15589
rect 7006 15580 7012 15592
rect 7064 15580 7070 15632
rect 9953 15623 10011 15629
rect 9953 15589 9965 15623
rect 9999 15620 10011 15623
rect 10318 15620 10324 15632
rect 9999 15592 10324 15620
rect 9999 15589 10011 15592
rect 9953 15583 10011 15589
rect 10318 15580 10324 15592
rect 10376 15580 10382 15632
rect 12799 15623 12857 15629
rect 12799 15589 12811 15623
rect 12845 15620 12857 15623
rect 14458 15620 14464 15632
rect 12845 15592 14464 15620
rect 12845 15589 12857 15592
rect 12799 15583 12857 15589
rect 14458 15580 14464 15592
rect 14516 15620 14522 15632
rect 16850 15620 16856 15632
rect 14516 15592 16856 15620
rect 14516 15580 14522 15592
rect 16850 15580 16856 15592
rect 16908 15620 16914 15632
rect 17310 15620 17316 15632
rect 16908 15592 17316 15620
rect 16908 15580 16914 15592
rect 17310 15580 17316 15592
rect 17368 15620 17374 15632
rect 17450 15623 17508 15629
rect 17450 15620 17462 15623
rect 17368 15592 17462 15620
rect 17368 15580 17374 15592
rect 17450 15589 17462 15592
rect 17496 15589 17508 15623
rect 17450 15583 17508 15589
rect 2317 15555 2375 15561
rect 2317 15521 2329 15555
rect 2363 15552 2375 15555
rect 2498 15552 2504 15564
rect 2363 15524 2504 15552
rect 2363 15521 2375 15524
rect 2317 15515 2375 15521
rect 2498 15512 2504 15524
rect 2556 15512 2562 15564
rect 8205 15555 8263 15561
rect 8205 15521 8217 15555
rect 8251 15552 8263 15555
rect 8294 15552 8300 15564
rect 8251 15524 8300 15552
rect 8251 15521 8263 15524
rect 8205 15515 8263 15521
rect 8294 15512 8300 15524
rect 8352 15512 8358 15564
rect 10045 15555 10103 15561
rect 10045 15521 10057 15555
rect 10091 15552 10103 15555
rect 11698 15552 11704 15564
rect 10091 15524 11704 15552
rect 10091 15521 10103 15524
rect 10045 15515 10103 15521
rect 11698 15512 11704 15524
rect 11756 15512 11762 15564
rect 12437 15555 12495 15561
rect 12437 15521 12449 15555
rect 12483 15552 12495 15555
rect 12526 15552 12532 15564
rect 12483 15524 12532 15552
rect 12483 15521 12495 15524
rect 12437 15515 12495 15521
rect 12526 15512 12532 15524
rect 12584 15512 12590 15564
rect 15102 15552 15108 15564
rect 13786 15524 15108 15552
rect 4246 15484 4252 15496
rect 4207 15456 4252 15484
rect 4246 15444 4252 15456
rect 4304 15444 4310 15496
rect 7374 15484 7380 15496
rect 7335 15456 7380 15484
rect 7374 15444 7380 15456
rect 7432 15444 7438 15496
rect 10778 15444 10784 15496
rect 10836 15484 10842 15496
rect 11333 15487 11391 15493
rect 11333 15484 11345 15487
rect 10836 15456 11345 15484
rect 10836 15444 10842 15456
rect 11333 15453 11345 15456
rect 11379 15484 11391 15487
rect 13786 15484 13814 15524
rect 15102 15512 15108 15524
rect 15160 15552 15166 15564
rect 15565 15555 15623 15561
rect 15565 15552 15577 15555
rect 15160 15524 15577 15552
rect 15160 15512 15166 15524
rect 15565 15521 15577 15524
rect 15611 15521 15623 15555
rect 15565 15515 15623 15521
rect 15746 15512 15752 15564
rect 15804 15552 15810 15564
rect 16025 15555 16083 15561
rect 16025 15552 16037 15555
rect 15804 15524 16037 15552
rect 15804 15512 15810 15524
rect 16025 15521 16037 15524
rect 16071 15521 16083 15555
rect 16025 15515 16083 15521
rect 20806 15512 20812 15564
rect 20864 15552 20870 15564
rect 20901 15555 20959 15561
rect 20901 15552 20913 15555
rect 20864 15524 20913 15552
rect 20864 15512 20870 15524
rect 20901 15521 20913 15524
rect 20947 15521 20959 15555
rect 20901 15515 20959 15521
rect 11379 15456 13814 15484
rect 16301 15487 16359 15493
rect 11379 15453 11391 15456
rect 11333 15447 11391 15453
rect 16301 15453 16313 15487
rect 16347 15484 16359 15487
rect 17129 15487 17187 15493
rect 17129 15484 17141 15487
rect 16347 15456 17141 15484
rect 16347 15453 16359 15456
rect 16301 15447 16359 15453
rect 17129 15453 17141 15456
rect 17175 15484 17187 15487
rect 17494 15484 17500 15496
rect 17175 15456 17500 15484
rect 17175 15453 17187 15456
rect 17129 15447 17187 15453
rect 17494 15444 17500 15456
rect 17552 15444 17558 15496
rect 4798 15416 4804 15428
rect 4759 15388 4804 15416
rect 4798 15376 4804 15388
rect 4856 15376 4862 15428
rect 6086 15376 6092 15428
rect 6144 15416 6150 15428
rect 10686 15416 10692 15428
rect 6144 15388 10692 15416
rect 6144 15376 6150 15388
rect 10686 15376 10692 15388
rect 10744 15376 10750 15428
rect 7926 15308 7932 15360
rect 7984 15348 7990 15360
rect 8343 15351 8401 15357
rect 8343 15348 8355 15351
rect 7984 15320 8355 15348
rect 7984 15308 7990 15320
rect 8343 15317 8355 15320
rect 8389 15317 8401 15351
rect 8754 15348 8760 15360
rect 8715 15320 8760 15348
rect 8343 15311 8401 15317
rect 8754 15308 8760 15320
rect 8812 15308 8818 15360
rect 10502 15308 10508 15360
rect 10560 15348 10566 15360
rect 10965 15351 11023 15357
rect 10965 15348 10977 15351
rect 10560 15320 10977 15348
rect 10560 15308 10566 15320
rect 10965 15317 10977 15320
rect 11011 15317 11023 15351
rect 10965 15311 11023 15317
rect 12434 15308 12440 15360
rect 12492 15348 12498 15360
rect 13357 15351 13415 15357
rect 13357 15348 13369 15351
rect 12492 15320 13369 15348
rect 12492 15308 12498 15320
rect 13357 15317 13369 15320
rect 13403 15348 13415 15351
rect 13446 15348 13452 15360
rect 13403 15320 13452 15348
rect 13403 15317 13415 15320
rect 13357 15311 13415 15317
rect 13446 15308 13452 15320
rect 13504 15308 13510 15360
rect 13725 15351 13783 15357
rect 13725 15317 13737 15351
rect 13771 15348 13783 15351
rect 13814 15348 13820 15360
rect 13771 15320 13820 15348
rect 13771 15317 13783 15320
rect 13725 15311 13783 15317
rect 13814 15308 13820 15320
rect 13872 15308 13878 15360
rect 1104 15258 22816 15280
rect 1104 15206 4982 15258
rect 5034 15206 5046 15258
rect 5098 15206 5110 15258
rect 5162 15206 5174 15258
rect 5226 15206 12982 15258
rect 13034 15206 13046 15258
rect 13098 15206 13110 15258
rect 13162 15206 13174 15258
rect 13226 15206 20982 15258
rect 21034 15206 21046 15258
rect 21098 15206 21110 15258
rect 21162 15206 21174 15258
rect 21226 15206 22816 15258
rect 1104 15184 22816 15206
rect 4249 15147 4307 15153
rect 4249 15113 4261 15147
rect 4295 15144 4307 15147
rect 4338 15144 4344 15156
rect 4295 15116 4344 15144
rect 4295 15113 4307 15116
rect 4249 15107 4307 15113
rect 4338 15104 4344 15116
rect 4396 15104 4402 15156
rect 4522 15104 4528 15156
rect 4580 15144 4586 15156
rect 4617 15147 4675 15153
rect 4617 15144 4629 15147
rect 4580 15116 4629 15144
rect 4580 15104 4586 15116
rect 4617 15113 4629 15116
rect 4663 15113 4675 15147
rect 6270 15144 6276 15156
rect 6231 15116 6276 15144
rect 4617 15107 4675 15113
rect 2406 15076 2412 15088
rect 2367 15048 2412 15076
rect 2406 15036 2412 15048
rect 2464 15036 2470 15088
rect 1857 15011 1915 15017
rect 1857 14977 1869 15011
rect 1903 15008 1915 15011
rect 3145 15011 3203 15017
rect 3145 15008 3157 15011
rect 1903 14980 3157 15008
rect 1903 14977 1915 14980
rect 1857 14971 1915 14977
rect 3145 14977 3157 14980
rect 3191 15008 3203 15011
rect 3467 15011 3525 15017
rect 3467 15008 3479 15011
rect 3191 14980 3479 15008
rect 3191 14977 3203 14980
rect 3145 14971 3203 14977
rect 3467 14977 3479 14980
rect 3513 14977 3525 15011
rect 4632 15008 4660 15107
rect 6270 15104 6276 15116
rect 6328 15104 6334 15156
rect 6641 15147 6699 15153
rect 6641 15113 6653 15147
rect 6687 15144 6699 15147
rect 7006 15144 7012 15156
rect 6687 15116 7012 15144
rect 6687 15113 6699 15116
rect 6641 15107 6699 15113
rect 7006 15104 7012 15116
rect 7064 15104 7070 15156
rect 11425 15147 11483 15153
rect 11425 15113 11437 15147
rect 11471 15144 11483 15147
rect 11698 15144 11704 15156
rect 11471 15116 11704 15144
rect 11471 15113 11483 15116
rect 11425 15107 11483 15113
rect 11698 15104 11704 15116
rect 11756 15104 11762 15156
rect 13449 15147 13507 15153
rect 13449 15113 13461 15147
rect 13495 15144 13507 15147
rect 13630 15144 13636 15156
rect 13495 15116 13636 15144
rect 13495 15113 13507 15116
rect 13449 15107 13507 15113
rect 13630 15104 13636 15116
rect 13688 15144 13694 15156
rect 14458 15144 14464 15156
rect 13688 15116 14464 15144
rect 13688 15104 13694 15116
rect 14458 15104 14464 15116
rect 14516 15104 14522 15156
rect 15102 15144 15108 15156
rect 15063 15116 15108 15144
rect 15102 15104 15108 15116
rect 15160 15104 15166 15156
rect 17494 15144 17500 15156
rect 17455 15116 17500 15144
rect 17494 15104 17500 15116
rect 17552 15104 17558 15156
rect 21085 15147 21143 15153
rect 21085 15113 21097 15147
rect 21131 15144 21143 15147
rect 21266 15144 21272 15156
rect 21131 15116 21272 15144
rect 21131 15113 21143 15116
rect 21085 15107 21143 15113
rect 21266 15104 21272 15116
rect 21324 15104 21330 15156
rect 4798 15036 4804 15088
rect 4856 15076 4862 15088
rect 4856 15048 5212 15076
rect 4856 15036 4862 15048
rect 5184 15017 5212 15048
rect 7374 15036 7380 15088
rect 7432 15076 7438 15088
rect 7745 15079 7803 15085
rect 7745 15076 7757 15079
rect 7432 15048 7757 15076
rect 7432 15036 7438 15048
rect 7745 15045 7757 15048
rect 7791 15045 7803 15079
rect 13262 15076 13268 15088
rect 7745 15039 7803 15045
rect 10060 15048 13268 15076
rect 4893 15011 4951 15017
rect 4893 15008 4905 15011
rect 4632 14980 4905 15008
rect 3467 14971 3525 14977
rect 4893 14977 4905 14980
rect 4939 14977 4951 15011
rect 4893 14971 4951 14977
rect 5169 15011 5227 15017
rect 5169 14977 5181 15011
rect 5215 14977 5227 15011
rect 5169 14971 5227 14977
rect 7193 15011 7251 15017
rect 7193 14977 7205 15011
rect 7239 15008 7251 15011
rect 7926 15008 7932 15020
rect 7239 14980 7932 15008
rect 7239 14977 7251 14980
rect 7193 14971 7251 14977
rect 7926 14968 7932 14980
rect 7984 14968 7990 15020
rect 8754 14968 8760 15020
rect 8812 15008 8818 15020
rect 10060 15008 10088 15048
rect 13262 15036 13268 15048
rect 13320 15036 13326 15088
rect 13814 15036 13820 15088
rect 13872 15076 13878 15088
rect 15381 15079 15439 15085
rect 15381 15076 15393 15079
rect 13872 15048 15393 15076
rect 13872 15036 13878 15048
rect 15381 15045 15393 15048
rect 15427 15076 15439 15079
rect 15746 15076 15752 15088
rect 15427 15048 15752 15076
rect 15427 15045 15439 15048
rect 15381 15039 15439 15045
rect 15746 15036 15752 15048
rect 15804 15036 15810 15088
rect 16206 15036 16212 15088
rect 16264 15076 16270 15088
rect 20717 15079 20775 15085
rect 20717 15076 20729 15079
rect 16264 15048 20729 15076
rect 16264 15036 16270 15048
rect 20717 15045 20729 15048
rect 20763 15045 20775 15079
rect 20717 15039 20775 15045
rect 8812 14980 10088 15008
rect 10413 15011 10471 15017
rect 8812 14968 8818 14980
rect 8956 14949 8984 14980
rect 10413 14977 10425 15011
rect 10459 15008 10471 15011
rect 11422 15008 11428 15020
rect 10459 14980 11428 15008
rect 10459 14977 10471 14980
rect 10413 14971 10471 14977
rect 11422 14968 11428 14980
rect 11480 15008 11486 15020
rect 11701 15011 11759 15017
rect 11701 15008 11713 15011
rect 11480 14980 11713 15008
rect 11480 14968 11486 14980
rect 11701 14977 11713 14980
rect 11747 14977 11759 15011
rect 11701 14971 11759 14977
rect 11974 14968 11980 15020
rect 12032 15008 12038 15020
rect 12032 14980 15608 15008
rect 12032 14968 12038 14980
rect 15580 14952 15608 14980
rect 3380 14943 3438 14949
rect 3380 14909 3392 14943
rect 3426 14940 3438 14943
rect 8941 14943 8999 14949
rect 3426 14912 3832 14940
rect 3426 14909 3438 14912
rect 3380 14903 3438 14909
rect 1949 14875 2007 14881
rect 1949 14841 1961 14875
rect 1995 14841 2007 14875
rect 1949 14835 2007 14841
rect 1673 14807 1731 14813
rect 1673 14773 1685 14807
rect 1719 14804 1731 14807
rect 1964 14804 1992 14835
rect 3804 14816 3832 14912
rect 8941 14909 8953 14943
rect 8987 14909 8999 14943
rect 8941 14903 8999 14909
rect 9217 14943 9275 14949
rect 9217 14909 9229 14943
rect 9263 14940 9275 14943
rect 9398 14940 9404 14952
rect 9263 14912 9404 14940
rect 9263 14909 9275 14912
rect 9217 14903 9275 14909
rect 9398 14900 9404 14912
rect 9456 14900 9462 14952
rect 12504 14943 12562 14949
rect 12504 14909 12516 14943
rect 12550 14940 12562 14943
rect 12550 14912 12848 14940
rect 12550 14909 12562 14912
rect 12504 14903 12562 14909
rect 4985 14875 5043 14881
rect 4985 14841 4997 14875
rect 5031 14872 5043 14875
rect 5350 14872 5356 14884
rect 5031 14844 5356 14872
rect 5031 14841 5043 14844
rect 4985 14835 5043 14841
rect 5350 14832 5356 14844
rect 5408 14872 5414 14884
rect 7282 14872 7288 14884
rect 5408 14844 7288 14872
rect 5408 14832 5414 14844
rect 7282 14832 7288 14844
rect 7340 14832 7346 14884
rect 8294 14872 8300 14884
rect 8207 14844 8300 14872
rect 8294 14832 8300 14844
rect 8352 14872 8358 14884
rect 8846 14872 8852 14884
rect 8352 14844 8852 14872
rect 8352 14832 8358 14844
rect 8846 14832 8852 14844
rect 8904 14832 8910 14884
rect 9769 14875 9827 14881
rect 9769 14841 9781 14875
rect 9815 14872 9827 14875
rect 10502 14872 10508 14884
rect 9815 14844 10508 14872
rect 9815 14841 9827 14844
rect 9769 14835 9827 14841
rect 10502 14832 10508 14844
rect 10560 14832 10566 14884
rect 10594 14832 10600 14884
rect 10652 14872 10658 14884
rect 11057 14875 11115 14881
rect 11057 14872 11069 14875
rect 10652 14844 11069 14872
rect 10652 14832 10658 14844
rect 11057 14841 11069 14844
rect 11103 14841 11115 14875
rect 11057 14835 11115 14841
rect 12820 14816 12848 14912
rect 13446 14900 13452 14952
rect 13504 14940 13510 14952
rect 13541 14943 13599 14949
rect 13541 14940 13553 14943
rect 13504 14912 13553 14940
rect 13504 14900 13510 14912
rect 13541 14909 13553 14912
rect 13587 14909 13599 14943
rect 15562 14940 15568 14952
rect 15475 14912 15568 14940
rect 13541 14903 13599 14909
rect 15562 14900 15568 14912
rect 15620 14900 15626 14952
rect 15764 14940 15792 15036
rect 16025 14943 16083 14949
rect 16025 14940 16037 14943
rect 15764 14912 16037 14940
rect 16025 14909 16037 14912
rect 16071 14909 16083 14943
rect 20732 14940 20760 15039
rect 20901 14943 20959 14949
rect 20901 14940 20913 14943
rect 20732 14912 20913 14940
rect 16025 14903 16083 14909
rect 20901 14909 20913 14912
rect 20947 14909 20959 14943
rect 20901 14903 20959 14909
rect 13630 14832 13636 14884
rect 13688 14872 13694 14884
rect 13862 14875 13920 14881
rect 13862 14872 13874 14875
rect 13688 14844 13874 14872
rect 13688 14832 13694 14844
rect 13862 14841 13874 14844
rect 13908 14841 13920 14875
rect 13862 14835 13920 14841
rect 16301 14875 16359 14881
rect 16301 14841 16313 14875
rect 16347 14872 16359 14875
rect 16482 14872 16488 14884
rect 16347 14844 16488 14872
rect 16347 14841 16359 14844
rect 16301 14835 16359 14841
rect 16482 14832 16488 14844
rect 16540 14832 16546 14884
rect 19334 14832 19340 14884
rect 19392 14872 19398 14884
rect 20806 14872 20812 14884
rect 19392 14844 20812 14872
rect 19392 14832 19398 14844
rect 20806 14832 20812 14844
rect 20864 14872 20870 14884
rect 21453 14875 21511 14881
rect 21453 14872 21465 14875
rect 20864 14844 21465 14872
rect 20864 14832 20870 14844
rect 21453 14841 21465 14844
rect 21499 14841 21511 14875
rect 21453 14835 21511 14841
rect 2498 14804 2504 14816
rect 1719 14776 2504 14804
rect 1719 14773 1731 14776
rect 1673 14767 1731 14773
rect 2498 14764 2504 14776
rect 2556 14804 2562 14816
rect 2777 14807 2835 14813
rect 2777 14804 2789 14807
rect 2556 14776 2789 14804
rect 2556 14764 2562 14776
rect 2777 14773 2789 14776
rect 2823 14773 2835 14807
rect 3786 14804 3792 14816
rect 3747 14776 3792 14804
rect 2777 14767 2835 14773
rect 3786 14764 3792 14776
rect 3844 14764 3850 14816
rect 8754 14804 8760 14816
rect 8715 14776 8760 14804
rect 8754 14764 8760 14776
rect 8812 14764 8818 14816
rect 10137 14807 10195 14813
rect 10137 14773 10149 14807
rect 10183 14804 10195 14807
rect 10410 14804 10416 14816
rect 10183 14776 10416 14804
rect 10183 14773 10195 14776
rect 10137 14767 10195 14773
rect 10410 14764 10416 14776
rect 10468 14804 10474 14816
rect 12161 14807 12219 14813
rect 12161 14804 12173 14807
rect 10468 14776 12173 14804
rect 10468 14764 10474 14776
rect 12161 14773 12173 14776
rect 12207 14773 12219 14807
rect 12161 14767 12219 14773
rect 12575 14807 12633 14813
rect 12575 14773 12587 14807
rect 12621 14804 12633 14807
rect 12710 14804 12716 14816
rect 12621 14776 12716 14804
rect 12621 14773 12633 14776
rect 12575 14767 12633 14773
rect 12710 14764 12716 14776
rect 12768 14764 12774 14816
rect 12802 14764 12808 14816
rect 12860 14804 12866 14816
rect 12897 14807 12955 14813
rect 12897 14804 12909 14807
rect 12860 14776 12909 14804
rect 12860 14764 12866 14776
rect 12897 14773 12909 14776
rect 12943 14773 12955 14807
rect 12897 14767 12955 14773
rect 14461 14807 14519 14813
rect 14461 14773 14473 14807
rect 14507 14804 14519 14807
rect 14734 14804 14740 14816
rect 14507 14776 14740 14804
rect 14507 14773 14519 14776
rect 14461 14767 14519 14773
rect 14734 14764 14740 14776
rect 14792 14764 14798 14816
rect 16850 14764 16856 14816
rect 16908 14804 16914 14816
rect 17129 14807 17187 14813
rect 17129 14804 17141 14807
rect 16908 14776 17141 14804
rect 16908 14764 16914 14776
rect 17129 14773 17141 14776
rect 17175 14773 17187 14807
rect 17129 14767 17187 14773
rect 1104 14714 22816 14736
rect 1104 14662 8982 14714
rect 9034 14662 9046 14714
rect 9098 14662 9110 14714
rect 9162 14662 9174 14714
rect 9226 14662 16982 14714
rect 17034 14662 17046 14714
rect 17098 14662 17110 14714
rect 17162 14662 17174 14714
rect 17226 14662 22816 14714
rect 1104 14640 22816 14662
rect 1946 14560 1952 14612
rect 2004 14600 2010 14612
rect 2041 14603 2099 14609
rect 2041 14600 2053 14603
rect 2004 14572 2053 14600
rect 2004 14560 2010 14572
rect 2041 14569 2053 14572
rect 2087 14569 2099 14603
rect 2590 14600 2596 14612
rect 2551 14572 2596 14600
rect 2041 14563 2099 14569
rect 2590 14560 2596 14572
rect 2648 14560 2654 14612
rect 4246 14560 4252 14612
rect 4304 14600 4310 14612
rect 4617 14603 4675 14609
rect 4617 14600 4629 14603
rect 4304 14572 4629 14600
rect 4304 14560 4310 14572
rect 4617 14569 4629 14572
rect 4663 14569 4675 14603
rect 4617 14563 4675 14569
rect 7282 14560 7288 14612
rect 7340 14600 7346 14612
rect 7469 14603 7527 14609
rect 7469 14600 7481 14603
rect 7340 14572 7481 14600
rect 7340 14560 7346 14572
rect 7469 14569 7481 14572
rect 7515 14569 7527 14603
rect 7926 14600 7932 14612
rect 7887 14572 7932 14600
rect 7469 14563 7527 14569
rect 7926 14560 7932 14572
rect 7984 14560 7990 14612
rect 9306 14560 9312 14612
rect 9364 14600 9370 14612
rect 11379 14603 11437 14609
rect 11379 14600 11391 14603
rect 9364 14572 11391 14600
rect 9364 14560 9370 14572
rect 11379 14569 11391 14572
rect 11425 14569 11437 14603
rect 12526 14600 12532 14612
rect 12487 14572 12532 14600
rect 11379 14563 11437 14569
rect 12526 14560 12532 14572
rect 12584 14560 12590 14612
rect 15562 14560 15568 14612
rect 15620 14600 15626 14612
rect 15933 14603 15991 14609
rect 15933 14600 15945 14603
rect 15620 14572 15945 14600
rect 15620 14560 15626 14572
rect 15933 14569 15945 14572
rect 15979 14569 15991 14603
rect 15933 14563 15991 14569
rect 4798 14492 4804 14544
rect 4856 14532 4862 14544
rect 4985 14535 5043 14541
rect 4985 14532 4997 14535
rect 4856 14504 4997 14532
rect 4856 14492 4862 14504
rect 4985 14501 4997 14504
rect 5031 14501 5043 14535
rect 4985 14495 5043 14501
rect 5077 14535 5135 14541
rect 5077 14501 5089 14535
rect 5123 14532 5135 14535
rect 5350 14532 5356 14544
rect 5123 14504 5356 14532
rect 5123 14501 5135 14504
rect 5077 14495 5135 14501
rect 5350 14492 5356 14504
rect 5408 14492 5414 14544
rect 6641 14535 6699 14541
rect 6641 14501 6653 14535
rect 6687 14532 6699 14535
rect 6730 14532 6736 14544
rect 6687 14504 6736 14532
rect 6687 14501 6699 14504
rect 6641 14495 6699 14501
rect 6730 14492 6736 14504
rect 6788 14532 6794 14544
rect 8205 14535 8263 14541
rect 8205 14532 8217 14535
rect 6788 14504 8217 14532
rect 6788 14492 6794 14504
rect 8205 14501 8217 14504
rect 8251 14501 8263 14535
rect 8205 14495 8263 14501
rect 9125 14535 9183 14541
rect 9125 14501 9137 14535
rect 9171 14532 9183 14535
rect 9398 14532 9404 14544
rect 9171 14504 9404 14532
rect 9171 14501 9183 14504
rect 9125 14495 9183 14501
rect 9398 14492 9404 14504
rect 9456 14492 9462 14544
rect 9858 14532 9864 14544
rect 9819 14504 9864 14532
rect 9858 14492 9864 14504
rect 9916 14492 9922 14544
rect 10778 14532 10784 14544
rect 10739 14504 10784 14532
rect 10778 14492 10784 14504
rect 10836 14492 10842 14544
rect 12434 14492 12440 14544
rect 12492 14532 12498 14544
rect 12805 14535 12863 14541
rect 12805 14532 12817 14535
rect 12492 14504 12817 14532
rect 12492 14492 12498 14504
rect 12805 14501 12817 14504
rect 12851 14501 12863 14535
rect 15657 14535 15715 14541
rect 15657 14532 15669 14535
rect 12805 14495 12863 14501
rect 15580 14504 15669 14532
rect 15580 14476 15608 14504
rect 15657 14501 15669 14504
rect 15703 14532 15715 14535
rect 15746 14532 15752 14544
rect 15703 14504 15752 14532
rect 15703 14501 15715 14504
rect 15657 14495 15715 14501
rect 15746 14492 15752 14504
rect 15804 14492 15810 14544
rect 16571 14535 16629 14541
rect 16571 14501 16583 14535
rect 16617 14532 16629 14535
rect 16850 14532 16856 14544
rect 16617 14504 16856 14532
rect 16617 14501 16629 14504
rect 16571 14495 16629 14501
rect 16850 14492 16856 14504
rect 16908 14492 16914 14544
rect 5629 14467 5687 14473
rect 5629 14433 5641 14467
rect 5675 14464 5687 14467
rect 6362 14464 6368 14476
rect 5675 14436 6368 14464
rect 5675 14433 5687 14436
rect 5629 14427 5687 14433
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14396 1731 14399
rect 3234 14396 3240 14408
rect 1719 14368 3240 14396
rect 1719 14365 1731 14368
rect 1673 14359 1731 14365
rect 3234 14356 3240 14368
rect 3292 14356 3298 14408
rect 3878 14356 3884 14408
rect 3936 14396 3942 14408
rect 5644 14396 5672 14427
rect 6362 14424 6368 14436
rect 6420 14424 6426 14476
rect 10686 14424 10692 14476
rect 10744 14464 10750 14476
rect 11308 14467 11366 14473
rect 11308 14464 11320 14467
rect 10744 14436 11320 14464
rect 10744 14424 10750 14436
rect 11308 14433 11320 14436
rect 11354 14464 11366 14467
rect 11790 14464 11796 14476
rect 11354 14436 11796 14464
rect 11354 14433 11366 14436
rect 11308 14427 11366 14433
rect 11790 14424 11796 14436
rect 11848 14424 11854 14476
rect 14090 14424 14096 14476
rect 14148 14464 14154 14476
rect 14220 14467 14278 14473
rect 14220 14464 14232 14467
rect 14148 14436 14232 14464
rect 14148 14424 14154 14436
rect 14220 14433 14232 14436
rect 14266 14433 14278 14467
rect 14220 14427 14278 14433
rect 15562 14424 15568 14476
rect 15620 14424 15626 14476
rect 6549 14399 6607 14405
rect 6549 14396 6561 14399
rect 3936 14368 5672 14396
rect 6288 14368 6561 14396
rect 3936 14356 3942 14368
rect 6288 14272 6316 14368
rect 6549 14365 6561 14368
rect 6595 14365 6607 14399
rect 6822 14396 6828 14408
rect 6783 14368 6828 14396
rect 6549 14359 6607 14365
rect 6822 14356 6828 14368
rect 6880 14356 6886 14408
rect 8110 14396 8116 14408
rect 8071 14368 8116 14396
rect 8110 14356 8116 14368
rect 8168 14356 8174 14408
rect 8389 14399 8447 14405
rect 8389 14365 8401 14399
rect 8435 14365 8447 14399
rect 9766 14396 9772 14408
rect 9727 14368 9772 14396
rect 8389 14359 8447 14365
rect 7374 14288 7380 14340
rect 7432 14328 7438 14340
rect 8404 14328 8432 14359
rect 9766 14356 9772 14368
rect 9824 14356 9830 14408
rect 9950 14356 9956 14408
rect 10008 14396 10014 14408
rect 10045 14399 10103 14405
rect 10045 14396 10057 14399
rect 10008 14368 10057 14396
rect 10008 14356 10014 14368
rect 10045 14365 10057 14368
rect 10091 14396 10103 14399
rect 10594 14396 10600 14408
rect 10091 14368 10600 14396
rect 10091 14365 10103 14368
rect 10045 14359 10103 14365
rect 10594 14356 10600 14368
rect 10652 14356 10658 14408
rect 12158 14356 12164 14408
rect 12216 14396 12222 14408
rect 12710 14396 12716 14408
rect 12216 14368 12716 14396
rect 12216 14356 12222 14368
rect 12710 14356 12716 14368
rect 12768 14356 12774 14408
rect 13357 14399 13415 14405
rect 13357 14365 13369 14399
rect 13403 14396 13415 14399
rect 13538 14396 13544 14408
rect 13403 14368 13544 14396
rect 13403 14365 13415 14368
rect 13357 14359 13415 14365
rect 13538 14356 13544 14368
rect 13596 14396 13602 14408
rect 14918 14396 14924 14408
rect 13596 14368 14924 14396
rect 13596 14356 13602 14368
rect 14918 14356 14924 14368
rect 14976 14356 14982 14408
rect 16209 14399 16267 14405
rect 16209 14365 16221 14399
rect 16255 14396 16267 14399
rect 16482 14396 16488 14408
rect 16255 14368 16488 14396
rect 16255 14365 16267 14368
rect 16209 14359 16267 14365
rect 16482 14356 16488 14368
rect 16540 14356 16546 14408
rect 7432 14300 8432 14328
rect 7432 14288 7438 14300
rect 4246 14260 4252 14272
rect 4207 14232 4252 14260
rect 4246 14220 4252 14232
rect 4304 14220 4310 14272
rect 6270 14260 6276 14272
rect 6231 14232 6276 14260
rect 6270 14220 6276 14232
rect 6328 14220 6334 14272
rect 6362 14220 6368 14272
rect 6420 14260 6426 14272
rect 7650 14260 7656 14272
rect 6420 14232 7656 14260
rect 6420 14220 6426 14232
rect 7650 14220 7656 14232
rect 7708 14220 7714 14272
rect 13446 14220 13452 14272
rect 13504 14260 13510 14272
rect 13633 14263 13691 14269
rect 13633 14260 13645 14263
rect 13504 14232 13645 14260
rect 13504 14220 13510 14232
rect 13633 14229 13645 14232
rect 13679 14229 13691 14263
rect 13633 14223 13691 14229
rect 14323 14263 14381 14269
rect 14323 14229 14335 14263
rect 14369 14260 14381 14263
rect 14642 14260 14648 14272
rect 14369 14232 14648 14260
rect 14369 14229 14381 14232
rect 14323 14223 14381 14229
rect 14642 14220 14648 14232
rect 14700 14220 14706 14272
rect 16574 14220 16580 14272
rect 16632 14260 16638 14272
rect 17129 14263 17187 14269
rect 17129 14260 17141 14263
rect 16632 14232 17141 14260
rect 16632 14220 16638 14232
rect 17129 14229 17141 14232
rect 17175 14260 17187 14263
rect 17586 14260 17592 14272
rect 17175 14232 17592 14260
rect 17175 14229 17187 14232
rect 17129 14223 17187 14229
rect 17586 14220 17592 14232
rect 17644 14220 17650 14272
rect 1104 14170 22816 14192
rect 1104 14118 4982 14170
rect 5034 14118 5046 14170
rect 5098 14118 5110 14170
rect 5162 14118 5174 14170
rect 5226 14118 12982 14170
rect 13034 14118 13046 14170
rect 13098 14118 13110 14170
rect 13162 14118 13174 14170
rect 13226 14118 20982 14170
rect 21034 14118 21046 14170
rect 21098 14118 21110 14170
rect 21162 14118 21174 14170
rect 21226 14118 22816 14170
rect 1104 14096 22816 14118
rect 2498 14056 2504 14068
rect 2459 14028 2504 14056
rect 2498 14016 2504 14028
rect 2556 14016 2562 14068
rect 5169 14059 5227 14065
rect 5169 14025 5181 14059
rect 5215 14056 5227 14059
rect 5350 14056 5356 14068
rect 5215 14028 5356 14056
rect 5215 14025 5227 14028
rect 5169 14019 5227 14025
rect 5350 14016 5356 14028
rect 5408 14056 5414 14068
rect 5445 14059 5503 14065
rect 5445 14056 5457 14059
rect 5408 14028 5457 14056
rect 5408 14016 5414 14028
rect 5445 14025 5457 14028
rect 5491 14025 5503 14059
rect 5445 14019 5503 14025
rect 6549 14059 6607 14065
rect 6549 14025 6561 14059
rect 6595 14056 6607 14059
rect 6730 14056 6736 14068
rect 6595 14028 6736 14056
rect 6595 14025 6607 14028
rect 6549 14019 6607 14025
rect 6730 14016 6736 14028
rect 6788 14056 6794 14068
rect 8021 14059 8079 14065
rect 8021 14056 8033 14059
rect 6788 14028 8033 14056
rect 6788 14016 6794 14028
rect 8021 14025 8033 14028
rect 8067 14025 8079 14059
rect 8021 14019 8079 14025
rect 8110 14016 8116 14068
rect 8168 14056 8174 14068
rect 8389 14059 8447 14065
rect 8389 14056 8401 14059
rect 8168 14028 8401 14056
rect 8168 14016 8174 14028
rect 8389 14025 8401 14028
rect 8435 14025 8447 14059
rect 8389 14019 8447 14025
rect 8478 14016 8484 14068
rect 8536 14056 8542 14068
rect 8665 14059 8723 14065
rect 8665 14056 8677 14059
rect 8536 14028 8677 14056
rect 8536 14016 8542 14028
rect 8665 14025 8677 14028
rect 8711 14056 8723 14059
rect 8757 14059 8815 14065
rect 8757 14056 8769 14059
rect 8711 14028 8769 14056
rect 8711 14025 8723 14028
rect 8665 14019 8723 14025
rect 8757 14025 8769 14028
rect 8803 14025 8815 14059
rect 9858 14056 9864 14068
rect 9771 14028 9864 14056
rect 8757 14019 8815 14025
rect 9858 14016 9864 14028
rect 9916 14056 9922 14068
rect 10137 14059 10195 14065
rect 10137 14056 10149 14059
rect 9916 14028 10149 14056
rect 9916 14016 9922 14028
rect 10137 14025 10149 14028
rect 10183 14025 10195 14059
rect 11790 14056 11796 14068
rect 11751 14028 11796 14056
rect 10137 14019 10195 14025
rect 11790 14016 11796 14028
rect 11848 14016 11854 14068
rect 12250 14056 12256 14068
rect 12211 14028 12256 14056
rect 12250 14016 12256 14028
rect 12308 14016 12314 14068
rect 6178 13948 6184 14000
rect 6236 13988 6242 14000
rect 9398 13988 9404 14000
rect 6236 13960 9404 13988
rect 6236 13948 6242 13960
rect 9398 13948 9404 13960
rect 9456 13948 9462 14000
rect 4246 13920 4252 13932
rect 4207 13892 4252 13920
rect 4246 13880 4252 13892
rect 4304 13880 4310 13932
rect 7009 13923 7067 13929
rect 7009 13889 7021 13923
rect 7055 13920 7067 13923
rect 7374 13920 7380 13932
rect 7055 13892 7380 13920
rect 7055 13889 7067 13892
rect 7009 13883 7067 13889
rect 7374 13880 7380 13892
rect 7432 13880 7438 13932
rect 7650 13920 7656 13932
rect 7611 13892 7656 13920
rect 7650 13880 7656 13892
rect 7708 13880 7714 13932
rect 8754 13880 8760 13932
rect 8812 13920 8818 13932
rect 8941 13923 8999 13929
rect 8941 13920 8953 13923
rect 8812 13892 8953 13920
rect 8812 13880 8818 13892
rect 8941 13889 8953 13892
rect 8987 13889 8999 13923
rect 8941 13883 8999 13889
rect 10778 13880 10784 13932
rect 10836 13920 10842 13932
rect 12268 13920 12296 14016
rect 16301 13991 16359 13997
rect 16301 13957 16313 13991
rect 16347 13988 16359 13991
rect 16850 13988 16856 14000
rect 16347 13960 16856 13988
rect 16347 13957 16359 13960
rect 16301 13951 16359 13957
rect 16850 13948 16856 13960
rect 16908 13948 16914 14000
rect 13446 13920 13452 13932
rect 10836 13892 10916 13920
rect 10836 13880 10842 13892
rect 1581 13855 1639 13861
rect 1581 13821 1593 13855
rect 1627 13852 1639 13855
rect 2038 13852 2044 13864
rect 1627 13824 2044 13852
rect 1627 13821 1639 13824
rect 1581 13815 1639 13821
rect 2038 13812 2044 13824
rect 2096 13812 2102 13864
rect 4065 13855 4123 13861
rect 4065 13852 4077 13855
rect 2792 13824 4077 13852
rect 1946 13793 1952 13796
rect 1922 13787 1952 13793
rect 1922 13784 1934 13787
rect 1859 13756 1934 13784
rect 1922 13753 1934 13756
rect 2004 13784 2010 13796
rect 2792 13793 2820 13824
rect 4065 13821 4077 13824
rect 4111 13852 4123 13855
rect 4430 13852 4436 13864
rect 4111 13824 4436 13852
rect 4111 13821 4123 13824
rect 4065 13815 4123 13821
rect 4430 13812 4436 13824
rect 4488 13852 4494 13864
rect 10888 13861 10916 13892
rect 11256 13892 13216 13920
rect 13407 13892 13452 13920
rect 10873 13855 10931 13861
rect 4488 13824 4613 13852
rect 4488 13812 4494 13824
rect 2777 13787 2835 13793
rect 2777 13784 2789 13787
rect 2004 13756 2789 13784
rect 1922 13747 1952 13753
rect 1946 13744 1952 13747
rect 2004 13744 2010 13756
rect 2777 13753 2789 13756
rect 2823 13753 2835 13787
rect 3234 13784 3240 13796
rect 3195 13756 3240 13784
rect 2777 13747 2835 13753
rect 3234 13744 3240 13756
rect 3292 13744 3298 13796
rect 4585 13793 4613 13824
rect 10873 13821 10885 13855
rect 10919 13852 10931 13855
rect 10962 13852 10968 13864
rect 10919 13824 10968 13852
rect 10919 13821 10931 13824
rect 10873 13815 10931 13821
rect 10962 13812 10968 13824
rect 11020 13812 11026 13864
rect 11256 13861 11284 13892
rect 11241 13855 11299 13861
rect 11241 13821 11253 13855
rect 11287 13821 11299 13855
rect 11241 13815 11299 13821
rect 4570 13787 4628 13793
rect 4570 13753 4582 13787
rect 4616 13753 4628 13787
rect 4570 13747 4628 13753
rect 6181 13787 6239 13793
rect 6181 13753 6193 13787
rect 6227 13784 6239 13787
rect 7101 13787 7159 13793
rect 7101 13784 7113 13787
rect 6227 13756 7113 13784
rect 6227 13753 6239 13756
rect 6181 13747 6239 13753
rect 7101 13753 7113 13756
rect 7147 13784 7159 13787
rect 7282 13784 7288 13796
rect 7147 13756 7288 13784
rect 7147 13753 7159 13756
rect 7101 13747 7159 13753
rect 7282 13744 7288 13756
rect 7340 13744 7346 13796
rect 8665 13787 8723 13793
rect 8665 13753 8677 13787
rect 8711 13784 8723 13787
rect 9262 13787 9320 13793
rect 9262 13784 9274 13787
rect 8711 13756 9274 13784
rect 8711 13753 8723 13756
rect 8665 13747 8723 13753
rect 9262 13753 9274 13756
rect 9308 13784 9320 13787
rect 10689 13787 10747 13793
rect 9308 13756 9674 13784
rect 9308 13753 9320 13756
rect 9262 13747 9320 13753
rect 4798 13676 4804 13728
rect 4856 13716 4862 13728
rect 5626 13716 5632 13728
rect 4856 13688 5632 13716
rect 4856 13676 4862 13688
rect 5626 13676 5632 13688
rect 5684 13716 5690 13728
rect 6822 13716 6828 13728
rect 5684 13688 6828 13716
rect 5684 13676 5690 13688
rect 6822 13676 6828 13688
rect 6880 13676 6886 13728
rect 9646 13716 9674 13756
rect 10689 13753 10701 13787
rect 10735 13784 10747 13787
rect 11256 13784 11284 13815
rect 12618 13812 12624 13864
rect 12676 13852 12682 13864
rect 13188 13861 13216 13892
rect 13446 13880 13452 13892
rect 13504 13880 13510 13932
rect 14642 13920 14648 13932
rect 14603 13892 14648 13920
rect 14642 13880 14648 13892
rect 14700 13880 14706 13932
rect 14918 13920 14924 13932
rect 14879 13892 14924 13920
rect 14918 13880 14924 13892
rect 14976 13880 14982 13932
rect 15933 13923 15991 13929
rect 15933 13889 15945 13923
rect 15979 13920 15991 13923
rect 16574 13920 16580 13932
rect 15979 13892 16580 13920
rect 15979 13889 15991 13892
rect 15933 13883 15991 13889
rect 16574 13880 16580 13892
rect 16632 13880 16638 13932
rect 16666 13880 16672 13932
rect 16724 13920 16730 13932
rect 16724 13892 17172 13920
rect 16724 13880 16730 13892
rect 17144 13861 17172 13892
rect 12713 13855 12771 13861
rect 12713 13852 12725 13855
rect 12676 13824 12725 13852
rect 12676 13812 12682 13824
rect 12713 13821 12725 13824
rect 12759 13852 12771 13855
rect 13173 13855 13231 13861
rect 12759 13824 13032 13852
rect 12759 13821 12771 13824
rect 12713 13815 12771 13821
rect 11514 13784 11520 13796
rect 10735 13756 11284 13784
rect 11475 13756 11520 13784
rect 10735 13753 10747 13756
rect 10689 13747 10747 13753
rect 11514 13744 11520 13756
rect 11572 13744 11578 13796
rect 13004 13784 13032 13824
rect 13173 13821 13185 13855
rect 13219 13821 13231 13855
rect 13173 13815 13231 13821
rect 17129 13855 17187 13861
rect 17129 13821 17141 13855
rect 17175 13852 17187 13855
rect 18322 13852 18328 13864
rect 17175 13824 18328 13852
rect 17175 13821 17187 13824
rect 17129 13815 17187 13821
rect 18322 13812 18328 13824
rect 18380 13812 18386 13864
rect 13817 13787 13875 13793
rect 13817 13784 13829 13787
rect 13004 13756 13829 13784
rect 13817 13753 13829 13756
rect 13863 13753 13875 13787
rect 13817 13747 13875 13753
rect 10410 13716 10416 13728
rect 9646 13688 10416 13716
rect 10410 13676 10416 13688
rect 10468 13676 10474 13728
rect 13832 13716 13860 13747
rect 14090 13744 14096 13796
rect 14148 13784 14154 13796
rect 14185 13787 14243 13793
rect 14185 13784 14197 13787
rect 14148 13756 14197 13784
rect 14148 13744 14154 13756
rect 14185 13753 14197 13756
rect 14231 13753 14243 13787
rect 14734 13784 14740 13796
rect 14695 13756 14740 13784
rect 14185 13747 14243 13753
rect 14734 13744 14740 13756
rect 14792 13744 14798 13796
rect 16485 13787 16543 13793
rect 16485 13753 16497 13787
rect 16531 13753 16543 13787
rect 16485 13747 16543 13753
rect 15930 13716 15936 13728
rect 13832 13688 15936 13716
rect 15930 13676 15936 13688
rect 15988 13676 15994 13728
rect 16500 13716 16528 13747
rect 16574 13744 16580 13796
rect 16632 13784 16638 13796
rect 16632 13756 16677 13784
rect 16632 13744 16638 13756
rect 17494 13716 17500 13728
rect 16500 13688 17500 13716
rect 17494 13676 17500 13688
rect 17552 13676 17558 13728
rect 1104 13626 22816 13648
rect 1104 13574 8982 13626
rect 9034 13574 9046 13626
rect 9098 13574 9110 13626
rect 9162 13574 9174 13626
rect 9226 13574 16982 13626
rect 17034 13574 17046 13626
rect 17098 13574 17110 13626
rect 17162 13574 17174 13626
rect 17226 13574 22816 13626
rect 1104 13552 22816 13574
rect 106 13472 112 13524
rect 164 13512 170 13524
rect 1581 13515 1639 13521
rect 1581 13512 1593 13515
rect 164 13484 1593 13512
rect 164 13472 170 13484
rect 1581 13481 1593 13484
rect 1627 13481 1639 13515
rect 1581 13475 1639 13481
rect 2639 13515 2697 13521
rect 2639 13481 2651 13515
rect 2685 13512 2697 13515
rect 2774 13512 2780 13524
rect 2685 13484 2780 13512
rect 2685 13481 2697 13484
rect 2639 13475 2697 13481
rect 2774 13472 2780 13484
rect 2832 13472 2838 13524
rect 4246 13512 4252 13524
rect 4207 13484 4252 13512
rect 4246 13472 4252 13484
rect 4304 13472 4310 13524
rect 5626 13512 5632 13524
rect 5587 13484 5632 13512
rect 5626 13472 5632 13484
rect 5684 13472 5690 13524
rect 6638 13472 6644 13524
rect 6696 13512 6702 13524
rect 6733 13515 6791 13521
rect 6733 13512 6745 13515
rect 6696 13484 6745 13512
rect 6696 13472 6702 13484
rect 6733 13481 6745 13484
rect 6779 13481 6791 13515
rect 7282 13512 7288 13524
rect 7243 13484 7288 13512
rect 6733 13475 6791 13481
rect 7282 13472 7288 13484
rect 7340 13472 7346 13524
rect 7374 13472 7380 13524
rect 7432 13512 7438 13524
rect 7561 13515 7619 13521
rect 7561 13512 7573 13515
rect 7432 13484 7573 13512
rect 7432 13472 7438 13484
rect 7561 13481 7573 13484
rect 7607 13481 7619 13515
rect 7561 13475 7619 13481
rect 8110 13472 8116 13524
rect 8168 13512 8174 13524
rect 8251 13515 8309 13521
rect 8251 13512 8263 13515
rect 8168 13484 8263 13512
rect 8168 13472 8174 13484
rect 8251 13481 8263 13484
rect 8297 13481 8309 13515
rect 8251 13475 8309 13481
rect 8754 13472 8760 13524
rect 8812 13512 8818 13524
rect 8941 13515 8999 13521
rect 8941 13512 8953 13515
rect 8812 13484 8953 13512
rect 8812 13472 8818 13484
rect 8941 13481 8953 13484
rect 8987 13481 8999 13515
rect 12158 13512 12164 13524
rect 12119 13484 12164 13512
rect 8941 13475 8999 13481
rect 12158 13472 12164 13484
rect 12216 13472 12222 13524
rect 12434 13512 12440 13524
rect 12395 13484 12440 13512
rect 12434 13472 12440 13484
rect 12492 13472 12498 13524
rect 13630 13512 13636 13524
rect 12998 13484 13636 13512
rect 10686 13444 10692 13456
rect 10647 13416 10692 13444
rect 10686 13404 10692 13416
rect 10744 13404 10750 13456
rect 11238 13444 11244 13456
rect 11199 13416 11244 13444
rect 11238 13404 11244 13416
rect 11296 13404 11302 13456
rect 12710 13404 12716 13456
rect 12768 13444 12774 13456
rect 12998 13453 13026 13484
rect 13630 13472 13636 13484
rect 13688 13472 13694 13524
rect 14645 13515 14703 13521
rect 14645 13481 14657 13515
rect 14691 13512 14703 13515
rect 14734 13512 14740 13524
rect 14691 13484 14740 13512
rect 14691 13481 14703 13484
rect 14645 13475 14703 13481
rect 14734 13472 14740 13484
rect 14792 13472 14798 13524
rect 16482 13512 16488 13524
rect 16443 13484 16488 13512
rect 16482 13472 16488 13484
rect 16540 13472 16546 13524
rect 17589 13515 17647 13521
rect 17589 13481 17601 13515
rect 17635 13512 17647 13515
rect 21082 13512 21088 13524
rect 17635 13484 18644 13512
rect 21043 13484 21088 13512
rect 17635 13481 17647 13484
rect 17589 13475 17647 13481
rect 12983 13447 13041 13453
rect 12983 13444 12995 13447
rect 12768 13416 12995 13444
rect 12768 13404 12774 13416
rect 12983 13413 12995 13416
rect 13029 13413 13041 13447
rect 12983 13407 13041 13413
rect 16850 13404 16856 13456
rect 16908 13444 16914 13456
rect 18616 13453 18644 13484
rect 21082 13472 21088 13484
rect 21140 13472 21146 13524
rect 16990 13447 17048 13453
rect 16990 13444 17002 13447
rect 16908 13416 17002 13444
rect 16908 13404 16914 13416
rect 16990 13413 17002 13416
rect 17036 13413 17048 13447
rect 16990 13407 17048 13413
rect 18601 13447 18659 13453
rect 18601 13413 18613 13447
rect 18647 13444 18659 13447
rect 18874 13444 18880 13456
rect 18647 13416 18880 13444
rect 18647 13413 18659 13416
rect 18601 13407 18659 13413
rect 18874 13404 18880 13416
rect 18932 13404 18938 13456
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 1670 13376 1676 13388
rect 1443 13348 1676 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 1670 13336 1676 13348
rect 1728 13336 1734 13388
rect 2568 13379 2626 13385
rect 2568 13345 2580 13379
rect 2614 13376 2626 13379
rect 3142 13376 3148 13388
rect 2614 13348 3148 13376
rect 2614 13345 2626 13348
rect 2568 13339 2626 13345
rect 3142 13336 3148 13348
rect 3200 13336 3206 13388
rect 3694 13336 3700 13388
rect 3752 13376 3758 13388
rect 4157 13379 4215 13385
rect 4157 13376 4169 13379
rect 3752 13348 4169 13376
rect 3752 13336 3758 13348
rect 4157 13345 4169 13348
rect 4203 13345 4215 13379
rect 4706 13376 4712 13388
rect 4667 13348 4712 13376
rect 4157 13339 4215 13345
rect 4706 13336 4712 13348
rect 4764 13336 4770 13388
rect 8113 13379 8171 13385
rect 8113 13345 8125 13379
rect 8159 13376 8171 13379
rect 8202 13376 8208 13388
rect 8159 13348 8208 13376
rect 8159 13345 8171 13348
rect 8113 13339 8171 13345
rect 8202 13336 8208 13348
rect 8260 13336 8266 13388
rect 11514 13336 11520 13388
rect 11572 13376 11578 13388
rect 12621 13379 12679 13385
rect 12621 13376 12633 13379
rect 11572 13348 12633 13376
rect 11572 13336 11578 13348
rect 12621 13345 12633 13348
rect 12667 13376 12679 13379
rect 13630 13376 13636 13388
rect 12667 13348 13636 13376
rect 12667 13345 12679 13348
rect 12621 13339 12679 13345
rect 13630 13336 13636 13348
rect 13688 13336 13694 13388
rect 15194 13376 15200 13388
rect 15155 13348 15200 13376
rect 15194 13336 15200 13348
rect 15252 13336 15258 13388
rect 20806 13336 20812 13388
rect 20864 13376 20870 13388
rect 20901 13379 20959 13385
rect 20901 13376 20913 13379
rect 20864 13348 20913 13376
rect 20864 13336 20870 13348
rect 20901 13345 20913 13348
rect 20947 13345 20959 13379
rect 20901 13339 20959 13345
rect 6362 13308 6368 13320
rect 6323 13280 6368 13308
rect 6362 13268 6368 13280
rect 6420 13268 6426 13320
rect 10594 13308 10600 13320
rect 10555 13280 10600 13308
rect 10594 13268 10600 13280
rect 10652 13268 10658 13320
rect 16666 13308 16672 13320
rect 16627 13280 16672 13308
rect 16666 13268 16672 13280
rect 16724 13268 16730 13320
rect 18506 13308 18512 13320
rect 18467 13280 18512 13308
rect 18506 13268 18512 13280
rect 18564 13268 18570 13320
rect 18690 13268 18696 13320
rect 18748 13308 18754 13320
rect 18785 13311 18843 13317
rect 18785 13308 18797 13311
rect 18748 13280 18797 13308
rect 18748 13268 18754 13280
rect 18785 13277 18797 13280
rect 18831 13277 18843 13311
rect 18785 13271 18843 13277
rect 10778 13200 10784 13252
rect 10836 13240 10842 13252
rect 10836 13212 15608 13240
rect 10836 13200 10842 13212
rect 15580 13184 15608 13212
rect 15746 13200 15752 13252
rect 15804 13240 15810 13252
rect 16117 13243 16175 13249
rect 16117 13240 16129 13243
rect 15804 13212 16129 13240
rect 15804 13200 15810 13212
rect 16117 13209 16129 13212
rect 16163 13209 16175 13243
rect 16117 13203 16175 13209
rect 1946 13172 1952 13184
rect 1907 13144 1952 13172
rect 1946 13132 1952 13144
rect 2004 13132 2010 13184
rect 2038 13132 2044 13184
rect 2096 13172 2102 13184
rect 2314 13172 2320 13184
rect 2096 13144 2320 13172
rect 2096 13132 2102 13144
rect 2314 13132 2320 13144
rect 2372 13132 2378 13184
rect 5261 13175 5319 13181
rect 5261 13141 5273 13175
rect 5307 13172 5319 13175
rect 5350 13172 5356 13184
rect 5307 13144 5356 13172
rect 5307 13141 5319 13144
rect 5261 13135 5319 13141
rect 5350 13132 5356 13144
rect 5408 13132 5414 13184
rect 9858 13172 9864 13184
rect 9819 13144 9864 13172
rect 9858 13132 9864 13144
rect 9916 13132 9922 13184
rect 13541 13175 13599 13181
rect 13541 13141 13553 13175
rect 13587 13172 13599 13175
rect 13998 13172 14004 13184
rect 13587 13144 14004 13172
rect 13587 13141 13599 13144
rect 13541 13135 13599 13141
rect 13998 13132 14004 13144
rect 14056 13132 14062 13184
rect 14274 13172 14280 13184
rect 14235 13144 14280 13172
rect 14274 13132 14280 13144
rect 14332 13132 14338 13184
rect 14734 13132 14740 13184
rect 14792 13172 14798 13184
rect 15427 13175 15485 13181
rect 15427 13172 15439 13175
rect 14792 13144 15439 13172
rect 14792 13132 14798 13144
rect 15427 13141 15439 13144
rect 15473 13141 15485 13175
rect 15427 13135 15485 13141
rect 15562 13132 15568 13184
rect 15620 13172 15626 13184
rect 15838 13172 15844 13184
rect 15620 13144 15844 13172
rect 15620 13132 15626 13144
rect 15838 13132 15844 13144
rect 15896 13132 15902 13184
rect 1104 13082 22816 13104
rect 1104 13030 4982 13082
rect 5034 13030 5046 13082
rect 5098 13030 5110 13082
rect 5162 13030 5174 13082
rect 5226 13030 12982 13082
rect 13034 13030 13046 13082
rect 13098 13030 13110 13082
rect 13162 13030 13174 13082
rect 13226 13030 20982 13082
rect 21034 13030 21046 13082
rect 21098 13030 21110 13082
rect 21162 13030 21174 13082
rect 21226 13030 22816 13082
rect 1104 13008 22816 13030
rect 4295 12971 4353 12977
rect 4295 12937 4307 12971
rect 4341 12968 4353 12971
rect 6270 12968 6276 12980
rect 4341 12940 6276 12968
rect 4341 12937 4353 12940
rect 4295 12931 4353 12937
rect 6270 12928 6276 12940
rect 6328 12928 6334 12980
rect 8711 12971 8769 12977
rect 8711 12937 8723 12971
rect 8757 12968 8769 12971
rect 9858 12968 9864 12980
rect 8757 12940 9864 12968
rect 8757 12937 8769 12940
rect 8711 12931 8769 12937
rect 9858 12928 9864 12940
rect 9916 12928 9922 12980
rect 10594 12928 10600 12980
rect 10652 12968 10658 12980
rect 10965 12971 11023 12977
rect 10965 12968 10977 12971
rect 10652 12940 10977 12968
rect 10652 12928 10658 12940
rect 10965 12937 10977 12940
rect 11011 12937 11023 12971
rect 10965 12931 11023 12937
rect 11287 12971 11345 12977
rect 11287 12937 11299 12971
rect 11333 12968 11345 12971
rect 11422 12968 11428 12980
rect 11333 12940 11428 12968
rect 11333 12937 11345 12940
rect 11287 12931 11345 12937
rect 11422 12928 11428 12940
rect 11480 12928 11486 12980
rect 13630 12968 13636 12980
rect 13591 12940 13636 12968
rect 13630 12928 13636 12940
rect 13688 12928 13694 12980
rect 13998 12968 14004 12980
rect 13959 12940 14004 12968
rect 13998 12928 14004 12940
rect 14056 12928 14062 12980
rect 17494 12928 17500 12980
rect 17552 12968 17558 12980
rect 18187 12971 18245 12977
rect 18187 12968 18199 12971
rect 17552 12940 18199 12968
rect 17552 12928 17558 12940
rect 18187 12937 18199 12940
rect 18233 12937 18245 12971
rect 18874 12968 18880 12980
rect 18835 12940 18880 12968
rect 18187 12931 18245 12937
rect 18874 12928 18880 12940
rect 18932 12928 18938 12980
rect 4430 12860 4436 12912
rect 4488 12900 4494 12912
rect 6365 12903 6423 12909
rect 6365 12900 6377 12903
rect 4488 12872 6377 12900
rect 4488 12860 4494 12872
rect 6365 12869 6377 12872
rect 6411 12900 6423 12903
rect 6638 12900 6644 12912
rect 6411 12872 6644 12900
rect 6411 12869 6423 12872
rect 6365 12863 6423 12869
rect 6638 12860 6644 12872
rect 6696 12860 6702 12912
rect 8846 12860 8852 12912
rect 8904 12900 8910 12912
rect 8904 12872 10818 12900
rect 8904 12860 8910 12872
rect 5368 12804 9628 12832
rect 5368 12776 5396 12804
rect 9600 12776 9628 12804
rect 1949 12767 2007 12773
rect 1949 12733 1961 12767
rect 1995 12764 2007 12767
rect 2133 12767 2191 12773
rect 2133 12764 2145 12767
rect 1995 12736 2145 12764
rect 1995 12733 2007 12736
rect 1949 12727 2007 12733
rect 2133 12733 2145 12736
rect 2179 12764 2191 12767
rect 2590 12764 2596 12776
rect 2179 12736 2596 12764
rect 2179 12733 2191 12736
rect 2133 12727 2191 12733
rect 2590 12724 2596 12736
rect 2648 12724 2654 12776
rect 3786 12724 3792 12776
rect 3844 12764 3850 12776
rect 4154 12764 4160 12776
rect 4212 12773 4218 12776
rect 4212 12767 4250 12773
rect 3844 12736 4160 12764
rect 3844 12724 3850 12736
rect 4154 12724 4160 12736
rect 4238 12764 4250 12767
rect 4617 12767 4675 12773
rect 4617 12764 4629 12767
rect 4238 12736 4629 12764
rect 4238 12733 4250 12736
rect 4212 12727 4250 12733
rect 4617 12733 4629 12736
rect 4663 12733 4675 12767
rect 5350 12764 5356 12776
rect 5311 12736 5356 12764
rect 4617 12727 4675 12733
rect 4212 12724 4218 12727
rect 5350 12724 5356 12736
rect 5408 12724 5414 12776
rect 5721 12767 5779 12773
rect 5721 12733 5733 12767
rect 5767 12733 5779 12767
rect 5721 12727 5779 12733
rect 5905 12767 5963 12773
rect 5905 12733 5917 12767
rect 5951 12764 5963 12767
rect 6362 12764 6368 12776
rect 5951 12736 6368 12764
rect 5951 12733 5963 12736
rect 5905 12727 5963 12733
rect 4065 12699 4123 12705
rect 4065 12665 4077 12699
rect 4111 12696 4123 12699
rect 4706 12696 4712 12708
rect 4111 12668 4712 12696
rect 4111 12665 4123 12668
rect 4065 12659 4123 12665
rect 4706 12656 4712 12668
rect 4764 12696 4770 12708
rect 5077 12699 5135 12705
rect 5077 12696 5089 12699
rect 4764 12668 5089 12696
rect 4764 12656 4770 12668
rect 5077 12665 5089 12668
rect 5123 12696 5135 12699
rect 5736 12696 5764 12727
rect 6362 12724 6368 12736
rect 6420 12724 6426 12776
rect 6638 12724 6644 12776
rect 6696 12764 6702 12776
rect 6917 12767 6975 12773
rect 6917 12764 6929 12767
rect 6696 12736 6929 12764
rect 6696 12724 6702 12736
rect 6917 12733 6929 12736
rect 6963 12733 6975 12767
rect 8202 12764 8208 12776
rect 8115 12736 8208 12764
rect 6917 12727 6975 12733
rect 8202 12724 8208 12736
rect 8260 12764 8266 12776
rect 8640 12767 8698 12773
rect 8640 12764 8652 12767
rect 8260 12736 8652 12764
rect 8260 12724 8266 12736
rect 8640 12733 8652 12736
rect 8686 12764 8698 12767
rect 9122 12764 9128 12776
rect 8686 12736 9128 12764
rect 8686 12733 8698 12736
rect 8640 12727 8698 12733
rect 9122 12724 9128 12736
rect 9180 12724 9186 12776
rect 9582 12764 9588 12776
rect 9495 12736 9588 12764
rect 9582 12724 9588 12736
rect 9640 12724 9646 12776
rect 10137 12767 10195 12773
rect 10137 12764 10149 12767
rect 10047 12736 10149 12764
rect 10137 12733 10149 12736
rect 10183 12764 10195 12767
rect 10318 12764 10324 12776
rect 10183 12736 10324 12764
rect 10183 12733 10195 12736
rect 10137 12727 10195 12733
rect 6822 12696 6828 12708
rect 5123 12668 5948 12696
rect 6783 12668 6828 12696
rect 5123 12665 5135 12668
rect 5077 12659 5135 12665
rect 2498 12628 2504 12640
rect 2459 12600 2504 12628
rect 2498 12588 2504 12600
rect 2556 12588 2562 12640
rect 3142 12628 3148 12640
rect 3103 12600 3148 12628
rect 3142 12588 3148 12600
rect 3200 12588 3206 12640
rect 3694 12628 3700 12640
rect 3655 12600 3700 12628
rect 3694 12588 3700 12600
rect 3752 12588 3758 12640
rect 5920 12628 5948 12668
rect 6822 12656 6828 12668
rect 6880 12656 6886 12708
rect 9306 12656 9312 12708
rect 9364 12696 9370 12708
rect 9493 12699 9551 12705
rect 9493 12696 9505 12699
rect 9364 12668 9505 12696
rect 9364 12656 9370 12668
rect 9493 12665 9505 12668
rect 9539 12696 9551 12699
rect 10152 12696 10180 12727
rect 10318 12724 10324 12736
rect 10376 12724 10382 12776
rect 10790 12764 10818 12872
rect 18506 12860 18512 12912
rect 18564 12900 18570 12912
rect 19245 12903 19303 12909
rect 19245 12900 19257 12903
rect 18564 12872 19257 12900
rect 18564 12860 18570 12872
rect 19245 12869 19257 12872
rect 19291 12869 19303 12903
rect 19245 12863 19303 12869
rect 20671 12903 20729 12909
rect 20671 12869 20683 12903
rect 20717 12900 20729 12903
rect 20806 12900 20812 12912
rect 20717 12872 20812 12900
rect 20717 12869 20729 12872
rect 20671 12863 20729 12869
rect 20806 12860 20812 12872
rect 20864 12900 20870 12912
rect 21361 12903 21419 12909
rect 21361 12900 21373 12903
rect 20864 12872 21373 12900
rect 20864 12860 20870 12872
rect 21361 12869 21373 12872
rect 21407 12869 21419 12903
rect 21361 12863 21419 12869
rect 12437 12835 12495 12841
rect 12437 12801 12449 12835
rect 12483 12832 12495 12835
rect 12802 12832 12808 12844
rect 12483 12804 12808 12832
rect 12483 12801 12495 12804
rect 12437 12795 12495 12801
rect 12802 12792 12808 12804
rect 12860 12792 12866 12844
rect 14550 12832 14556 12844
rect 14511 12804 14556 12832
rect 14550 12792 14556 12804
rect 14608 12792 14614 12844
rect 16485 12835 16543 12841
rect 16485 12801 16497 12835
rect 16531 12832 16543 12835
rect 16666 12832 16672 12844
rect 16531 12804 16672 12832
rect 16531 12801 16543 12804
rect 16485 12795 16543 12801
rect 16666 12792 16672 12804
rect 16724 12832 16730 12844
rect 17129 12835 17187 12841
rect 17129 12832 17141 12835
rect 16724 12804 17141 12832
rect 16724 12792 16730 12804
rect 17129 12801 17141 12804
rect 17175 12801 17187 12835
rect 17129 12795 17187 12801
rect 11184 12767 11242 12773
rect 11184 12764 11196 12767
rect 10790 12736 11196 12764
rect 11184 12733 11196 12736
rect 11230 12764 11242 12767
rect 11609 12767 11667 12773
rect 11609 12764 11621 12767
rect 11230 12736 11621 12764
rect 11230 12733 11242 12736
rect 11184 12727 11242 12733
rect 11609 12733 11621 12736
rect 11655 12764 11667 12767
rect 11790 12764 11796 12776
rect 11655 12736 11796 12764
rect 11655 12733 11667 12736
rect 11609 12727 11667 12733
rect 11790 12724 11796 12736
rect 11848 12724 11854 12776
rect 15378 12724 15384 12776
rect 15436 12764 15442 12776
rect 15746 12764 15752 12776
rect 15436 12736 15752 12764
rect 15436 12724 15442 12736
rect 15746 12724 15752 12736
rect 15804 12724 15810 12776
rect 15838 12724 15844 12776
rect 15896 12764 15902 12776
rect 16209 12767 16267 12773
rect 16209 12764 16221 12767
rect 15896 12736 16221 12764
rect 15896 12724 15902 12736
rect 16209 12733 16221 12736
rect 16255 12733 16267 12767
rect 16209 12727 16267 12733
rect 18084 12767 18142 12773
rect 18084 12733 18096 12767
rect 18130 12733 18142 12767
rect 18084 12727 18142 12733
rect 14274 12696 14280 12708
rect 9539 12668 10180 12696
rect 14235 12668 14280 12696
rect 9539 12665 9551 12668
rect 9493 12659 9551 12665
rect 14274 12656 14280 12668
rect 14332 12656 14338 12708
rect 14369 12699 14427 12705
rect 14369 12665 14381 12699
rect 14415 12665 14427 12699
rect 18099 12696 18127 12727
rect 18690 12724 18696 12776
rect 18748 12764 18754 12776
rect 19556 12767 19614 12773
rect 19556 12764 19568 12767
rect 18748 12736 19568 12764
rect 18748 12724 18754 12736
rect 19556 12733 19568 12736
rect 19602 12764 19614 12767
rect 19981 12767 20039 12773
rect 19981 12764 19993 12767
rect 19602 12736 19993 12764
rect 19602 12733 19614 12736
rect 19556 12727 19614 12733
rect 19981 12733 19993 12736
rect 20027 12733 20039 12767
rect 19981 12727 20039 12733
rect 20600 12767 20658 12773
rect 20600 12733 20612 12767
rect 20646 12764 20658 12767
rect 20714 12764 20720 12776
rect 20646 12736 20720 12764
rect 20646 12733 20658 12736
rect 20600 12727 20658 12733
rect 20714 12724 20720 12736
rect 20772 12764 20778 12776
rect 20993 12767 21051 12773
rect 20993 12764 21005 12767
rect 20772 12736 21005 12764
rect 20772 12724 20778 12736
rect 20993 12733 21005 12736
rect 21039 12733 21051 12767
rect 20993 12727 21051 12733
rect 18509 12699 18567 12705
rect 18509 12696 18521 12699
rect 14369 12659 14427 12665
rect 15304 12668 18521 12696
rect 9674 12628 9680 12640
rect 5920 12600 9680 12628
rect 9674 12588 9680 12600
rect 9732 12588 9738 12640
rect 9858 12628 9864 12640
rect 9819 12600 9864 12628
rect 9858 12588 9864 12600
rect 9916 12588 9922 12640
rect 10686 12628 10692 12640
rect 10647 12600 10692 12628
rect 10686 12588 10692 12600
rect 10744 12588 10750 12640
rect 12253 12631 12311 12637
rect 12253 12597 12265 12631
rect 12299 12628 12311 12631
rect 12710 12628 12716 12640
rect 12299 12600 12716 12628
rect 12299 12597 12311 12600
rect 12253 12591 12311 12597
rect 12710 12588 12716 12600
rect 12768 12628 12774 12640
rect 12805 12631 12863 12637
rect 12805 12628 12817 12631
rect 12768 12600 12817 12628
rect 12768 12588 12774 12600
rect 12805 12597 12817 12600
rect 12851 12597 12863 12631
rect 13354 12628 13360 12640
rect 13315 12600 13360 12628
rect 12805 12591 12863 12597
rect 13354 12588 13360 12600
rect 13412 12588 13418 12640
rect 13998 12588 14004 12640
rect 14056 12628 14062 12640
rect 14384 12628 14412 12659
rect 14056 12600 14412 12628
rect 14056 12588 14062 12600
rect 14458 12588 14464 12640
rect 14516 12628 14522 12640
rect 15194 12628 15200 12640
rect 14516 12600 15200 12628
rect 14516 12588 14522 12600
rect 15194 12588 15200 12600
rect 15252 12628 15258 12640
rect 15304 12637 15332 12668
rect 18509 12665 18521 12668
rect 18555 12665 18567 12699
rect 18509 12659 18567 12665
rect 15289 12631 15347 12637
rect 15289 12628 15301 12631
rect 15252 12600 15301 12628
rect 15252 12588 15258 12600
rect 15289 12597 15301 12600
rect 15335 12597 15347 12631
rect 16850 12628 16856 12640
rect 16811 12600 16856 12628
rect 15289 12591 15347 12597
rect 16850 12588 16856 12600
rect 16908 12588 16914 12640
rect 19659 12631 19717 12637
rect 19659 12597 19671 12631
rect 19705 12628 19717 12631
rect 19886 12628 19892 12640
rect 19705 12600 19892 12628
rect 19705 12597 19717 12600
rect 19659 12591 19717 12597
rect 19886 12588 19892 12600
rect 19944 12588 19950 12640
rect 1104 12538 22816 12560
rect 1104 12486 8982 12538
rect 9034 12486 9046 12538
rect 9098 12486 9110 12538
rect 9162 12486 9174 12538
rect 9226 12486 16982 12538
rect 17034 12486 17046 12538
rect 17098 12486 17110 12538
rect 17162 12486 17174 12538
rect 17226 12486 22816 12538
rect 1104 12464 22816 12486
rect 6362 12424 6368 12436
rect 6323 12396 6368 12424
rect 6362 12384 6368 12396
rect 6420 12384 6426 12436
rect 7742 12384 7748 12436
rect 7800 12424 7806 12436
rect 8662 12424 8668 12436
rect 7800 12396 8668 12424
rect 7800 12384 7806 12396
rect 8662 12384 8668 12396
rect 8720 12424 8726 12436
rect 8757 12427 8815 12433
rect 8757 12424 8769 12427
rect 8720 12396 8769 12424
rect 8720 12384 8726 12396
rect 8757 12393 8769 12396
rect 8803 12393 8815 12427
rect 8757 12387 8815 12393
rect 9582 12384 9588 12436
rect 9640 12424 9646 12436
rect 9861 12427 9919 12433
rect 9861 12424 9873 12427
rect 9640 12396 9873 12424
rect 9640 12384 9646 12396
rect 9861 12393 9873 12396
rect 9907 12393 9919 12427
rect 10410 12424 10416 12436
rect 10371 12396 10416 12424
rect 9861 12387 9919 12393
rect 10410 12384 10416 12396
rect 10468 12384 10474 12436
rect 10686 12384 10692 12436
rect 10744 12424 10750 12436
rect 10965 12427 11023 12433
rect 10965 12424 10977 12427
rect 10744 12396 10977 12424
rect 10744 12384 10750 12396
rect 10965 12393 10977 12396
rect 11011 12393 11023 12427
rect 10965 12387 11023 12393
rect 12529 12427 12587 12433
rect 12529 12393 12541 12427
rect 12575 12424 12587 12427
rect 12710 12424 12716 12436
rect 12575 12396 12716 12424
rect 12575 12393 12587 12396
rect 12529 12387 12587 12393
rect 12710 12384 12716 12396
rect 12768 12384 12774 12436
rect 14734 12424 14740 12436
rect 14695 12396 14740 12424
rect 14734 12384 14740 12396
rect 14792 12384 14798 12436
rect 2498 12356 2504 12368
rect 2459 12328 2504 12356
rect 2498 12316 2504 12328
rect 2556 12316 2562 12368
rect 4985 12359 5043 12365
rect 4985 12325 4997 12359
rect 5031 12356 5043 12359
rect 5350 12356 5356 12368
rect 5031 12328 5356 12356
rect 5031 12325 5043 12328
rect 4985 12319 5043 12325
rect 5350 12316 5356 12328
rect 5408 12316 5414 12368
rect 13354 12316 13360 12368
rect 13412 12356 13418 12368
rect 13449 12359 13507 12365
rect 13449 12356 13461 12359
rect 13412 12328 13461 12356
rect 13412 12316 13418 12328
rect 13449 12325 13461 12328
rect 13495 12325 13507 12359
rect 13998 12356 14004 12368
rect 13911 12328 14004 12356
rect 13449 12319 13507 12325
rect 13998 12316 14004 12328
rect 14056 12356 14062 12368
rect 14550 12356 14556 12368
rect 14056 12328 14556 12356
rect 14056 12316 14062 12328
rect 14550 12316 14556 12328
rect 14608 12316 14614 12368
rect 15470 12356 15476 12368
rect 15431 12328 15476 12356
rect 15470 12316 15476 12328
rect 15528 12316 15534 12368
rect 8018 12288 8024 12300
rect 7979 12260 8024 12288
rect 8018 12248 8024 12260
rect 8076 12248 8082 12300
rect 9858 12248 9864 12300
rect 9916 12288 9922 12300
rect 10045 12291 10103 12297
rect 10045 12288 10057 12291
rect 9916 12260 10057 12288
rect 9916 12248 9922 12260
rect 10045 12257 10057 12260
rect 10091 12257 10103 12291
rect 10045 12251 10103 12257
rect 19886 12248 19892 12300
rect 19944 12288 19950 12300
rect 20806 12288 20812 12300
rect 19944 12260 20812 12288
rect 19944 12248 19950 12260
rect 20806 12248 20812 12260
rect 20864 12288 20870 12300
rect 20901 12291 20959 12297
rect 20901 12288 20913 12291
rect 20864 12260 20913 12288
rect 20864 12248 20870 12260
rect 20901 12257 20913 12260
rect 20947 12257 20959 12291
rect 20901 12251 20959 12257
rect 2409 12223 2467 12229
rect 2409 12220 2421 12223
rect 2148 12192 2421 12220
rect 2148 12096 2176 12192
rect 2409 12189 2421 12192
rect 2455 12189 2467 12223
rect 2409 12183 2467 12189
rect 4893 12223 4951 12229
rect 4893 12189 4905 12223
rect 4939 12220 4951 12223
rect 5626 12220 5632 12232
rect 4939 12192 5632 12220
rect 4939 12189 4951 12192
rect 4893 12183 4951 12189
rect 5626 12180 5632 12192
rect 5684 12180 5690 12232
rect 7742 12220 7748 12232
rect 7703 12192 7748 12220
rect 7742 12180 7748 12192
rect 7800 12180 7806 12232
rect 13357 12223 13415 12229
rect 13357 12189 13369 12223
rect 13403 12220 13415 12223
rect 13722 12220 13728 12232
rect 13403 12192 13728 12220
rect 13403 12189 13415 12192
rect 13357 12183 13415 12189
rect 13722 12180 13728 12192
rect 13780 12180 13786 12232
rect 14550 12180 14556 12232
rect 14608 12220 14614 12232
rect 15381 12223 15439 12229
rect 15381 12220 15393 12223
rect 14608 12192 15393 12220
rect 14608 12180 14614 12192
rect 15381 12189 15393 12192
rect 15427 12220 15439 12223
rect 16853 12223 16911 12229
rect 16853 12220 16865 12223
rect 15427 12192 16865 12220
rect 15427 12189 15439 12192
rect 15381 12183 15439 12189
rect 16853 12189 16865 12192
rect 16899 12189 16911 12223
rect 16853 12183 16911 12189
rect 2961 12155 3019 12161
rect 2961 12121 2973 12155
rect 3007 12152 3019 12155
rect 3050 12152 3056 12164
rect 3007 12124 3056 12152
rect 3007 12121 3019 12124
rect 2961 12115 3019 12121
rect 3050 12112 3056 12124
rect 3108 12152 3114 12164
rect 4249 12155 4307 12161
rect 4249 12152 4261 12155
rect 3108 12124 4261 12152
rect 3108 12112 3114 12124
rect 4249 12121 4261 12124
rect 4295 12152 4307 12155
rect 4338 12152 4344 12164
rect 4295 12124 4344 12152
rect 4295 12121 4307 12124
rect 4249 12115 4307 12121
rect 4338 12112 4344 12124
rect 4396 12112 4402 12164
rect 5442 12152 5448 12164
rect 5403 12124 5448 12152
rect 5442 12112 5448 12124
rect 5500 12112 5506 12164
rect 14274 12112 14280 12164
rect 14332 12152 14338 12164
rect 15933 12155 15991 12161
rect 15933 12152 15945 12155
rect 14332 12124 15945 12152
rect 14332 12112 14338 12124
rect 15933 12121 15945 12124
rect 15979 12121 15991 12155
rect 15933 12115 15991 12121
rect 1670 12084 1676 12096
rect 1631 12056 1676 12084
rect 1670 12044 1676 12056
rect 1728 12044 1734 12096
rect 2130 12084 2136 12096
rect 2091 12056 2136 12084
rect 2130 12044 2136 12056
rect 2188 12044 2194 12096
rect 6638 12044 6644 12096
rect 6696 12084 6702 12096
rect 6825 12087 6883 12093
rect 6825 12084 6837 12087
rect 6696 12056 6837 12084
rect 6696 12044 6702 12056
rect 6825 12053 6837 12056
rect 6871 12053 6883 12087
rect 7190 12084 7196 12096
rect 7151 12056 7196 12084
rect 6825 12047 6883 12053
rect 7190 12044 7196 12056
rect 7248 12044 7254 12096
rect 12802 12084 12808 12096
rect 12763 12056 12808 12084
rect 12802 12044 12808 12056
rect 12860 12044 12866 12096
rect 21085 12087 21143 12093
rect 21085 12053 21097 12087
rect 21131 12084 21143 12087
rect 23566 12084 23572 12096
rect 21131 12056 23572 12084
rect 21131 12053 21143 12056
rect 21085 12047 21143 12053
rect 23566 12044 23572 12056
rect 23624 12044 23630 12096
rect 1104 11994 22816 12016
rect 1104 11942 4982 11994
rect 5034 11942 5046 11994
rect 5098 11942 5110 11994
rect 5162 11942 5174 11994
rect 5226 11942 12982 11994
rect 13034 11942 13046 11994
rect 13098 11942 13110 11994
rect 13162 11942 13174 11994
rect 13226 11942 20982 11994
rect 21034 11942 21046 11994
rect 21098 11942 21110 11994
rect 21162 11942 21174 11994
rect 21226 11942 22816 11994
rect 1104 11920 22816 11942
rect 1535 11883 1593 11889
rect 1535 11849 1547 11883
rect 1581 11880 1593 11883
rect 2130 11880 2136 11892
rect 1581 11852 2136 11880
rect 1581 11849 1593 11852
rect 1535 11843 1593 11849
rect 2130 11840 2136 11852
rect 2188 11840 2194 11892
rect 2317 11883 2375 11889
rect 2317 11849 2329 11883
rect 2363 11880 2375 11883
rect 2498 11880 2504 11892
rect 2363 11852 2504 11880
rect 2363 11849 2375 11852
rect 2317 11843 2375 11849
rect 2498 11840 2504 11852
rect 2556 11840 2562 11892
rect 5626 11880 5632 11892
rect 5587 11852 5632 11880
rect 5626 11840 5632 11852
rect 5684 11840 5690 11892
rect 6641 11883 6699 11889
rect 6641 11849 6653 11883
rect 6687 11880 6699 11883
rect 6822 11880 6828 11892
rect 6687 11852 6828 11880
rect 6687 11849 6699 11852
rect 6641 11843 6699 11849
rect 6822 11840 6828 11852
rect 6880 11840 6886 11892
rect 7190 11840 7196 11892
rect 7248 11880 7254 11892
rect 7248 11852 8432 11880
rect 7248 11840 7254 11852
rect 8404 11824 8432 11852
rect 9858 11840 9864 11892
rect 9916 11880 9922 11892
rect 9953 11883 10011 11889
rect 9953 11880 9965 11883
rect 9916 11852 9965 11880
rect 9916 11840 9922 11852
rect 9953 11849 9965 11852
rect 9999 11849 10011 11883
rect 9953 11843 10011 11849
rect 11057 11883 11115 11889
rect 11057 11849 11069 11883
rect 11103 11880 11115 11883
rect 11238 11880 11244 11892
rect 11103 11852 11244 11880
rect 11103 11849 11115 11852
rect 11057 11843 11115 11849
rect 3050 11812 3056 11824
rect 3011 11784 3056 11812
rect 3050 11772 3056 11784
rect 3108 11772 3114 11824
rect 3142 11772 3148 11824
rect 3200 11812 3206 11824
rect 8386 11812 8392 11824
rect 3200 11784 7420 11812
rect 8299 11784 8392 11812
rect 3200 11772 3206 11784
rect 7392 11756 7420 11784
rect 8386 11772 8392 11784
rect 8444 11812 8450 11824
rect 8444 11784 8984 11812
rect 8444 11772 8450 11784
rect 4338 11744 4344 11756
rect 4299 11716 4344 11744
rect 4338 11704 4344 11716
rect 4396 11704 4402 11756
rect 4985 11747 5043 11753
rect 4985 11713 4997 11747
rect 5031 11744 5043 11747
rect 5442 11744 5448 11756
rect 5031 11716 5448 11744
rect 5031 11713 5043 11716
rect 4985 11707 5043 11713
rect 5442 11704 5448 11716
rect 5500 11704 5506 11756
rect 7101 11747 7159 11753
rect 7101 11713 7113 11747
rect 7147 11744 7159 11747
rect 7190 11744 7196 11756
rect 7147 11716 7196 11744
rect 7147 11713 7159 11716
rect 7101 11707 7159 11713
rect 7190 11704 7196 11716
rect 7248 11704 7254 11756
rect 7374 11744 7380 11756
rect 7287 11716 7380 11744
rect 7374 11704 7380 11716
rect 7432 11704 7438 11756
rect 8662 11744 8668 11756
rect 8623 11716 8668 11744
rect 8662 11704 8668 11716
rect 8720 11704 8726 11756
rect 8956 11753 8984 11784
rect 8941 11747 8999 11753
rect 8941 11713 8953 11747
rect 8987 11713 8999 11747
rect 8941 11707 8999 11713
rect 1464 11679 1522 11685
rect 1464 11645 1476 11679
rect 1510 11676 1522 11679
rect 10204 11679 10262 11685
rect 1510 11648 1992 11676
rect 1510 11645 1522 11648
rect 1464 11639 1522 11645
rect 1964 11549 1992 11648
rect 10204 11645 10216 11679
rect 10250 11676 10262 11679
rect 11072 11676 11100 11843
rect 11238 11840 11244 11852
rect 11296 11840 11302 11892
rect 12250 11880 12256 11892
rect 12211 11852 12256 11880
rect 12250 11840 12256 11852
rect 12308 11840 12314 11892
rect 13354 11840 13360 11892
rect 13412 11880 13418 11892
rect 13449 11883 13507 11889
rect 13449 11880 13461 11883
rect 13412 11852 13461 11880
rect 13412 11840 13418 11852
rect 13449 11849 13461 11852
rect 13495 11849 13507 11883
rect 13449 11843 13507 11849
rect 13722 11840 13728 11892
rect 13780 11880 13786 11892
rect 14550 11880 14556 11892
rect 13780 11840 13814 11880
rect 14511 11852 14556 11880
rect 14550 11840 14556 11852
rect 14608 11840 14614 11892
rect 15654 11880 15660 11892
rect 15615 11852 15660 11880
rect 15654 11840 15660 11852
rect 15712 11840 15718 11892
rect 20806 11840 20812 11892
rect 20864 11880 20870 11892
rect 20901 11883 20959 11889
rect 20901 11880 20913 11883
rect 20864 11852 20913 11880
rect 20864 11840 20870 11852
rect 20901 11849 20913 11852
rect 20947 11849 20959 11883
rect 20901 11843 20959 11849
rect 12268 11744 12296 11840
rect 12268 11716 12572 11744
rect 12437 11679 12495 11685
rect 12437 11676 12449 11679
rect 10250 11648 11100 11676
rect 11808 11648 12449 11676
rect 10250 11645 10262 11648
rect 10204 11639 10262 11645
rect 2498 11608 2504 11620
rect 2459 11580 2504 11608
rect 2498 11568 2504 11580
rect 2556 11568 2562 11620
rect 2590 11568 2596 11620
rect 2648 11608 2654 11620
rect 3421 11611 3479 11617
rect 3421 11608 3433 11611
rect 2648 11580 3433 11608
rect 2648 11568 2654 11580
rect 3421 11577 3433 11580
rect 3467 11577 3479 11611
rect 3421 11571 3479 11577
rect 4157 11611 4215 11617
rect 4157 11577 4169 11611
rect 4203 11608 4215 11611
rect 4433 11611 4491 11617
rect 4433 11608 4445 11611
rect 4203 11580 4445 11608
rect 4203 11577 4215 11580
rect 4157 11571 4215 11577
rect 4433 11577 4445 11580
rect 4479 11608 4491 11611
rect 4798 11608 4804 11620
rect 4479 11580 4804 11608
rect 4479 11577 4491 11580
rect 4433 11571 4491 11577
rect 4798 11568 4804 11580
rect 4856 11568 4862 11620
rect 7193 11611 7251 11617
rect 7193 11577 7205 11611
rect 7239 11577 7251 11611
rect 7193 11571 7251 11577
rect 8757 11611 8815 11617
rect 8757 11577 8769 11611
rect 8803 11577 8815 11611
rect 8757 11571 8815 11577
rect 1949 11543 2007 11549
rect 1949 11509 1961 11543
rect 1995 11540 2007 11543
rect 2038 11540 2044 11552
rect 1995 11512 2044 11540
rect 1995 11509 2007 11512
rect 1949 11503 2007 11509
rect 2038 11500 2044 11512
rect 2096 11540 2102 11552
rect 2866 11540 2872 11552
rect 2096 11512 2872 11540
rect 2096 11500 2102 11512
rect 2866 11500 2872 11512
rect 2924 11500 2930 11552
rect 5350 11540 5356 11552
rect 5311 11512 5356 11540
rect 5350 11500 5356 11512
rect 5408 11500 5414 11552
rect 6822 11500 6828 11552
rect 6880 11540 6886 11552
rect 7208 11540 7236 11571
rect 8018 11540 8024 11552
rect 6880 11512 7236 11540
rect 7979 11512 8024 11540
rect 6880 11500 6886 11512
rect 8018 11500 8024 11512
rect 8076 11540 8082 11552
rect 8389 11543 8447 11549
rect 8389 11540 8401 11543
rect 8076 11512 8401 11540
rect 8076 11500 8082 11512
rect 8389 11509 8401 11512
rect 8435 11540 8447 11543
rect 8772 11540 8800 11571
rect 9582 11568 9588 11620
rect 9640 11608 9646 11620
rect 11808 11617 11836 11648
rect 12437 11645 12449 11648
rect 12483 11645 12495 11679
rect 12544 11676 12572 11716
rect 12802 11704 12808 11756
rect 12860 11744 12866 11756
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 12860 11716 13001 11744
rect 12860 11704 12866 11716
rect 12989 11713 13001 11716
rect 13035 11713 13047 11747
rect 13786 11744 13814 11840
rect 13909 11747 13967 11753
rect 13909 11744 13921 11747
rect 13786 11716 13921 11744
rect 12989 11707 13047 11713
rect 13909 11713 13921 11716
rect 13955 11744 13967 11747
rect 15013 11747 15071 11753
rect 15013 11744 15025 11747
rect 13955 11716 15025 11744
rect 13955 11713 13967 11716
rect 13909 11707 13967 11713
rect 15013 11713 15025 11716
rect 15059 11713 15071 11747
rect 15672 11744 15700 11840
rect 15672 11716 16712 11744
rect 15013 11707 15071 11713
rect 12897 11679 12955 11685
rect 12897 11676 12909 11679
rect 12544 11648 12909 11676
rect 12437 11639 12495 11645
rect 12897 11645 12909 11648
rect 12943 11645 12955 11679
rect 12897 11639 12955 11645
rect 16117 11679 16175 11685
rect 16117 11645 16129 11679
rect 16163 11676 16175 11679
rect 16206 11676 16212 11688
rect 16163 11648 16212 11676
rect 16163 11645 16175 11648
rect 16117 11639 16175 11645
rect 11793 11611 11851 11617
rect 11793 11608 11805 11611
rect 9640 11580 11805 11608
rect 9640 11568 9646 11580
rect 11793 11577 11805 11580
rect 11839 11577 11851 11611
rect 11793 11571 11851 11577
rect 8435 11512 8800 11540
rect 8435 11509 8447 11512
rect 8389 11503 8447 11509
rect 9398 11500 9404 11552
rect 9456 11540 9462 11552
rect 10275 11543 10333 11549
rect 10275 11540 10287 11543
rect 9456 11512 10287 11540
rect 9456 11500 9462 11512
rect 10275 11509 10287 11512
rect 10321 11509 10333 11543
rect 10275 11503 10333 11509
rect 10410 11500 10416 11552
rect 10468 11540 10474 11552
rect 10689 11543 10747 11549
rect 10689 11540 10701 11543
rect 10468 11512 10701 11540
rect 10468 11500 10474 11512
rect 10689 11509 10701 11512
rect 10735 11540 10747 11543
rect 11698 11540 11704 11552
rect 10735 11512 11704 11540
rect 10735 11509 10747 11512
rect 10689 11503 10747 11509
rect 11698 11500 11704 11512
rect 11756 11500 11762 11552
rect 12452 11540 12480 11639
rect 16206 11636 16212 11648
rect 16264 11636 16270 11688
rect 16684 11685 16712 11716
rect 16669 11679 16727 11685
rect 16669 11645 16681 11679
rect 16715 11645 16727 11679
rect 16669 11639 16727 11645
rect 14734 11608 14740 11620
rect 14695 11580 14740 11608
rect 14734 11568 14740 11580
rect 14792 11568 14798 11620
rect 14829 11611 14887 11617
rect 14829 11577 14841 11611
rect 14875 11608 14887 11611
rect 15470 11608 15476 11620
rect 14875 11580 15476 11608
rect 14875 11577 14887 11580
rect 14829 11571 14887 11577
rect 15470 11568 15476 11580
rect 15528 11568 15534 11620
rect 14274 11540 14280 11552
rect 12452 11512 14280 11540
rect 14274 11500 14280 11512
rect 14332 11540 14338 11552
rect 15378 11540 15384 11552
rect 14332 11512 15384 11540
rect 14332 11500 14338 11512
rect 15378 11500 15384 11512
rect 15436 11500 15442 11552
rect 16482 11540 16488 11552
rect 16443 11512 16488 11540
rect 16482 11500 16488 11512
rect 16540 11500 16546 11552
rect 1104 11450 22816 11472
rect 1104 11398 8982 11450
rect 9034 11398 9046 11450
rect 9098 11398 9110 11450
rect 9162 11398 9174 11450
rect 9226 11398 16982 11450
rect 17034 11398 17046 11450
rect 17098 11398 17110 11450
rect 17162 11398 17174 11450
rect 17226 11398 22816 11450
rect 1104 11376 22816 11398
rect 2130 11336 2136 11348
rect 2091 11308 2136 11336
rect 2130 11296 2136 11308
rect 2188 11296 2194 11348
rect 2498 11296 2504 11348
rect 2556 11336 2562 11348
rect 2961 11339 3019 11345
rect 2961 11336 2973 11339
rect 2556 11308 2973 11336
rect 2556 11296 2562 11308
rect 2961 11305 2973 11308
rect 3007 11305 3019 11339
rect 4430 11336 4436 11348
rect 4391 11308 4436 11336
rect 2961 11299 3019 11305
rect 4430 11296 4436 11308
rect 4488 11296 4494 11348
rect 4798 11296 4804 11348
rect 4856 11336 4862 11348
rect 4985 11339 5043 11345
rect 4985 11336 4997 11339
rect 4856 11308 4997 11336
rect 4856 11296 4862 11308
rect 4985 11305 4997 11308
rect 5031 11305 5043 11339
rect 4985 11299 5043 11305
rect 5626 11296 5632 11348
rect 5684 11336 5690 11348
rect 5813 11339 5871 11345
rect 5813 11336 5825 11339
rect 5684 11308 5825 11336
rect 5684 11296 5690 11308
rect 5813 11305 5825 11308
rect 5859 11305 5871 11339
rect 5813 11299 5871 11305
rect 12437 11339 12495 11345
rect 12437 11305 12449 11339
rect 12483 11336 12495 11339
rect 13354 11336 13360 11348
rect 12483 11308 13360 11336
rect 12483 11305 12495 11308
rect 12437 11299 12495 11305
rect 13354 11296 13360 11308
rect 13412 11336 13418 11348
rect 13412 11308 13492 11336
rect 13412 11296 13418 11308
rect 6638 11228 6644 11280
rect 6696 11268 6702 11280
rect 7101 11271 7159 11277
rect 7101 11268 7113 11271
rect 6696 11240 7113 11268
rect 6696 11228 6702 11240
rect 7101 11237 7113 11240
rect 7147 11237 7159 11271
rect 7101 11231 7159 11237
rect 10689 11271 10747 11277
rect 10689 11237 10701 11271
rect 10735 11268 10747 11271
rect 10778 11268 10784 11280
rect 10735 11240 10784 11268
rect 10735 11237 10747 11240
rect 10689 11231 10747 11237
rect 10778 11228 10784 11240
rect 10836 11228 10842 11280
rect 11698 11228 11704 11280
rect 11756 11268 11762 11280
rect 11879 11271 11937 11277
rect 11879 11268 11891 11271
rect 11756 11240 11891 11268
rect 11756 11228 11762 11240
rect 11879 11237 11891 11240
rect 11925 11268 11937 11271
rect 12710 11268 12716 11280
rect 11925 11240 12716 11268
rect 11925 11237 11937 11240
rect 11879 11231 11937 11237
rect 12710 11228 12716 11240
rect 12768 11228 12774 11280
rect 13464 11277 13492 11308
rect 13449 11271 13507 11277
rect 13449 11237 13461 11271
rect 13495 11237 13507 11271
rect 13998 11268 14004 11280
rect 13959 11240 14004 11268
rect 13449 11231 13507 11237
rect 13998 11228 14004 11240
rect 14056 11228 14062 11280
rect 14737 11271 14795 11277
rect 14737 11237 14749 11271
rect 14783 11268 14795 11271
rect 14826 11268 14832 11280
rect 14783 11240 14832 11268
rect 14783 11237 14795 11240
rect 14737 11231 14795 11237
rect 14826 11228 14832 11240
rect 14884 11268 14890 11280
rect 15105 11271 15163 11277
rect 15105 11268 15117 11271
rect 14884 11240 15117 11268
rect 14884 11228 14890 11240
rect 15105 11237 15117 11240
rect 15151 11268 15163 11271
rect 15470 11268 15476 11280
rect 15151 11240 15476 11268
rect 15151 11237 15163 11240
rect 15105 11231 15163 11237
rect 15470 11228 15476 11240
rect 15528 11228 15534 11280
rect 18690 11268 18696 11280
rect 18651 11240 18696 11268
rect 18690 11228 18696 11240
rect 18748 11228 18754 11280
rect 2590 11160 2596 11212
rect 2648 11200 2654 11212
rect 2685 11203 2743 11209
rect 2685 11200 2697 11203
rect 2648 11172 2697 11200
rect 2648 11160 2654 11172
rect 2685 11169 2697 11172
rect 2731 11169 2743 11203
rect 9950 11200 9956 11212
rect 9911 11172 9956 11200
rect 2685 11163 2743 11169
rect 9950 11160 9956 11172
rect 10008 11160 10014 11212
rect 10229 11203 10287 11209
rect 10229 11169 10241 11203
rect 10275 11169 10287 11203
rect 10229 11163 10287 11169
rect 1765 11135 1823 11141
rect 1765 11101 1777 11135
rect 1811 11132 1823 11135
rect 3326 11132 3332 11144
rect 1811 11104 3332 11132
rect 1811 11101 1823 11104
rect 1765 11095 1823 11101
rect 3326 11092 3332 11104
rect 3384 11092 3390 11144
rect 4062 11132 4068 11144
rect 4023 11104 4068 11132
rect 4062 11092 4068 11104
rect 4120 11092 4126 11144
rect 7009 11135 7067 11141
rect 7009 11101 7021 11135
rect 7055 11101 7067 11135
rect 7374 11132 7380 11144
rect 7335 11104 7380 11132
rect 7009 11095 7067 11101
rect 6270 11024 6276 11076
rect 6328 11064 6334 11076
rect 7024 11064 7052 11095
rect 7374 11092 7380 11104
rect 7432 11092 7438 11144
rect 7926 11092 7932 11144
rect 7984 11132 7990 11144
rect 8021 11135 8079 11141
rect 8021 11132 8033 11135
rect 7984 11104 8033 11132
rect 7984 11092 7990 11104
rect 8021 11101 8033 11104
rect 8067 11132 8079 11135
rect 8481 11135 8539 11141
rect 8481 11132 8493 11135
rect 8067 11104 8493 11132
rect 8067 11101 8079 11104
rect 8021 11095 8079 11101
rect 8481 11101 8493 11104
rect 8527 11101 8539 11135
rect 10244 11132 10272 11163
rect 20806 11160 20812 11212
rect 20864 11200 20870 11212
rect 20968 11203 21026 11209
rect 20968 11200 20980 11203
rect 20864 11172 20980 11200
rect 20864 11160 20870 11172
rect 20968 11169 20980 11172
rect 21014 11200 21026 11203
rect 22094 11200 22100 11212
rect 21014 11172 22100 11200
rect 21014 11169 21026 11172
rect 20968 11163 21026 11169
rect 22094 11160 22100 11172
rect 22152 11160 22158 11212
rect 10686 11132 10692 11144
rect 10244 11104 10692 11132
rect 8481 11095 8539 11101
rect 10686 11092 10692 11104
rect 10744 11092 10750 11144
rect 11517 11135 11575 11141
rect 11517 11101 11529 11135
rect 11563 11132 11575 11135
rect 11606 11132 11612 11144
rect 11563 11104 11612 11132
rect 11563 11101 11575 11104
rect 11517 11095 11575 11101
rect 11606 11092 11612 11104
rect 11664 11092 11670 11144
rect 13357 11135 13415 11141
rect 13357 11101 13369 11135
rect 13403 11101 13415 11135
rect 15378 11132 15384 11144
rect 13357 11095 13415 11101
rect 13786 11104 14044 11132
rect 15339 11104 15384 11132
rect 9766 11064 9772 11076
rect 6328 11036 9772 11064
rect 6328 11024 6334 11036
rect 9766 11024 9772 11036
rect 9824 11024 9830 11076
rect 10045 11067 10103 11073
rect 10045 11033 10057 11067
rect 10091 11064 10103 11067
rect 10410 11064 10416 11076
rect 10091 11036 10416 11064
rect 10091 11033 10103 11036
rect 10045 11027 10103 11033
rect 10410 11024 10416 11036
rect 10468 11024 10474 11076
rect 13372 11064 13400 11095
rect 13538 11064 13544 11076
rect 13372 11036 13544 11064
rect 13538 11024 13544 11036
rect 13596 11064 13602 11076
rect 13786 11064 13814 11104
rect 13596 11036 13814 11064
rect 14016 11064 14044 11104
rect 15378 11092 15384 11104
rect 15436 11092 15442 11144
rect 15657 11135 15715 11141
rect 15657 11101 15669 11135
rect 15703 11101 15715 11135
rect 15657 11095 15715 11101
rect 18601 11135 18659 11141
rect 18601 11101 18613 11135
rect 18647 11132 18659 11135
rect 18782 11132 18788 11144
rect 18647 11104 18788 11132
rect 18647 11101 18659 11104
rect 18601 11095 18659 11101
rect 15672 11064 15700 11095
rect 18782 11092 18788 11104
rect 18840 11092 18846 11144
rect 19150 11064 19156 11076
rect 14016 11036 15700 11064
rect 19111 11036 19156 11064
rect 13596 11024 13602 11036
rect 19150 11024 19156 11036
rect 19208 11024 19214 11076
rect 11790 10956 11796 11008
rect 11848 10996 11854 11008
rect 15194 10996 15200 11008
rect 11848 10968 15200 10996
rect 11848 10956 11854 10968
rect 15194 10956 15200 10968
rect 15252 10956 15258 11008
rect 16390 10956 16396 11008
rect 16448 10996 16454 11008
rect 16485 10999 16543 11005
rect 16485 10996 16497 10999
rect 16448 10968 16497 10996
rect 16448 10956 16454 10968
rect 16485 10965 16497 10968
rect 16531 10996 16543 10999
rect 17310 10996 17316 11008
rect 16531 10968 17316 10996
rect 16531 10965 16543 10968
rect 16485 10959 16543 10965
rect 17310 10956 17316 10968
rect 17368 10956 17374 11008
rect 19242 10956 19248 11008
rect 19300 10996 19306 11008
rect 21039 10999 21097 11005
rect 21039 10996 21051 10999
rect 19300 10968 21051 10996
rect 19300 10956 19306 10968
rect 21039 10965 21051 10968
rect 21085 10965 21097 10999
rect 21039 10959 21097 10965
rect 1104 10906 22816 10928
rect 1104 10854 4982 10906
rect 5034 10854 5046 10906
rect 5098 10854 5110 10906
rect 5162 10854 5174 10906
rect 5226 10854 12982 10906
rect 13034 10854 13046 10906
rect 13098 10854 13110 10906
rect 13162 10854 13174 10906
rect 13226 10854 20982 10906
rect 21034 10854 21046 10906
rect 21098 10854 21110 10906
rect 21162 10854 21174 10906
rect 21226 10854 22816 10906
rect 1104 10832 22816 10854
rect 1578 10792 1584 10804
rect 1539 10764 1584 10792
rect 1578 10752 1584 10764
rect 1636 10752 1642 10804
rect 2130 10752 2136 10804
rect 2188 10792 2194 10804
rect 2317 10795 2375 10801
rect 2317 10792 2329 10795
rect 2188 10764 2329 10792
rect 2188 10752 2194 10764
rect 2317 10761 2329 10764
rect 2363 10761 2375 10795
rect 2317 10755 2375 10761
rect 2332 10724 2360 10755
rect 2498 10752 2504 10804
rect 2556 10792 2562 10804
rect 2639 10795 2697 10801
rect 2639 10792 2651 10795
rect 2556 10764 2651 10792
rect 2556 10752 2562 10764
rect 2639 10761 2651 10764
rect 2685 10761 2697 10795
rect 2639 10755 2697 10761
rect 4062 10752 4068 10804
rect 4120 10792 4126 10804
rect 5442 10792 5448 10804
rect 4120 10764 5448 10792
rect 4120 10752 4126 10764
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 6270 10792 6276 10804
rect 6231 10764 6276 10792
rect 6270 10752 6276 10764
rect 6328 10752 6334 10804
rect 7742 10792 7748 10804
rect 7703 10764 7748 10792
rect 7742 10752 7748 10764
rect 7800 10752 7806 10804
rect 9950 10752 9956 10804
rect 10008 10792 10014 10804
rect 11149 10795 11207 10801
rect 11149 10792 11161 10795
rect 10008 10764 11161 10792
rect 10008 10752 10014 10764
rect 11149 10761 11161 10764
rect 11195 10792 11207 10795
rect 11238 10792 11244 10804
rect 11195 10764 11244 10792
rect 11195 10761 11207 10764
rect 11149 10755 11207 10761
rect 11238 10752 11244 10764
rect 11296 10752 11302 10804
rect 11609 10795 11667 10801
rect 11609 10761 11621 10795
rect 11655 10792 11667 10795
rect 11698 10792 11704 10804
rect 11655 10764 11704 10792
rect 11655 10761 11667 10764
rect 11609 10755 11667 10761
rect 11698 10752 11704 10764
rect 11756 10752 11762 10804
rect 13354 10792 13360 10804
rect 13315 10764 13360 10792
rect 13354 10752 13360 10764
rect 13412 10752 13418 10804
rect 14826 10792 14832 10804
rect 14787 10764 14832 10792
rect 14826 10752 14832 10764
rect 14884 10792 14890 10804
rect 15289 10795 15347 10801
rect 15289 10792 15301 10795
rect 14884 10764 15301 10792
rect 14884 10752 14890 10764
rect 15289 10761 15301 10764
rect 15335 10761 15347 10795
rect 16206 10792 16212 10804
rect 16167 10764 16212 10792
rect 15289 10755 15347 10761
rect 16206 10752 16212 10764
rect 16264 10752 16270 10804
rect 20806 10752 20812 10804
rect 20864 10792 20870 10804
rect 20901 10795 20959 10801
rect 20901 10792 20913 10795
rect 20864 10764 20913 10792
rect 20864 10752 20870 10764
rect 20901 10761 20913 10764
rect 20947 10761 20959 10795
rect 20901 10755 20959 10761
rect 4157 10727 4215 10733
rect 4157 10724 4169 10727
rect 2332 10696 4169 10724
rect 4157 10693 4169 10696
rect 4203 10693 4215 10727
rect 4157 10687 4215 10693
rect 6963 10727 7021 10733
rect 6963 10693 6975 10727
rect 7009 10724 7021 10727
rect 12989 10727 13047 10733
rect 7009 10696 9536 10724
rect 7009 10693 7021 10696
rect 6963 10687 7021 10693
rect 9508 10668 9536 10696
rect 12989 10693 13001 10727
rect 13035 10724 13047 10727
rect 13538 10724 13544 10736
rect 13035 10696 13544 10724
rect 13035 10693 13047 10696
rect 12989 10687 13047 10693
rect 13538 10684 13544 10696
rect 13596 10684 13602 10736
rect 13814 10684 13820 10736
rect 13872 10724 13878 10736
rect 17954 10724 17960 10736
rect 13872 10696 17960 10724
rect 13872 10684 13878 10696
rect 17954 10684 17960 10696
rect 18012 10684 18018 10736
rect 18598 10684 18604 10736
rect 18656 10724 18662 10736
rect 18874 10724 18880 10736
rect 18656 10696 18880 10724
rect 18656 10684 18662 10696
rect 18874 10684 18880 10696
rect 18932 10684 18938 10736
rect 5077 10659 5135 10665
rect 5077 10625 5089 10659
rect 5123 10656 5135 10659
rect 5350 10656 5356 10668
rect 5123 10628 5356 10656
rect 5123 10625 5135 10628
rect 5077 10619 5135 10625
rect 5350 10616 5356 10628
rect 5408 10616 5414 10668
rect 7926 10656 7932 10668
rect 7887 10628 7932 10656
rect 7926 10616 7932 10628
rect 7984 10616 7990 10668
rect 8386 10656 8392 10668
rect 8347 10628 8392 10656
rect 8386 10616 8392 10628
rect 8444 10616 8450 10668
rect 9490 10656 9496 10668
rect 9403 10628 9496 10656
rect 9490 10616 9496 10628
rect 9548 10616 9554 10668
rect 9766 10656 9772 10668
rect 9727 10628 9772 10656
rect 9766 10616 9772 10628
rect 9824 10616 9830 10668
rect 13998 10656 14004 10668
rect 12519 10628 14004 10656
rect 12519 10600 12547 10628
rect 13998 10616 14004 10628
rect 14056 10616 14062 10668
rect 17865 10659 17923 10665
rect 17865 10625 17877 10659
rect 17911 10656 17923 10659
rect 18690 10656 18696 10668
rect 17911 10628 18696 10656
rect 17911 10625 17923 10628
rect 17865 10619 17923 10625
rect 18690 10616 18696 10628
rect 18748 10616 18754 10668
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10588 1455 10591
rect 1443 10560 2084 10588
rect 1443 10557 1455 10560
rect 1397 10551 1455 10557
rect 2056 10464 2084 10560
rect 2222 10548 2228 10600
rect 2280 10588 2286 10600
rect 2536 10591 2594 10597
rect 2536 10588 2548 10591
rect 2280 10560 2548 10588
rect 2280 10548 2286 10560
rect 2536 10557 2548 10560
rect 2582 10588 2594 10591
rect 2961 10591 3019 10597
rect 2961 10588 2973 10591
rect 2582 10560 2973 10588
rect 2582 10557 2594 10560
rect 2536 10551 2594 10557
rect 2961 10557 2973 10560
rect 3007 10588 3019 10591
rect 3602 10588 3608 10600
rect 3007 10560 3608 10588
rect 3007 10557 3019 10560
rect 2961 10551 3019 10557
rect 3602 10548 3608 10560
rect 3660 10548 3666 10600
rect 3789 10591 3847 10597
rect 3789 10557 3801 10591
rect 3835 10588 3847 10591
rect 4798 10588 4804 10600
rect 3835 10560 4804 10588
rect 3835 10557 3847 10560
rect 3789 10551 3847 10557
rect 4798 10548 4804 10560
rect 4856 10548 4862 10600
rect 12519 10597 12532 10600
rect 6892 10591 6950 10597
rect 6892 10557 6904 10591
rect 6938 10588 6950 10591
rect 12504 10591 12532 10597
rect 12504 10588 12516 10591
rect 6938 10557 6960 10588
rect 12439 10560 12516 10588
rect 6892 10551 6960 10557
rect 12504 10557 12516 10560
rect 12504 10551 12532 10557
rect 4706 10480 4712 10532
rect 4764 10520 4770 10532
rect 6932 10520 6960 10551
rect 12526 10548 12532 10551
rect 12584 10548 12590 10600
rect 13906 10588 13912 10600
rect 13867 10560 13912 10588
rect 13906 10548 13912 10560
rect 13964 10548 13970 10600
rect 16206 10548 16212 10600
rect 16264 10588 16270 10600
rect 16393 10591 16451 10597
rect 16393 10588 16405 10591
rect 16264 10560 16405 10588
rect 16264 10548 16270 10560
rect 16393 10557 16405 10560
rect 16439 10588 16451 10591
rect 16758 10588 16764 10600
rect 16439 10560 16764 10588
rect 16439 10557 16451 10560
rect 16393 10551 16451 10557
rect 16758 10548 16764 10560
rect 16816 10548 16822 10600
rect 16945 10591 17003 10597
rect 16945 10557 16957 10591
rect 16991 10588 17003 10591
rect 17310 10588 17316 10600
rect 16991 10560 17316 10588
rect 16991 10557 17003 10560
rect 16945 10551 17003 10557
rect 17310 10548 17316 10560
rect 17368 10548 17374 10600
rect 7285 10523 7343 10529
rect 7285 10520 7297 10523
rect 4764 10492 7297 10520
rect 4764 10480 4770 10492
rect 7285 10489 7297 10492
rect 7331 10520 7343 10523
rect 7558 10520 7564 10532
rect 7331 10492 7564 10520
rect 7331 10489 7343 10492
rect 7285 10483 7343 10489
rect 7558 10480 7564 10492
rect 7616 10480 7622 10532
rect 7742 10480 7748 10532
rect 7800 10520 7806 10532
rect 8021 10523 8079 10529
rect 8021 10520 8033 10523
rect 7800 10492 8033 10520
rect 7800 10480 7806 10492
rect 8021 10489 8033 10492
rect 8067 10489 8079 10523
rect 8021 10483 8079 10489
rect 9585 10523 9643 10529
rect 9585 10489 9597 10523
rect 9631 10489 9643 10523
rect 9585 10483 9643 10489
rect 13817 10523 13875 10529
rect 13817 10489 13829 10523
rect 13863 10520 13875 10523
rect 13998 10520 14004 10532
rect 13863 10492 14004 10520
rect 13863 10489 13875 10492
rect 13817 10483 13875 10489
rect 2038 10452 2044 10464
rect 1999 10424 2044 10452
rect 2038 10412 2044 10424
rect 2096 10412 2102 10464
rect 3326 10452 3332 10464
rect 3287 10424 3332 10452
rect 3326 10412 3332 10424
rect 3384 10412 3390 10464
rect 5442 10452 5448 10464
rect 5403 10424 5448 10452
rect 5442 10412 5448 10424
rect 5500 10412 5506 10464
rect 6638 10452 6644 10464
rect 6599 10424 6644 10452
rect 6638 10412 6644 10424
rect 6696 10412 6702 10464
rect 8036 10452 8064 10483
rect 9217 10455 9275 10461
rect 9217 10452 9229 10455
rect 8036 10424 9229 10452
rect 9217 10421 9229 10424
rect 9263 10452 9275 10455
rect 9600 10452 9628 10483
rect 13998 10480 14004 10492
rect 14056 10520 14062 10532
rect 14271 10523 14329 10529
rect 14271 10520 14283 10523
rect 14056 10492 14283 10520
rect 14056 10480 14062 10492
rect 14271 10489 14283 10492
rect 14317 10520 14329 10523
rect 16850 10520 16856 10532
rect 14317 10492 16856 10520
rect 14317 10489 14329 10492
rect 14271 10483 14329 10489
rect 16850 10480 16856 10492
rect 16908 10480 16914 10532
rect 17129 10523 17187 10529
rect 17129 10489 17141 10523
rect 17175 10520 17187 10523
rect 17770 10520 17776 10532
rect 17175 10492 17776 10520
rect 17175 10489 17187 10492
rect 17129 10483 17187 10489
rect 17770 10480 17776 10492
rect 17828 10480 17834 10532
rect 18598 10520 18604 10532
rect 18559 10492 18604 10520
rect 18598 10480 18604 10492
rect 18656 10480 18662 10532
rect 18693 10523 18751 10529
rect 18693 10489 18705 10523
rect 18739 10489 18751 10523
rect 18693 10483 18751 10489
rect 10410 10452 10416 10464
rect 9263 10424 9628 10452
rect 10371 10424 10416 10452
rect 9263 10421 9275 10424
rect 9217 10415 9275 10421
rect 10410 10412 10416 10424
rect 10468 10412 10474 10464
rect 10686 10412 10692 10464
rect 10744 10452 10750 10464
rect 10781 10455 10839 10461
rect 10781 10452 10793 10455
rect 10744 10424 10793 10452
rect 10744 10412 10750 10424
rect 10781 10421 10793 10424
rect 10827 10421 10839 10455
rect 10781 10415 10839 10421
rect 11606 10412 11612 10464
rect 11664 10452 11670 10464
rect 11885 10455 11943 10461
rect 11885 10452 11897 10455
rect 11664 10424 11897 10452
rect 11664 10412 11670 10424
rect 11885 10421 11897 10424
rect 11931 10421 11943 10455
rect 11885 10415 11943 10421
rect 12250 10412 12256 10464
rect 12308 10452 12314 10464
rect 12575 10455 12633 10461
rect 12575 10452 12587 10455
rect 12308 10424 12587 10452
rect 12308 10412 12314 10424
rect 12575 10421 12587 10424
rect 12621 10421 12633 10455
rect 12575 10415 12633 10421
rect 15378 10412 15384 10464
rect 15436 10452 15442 10464
rect 15746 10452 15752 10464
rect 15436 10424 15752 10452
rect 15436 10412 15442 10424
rect 15746 10412 15752 10424
rect 15804 10412 15810 10464
rect 17402 10412 17408 10464
rect 17460 10452 17466 10464
rect 18325 10455 18383 10461
rect 18325 10452 18337 10455
rect 17460 10424 18337 10452
rect 17460 10412 17466 10424
rect 18325 10421 18337 10424
rect 18371 10452 18383 10455
rect 18708 10452 18736 10483
rect 18782 10480 18788 10532
rect 18840 10520 18846 10532
rect 19245 10523 19303 10529
rect 19245 10520 19257 10523
rect 18840 10492 19257 10520
rect 18840 10480 18846 10492
rect 19245 10489 19257 10492
rect 19291 10520 19303 10523
rect 19291 10492 19932 10520
rect 19291 10489 19303 10492
rect 19245 10483 19303 10489
rect 19904 10464 19932 10492
rect 18371 10424 18736 10452
rect 18371 10421 18383 10424
rect 18325 10415 18383 10421
rect 18874 10412 18880 10464
rect 18932 10452 18938 10464
rect 19521 10455 19579 10461
rect 19521 10452 19533 10455
rect 18932 10424 19533 10452
rect 18932 10412 18938 10424
rect 19521 10421 19533 10424
rect 19567 10421 19579 10455
rect 19886 10452 19892 10464
rect 19847 10424 19892 10452
rect 19521 10415 19579 10421
rect 19886 10412 19892 10424
rect 19944 10412 19950 10464
rect 1104 10362 22816 10384
rect 1104 10310 8982 10362
rect 9034 10310 9046 10362
rect 9098 10310 9110 10362
rect 9162 10310 9174 10362
rect 9226 10310 16982 10362
rect 17034 10310 17046 10362
rect 17098 10310 17110 10362
rect 17162 10310 17174 10362
rect 17226 10310 22816 10362
rect 1104 10288 22816 10310
rect 1670 10208 1676 10260
rect 1728 10248 1734 10260
rect 2639 10251 2697 10257
rect 2639 10248 2651 10251
rect 1728 10220 2651 10248
rect 1728 10208 1734 10220
rect 2639 10217 2651 10220
rect 2685 10217 2697 10251
rect 2639 10211 2697 10217
rect 3789 10251 3847 10257
rect 3789 10217 3801 10251
rect 3835 10248 3847 10251
rect 3878 10248 3884 10260
rect 3835 10220 3884 10248
rect 3835 10217 3847 10220
rect 3789 10211 3847 10217
rect 3804 10180 3832 10211
rect 3878 10208 3884 10220
rect 3936 10208 3942 10260
rect 4246 10248 4252 10260
rect 4159 10220 4252 10248
rect 4246 10208 4252 10220
rect 4304 10208 4310 10260
rect 4430 10208 4436 10260
rect 4488 10248 4494 10260
rect 4488 10220 5488 10248
rect 4488 10208 4494 10220
rect 2583 10152 3832 10180
rect 2583 10121 2611 10152
rect 3970 10140 3976 10192
rect 4028 10180 4034 10192
rect 5460 10180 5488 10220
rect 6638 10208 6644 10260
rect 6696 10248 6702 10260
rect 7929 10251 7987 10257
rect 7929 10248 7941 10251
rect 6696 10220 7941 10248
rect 6696 10208 6702 10220
rect 7929 10217 7941 10220
rect 7975 10217 7987 10251
rect 9490 10248 9496 10260
rect 9451 10220 9496 10248
rect 7929 10211 7987 10217
rect 9490 10208 9496 10220
rect 9548 10208 9554 10260
rect 12526 10248 12532 10260
rect 12487 10220 12532 10248
rect 12526 10208 12532 10220
rect 12584 10208 12590 10260
rect 15654 10248 15660 10260
rect 13188 10220 15660 10248
rect 7098 10180 7104 10192
rect 4028 10152 4936 10180
rect 5460 10152 7104 10180
rect 4028 10140 4034 10152
rect 1397 10115 1455 10121
rect 1397 10081 1409 10115
rect 1443 10112 1455 10115
rect 2568 10115 2626 10121
rect 1443 10084 2084 10112
rect 1443 10081 1455 10084
rect 1397 10075 1455 10081
rect 2056 10053 2084 10084
rect 2568 10081 2580 10115
rect 2614 10081 2626 10115
rect 2568 10075 2626 10081
rect 4062 10072 4068 10124
rect 4120 10112 4126 10124
rect 4154 10112 4160 10124
rect 4120 10084 4160 10112
rect 4120 10072 4126 10084
rect 4154 10072 4160 10084
rect 4212 10112 4218 10124
rect 4798 10112 4804 10124
rect 4212 10084 4305 10112
rect 4759 10084 4804 10112
rect 4212 10072 4218 10084
rect 4798 10072 4804 10084
rect 4856 10072 4862 10124
rect 4908 10112 4936 10152
rect 7098 10140 7104 10152
rect 7156 10180 7162 10192
rect 7330 10183 7388 10189
rect 7330 10180 7342 10183
rect 7156 10152 7342 10180
rect 7156 10140 7162 10152
rect 7330 10149 7342 10152
rect 7376 10149 7388 10183
rect 11606 10180 11612 10192
rect 11567 10152 11612 10180
rect 7330 10143 7388 10149
rect 11606 10140 11612 10152
rect 11664 10140 11670 10192
rect 5169 10115 5227 10121
rect 5169 10112 5181 10115
rect 4908 10084 5181 10112
rect 5169 10081 5181 10084
rect 5215 10081 5227 10115
rect 5534 10112 5540 10124
rect 5495 10084 5540 10112
rect 5169 10075 5227 10081
rect 5534 10072 5540 10084
rect 5592 10072 5598 10124
rect 6086 10112 6092 10124
rect 6047 10084 6092 10112
rect 6086 10072 6092 10084
rect 6144 10072 6150 10124
rect 10962 10112 10968 10124
rect 10923 10084 10968 10112
rect 10962 10072 10968 10084
rect 11020 10072 11026 10124
rect 11330 10072 11336 10124
rect 11388 10112 11394 10124
rect 11425 10115 11483 10121
rect 11425 10112 11437 10115
rect 11388 10084 11437 10112
rect 11388 10072 11394 10084
rect 11425 10081 11437 10084
rect 11471 10112 11483 10115
rect 12158 10112 12164 10124
rect 11471 10084 12164 10112
rect 11471 10081 11483 10084
rect 11425 10075 11483 10081
rect 12158 10072 12164 10084
rect 12216 10072 12222 10124
rect 12342 10072 12348 10124
rect 12400 10112 12406 10124
rect 13188 10121 13216 10220
rect 15654 10208 15660 10220
rect 15712 10208 15718 10260
rect 16850 10248 16856 10260
rect 16811 10220 16856 10248
rect 16850 10208 16856 10220
rect 16908 10208 16914 10260
rect 18690 10208 18696 10260
rect 18748 10248 18754 10260
rect 19153 10251 19211 10257
rect 19153 10248 19165 10251
rect 18748 10220 19165 10248
rect 18748 10208 18754 10220
rect 19153 10217 19165 10220
rect 19199 10217 19211 10251
rect 19153 10211 19211 10217
rect 16114 10140 16120 10192
rect 16172 10180 16178 10192
rect 16172 10152 16620 10180
rect 16172 10140 16178 10152
rect 13173 10115 13231 10121
rect 13173 10112 13185 10115
rect 12400 10084 13185 10112
rect 12400 10072 12406 10084
rect 13173 10081 13185 10084
rect 13219 10081 13231 10115
rect 13173 10075 13231 10081
rect 13357 10115 13415 10121
rect 13357 10081 13369 10115
rect 13403 10081 13415 10115
rect 13357 10075 13415 10081
rect 13633 10115 13691 10121
rect 13633 10081 13645 10115
rect 13679 10112 13691 10115
rect 13906 10112 13912 10124
rect 13679 10084 13912 10112
rect 13679 10081 13691 10084
rect 13633 10075 13691 10081
rect 2041 10047 2099 10053
rect 2041 10013 2053 10047
rect 2087 10044 2099 10047
rect 4080 10044 4108 10072
rect 2087 10016 4108 10044
rect 6181 10047 6239 10053
rect 2087 10013 2099 10016
rect 2041 10007 2099 10013
rect 6181 10013 6193 10047
rect 6227 10044 6239 10047
rect 7009 10047 7067 10053
rect 7009 10044 7021 10047
rect 6227 10016 7021 10044
rect 6227 10013 6239 10016
rect 6181 10007 6239 10013
rect 7009 10013 7021 10016
rect 7055 10044 7067 10047
rect 7374 10044 7380 10056
rect 7055 10016 7380 10044
rect 7055 10013 7067 10016
rect 7009 10007 7067 10013
rect 7374 10004 7380 10016
rect 7432 10004 7438 10056
rect 12176 10044 12204 10072
rect 12802 10044 12808 10056
rect 12176 10016 12808 10044
rect 12802 10004 12808 10016
rect 12860 10044 12866 10056
rect 13372 10044 13400 10075
rect 13906 10072 13912 10084
rect 13964 10072 13970 10124
rect 15356 10115 15414 10121
rect 15356 10081 15368 10115
rect 15402 10112 15414 10115
rect 15838 10112 15844 10124
rect 15402 10084 15844 10112
rect 15402 10081 15414 10084
rect 15356 10075 15414 10081
rect 15838 10072 15844 10084
rect 15896 10072 15902 10124
rect 16482 10112 16488 10124
rect 16443 10084 16488 10112
rect 16482 10072 16488 10084
rect 16540 10072 16546 10124
rect 16592 10112 16620 10152
rect 18322 10140 18328 10192
rect 18380 10180 18386 10192
rect 18554 10183 18612 10189
rect 18554 10180 18566 10183
rect 18380 10152 18566 10180
rect 18380 10140 18386 10152
rect 18554 10149 18566 10152
rect 18600 10149 18612 10183
rect 18554 10143 18612 10149
rect 20714 10112 20720 10124
rect 16592 10084 20720 10112
rect 20714 10072 20720 10084
rect 20772 10112 20778 10124
rect 20901 10115 20959 10121
rect 20901 10112 20913 10115
rect 20772 10084 20913 10112
rect 20772 10072 20778 10084
rect 20901 10081 20913 10084
rect 20947 10081 20959 10115
rect 20901 10075 20959 10081
rect 12860 10016 13400 10044
rect 12860 10004 12866 10016
rect 13538 10004 13544 10056
rect 13596 10044 13602 10056
rect 14277 10047 14335 10053
rect 14277 10044 14289 10047
rect 13596 10016 14289 10044
rect 13596 10004 13602 10016
rect 14277 10013 14289 10016
rect 14323 10013 14335 10047
rect 14277 10007 14335 10013
rect 17770 10004 17776 10056
rect 17828 10044 17834 10056
rect 18233 10047 18291 10053
rect 18233 10044 18245 10047
rect 17828 10016 18245 10044
rect 17828 10004 17834 10016
rect 18233 10013 18245 10016
rect 18279 10013 18291 10047
rect 18233 10007 18291 10013
rect 1578 9976 1584 9988
rect 1539 9948 1584 9976
rect 1578 9936 1584 9948
rect 1636 9936 1642 9988
rect 2406 9936 2412 9988
rect 2464 9976 2470 9988
rect 3329 9979 3387 9985
rect 3329 9976 3341 9979
rect 2464 9948 3341 9976
rect 2464 9936 2470 9948
rect 3329 9945 3341 9948
rect 3375 9976 3387 9979
rect 3970 9976 3976 9988
rect 3375 9948 3976 9976
rect 3375 9945 3387 9948
rect 3329 9939 3387 9945
rect 3970 9936 3976 9948
rect 4028 9936 4034 9988
rect 10321 9979 10379 9985
rect 10321 9945 10333 9979
rect 10367 9976 10379 9979
rect 10778 9976 10784 9988
rect 10367 9948 10784 9976
rect 10367 9945 10379 9948
rect 10321 9939 10379 9945
rect 10778 9936 10784 9948
rect 10836 9936 10842 9988
rect 15746 9936 15752 9988
rect 15804 9976 15810 9988
rect 20162 9976 20168 9988
rect 15804 9948 20168 9976
rect 15804 9936 15810 9948
rect 20162 9936 20168 9948
rect 20220 9936 20226 9988
rect 21082 9976 21088 9988
rect 21043 9948 21088 9976
rect 21082 9936 21088 9948
rect 21140 9936 21146 9988
rect 2317 9911 2375 9917
rect 2317 9877 2329 9911
rect 2363 9908 2375 9911
rect 2498 9908 2504 9920
rect 2363 9880 2504 9908
rect 2363 9877 2375 9880
rect 2317 9871 2375 9877
rect 2498 9868 2504 9880
rect 2556 9868 2562 9920
rect 2590 9868 2596 9920
rect 2648 9908 2654 9920
rect 3053 9911 3111 9917
rect 3053 9908 3065 9911
rect 2648 9880 3065 9908
rect 2648 9868 2654 9880
rect 3053 9877 3065 9880
rect 3099 9908 3111 9911
rect 3786 9908 3792 9920
rect 3099 9880 3792 9908
rect 3099 9877 3111 9880
rect 3053 9871 3111 9877
rect 3786 9868 3792 9880
rect 3844 9868 3850 9920
rect 8110 9868 8116 9920
rect 8168 9908 8174 9920
rect 8205 9911 8263 9917
rect 8205 9908 8217 9911
rect 8168 9880 8217 9908
rect 8168 9868 8174 9880
rect 8205 9877 8217 9880
rect 8251 9877 8263 9911
rect 10594 9908 10600 9920
rect 10555 9880 10600 9908
rect 8205 9871 8263 9877
rect 10594 9868 10600 9880
rect 10652 9868 10658 9920
rect 14550 9868 14556 9920
rect 14608 9908 14614 9920
rect 15427 9911 15485 9917
rect 15427 9908 15439 9911
rect 14608 9880 15439 9908
rect 14608 9868 14614 9880
rect 15427 9877 15439 9880
rect 15473 9877 15485 9911
rect 15838 9908 15844 9920
rect 15799 9880 15844 9908
rect 15427 9871 15485 9877
rect 15838 9868 15844 9880
rect 15896 9868 15902 9920
rect 17402 9908 17408 9920
rect 17363 9880 17408 9908
rect 17402 9868 17408 9880
rect 17460 9868 17466 9920
rect 1104 9818 22816 9840
rect 1104 9766 4982 9818
rect 5034 9766 5046 9818
rect 5098 9766 5110 9818
rect 5162 9766 5174 9818
rect 5226 9766 12982 9818
rect 13034 9766 13046 9818
rect 13098 9766 13110 9818
rect 13162 9766 13174 9818
rect 13226 9766 20982 9818
rect 21034 9766 21046 9818
rect 21098 9766 21110 9818
rect 21162 9766 21174 9818
rect 21226 9766 22816 9818
rect 1104 9744 22816 9766
rect 6086 9664 6092 9716
rect 6144 9704 6150 9716
rect 6273 9707 6331 9713
rect 6273 9704 6285 9707
rect 6144 9676 6285 9704
rect 6144 9664 6150 9676
rect 6273 9673 6285 9676
rect 6319 9673 6331 9707
rect 7098 9704 7104 9716
rect 7059 9676 7104 9704
rect 6273 9667 6331 9673
rect 7098 9664 7104 9676
rect 7156 9664 7162 9716
rect 7374 9704 7380 9716
rect 7335 9676 7380 9704
rect 7374 9664 7380 9676
rect 7432 9664 7438 9716
rect 10394 9707 10452 9713
rect 10394 9673 10406 9707
rect 10440 9704 10452 9707
rect 10594 9704 10600 9716
rect 10440 9676 10600 9704
rect 10440 9673 10452 9676
rect 10394 9667 10452 9673
rect 10594 9664 10600 9676
rect 10652 9664 10658 9716
rect 10873 9707 10931 9713
rect 10873 9673 10885 9707
rect 10919 9704 10931 9707
rect 11330 9704 11336 9716
rect 10919 9676 11336 9704
rect 10919 9673 10931 9676
rect 10873 9667 10931 9673
rect 11330 9664 11336 9676
rect 11388 9664 11394 9716
rect 13541 9707 13599 9713
rect 13541 9673 13553 9707
rect 13587 9704 13599 9707
rect 13998 9704 14004 9716
rect 13587 9676 14004 9704
rect 13587 9673 13599 9676
rect 13541 9667 13599 9673
rect 13998 9664 14004 9676
rect 14056 9664 14062 9716
rect 16482 9664 16488 9716
rect 16540 9704 16546 9716
rect 17037 9707 17095 9713
rect 17037 9704 17049 9707
rect 16540 9676 17049 9704
rect 16540 9664 16546 9676
rect 17037 9673 17049 9676
rect 17083 9673 17095 9707
rect 17770 9704 17776 9716
rect 17731 9676 17776 9704
rect 17037 9667 17095 9673
rect 17770 9664 17776 9676
rect 17828 9664 17834 9716
rect 5442 9596 5448 9648
rect 5500 9636 5506 9648
rect 5537 9639 5595 9645
rect 5537 9636 5549 9639
rect 5500 9608 5549 9636
rect 5500 9596 5506 9608
rect 5537 9605 5549 9608
rect 5583 9605 5595 9639
rect 5537 9599 5595 9605
rect 10505 9639 10563 9645
rect 10505 9605 10517 9639
rect 10551 9605 10563 9639
rect 10505 9599 10563 9605
rect 11624 9608 13814 9636
rect 2590 9568 2596 9580
rect 2148 9540 2596 9568
rect 1946 9460 1952 9512
rect 2004 9500 2010 9512
rect 2148 9509 2176 9540
rect 2590 9528 2596 9540
rect 2648 9528 2654 9580
rect 3605 9571 3663 9577
rect 3605 9568 3617 9571
rect 2700 9540 3617 9568
rect 2133 9503 2191 9509
rect 2133 9500 2145 9503
rect 2004 9472 2145 9500
rect 2004 9460 2010 9472
rect 2133 9469 2145 9472
rect 2179 9469 2191 9503
rect 2406 9500 2412 9512
rect 2367 9472 2412 9500
rect 2133 9463 2191 9469
rect 2406 9460 2412 9472
rect 2464 9460 2470 9512
rect 2498 9460 2504 9512
rect 2556 9500 2562 9512
rect 2700 9509 2728 9540
rect 3605 9537 3617 9540
rect 3651 9568 3663 9571
rect 8757 9571 8815 9577
rect 3651 9540 5212 9568
rect 3651 9537 3663 9540
rect 3605 9531 3663 9537
rect 2685 9503 2743 9509
rect 2685 9500 2697 9503
rect 2556 9472 2697 9500
rect 2556 9460 2562 9472
rect 2685 9469 2697 9472
rect 2731 9469 2743 9503
rect 3142 9500 3148 9512
rect 3103 9472 3148 9500
rect 2685 9463 2743 9469
rect 3142 9460 3148 9472
rect 3200 9460 3206 9512
rect 3786 9460 3792 9512
rect 3844 9500 3850 9512
rect 5184 9509 5212 9540
rect 8757 9537 8769 9571
rect 8803 9568 8815 9571
rect 9766 9568 9772 9580
rect 8803 9540 9772 9568
rect 8803 9537 8815 9540
rect 8757 9531 8815 9537
rect 9766 9528 9772 9540
rect 9824 9528 9830 9580
rect 10410 9528 10416 9580
rect 10468 9568 10474 9580
rect 10520 9568 10548 9599
rect 10468 9540 10548 9568
rect 10597 9571 10655 9577
rect 10468 9528 10474 9540
rect 10597 9537 10609 9571
rect 10643 9568 10655 9571
rect 10778 9568 10784 9580
rect 10643 9540 10784 9568
rect 10643 9537 10655 9540
rect 10597 9531 10655 9537
rect 10778 9528 10784 9540
rect 10836 9568 10842 9580
rect 11514 9568 11520 9580
rect 10836 9540 11520 9568
rect 10836 9528 10842 9540
rect 11514 9528 11520 9540
rect 11572 9528 11578 9580
rect 4157 9503 4215 9509
rect 4157 9500 4169 9503
rect 3844 9472 4169 9500
rect 3844 9460 3850 9472
rect 4157 9469 4169 9472
rect 4203 9469 4215 9503
rect 4617 9503 4675 9509
rect 4617 9500 4629 9503
rect 4157 9463 4215 9469
rect 4356 9472 4629 9500
rect 4356 9432 4384 9472
rect 4617 9469 4629 9472
rect 4663 9469 4675 9503
rect 4617 9463 4675 9469
rect 5169 9503 5227 9509
rect 5169 9469 5181 9503
rect 5215 9469 5227 9503
rect 5169 9463 5227 9469
rect 4172 9404 4384 9432
rect 1762 9364 1768 9376
rect 1723 9336 1768 9364
rect 1762 9324 1768 9336
rect 1820 9324 1826 9376
rect 2133 9367 2191 9373
rect 2133 9333 2145 9367
rect 2179 9364 2191 9367
rect 2314 9364 2320 9376
rect 2179 9336 2320 9364
rect 2179 9333 2191 9336
rect 2133 9327 2191 9333
rect 2314 9324 2320 9336
rect 2372 9324 2378 9376
rect 4062 9364 4068 9376
rect 4023 9336 4068 9364
rect 4062 9324 4068 9336
rect 4120 9364 4126 9376
rect 4172 9364 4200 9404
rect 4120 9336 4200 9364
rect 5184 9364 5212 9463
rect 5258 9460 5264 9512
rect 5316 9500 5322 9512
rect 5537 9503 5595 9509
rect 5537 9500 5549 9503
rect 5316 9472 5549 9500
rect 5316 9460 5322 9472
rect 5537 9469 5549 9472
rect 5583 9500 5595 9503
rect 6086 9500 6092 9512
rect 5583 9472 6092 9500
rect 5583 9469 5595 9472
rect 5537 9463 5595 9469
rect 6086 9460 6092 9472
rect 6144 9460 6150 9512
rect 8110 9432 8116 9444
rect 8071 9404 8116 9432
rect 8110 9392 8116 9404
rect 8168 9392 8174 9444
rect 8205 9435 8263 9441
rect 8205 9401 8217 9435
rect 8251 9432 8263 9435
rect 8386 9432 8392 9444
rect 8251 9404 8392 9432
rect 8251 9401 8263 9404
rect 8205 9395 8263 9401
rect 5534 9364 5540 9376
rect 5184 9336 5540 9364
rect 4120 9324 4126 9336
rect 5534 9324 5540 9336
rect 5592 9364 5598 9376
rect 5994 9364 6000 9376
rect 5592 9336 6000 9364
rect 5592 9324 5598 9336
rect 5994 9324 6000 9336
rect 6052 9324 6058 9376
rect 7929 9367 7987 9373
rect 7929 9333 7941 9367
rect 7975 9364 7987 9367
rect 8018 9364 8024 9376
rect 7975 9336 8024 9364
rect 7975 9333 7987 9336
rect 7929 9327 7987 9333
rect 8018 9324 8024 9336
rect 8076 9364 8082 9376
rect 8220 9364 8248 9395
rect 8386 9392 8392 9404
rect 8444 9392 8450 9444
rect 10229 9435 10287 9441
rect 10229 9432 10241 9435
rect 9692 9404 10241 9432
rect 9692 9376 9720 9404
rect 10229 9401 10241 9404
rect 10275 9401 10287 9435
rect 10229 9395 10287 9401
rect 9674 9364 9680 9376
rect 8076 9336 8248 9364
rect 9635 9336 9680 9364
rect 8076 9324 8082 9336
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 10137 9367 10195 9373
rect 10137 9333 10149 9367
rect 10183 9364 10195 9367
rect 10410 9364 10416 9376
rect 10183 9336 10416 9364
rect 10183 9333 10195 9336
rect 10137 9327 10195 9333
rect 10410 9324 10416 9336
rect 10468 9324 10474 9376
rect 10962 9324 10968 9376
rect 11020 9364 11026 9376
rect 11624 9373 11652 9608
rect 13786 9568 13814 9608
rect 15838 9596 15844 9648
rect 15896 9636 15902 9648
rect 16301 9639 16359 9645
rect 16301 9636 16313 9639
rect 15896 9608 16313 9636
rect 15896 9596 15902 9608
rect 16301 9605 16313 9608
rect 16347 9636 16359 9639
rect 19058 9636 19064 9648
rect 16347 9608 19064 9636
rect 16347 9605 16359 9608
rect 16301 9599 16359 9605
rect 19058 9596 19064 9608
rect 19116 9596 19122 9648
rect 17310 9568 17316 9580
rect 13786 9540 17316 9568
rect 17310 9528 17316 9540
rect 17368 9528 17374 9580
rect 19153 9571 19211 9577
rect 19153 9537 19165 9571
rect 19199 9568 19211 9571
rect 19242 9568 19248 9580
rect 19199 9540 19248 9568
rect 19199 9537 19211 9540
rect 19153 9531 19211 9537
rect 19242 9528 19248 9540
rect 19300 9528 19306 9580
rect 12688 9503 12746 9509
rect 12688 9469 12700 9503
rect 12734 9500 12746 9503
rect 12734 9472 13216 9500
rect 12734 9469 12746 9472
rect 12688 9463 12746 9469
rect 11609 9367 11667 9373
rect 11609 9364 11621 9367
rect 11020 9336 11621 9364
rect 11020 9324 11026 9336
rect 11609 9333 11621 9336
rect 11655 9333 11667 9367
rect 11609 9327 11667 9333
rect 12253 9367 12311 9373
rect 12253 9333 12265 9367
rect 12299 9364 12311 9367
rect 12342 9364 12348 9376
rect 12299 9336 12348 9364
rect 12299 9333 12311 9336
rect 12253 9327 12311 9333
rect 12342 9324 12348 9336
rect 12400 9324 12406 9376
rect 12759 9367 12817 9373
rect 12759 9333 12771 9367
rect 12805 9364 12817 9367
rect 12986 9364 12992 9376
rect 12805 9336 12992 9364
rect 12805 9333 12817 9336
rect 12759 9327 12817 9333
rect 12986 9324 12992 9336
rect 13044 9324 13050 9376
rect 13188 9373 13216 9472
rect 13538 9460 13544 9512
rect 13596 9500 13602 9512
rect 13633 9503 13691 9509
rect 13633 9500 13645 9503
rect 13596 9472 13645 9500
rect 13596 9460 13602 9472
rect 13633 9469 13645 9472
rect 13679 9469 13691 9503
rect 13633 9463 13691 9469
rect 15197 9503 15255 9509
rect 15197 9469 15209 9503
rect 15243 9500 15255 9503
rect 15562 9500 15568 9512
rect 15243 9472 15568 9500
rect 15243 9469 15255 9472
rect 15197 9463 15255 9469
rect 15562 9460 15568 9472
rect 15620 9460 15626 9512
rect 15580 9432 15608 9460
rect 15749 9435 15807 9441
rect 15749 9432 15761 9435
rect 15580 9404 15761 9432
rect 15749 9401 15761 9404
rect 15795 9401 15807 9435
rect 15749 9395 15807 9401
rect 15841 9435 15899 9441
rect 15841 9401 15853 9435
rect 15887 9401 15899 9435
rect 15841 9395 15899 9401
rect 13173 9367 13231 9373
rect 13173 9333 13185 9367
rect 13219 9364 13231 9367
rect 13262 9364 13268 9376
rect 13219 9336 13268 9364
rect 13219 9333 13231 9336
rect 13173 9327 13231 9333
rect 13262 9324 13268 9336
rect 13320 9324 13326 9376
rect 13998 9364 14004 9376
rect 13959 9336 14004 9364
rect 13998 9324 14004 9336
rect 14056 9324 14062 9376
rect 14553 9367 14611 9373
rect 14553 9333 14565 9367
rect 14599 9364 14611 9367
rect 14642 9364 14648 9376
rect 14599 9336 14648 9364
rect 14599 9333 14611 9336
rect 14553 9327 14611 9333
rect 14642 9324 14648 9336
rect 14700 9324 14706 9376
rect 15565 9367 15623 9373
rect 15565 9333 15577 9367
rect 15611 9364 15623 9367
rect 15856 9364 15884 9395
rect 18046 9392 18052 9444
rect 18104 9432 18110 9444
rect 18877 9435 18935 9441
rect 18877 9432 18889 9435
rect 18104 9404 18889 9432
rect 18104 9392 18110 9404
rect 18877 9401 18889 9404
rect 18923 9432 18935 9435
rect 19245 9435 19303 9441
rect 19245 9432 19257 9435
rect 18923 9404 19257 9432
rect 18923 9401 18935 9404
rect 18877 9395 18935 9401
rect 19245 9401 19257 9404
rect 19291 9401 19303 9435
rect 19245 9395 19303 9401
rect 19797 9435 19855 9441
rect 19797 9401 19809 9435
rect 19843 9432 19855 9435
rect 19886 9432 19892 9444
rect 19843 9404 19892 9432
rect 19843 9401 19855 9404
rect 19797 9395 19855 9401
rect 19886 9392 19892 9404
rect 19944 9392 19950 9444
rect 16206 9364 16212 9376
rect 15611 9336 16212 9364
rect 15611 9333 15623 9336
rect 15565 9327 15623 9333
rect 16206 9324 16212 9336
rect 16264 9324 16270 9376
rect 16761 9367 16819 9373
rect 16761 9333 16773 9367
rect 16807 9364 16819 9367
rect 16850 9364 16856 9376
rect 16807 9336 16856 9364
rect 16807 9333 16819 9336
rect 16761 9327 16819 9333
rect 16850 9324 16856 9336
rect 16908 9364 16914 9376
rect 18322 9364 18328 9376
rect 16908 9336 18328 9364
rect 16908 9324 16914 9336
rect 18322 9324 18328 9336
rect 18380 9324 18386 9376
rect 20714 9324 20720 9376
rect 20772 9364 20778 9376
rect 20901 9367 20959 9373
rect 20901 9364 20913 9367
rect 20772 9336 20913 9364
rect 20772 9324 20778 9336
rect 20901 9333 20913 9336
rect 20947 9333 20959 9367
rect 20901 9327 20959 9333
rect 1104 9274 22816 9296
rect 1104 9222 8982 9274
rect 9034 9222 9046 9274
rect 9098 9222 9110 9274
rect 9162 9222 9174 9274
rect 9226 9222 16982 9274
rect 17034 9222 17046 9274
rect 17098 9222 17110 9274
rect 17162 9222 17174 9274
rect 17226 9222 22816 9274
rect 1104 9200 22816 9222
rect 3513 9163 3571 9169
rect 3513 9129 3525 9163
rect 3559 9160 3571 9163
rect 3786 9160 3792 9172
rect 3559 9132 3792 9160
rect 3559 9129 3571 9132
rect 3513 9123 3571 9129
rect 3786 9120 3792 9132
rect 3844 9120 3850 9172
rect 4341 9163 4399 9169
rect 4341 9129 4353 9163
rect 4387 9160 4399 9163
rect 5258 9160 5264 9172
rect 4387 9132 5264 9160
rect 4387 9129 4399 9132
rect 4341 9123 4399 9129
rect 3145 9095 3203 9101
rect 3145 9061 3157 9095
rect 3191 9092 3203 9095
rect 3234 9092 3240 9104
rect 3191 9064 3240 9092
rect 3191 9061 3203 9064
rect 3145 9055 3203 9061
rect 3234 9052 3240 9064
rect 3292 9052 3298 9104
rect 1946 9024 1952 9036
rect 1907 8996 1952 9024
rect 1946 8984 1952 8996
rect 2004 8984 2010 9036
rect 2314 9024 2320 9036
rect 2275 8996 2320 9024
rect 2314 8984 2320 8996
rect 2372 8984 2378 9036
rect 2498 9024 2504 9036
rect 2459 8996 2504 9024
rect 2498 8984 2504 8996
rect 2556 8984 2562 9036
rect 2958 9024 2964 9036
rect 2919 8996 2964 9024
rect 2958 8984 2964 8996
rect 3016 9024 3022 9036
rect 4356 9024 4384 9123
rect 5258 9120 5264 9132
rect 5316 9120 5322 9172
rect 8386 9160 8392 9172
rect 8347 9132 8392 9160
rect 8386 9120 8392 9132
rect 8444 9120 8450 9172
rect 10318 9160 10324 9172
rect 10279 9132 10324 9160
rect 10318 9120 10324 9132
rect 10376 9120 10382 9172
rect 12802 9120 12808 9172
rect 12860 9160 12866 9172
rect 12897 9163 12955 9169
rect 12897 9160 12909 9163
rect 12860 9132 12909 9160
rect 12860 9120 12866 9132
rect 12897 9129 12909 9132
rect 12943 9129 12955 9163
rect 12897 9123 12955 9129
rect 12986 9120 12992 9172
rect 13044 9160 13050 9172
rect 14829 9163 14887 9169
rect 14829 9160 14841 9163
rect 13044 9132 14841 9160
rect 13044 9120 13050 9132
rect 14829 9129 14841 9132
rect 14875 9160 14887 9163
rect 14918 9160 14924 9172
rect 14875 9132 14924 9160
rect 14875 9129 14887 9132
rect 14829 9123 14887 9129
rect 14918 9120 14924 9132
rect 14976 9120 14982 9172
rect 15654 9160 15660 9172
rect 15615 9132 15660 9160
rect 15654 9120 15660 9132
rect 15712 9120 15718 9172
rect 16206 9160 16212 9172
rect 16167 9132 16212 9160
rect 16206 9120 16212 9132
rect 16264 9120 16270 9172
rect 19153 9163 19211 9169
rect 19153 9129 19165 9163
rect 19199 9160 19211 9163
rect 19242 9160 19248 9172
rect 19199 9132 19248 9160
rect 19199 9129 19211 9132
rect 19153 9123 19211 9129
rect 19242 9120 19248 9132
rect 19300 9120 19306 9172
rect 21039 9163 21097 9169
rect 21039 9129 21051 9163
rect 21085 9129 21097 9163
rect 21039 9123 21097 9129
rect 4798 9092 4804 9104
rect 4711 9064 4804 9092
rect 4798 9052 4804 9064
rect 4856 9092 4862 9104
rect 5902 9092 5908 9104
rect 4856 9064 5908 9092
rect 4856 9052 4862 9064
rect 5460 9033 5488 9064
rect 5902 9052 5908 9064
rect 5960 9052 5966 9104
rect 7098 9052 7104 9104
rect 7156 9092 7162 9104
rect 7790 9095 7848 9101
rect 7790 9092 7802 9095
rect 7156 9064 7802 9092
rect 7156 9052 7162 9064
rect 7790 9061 7802 9064
rect 7836 9061 7848 9095
rect 7790 9055 7848 9061
rect 9125 9095 9183 9101
rect 9125 9061 9137 9095
rect 9171 9092 9183 9095
rect 9306 9092 9312 9104
rect 9171 9064 9312 9092
rect 9171 9061 9183 9064
rect 9125 9055 9183 9061
rect 9306 9052 9312 9064
rect 9364 9092 9370 9104
rect 18046 9092 18052 9104
rect 9364 9064 11284 9092
rect 18007 9064 18052 9092
rect 9364 9052 9370 9064
rect 11256 9036 11284 9064
rect 18046 9052 18052 9064
rect 18104 9052 18110 9104
rect 20806 9052 20812 9104
rect 20864 9092 20870 9104
rect 21054 9092 21082 9123
rect 20864 9064 21082 9092
rect 20864 9052 20870 9064
rect 3016 8996 4384 9024
rect 5445 9027 5503 9033
rect 3016 8984 3022 8996
rect 5445 8993 5457 9027
rect 5491 8993 5503 9027
rect 5445 8987 5503 8993
rect 5629 9027 5687 9033
rect 5629 8993 5641 9027
rect 5675 8993 5687 9027
rect 5994 9024 6000 9036
rect 5955 8996 6000 9024
rect 5629 8987 5687 8993
rect 2332 8956 2360 8984
rect 3789 8959 3847 8965
rect 3789 8956 3801 8959
rect 2332 8928 3801 8956
rect 3789 8925 3801 8928
rect 3835 8956 3847 8959
rect 3970 8956 3976 8968
rect 3835 8928 3976 8956
rect 3835 8925 3847 8928
rect 3789 8919 3847 8925
rect 3970 8916 3976 8928
rect 4028 8916 4034 8968
rect 4338 8916 4344 8968
rect 4396 8956 4402 8968
rect 5644 8956 5672 8987
rect 5994 8984 6000 8996
rect 6052 8984 6058 9036
rect 6362 9024 6368 9036
rect 6323 8996 6368 9024
rect 6362 8984 6368 8996
rect 6420 8984 6426 9036
rect 9674 9024 9680 9036
rect 9635 8996 9680 9024
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 9858 9033 9864 9036
rect 9824 9027 9864 9033
rect 9824 9024 9836 9027
rect 9771 8996 9836 9024
rect 9824 8993 9836 8996
rect 9916 9024 9922 9036
rect 10594 9024 10600 9036
rect 9916 8996 10600 9024
rect 9824 8987 9864 8993
rect 9858 8984 9864 8987
rect 9916 8984 9922 8996
rect 10594 8984 10600 8996
rect 10652 8984 10658 9036
rect 11238 9024 11244 9036
rect 11199 8996 11244 9024
rect 11238 8984 11244 8996
rect 11296 8984 11302 9036
rect 11514 9024 11520 9036
rect 11475 8996 11520 9024
rect 11514 8984 11520 8996
rect 11572 8984 11578 9036
rect 11977 9027 12035 9033
rect 11977 8993 11989 9027
rect 12023 9024 12035 9027
rect 13906 9024 13912 9036
rect 12023 8996 13912 9024
rect 12023 8993 12035 8996
rect 11977 8987 12035 8993
rect 13906 8984 13912 8996
rect 13964 8984 13970 9036
rect 14185 9027 14243 9033
rect 14185 8993 14197 9027
rect 14231 9024 14243 9027
rect 14274 9024 14280 9036
rect 14231 8996 14280 9024
rect 14231 8993 14243 8996
rect 14185 8987 14243 8993
rect 14274 8984 14280 8996
rect 14332 8984 14338 9036
rect 20968 9027 21026 9033
rect 20968 8993 20980 9027
rect 21014 9024 21026 9027
rect 21266 9024 21272 9036
rect 21014 8996 21272 9024
rect 21014 8993 21026 8996
rect 20968 8987 21026 8993
rect 21266 8984 21272 8996
rect 21324 8984 21330 9036
rect 6454 8956 6460 8968
rect 4396 8928 6460 8956
rect 4396 8916 4402 8928
rect 6454 8916 6460 8928
rect 6512 8916 6518 8968
rect 6641 8959 6699 8965
rect 6641 8925 6653 8959
rect 6687 8956 6699 8959
rect 7466 8956 7472 8968
rect 6687 8928 7472 8956
rect 6687 8925 6699 8928
rect 6641 8919 6699 8925
rect 7466 8916 7472 8928
rect 7524 8916 7530 8968
rect 10045 8959 10103 8965
rect 10045 8956 10057 8959
rect 9600 8928 10057 8956
rect 9600 8832 9628 8928
rect 10045 8925 10057 8928
rect 10091 8956 10103 8959
rect 10686 8956 10692 8968
rect 10091 8928 10692 8956
rect 10091 8925 10103 8928
rect 10045 8919 10103 8925
rect 10686 8916 10692 8928
rect 10744 8916 10750 8968
rect 14369 8959 14427 8965
rect 14369 8925 14381 8959
rect 14415 8956 14427 8959
rect 15010 8956 15016 8968
rect 14415 8928 15016 8956
rect 14415 8925 14427 8928
rect 14369 8919 14427 8925
rect 15010 8916 15016 8928
rect 15068 8956 15074 8968
rect 15289 8959 15347 8965
rect 15289 8956 15301 8959
rect 15068 8928 15301 8956
rect 15068 8916 15074 8928
rect 15289 8925 15301 8928
rect 15335 8925 15347 8959
rect 17954 8956 17960 8968
rect 17915 8928 17960 8956
rect 15289 8919 15347 8925
rect 17954 8916 17960 8928
rect 18012 8916 18018 8968
rect 18598 8956 18604 8968
rect 18559 8928 18604 8956
rect 18598 8916 18604 8928
rect 18656 8916 18662 8968
rect 10778 8848 10784 8900
rect 10836 8888 10842 8900
rect 11333 8891 11391 8897
rect 11333 8888 11345 8891
rect 10836 8860 11345 8888
rect 10836 8848 10842 8860
rect 11333 8857 11345 8860
rect 11379 8857 11391 8891
rect 11333 8851 11391 8857
rect 9493 8823 9551 8829
rect 9493 8789 9505 8823
rect 9539 8820 9551 8823
rect 9582 8820 9588 8832
rect 9539 8792 9588 8820
rect 9539 8789 9551 8792
rect 9493 8783 9551 8789
rect 9582 8780 9588 8792
rect 9640 8780 9646 8832
rect 9953 8823 10011 8829
rect 9953 8789 9965 8823
rect 9999 8820 10011 8823
rect 10410 8820 10416 8832
rect 9999 8792 10416 8820
rect 9999 8789 10011 8792
rect 9953 8783 10011 8789
rect 10410 8780 10416 8792
rect 10468 8780 10474 8832
rect 1104 8730 22816 8752
rect 1104 8678 4982 8730
rect 5034 8678 5046 8730
rect 5098 8678 5110 8730
rect 5162 8678 5174 8730
rect 5226 8678 12982 8730
rect 13034 8678 13046 8730
rect 13098 8678 13110 8730
rect 13162 8678 13174 8730
rect 13226 8678 20982 8730
rect 21034 8678 21046 8730
rect 21098 8678 21110 8730
rect 21162 8678 21174 8730
rect 21226 8678 22816 8730
rect 1104 8656 22816 8678
rect 3970 8616 3976 8628
rect 3931 8588 3976 8616
rect 3970 8576 3976 8588
rect 4028 8616 4034 8628
rect 4338 8616 4344 8628
rect 4028 8588 4344 8616
rect 4028 8576 4034 8588
rect 4338 8576 4344 8588
rect 4396 8576 4402 8628
rect 4433 8619 4491 8625
rect 4433 8585 4445 8619
rect 4479 8616 4491 8619
rect 5537 8619 5595 8625
rect 5537 8616 5549 8619
rect 4479 8588 5549 8616
rect 4479 8585 4491 8588
rect 4433 8579 4491 8585
rect 5537 8585 5549 8588
rect 5583 8585 5595 8619
rect 6454 8616 6460 8628
rect 6415 8588 6460 8616
rect 5537 8579 5595 8585
rect 1762 8480 1768 8492
rect 1675 8452 1768 8480
rect 1762 8440 1768 8452
rect 1820 8480 1826 8492
rect 3142 8480 3148 8492
rect 1820 8452 3148 8480
rect 1820 8440 1826 8452
rect 3142 8440 3148 8452
rect 3200 8440 3206 8492
rect 3326 8480 3332 8492
rect 3287 8452 3332 8480
rect 3326 8440 3332 8452
rect 3384 8440 3390 8492
rect 3789 8483 3847 8489
rect 3789 8449 3801 8483
rect 3835 8480 3847 8483
rect 4448 8480 4476 8579
rect 6454 8576 6460 8588
rect 6512 8616 6518 8628
rect 14642 8616 14648 8628
rect 6512 8588 9536 8616
rect 14603 8588 14648 8616
rect 6512 8576 6518 8588
rect 4798 8548 4804 8560
rect 4759 8520 4804 8548
rect 4798 8508 4804 8520
rect 4856 8508 4862 8560
rect 6730 8508 6736 8560
rect 6788 8548 6794 8560
rect 9508 8557 9536 8588
rect 14642 8576 14648 8588
rect 14700 8616 14706 8628
rect 17405 8619 17463 8625
rect 17405 8616 17417 8619
rect 14700 8588 17417 8616
rect 14700 8576 14706 8588
rect 17405 8585 17417 8588
rect 17451 8616 17463 8619
rect 18046 8616 18052 8628
rect 17451 8588 18052 8616
rect 17451 8585 17463 8588
rect 17405 8579 17463 8585
rect 18046 8576 18052 8588
rect 18104 8576 18110 8628
rect 9125 8551 9183 8557
rect 9125 8548 9137 8551
rect 6788 8520 9137 8548
rect 6788 8508 6794 8520
rect 9125 8517 9137 8520
rect 9171 8517 9183 8551
rect 9125 8511 9183 8517
rect 9493 8551 9551 8557
rect 9493 8517 9505 8551
rect 9539 8548 9551 8551
rect 10778 8548 10784 8560
rect 9539 8520 10784 8548
rect 9539 8517 9551 8520
rect 9493 8511 9551 8517
rect 10778 8508 10784 8520
rect 10836 8508 10842 8560
rect 11103 8551 11161 8557
rect 11103 8517 11115 8551
rect 11149 8548 11161 8551
rect 17954 8548 17960 8560
rect 11149 8520 17960 8548
rect 11149 8517 11161 8520
rect 11103 8511 11161 8517
rect 17954 8508 17960 8520
rect 18012 8548 18018 8560
rect 19245 8551 19303 8557
rect 19245 8548 19257 8551
rect 18012 8520 19257 8548
rect 18012 8508 18018 8520
rect 19245 8517 19257 8520
rect 19291 8517 19303 8551
rect 19245 8511 19303 8517
rect 3835 8452 4476 8480
rect 5169 8483 5227 8489
rect 3835 8449 3847 8452
rect 3789 8443 3847 8449
rect 5169 8449 5181 8483
rect 5215 8480 5227 8483
rect 5626 8480 5632 8492
rect 5215 8452 5632 8480
rect 5215 8449 5227 8452
rect 5169 8443 5227 8449
rect 1946 8412 1952 8424
rect 1907 8384 1952 8412
rect 1946 8372 1952 8384
rect 2004 8372 2010 8424
rect 2130 8372 2136 8424
rect 2188 8412 2194 8424
rect 2317 8415 2375 8421
rect 2317 8412 2329 8415
rect 2188 8384 2329 8412
rect 2188 8372 2194 8384
rect 2317 8381 2329 8384
rect 2363 8381 2375 8415
rect 2317 8375 2375 8381
rect 2498 8372 2504 8424
rect 2556 8412 2562 8424
rect 2685 8415 2743 8421
rect 2685 8412 2697 8415
rect 2556 8384 2697 8412
rect 2556 8372 2562 8384
rect 2685 8381 2697 8384
rect 2731 8381 2743 8415
rect 3160 8412 3188 8440
rect 3237 8415 3295 8421
rect 3237 8412 3249 8415
rect 3160 8384 3249 8412
rect 2685 8375 2743 8381
rect 3237 8381 3249 8384
rect 3283 8412 3295 8415
rect 5184 8412 5212 8443
rect 5626 8440 5632 8452
rect 5684 8480 5690 8492
rect 6362 8480 6368 8492
rect 5684 8452 6368 8480
rect 5684 8440 5690 8452
rect 6362 8440 6368 8452
rect 6420 8440 6426 8492
rect 7098 8480 7104 8492
rect 7059 8452 7104 8480
rect 7098 8440 7104 8452
rect 7156 8440 7162 8492
rect 8849 8483 8907 8489
rect 8849 8480 8861 8483
rect 7576 8452 8861 8480
rect 3283 8384 5212 8412
rect 5445 8415 5503 8421
rect 3283 8381 3295 8384
rect 3237 8375 3295 8381
rect 5445 8381 5457 8415
rect 5491 8381 5503 8415
rect 5445 8375 5503 8381
rect 2700 8344 2728 8375
rect 3605 8347 3663 8353
rect 3605 8344 3617 8347
rect 2700 8316 3617 8344
rect 3605 8313 3617 8316
rect 3651 8344 3663 8347
rect 3789 8347 3847 8353
rect 3789 8344 3801 8347
rect 3651 8316 3801 8344
rect 3651 8313 3663 8316
rect 3605 8307 3663 8313
rect 3789 8313 3801 8316
rect 3835 8313 3847 8347
rect 3789 8307 3847 8313
rect 5261 8347 5319 8353
rect 5261 8313 5273 8347
rect 5307 8313 5319 8347
rect 5261 8307 5319 8313
rect 5276 8276 5304 8307
rect 5350 8304 5356 8356
rect 5408 8344 5414 8356
rect 5460 8344 5488 8375
rect 7282 8372 7288 8424
rect 7340 8412 7346 8424
rect 7576 8421 7604 8452
rect 8849 8449 8861 8452
rect 8895 8480 8907 8483
rect 9582 8480 9588 8492
rect 8895 8452 9588 8480
rect 8895 8449 8907 8452
rect 8849 8443 8907 8449
rect 9582 8440 9588 8452
rect 9640 8480 9646 8492
rect 9640 8452 9720 8480
rect 9640 8440 9646 8452
rect 7561 8415 7619 8421
rect 7561 8412 7573 8415
rect 7340 8384 7573 8412
rect 7340 8372 7346 8384
rect 7561 8381 7573 8384
rect 7607 8381 7619 8415
rect 8202 8412 8208 8424
rect 8163 8384 8208 8412
rect 7561 8375 7619 8381
rect 8202 8372 8208 8384
rect 8260 8372 8266 8424
rect 9306 8372 9312 8424
rect 9364 8412 9370 8424
rect 9692 8421 9720 8452
rect 9766 8440 9772 8492
rect 9824 8480 9830 8492
rect 9861 8483 9919 8489
rect 9861 8480 9873 8483
rect 9824 8452 9873 8480
rect 9824 8440 9830 8452
rect 9861 8449 9873 8452
rect 9907 8449 9919 8483
rect 9861 8443 9919 8449
rect 12713 8483 12771 8489
rect 12713 8449 12725 8483
rect 12759 8480 12771 8483
rect 13538 8480 13544 8492
rect 12759 8452 13400 8480
rect 13499 8452 13544 8480
rect 12759 8449 12771 8452
rect 12713 8443 12771 8449
rect 9401 8415 9459 8421
rect 9401 8412 9413 8415
rect 9364 8384 9413 8412
rect 9364 8372 9370 8384
rect 9401 8381 9413 8384
rect 9447 8381 9459 8415
rect 9401 8375 9459 8381
rect 9677 8415 9735 8421
rect 9677 8381 9689 8415
rect 9723 8381 9735 8415
rect 11000 8415 11058 8421
rect 11000 8412 11012 8415
rect 9677 8375 9735 8381
rect 9784 8384 11012 8412
rect 6181 8347 6239 8353
rect 6181 8344 6193 8347
rect 5408 8316 6193 8344
rect 5408 8304 5414 8316
rect 6181 8313 6193 8316
rect 6227 8344 6239 8347
rect 8478 8344 8484 8356
rect 6227 8316 8484 8344
rect 6227 8313 6239 8316
rect 6181 8307 6239 8313
rect 8478 8304 8484 8316
rect 8536 8304 8542 8356
rect 8846 8304 8852 8356
rect 8904 8344 8910 8356
rect 9217 8347 9275 8353
rect 9217 8344 9229 8347
rect 8904 8316 9229 8344
rect 8904 8304 8910 8316
rect 9217 8313 9229 8316
rect 9263 8313 9275 8347
rect 9217 8307 9275 8313
rect 5534 8276 5540 8288
rect 5276 8248 5540 8276
rect 5534 8236 5540 8248
rect 5592 8236 5598 8288
rect 7469 8279 7527 8285
rect 7469 8245 7481 8279
rect 7515 8276 7527 8279
rect 8202 8276 8208 8288
rect 7515 8248 8208 8276
rect 7515 8245 7527 8248
rect 7469 8239 7527 8245
rect 8202 8236 8208 8248
rect 8260 8236 8266 8288
rect 9125 8279 9183 8285
rect 9125 8245 9137 8279
rect 9171 8276 9183 8279
rect 9784 8276 9812 8384
rect 11000 8381 11012 8384
rect 11046 8412 11058 8415
rect 11793 8415 11851 8421
rect 11793 8412 11805 8415
rect 11046 8384 11805 8412
rect 11046 8381 11058 8384
rect 11000 8375 11058 8381
rect 11793 8381 11805 8384
rect 11839 8381 11851 8415
rect 11793 8375 11851 8381
rect 12989 8415 13047 8421
rect 12989 8381 13001 8415
rect 13035 8381 13047 8415
rect 12989 8375 13047 8381
rect 10410 8276 10416 8288
rect 9171 8248 9812 8276
rect 10371 8248 10416 8276
rect 9171 8245 9183 8248
rect 9125 8239 9183 8245
rect 10410 8236 10416 8248
rect 10468 8236 10474 8288
rect 10686 8236 10692 8288
rect 10744 8276 10750 8288
rect 11425 8279 11483 8285
rect 11425 8276 11437 8279
rect 10744 8248 11437 8276
rect 10744 8236 10750 8248
rect 11425 8245 11437 8248
rect 11471 8276 11483 8279
rect 11514 8276 11520 8288
rect 11471 8248 11520 8276
rect 11471 8245 11483 8248
rect 11425 8239 11483 8245
rect 11514 8236 11520 8248
rect 11572 8236 11578 8288
rect 13004 8276 13032 8375
rect 13262 8372 13268 8424
rect 13320 8412 13326 8424
rect 13372 8421 13400 8452
rect 13538 8440 13544 8452
rect 13596 8440 13602 8492
rect 14918 8480 14924 8492
rect 14879 8452 14924 8480
rect 14918 8440 14924 8452
rect 14976 8440 14982 8492
rect 15654 8440 15660 8492
rect 15712 8480 15718 8492
rect 15933 8483 15991 8489
rect 15933 8480 15945 8483
rect 15712 8452 15945 8480
rect 15712 8440 15718 8452
rect 15933 8449 15945 8452
rect 15979 8480 15991 8483
rect 17494 8480 17500 8492
rect 15979 8452 17500 8480
rect 15979 8449 15991 8452
rect 15933 8443 15991 8449
rect 17494 8440 17500 8452
rect 17552 8440 17558 8492
rect 18598 8440 18604 8492
rect 18656 8480 18662 8492
rect 20165 8483 20223 8489
rect 20165 8480 20177 8483
rect 18656 8452 20177 8480
rect 18656 8440 18662 8452
rect 20165 8449 20177 8452
rect 20211 8449 20223 8483
rect 20165 8443 20223 8449
rect 13357 8415 13415 8421
rect 13357 8412 13369 8415
rect 13320 8384 13369 8412
rect 13320 8372 13326 8384
rect 13357 8381 13369 8384
rect 13403 8412 13415 8415
rect 13446 8412 13452 8424
rect 13403 8384 13452 8412
rect 13403 8381 13415 8384
rect 13357 8375 13415 8381
rect 13446 8372 13452 8384
rect 13504 8372 13510 8424
rect 16393 8415 16451 8421
rect 16393 8412 16405 8415
rect 16224 8384 16405 8412
rect 14642 8304 14648 8356
rect 14700 8344 14706 8356
rect 15013 8347 15071 8353
rect 15013 8344 15025 8347
rect 14700 8316 15025 8344
rect 14700 8304 14706 8316
rect 15013 8313 15025 8316
rect 15059 8313 15071 8347
rect 15562 8344 15568 8356
rect 15523 8316 15568 8344
rect 15013 8307 15071 8313
rect 15562 8304 15568 8316
rect 15620 8304 15626 8356
rect 16224 8288 16252 8384
rect 16393 8381 16405 8384
rect 16439 8381 16451 8415
rect 16393 8375 16451 8381
rect 16758 8372 16764 8424
rect 16816 8412 16822 8424
rect 16853 8415 16911 8421
rect 16853 8412 16865 8415
rect 16816 8384 16865 8412
rect 16816 8372 16822 8384
rect 16853 8381 16865 8384
rect 16899 8381 16911 8415
rect 16853 8375 16911 8381
rect 17129 8415 17187 8421
rect 17129 8381 17141 8415
rect 17175 8412 17187 8415
rect 18046 8412 18052 8424
rect 17175 8384 18052 8412
rect 17175 8381 17187 8384
rect 17129 8375 17187 8381
rect 18046 8372 18052 8384
rect 18104 8372 18110 8424
rect 18322 8344 18328 8356
rect 18280 8316 18328 8344
rect 18322 8304 18328 8316
rect 18380 8353 18386 8356
rect 18380 8347 18428 8353
rect 18380 8313 18382 8347
rect 18416 8313 18428 8347
rect 18380 8307 18428 8313
rect 19889 8347 19947 8353
rect 19889 8313 19901 8347
rect 19935 8313 19947 8347
rect 19889 8307 19947 8313
rect 18380 8304 18413 8307
rect 13906 8276 13912 8288
rect 13004 8248 13912 8276
rect 13906 8236 13912 8248
rect 13964 8236 13970 8288
rect 14274 8276 14280 8288
rect 14235 8248 14280 8276
rect 14274 8236 14280 8248
rect 14332 8236 14338 8288
rect 16206 8276 16212 8288
rect 16167 8248 16212 8276
rect 16206 8236 16212 8248
rect 16264 8236 16270 8288
rect 17494 8236 17500 8288
rect 17552 8276 17558 8288
rect 17773 8279 17831 8285
rect 17773 8276 17785 8279
rect 17552 8248 17785 8276
rect 17552 8236 17558 8248
rect 17773 8245 17785 8248
rect 17819 8276 17831 8279
rect 18385 8276 18413 8304
rect 18966 8276 18972 8288
rect 17819 8248 18413 8276
rect 18927 8248 18972 8276
rect 17819 8245 17831 8248
rect 17773 8239 17831 8245
rect 18966 8236 18972 8248
rect 19024 8236 19030 8288
rect 19518 8236 19524 8288
rect 19576 8276 19582 8288
rect 19613 8279 19671 8285
rect 19613 8276 19625 8279
rect 19576 8248 19625 8276
rect 19576 8236 19582 8248
rect 19613 8245 19625 8248
rect 19659 8245 19671 8279
rect 19613 8239 19671 8245
rect 19794 8236 19800 8288
rect 19852 8276 19858 8288
rect 19904 8276 19932 8307
rect 19978 8304 19984 8356
rect 20036 8344 20042 8356
rect 20036 8316 20081 8344
rect 20036 8304 20042 8316
rect 19852 8248 19932 8276
rect 20993 8279 21051 8285
rect 19852 8236 19858 8248
rect 20993 8245 21005 8279
rect 21039 8276 21051 8279
rect 21266 8276 21272 8288
rect 21039 8248 21272 8276
rect 21039 8245 21051 8248
rect 20993 8239 21051 8245
rect 21266 8236 21272 8248
rect 21324 8276 21330 8288
rect 23198 8276 23204 8288
rect 21324 8248 23204 8276
rect 21324 8236 21330 8248
rect 23198 8236 23204 8248
rect 23256 8236 23262 8288
rect 1104 8186 22816 8208
rect 1104 8134 8982 8186
rect 9034 8134 9046 8186
rect 9098 8134 9110 8186
rect 9162 8134 9174 8186
rect 9226 8134 16982 8186
rect 17034 8134 17046 8186
rect 17098 8134 17110 8186
rect 17162 8134 17174 8186
rect 17226 8134 22816 8186
rect 1104 8112 22816 8134
rect 2314 8072 2320 8084
rect 2275 8044 2320 8072
rect 2314 8032 2320 8044
rect 2372 8032 2378 8084
rect 2958 8032 2964 8084
rect 3016 8072 3022 8084
rect 3053 8075 3111 8081
rect 3053 8072 3065 8075
rect 3016 8044 3065 8072
rect 3016 8032 3022 8044
rect 3053 8041 3065 8044
rect 3099 8072 3111 8075
rect 3418 8072 3424 8084
rect 3099 8044 3424 8072
rect 3099 8041 3111 8044
rect 3053 8035 3111 8041
rect 3418 8032 3424 8044
rect 3476 8032 3482 8084
rect 3513 8075 3571 8081
rect 3513 8041 3525 8075
rect 3559 8072 3571 8075
rect 3786 8072 3792 8084
rect 3559 8044 3792 8072
rect 3559 8041 3571 8044
rect 3513 8035 3571 8041
rect 3786 8032 3792 8044
rect 3844 8072 3850 8084
rect 4246 8072 4252 8084
rect 3844 8044 4252 8072
rect 3844 8032 3850 8044
rect 4246 8032 4252 8044
rect 4304 8072 4310 8084
rect 7282 8072 7288 8084
rect 4304 8044 7288 8072
rect 4304 8032 4310 8044
rect 7282 8032 7288 8044
rect 7340 8032 7346 8084
rect 7466 8072 7472 8084
rect 7427 8044 7472 8072
rect 7466 8032 7472 8044
rect 7524 8032 7530 8084
rect 9401 8075 9459 8081
rect 9401 8072 9413 8075
rect 8588 8044 9413 8072
rect 5353 8007 5411 8013
rect 5353 7973 5365 8007
rect 5399 8004 5411 8007
rect 5534 8004 5540 8016
rect 5399 7976 5540 8004
rect 5399 7973 5411 7976
rect 5353 7967 5411 7973
rect 5534 7964 5540 7976
rect 5592 7964 5598 8016
rect 8588 8013 8616 8044
rect 9401 8041 9413 8044
rect 9447 8072 9459 8075
rect 9582 8072 9588 8084
rect 9447 8044 9588 8072
rect 9447 8041 9459 8044
rect 9401 8035 9459 8041
rect 9582 8032 9588 8044
rect 9640 8072 9646 8084
rect 9858 8072 9864 8084
rect 9640 8044 9864 8072
rect 9640 8032 9646 8044
rect 9858 8032 9864 8044
rect 9916 8032 9922 8084
rect 11238 8032 11244 8084
rect 11296 8072 11302 8084
rect 11609 8075 11667 8081
rect 11609 8072 11621 8075
rect 11296 8044 11621 8072
rect 11296 8032 11302 8044
rect 11609 8041 11621 8044
rect 11655 8041 11667 8075
rect 11609 8035 11667 8041
rect 13817 8075 13875 8081
rect 13817 8041 13829 8075
rect 13863 8072 13875 8075
rect 13998 8072 14004 8084
rect 13863 8044 14004 8072
rect 13863 8041 13875 8044
rect 13817 8035 13875 8041
rect 13998 8032 14004 8044
rect 14056 8032 14062 8084
rect 15010 8072 15016 8084
rect 14971 8044 15016 8072
rect 15010 8032 15016 8044
rect 15068 8032 15074 8084
rect 15378 8072 15384 8084
rect 15339 8044 15384 8072
rect 15378 8032 15384 8044
rect 15436 8032 15442 8084
rect 16485 8075 16543 8081
rect 16485 8041 16497 8075
rect 16531 8072 16543 8075
rect 16758 8072 16764 8084
rect 16531 8044 16764 8072
rect 16531 8041 16543 8044
rect 16485 8035 16543 8041
rect 8573 8007 8631 8013
rect 8573 7973 8585 8007
rect 8619 7973 8631 8007
rect 9876 8004 9904 8032
rect 9876 7976 10410 8004
rect 8573 7967 8631 7973
rect 1946 7896 1952 7948
rect 2004 7936 2010 7948
rect 2130 7936 2136 7948
rect 2004 7908 2136 7936
rect 2004 7896 2010 7908
rect 2130 7896 2136 7908
rect 2188 7896 2194 7948
rect 8478 7936 8484 7948
rect 8439 7908 8484 7936
rect 8478 7896 8484 7908
rect 8536 7896 8542 7948
rect 8846 7896 8852 7948
rect 8904 7936 8910 7948
rect 9674 7936 9680 7948
rect 8904 7908 9680 7936
rect 8904 7896 8910 7908
rect 9674 7896 9680 7908
rect 9732 7936 9738 7948
rect 10226 7936 10232 7948
rect 9732 7908 10232 7936
rect 9732 7896 9738 7908
rect 10226 7896 10232 7908
rect 10284 7896 10290 7948
rect 10382 7945 10410 7976
rect 11054 7964 11060 8016
rect 11112 8004 11118 8016
rect 16206 8004 16212 8016
rect 11112 7976 16212 8004
rect 11112 7964 11118 7976
rect 11808 7948 11836 7976
rect 16206 7964 16212 7976
rect 16264 7964 16270 8016
rect 10376 7939 10434 7945
rect 10376 7905 10388 7939
rect 10422 7905 10434 7939
rect 10778 7936 10784 7948
rect 10376 7899 10434 7905
rect 10520 7908 10784 7936
rect 5902 7868 5908 7880
rect 5863 7840 5908 7868
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 5442 7760 5448 7812
rect 5500 7800 5506 7812
rect 10520 7809 10548 7908
rect 10778 7896 10784 7908
rect 10836 7936 10842 7948
rect 11146 7936 11152 7948
rect 10836 7908 11152 7936
rect 10836 7896 10842 7908
rect 11146 7896 11152 7908
rect 11204 7936 11210 7948
rect 11241 7939 11299 7945
rect 11241 7936 11253 7939
rect 11204 7908 11253 7936
rect 11204 7896 11210 7908
rect 11241 7905 11253 7908
rect 11287 7905 11299 7939
rect 11790 7936 11796 7948
rect 11703 7908 11796 7936
rect 11241 7899 11299 7905
rect 11790 7896 11796 7908
rect 11848 7896 11854 7948
rect 11882 7896 11888 7948
rect 11940 7936 11946 7948
rect 12253 7939 12311 7945
rect 12253 7936 12265 7939
rect 11940 7908 12265 7936
rect 11940 7896 11946 7908
rect 12253 7905 12265 7908
rect 12299 7905 12311 7939
rect 12253 7899 12311 7905
rect 12897 7939 12955 7945
rect 12897 7905 12909 7939
rect 12943 7936 12955 7939
rect 13906 7936 13912 7948
rect 12943 7908 13912 7936
rect 12943 7905 12955 7908
rect 12897 7899 12955 7905
rect 13906 7896 13912 7908
rect 13964 7936 13970 7948
rect 15565 7939 15623 7945
rect 15565 7936 15577 7939
rect 13964 7908 15577 7936
rect 13964 7896 13970 7908
rect 15565 7905 15577 7908
rect 15611 7905 15623 7939
rect 15565 7899 15623 7905
rect 15841 7939 15899 7945
rect 15841 7905 15853 7939
rect 15887 7936 15899 7939
rect 15930 7936 15936 7948
rect 15887 7908 15936 7936
rect 15887 7905 15899 7908
rect 15841 7899 15899 7905
rect 10597 7871 10655 7877
rect 10597 7837 10609 7871
rect 10643 7837 10655 7871
rect 12434 7868 12440 7880
rect 12395 7840 12440 7868
rect 10597 7831 10655 7837
rect 5813 7803 5871 7809
rect 5813 7800 5825 7803
rect 5500 7772 5825 7800
rect 5500 7760 5506 7772
rect 5813 7769 5825 7772
rect 5859 7769 5871 7803
rect 5813 7763 5871 7769
rect 10505 7803 10563 7809
rect 10505 7769 10517 7803
rect 10551 7769 10563 7803
rect 10505 7763 10563 7769
rect 10612 7800 10640 7831
rect 12434 7828 12440 7840
rect 12492 7828 12498 7880
rect 13446 7868 13452 7880
rect 13407 7840 13452 7868
rect 13446 7828 13452 7840
rect 13504 7828 13510 7880
rect 15580 7868 15608 7899
rect 15930 7896 15936 7908
rect 15988 7896 15994 7948
rect 15654 7868 15660 7880
rect 15567 7840 15660 7868
rect 15654 7828 15660 7840
rect 15712 7868 15718 7880
rect 16500 7868 16528 8035
rect 16758 8032 16764 8044
rect 16816 8032 16822 8084
rect 18046 8072 18052 8084
rect 18007 8044 18052 8072
rect 18046 8032 18052 8044
rect 18104 8032 18110 8084
rect 19518 8032 19524 8084
rect 19576 8072 19582 8084
rect 19978 8072 19984 8084
rect 19576 8044 19984 8072
rect 19576 8032 19582 8044
rect 19978 8032 19984 8044
rect 20036 8032 20042 8084
rect 17862 7964 17868 8016
rect 17920 8004 17926 8016
rect 18601 8007 18659 8013
rect 18601 8004 18613 8007
rect 17920 7976 18613 8004
rect 17920 7964 17926 7976
rect 18601 7973 18613 7976
rect 18647 8004 18659 8007
rect 18966 8004 18972 8016
rect 18647 7976 18972 8004
rect 18647 7973 18659 7976
rect 18601 7967 18659 7973
rect 18966 7964 18972 7976
rect 19024 7964 19030 8016
rect 19150 8004 19156 8016
rect 19111 7976 19156 8004
rect 19150 7964 19156 7976
rect 19208 7964 19214 8016
rect 16850 7936 16856 7948
rect 16811 7908 16856 7936
rect 16850 7896 16856 7908
rect 16908 7896 16914 7948
rect 18506 7868 18512 7880
rect 15712 7840 16528 7868
rect 18467 7840 18512 7868
rect 15712 7828 15718 7840
rect 18506 7828 18512 7840
rect 18564 7828 18570 7880
rect 18598 7828 18604 7880
rect 18656 7868 18662 7880
rect 20901 7871 20959 7877
rect 20901 7868 20913 7871
rect 18656 7840 20913 7868
rect 18656 7828 18662 7840
rect 20901 7837 20913 7840
rect 20947 7837 20959 7871
rect 20901 7831 20959 7837
rect 10778 7800 10784 7812
rect 10612 7772 10784 7800
rect 1946 7732 1952 7744
rect 1907 7704 1952 7732
rect 1946 7692 1952 7704
rect 2004 7692 2010 7744
rect 5350 7692 5356 7744
rect 5408 7732 5414 7744
rect 5675 7735 5733 7741
rect 5675 7732 5687 7735
rect 5408 7704 5687 7732
rect 5408 7692 5414 7704
rect 5675 7701 5687 7704
rect 5721 7701 5733 7735
rect 6178 7732 6184 7744
rect 6139 7704 6184 7732
rect 5675 7695 5733 7701
rect 6178 7692 6184 7704
rect 6236 7692 6242 7744
rect 8202 7692 8208 7744
rect 8260 7732 8266 7744
rect 10612 7732 10640 7772
rect 10778 7760 10784 7772
rect 10836 7760 10842 7812
rect 10873 7803 10931 7809
rect 10873 7769 10885 7803
rect 10919 7800 10931 7803
rect 12710 7800 12716 7812
rect 10919 7772 12716 7800
rect 10919 7769 10931 7772
rect 10873 7763 10931 7769
rect 12710 7760 12716 7772
rect 12768 7760 12774 7812
rect 14366 7732 14372 7744
rect 8260 7704 10640 7732
rect 14327 7704 14372 7732
rect 8260 7692 8266 7704
rect 14366 7692 14372 7704
rect 14424 7692 14430 7744
rect 16482 7692 16488 7744
rect 16540 7732 16546 7744
rect 16991 7735 17049 7741
rect 16991 7732 17003 7735
rect 16540 7704 17003 7732
rect 16540 7692 16546 7704
rect 16991 7701 17003 7704
rect 17037 7701 17049 7735
rect 19426 7732 19432 7744
rect 19387 7704 19432 7732
rect 16991 7695 17049 7701
rect 19426 7692 19432 7704
rect 19484 7692 19490 7744
rect 19794 7732 19800 7744
rect 19755 7704 19800 7732
rect 19794 7692 19800 7704
rect 19852 7692 19858 7744
rect 1104 7642 22816 7664
rect 1104 7590 4982 7642
rect 5034 7590 5046 7642
rect 5098 7590 5110 7642
rect 5162 7590 5174 7642
rect 5226 7590 12982 7642
rect 13034 7590 13046 7642
rect 13098 7590 13110 7642
rect 13162 7590 13174 7642
rect 13226 7590 20982 7642
rect 21034 7590 21046 7642
rect 21098 7590 21110 7642
rect 21162 7590 21174 7642
rect 21226 7590 22816 7642
rect 1104 7568 22816 7590
rect 1578 7528 1584 7540
rect 1539 7500 1584 7528
rect 1578 7488 1584 7500
rect 1636 7488 1642 7540
rect 2498 7528 2504 7540
rect 2459 7500 2504 7528
rect 2498 7488 2504 7500
rect 2556 7488 2562 7540
rect 2682 7488 2688 7540
rect 2740 7528 2746 7540
rect 3605 7531 3663 7537
rect 3605 7528 3617 7531
rect 2740 7500 3617 7528
rect 2740 7488 2746 7500
rect 3605 7497 3617 7500
rect 3651 7497 3663 7531
rect 3605 7491 3663 7497
rect 3789 7531 3847 7537
rect 3789 7497 3801 7531
rect 3835 7528 3847 7531
rect 4062 7528 4068 7540
rect 3835 7500 4068 7528
rect 3835 7497 3847 7500
rect 3789 7491 3847 7497
rect 1486 7392 1492 7404
rect 1412 7364 1492 7392
rect 1412 7333 1440 7364
rect 1486 7352 1492 7364
rect 1544 7352 1550 7404
rect 3620 7392 3648 7491
rect 4062 7488 4068 7500
rect 4120 7528 4126 7540
rect 5077 7531 5135 7537
rect 5077 7528 5089 7531
rect 4120 7500 5089 7528
rect 4120 7488 4126 7500
rect 5077 7497 5089 7500
rect 5123 7497 5135 7531
rect 5077 7491 5135 7497
rect 5261 7531 5319 7537
rect 5261 7497 5273 7531
rect 5307 7528 5319 7531
rect 5350 7528 5356 7540
rect 5307 7500 5356 7528
rect 5307 7497 5319 7500
rect 5261 7491 5319 7497
rect 3878 7420 3884 7472
rect 3936 7460 3942 7472
rect 5276 7460 5304 7491
rect 5350 7488 5356 7500
rect 5408 7488 5414 7540
rect 6641 7531 6699 7537
rect 6641 7497 6653 7531
rect 6687 7528 6699 7531
rect 6730 7528 6736 7540
rect 6687 7500 6736 7528
rect 6687 7497 6699 7500
rect 6641 7491 6699 7497
rect 6730 7488 6736 7500
rect 6788 7488 6794 7540
rect 7469 7531 7527 7537
rect 7469 7497 7481 7531
rect 7515 7528 7527 7531
rect 7742 7528 7748 7540
rect 7515 7500 7748 7528
rect 7515 7497 7527 7500
rect 7469 7491 7527 7497
rect 7742 7488 7748 7500
rect 7800 7488 7806 7540
rect 8478 7488 8484 7540
rect 8536 7528 8542 7540
rect 8573 7531 8631 7537
rect 8573 7528 8585 7531
rect 8536 7500 8585 7528
rect 8536 7488 8542 7500
rect 8573 7497 8585 7500
rect 8619 7497 8631 7531
rect 8573 7491 8631 7497
rect 9306 7488 9312 7540
rect 9364 7528 9370 7540
rect 9401 7531 9459 7537
rect 9401 7528 9413 7531
rect 9364 7500 9413 7528
rect 9364 7488 9370 7500
rect 9401 7497 9413 7500
rect 9447 7528 9459 7531
rect 10134 7528 10140 7540
rect 9447 7500 10140 7528
rect 9447 7497 9459 7500
rect 9401 7491 9459 7497
rect 10134 7488 10140 7500
rect 10192 7488 10198 7540
rect 10226 7488 10232 7540
rect 10284 7528 10290 7540
rect 11149 7531 11207 7537
rect 11149 7528 11161 7531
rect 10284 7500 11161 7528
rect 10284 7488 10290 7500
rect 11149 7497 11161 7500
rect 11195 7497 11207 7531
rect 11882 7528 11888 7540
rect 11843 7500 11888 7528
rect 11149 7491 11207 7497
rect 11882 7488 11888 7500
rect 11940 7488 11946 7540
rect 13446 7488 13452 7540
rect 13504 7528 13510 7540
rect 14093 7531 14151 7537
rect 14093 7528 14105 7531
rect 13504 7500 14105 7528
rect 13504 7488 13510 7500
rect 14093 7497 14105 7500
rect 14139 7528 14151 7531
rect 15378 7528 15384 7540
rect 14139 7500 15384 7528
rect 14139 7497 14151 7500
rect 14093 7491 14151 7497
rect 15378 7488 15384 7500
rect 15436 7488 15442 7540
rect 15654 7528 15660 7540
rect 15615 7500 15660 7528
rect 15654 7488 15660 7500
rect 15712 7488 15718 7540
rect 15841 7531 15899 7537
rect 15841 7497 15853 7531
rect 15887 7528 15899 7531
rect 17862 7528 17868 7540
rect 15887 7500 17033 7528
rect 17823 7500 17868 7528
rect 15887 7497 15899 7500
rect 15841 7491 15899 7497
rect 3936 7432 5304 7460
rect 3936 7420 3942 7432
rect 5902 7420 5908 7472
rect 5960 7460 5966 7472
rect 6273 7463 6331 7469
rect 6273 7460 6285 7463
rect 5960 7432 6285 7460
rect 5960 7420 5966 7432
rect 6273 7429 6285 7432
rect 6319 7460 6331 7463
rect 8202 7460 8208 7472
rect 6319 7432 8208 7460
rect 6319 7429 6331 7432
rect 6273 7423 6331 7429
rect 8202 7420 8208 7432
rect 8260 7420 8266 7472
rect 13725 7463 13783 7469
rect 13725 7429 13737 7463
rect 13771 7460 13783 7463
rect 13998 7460 14004 7472
rect 13771 7432 14004 7460
rect 13771 7429 13783 7432
rect 13725 7423 13783 7429
rect 4249 7395 4307 7401
rect 4249 7392 4261 7395
rect 3620 7364 4261 7392
rect 4249 7361 4261 7364
rect 4295 7361 4307 7395
rect 4249 7355 4307 7361
rect 4893 7395 4951 7401
rect 4893 7361 4905 7395
rect 4939 7392 4951 7395
rect 7650 7392 7656 7404
rect 4939 7364 7656 7392
rect 4939 7361 4951 7364
rect 4893 7355 4951 7361
rect 7650 7352 7656 7364
rect 7708 7392 7714 7404
rect 7929 7395 7987 7401
rect 7929 7392 7941 7395
rect 7708 7364 7941 7392
rect 7708 7352 7714 7364
rect 7929 7361 7941 7364
rect 7975 7361 7987 7395
rect 7929 7355 7987 7361
rect 9217 7395 9275 7401
rect 9217 7361 9229 7395
rect 9263 7392 9275 7395
rect 12434 7392 12440 7404
rect 9263 7364 9996 7392
rect 12395 7364 12440 7392
rect 9263 7361 9275 7364
rect 9217 7355 9275 7361
rect 9968 7336 9996 7364
rect 12434 7352 12440 7364
rect 12492 7352 12498 7404
rect 1397 7327 1455 7333
rect 1397 7293 1409 7327
rect 1443 7293 1455 7327
rect 1397 7287 1455 7293
rect 5077 7327 5135 7333
rect 5077 7293 5089 7327
rect 5123 7324 5135 7327
rect 5442 7324 5448 7336
rect 5123 7296 5448 7324
rect 5123 7293 5135 7296
rect 5077 7287 5135 7293
rect 5442 7284 5448 7296
rect 5500 7324 5506 7336
rect 5537 7327 5595 7333
rect 5537 7324 5549 7327
rect 5500 7296 5549 7324
rect 5500 7284 5506 7296
rect 5537 7293 5549 7296
rect 5583 7293 5595 7327
rect 5537 7287 5595 7293
rect 5772 7327 5830 7333
rect 5772 7293 5784 7327
rect 5818 7324 5830 7327
rect 6730 7324 6736 7336
rect 5818 7296 6736 7324
rect 5818 7293 5830 7296
rect 5772 7287 5830 7293
rect 6730 7284 6736 7296
rect 6788 7284 6794 7336
rect 9582 7324 9588 7336
rect 9543 7296 9588 7324
rect 9582 7284 9588 7296
rect 9640 7284 9646 7336
rect 9950 7324 9956 7336
rect 9911 7296 9956 7324
rect 9950 7284 9956 7296
rect 10008 7284 10014 7336
rect 10045 7327 10103 7333
rect 10045 7293 10057 7327
rect 10091 7293 10103 7327
rect 10045 7287 10103 7293
rect 4341 7259 4399 7265
rect 4341 7225 4353 7259
rect 4387 7225 4399 7259
rect 4341 7219 4399 7225
rect 5859 7259 5917 7265
rect 5859 7225 5871 7259
rect 5905 7256 5917 7259
rect 7009 7259 7067 7265
rect 7009 7256 7021 7259
rect 5905 7228 7021 7256
rect 5905 7225 5917 7228
rect 5859 7219 5917 7225
rect 7009 7225 7021 7228
rect 7055 7256 7067 7259
rect 7653 7259 7711 7265
rect 7653 7256 7665 7259
rect 7055 7228 7665 7256
rect 7055 7225 7067 7228
rect 7009 7219 7067 7225
rect 7653 7225 7665 7228
rect 7699 7225 7711 7259
rect 7653 7219 7711 7225
rect 1946 7148 1952 7200
rect 2004 7188 2010 7200
rect 2133 7191 2191 7197
rect 2133 7188 2145 7191
rect 2004 7160 2145 7188
rect 2004 7148 2010 7160
rect 2133 7157 2145 7160
rect 2179 7188 2191 7191
rect 2590 7188 2596 7200
rect 2179 7160 2596 7188
rect 2179 7157 2191 7160
rect 2133 7151 2191 7157
rect 2590 7148 2596 7160
rect 2648 7188 2654 7200
rect 3789 7191 3847 7197
rect 3789 7188 3801 7191
rect 2648 7160 3801 7188
rect 2648 7148 2654 7160
rect 3789 7157 3801 7160
rect 3835 7157 3847 7191
rect 3789 7151 3847 7157
rect 4065 7191 4123 7197
rect 4065 7157 4077 7191
rect 4111 7188 4123 7191
rect 4356 7188 4384 7219
rect 7742 7216 7748 7268
rect 7800 7256 7806 7268
rect 7800 7228 7845 7256
rect 7800 7216 7806 7228
rect 9306 7216 9312 7268
rect 9364 7256 9370 7268
rect 10060 7256 10088 7287
rect 9364 7228 10088 7256
rect 12253 7259 12311 7265
rect 9364 7216 9370 7228
rect 12253 7225 12265 7259
rect 12299 7256 12311 7259
rect 12526 7256 12532 7268
rect 12299 7228 12532 7256
rect 12299 7225 12311 7228
rect 12253 7219 12311 7225
rect 12526 7216 12532 7228
rect 12584 7256 12590 7268
rect 12799 7259 12857 7265
rect 12799 7256 12811 7259
rect 12584 7228 12811 7256
rect 12584 7216 12590 7228
rect 12799 7225 12811 7228
rect 12845 7256 12857 7259
rect 13740 7256 13768 7423
rect 13998 7420 14004 7432
rect 14056 7420 14062 7472
rect 14366 7460 14372 7472
rect 14327 7432 14372 7460
rect 14366 7420 14372 7432
rect 14424 7460 14430 7472
rect 14734 7460 14740 7472
rect 14424 7432 14740 7460
rect 14424 7420 14430 7432
rect 14734 7420 14740 7432
rect 14792 7420 14798 7472
rect 15197 7463 15255 7469
rect 15197 7429 15209 7463
rect 15243 7460 15255 7463
rect 15562 7460 15568 7472
rect 15243 7432 15568 7460
rect 15243 7429 15255 7432
rect 15197 7423 15255 7429
rect 15562 7420 15568 7432
rect 15620 7460 15626 7472
rect 16761 7463 16819 7469
rect 16761 7460 16773 7463
rect 15620 7432 16773 7460
rect 15620 7420 15626 7432
rect 16761 7429 16773 7432
rect 16807 7429 16819 7463
rect 17005 7460 17033 7500
rect 17862 7488 17868 7500
rect 17920 7488 17926 7540
rect 18463 7531 18521 7537
rect 18463 7497 18475 7531
rect 18509 7528 18521 7531
rect 19794 7528 19800 7540
rect 18509 7500 19800 7528
rect 18509 7497 18521 7500
rect 18463 7491 18521 7497
rect 19794 7488 19800 7500
rect 19852 7488 19858 7540
rect 19153 7463 19211 7469
rect 19153 7460 19165 7463
rect 17005 7432 19165 7460
rect 16761 7423 16819 7429
rect 19153 7429 19165 7432
rect 19199 7460 19211 7463
rect 19518 7460 19524 7472
rect 19199 7432 19524 7460
rect 19199 7429 19211 7432
rect 19153 7423 19211 7429
rect 19518 7420 19524 7432
rect 19576 7420 19582 7472
rect 15930 7392 15936 7404
rect 15891 7364 15936 7392
rect 15930 7352 15936 7364
rect 15988 7352 15994 7404
rect 16209 7395 16267 7401
rect 16209 7361 16221 7395
rect 16255 7392 16267 7395
rect 16482 7392 16488 7404
rect 16255 7364 16488 7392
rect 16255 7361 16267 7364
rect 16209 7355 16267 7361
rect 16482 7352 16488 7364
rect 16540 7352 16546 7404
rect 18877 7395 18935 7401
rect 18877 7361 18889 7395
rect 18923 7392 18935 7395
rect 19242 7392 19248 7404
rect 18923 7364 19248 7392
rect 18923 7361 18935 7364
rect 18877 7355 18935 7361
rect 18230 7284 18236 7336
rect 18288 7324 18294 7336
rect 18392 7327 18450 7333
rect 18392 7324 18404 7327
rect 18288 7296 18404 7324
rect 18288 7284 18294 7296
rect 18392 7293 18404 7296
rect 18438 7324 18450 7327
rect 18892 7324 18920 7355
rect 19242 7352 19248 7364
rect 19300 7352 19306 7404
rect 19886 7392 19892 7404
rect 19847 7364 19892 7392
rect 19886 7352 19892 7364
rect 19944 7352 19950 7404
rect 18438 7296 18920 7324
rect 18438 7293 18450 7296
rect 18392 7287 18450 7293
rect 12845 7228 13768 7256
rect 14645 7259 14703 7265
rect 12845 7225 12857 7228
rect 12799 7219 12857 7225
rect 14645 7225 14657 7259
rect 14691 7225 14703 7259
rect 14645 7219 14703 7225
rect 4614 7188 4620 7200
rect 4111 7160 4620 7188
rect 4111 7157 4123 7160
rect 4065 7151 4123 7157
rect 4614 7148 4620 7160
rect 4672 7188 4678 7200
rect 4982 7188 4988 7200
rect 4672 7160 4988 7188
rect 4672 7148 4678 7160
rect 4982 7148 4988 7160
rect 5040 7148 5046 7200
rect 10778 7188 10784 7200
rect 10739 7160 10784 7188
rect 10778 7148 10784 7160
rect 10836 7148 10842 7200
rect 11330 7188 11336 7200
rect 11291 7160 11336 7188
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 13354 7188 13360 7200
rect 13315 7160 13360 7188
rect 13354 7148 13360 7160
rect 13412 7148 13418 7200
rect 14550 7148 14556 7200
rect 14608 7188 14614 7200
rect 14660 7188 14688 7219
rect 14734 7216 14740 7268
rect 14792 7256 14798 7268
rect 15841 7259 15899 7265
rect 15841 7256 15853 7259
rect 14792 7228 15853 7256
rect 14792 7216 14798 7228
rect 15841 7225 15853 7228
rect 15887 7225 15899 7259
rect 16298 7256 16304 7268
rect 16259 7228 16304 7256
rect 15841 7219 15899 7225
rect 16298 7216 16304 7228
rect 16356 7216 16362 7268
rect 19426 7256 19432 7268
rect 19387 7228 19432 7256
rect 19426 7216 19432 7228
rect 19484 7216 19490 7268
rect 19518 7216 19524 7268
rect 19576 7256 19582 7268
rect 19576 7228 19621 7256
rect 19576 7216 19582 7228
rect 14608 7160 14688 7188
rect 14608 7148 14614 7160
rect 16022 7148 16028 7200
rect 16080 7188 16086 7200
rect 16850 7188 16856 7200
rect 16080 7160 16856 7188
rect 16080 7148 16086 7160
rect 16850 7148 16856 7160
rect 16908 7188 16914 7200
rect 17129 7191 17187 7197
rect 17129 7188 17141 7191
rect 16908 7160 17141 7188
rect 16908 7148 16914 7160
rect 17129 7157 17141 7160
rect 17175 7157 17187 7191
rect 17129 7151 17187 7157
rect 19610 7148 19616 7200
rect 19668 7188 19674 7200
rect 20901 7191 20959 7197
rect 20901 7188 20913 7191
rect 19668 7160 20913 7188
rect 19668 7148 19674 7160
rect 20901 7157 20913 7160
rect 20947 7157 20959 7191
rect 20901 7151 20959 7157
rect 1104 7098 22816 7120
rect 1104 7046 8982 7098
rect 9034 7046 9046 7098
rect 9098 7046 9110 7098
rect 9162 7046 9174 7098
rect 9226 7046 16982 7098
rect 17034 7046 17046 7098
rect 17098 7046 17110 7098
rect 17162 7046 17174 7098
rect 17226 7046 22816 7098
rect 1104 7024 22816 7046
rect 1486 6944 1492 6996
rect 1544 6984 1550 6996
rect 1581 6987 1639 6993
rect 1581 6984 1593 6987
rect 1544 6956 1593 6984
rect 1544 6944 1550 6956
rect 1581 6953 1593 6956
rect 1627 6953 1639 6987
rect 4982 6984 4988 6996
rect 4943 6956 4988 6984
rect 1581 6947 1639 6953
rect 4982 6944 4988 6956
rect 5040 6944 5046 6996
rect 5534 6944 5540 6996
rect 5592 6984 5598 6996
rect 5629 6987 5687 6993
rect 5629 6984 5641 6987
rect 5592 6956 5641 6984
rect 5592 6944 5598 6956
rect 5629 6953 5641 6956
rect 5675 6984 5687 6987
rect 5675 6956 8800 6984
rect 5675 6953 5687 6956
rect 5629 6947 5687 6953
rect 4062 6876 4068 6928
rect 4120 6916 4126 6928
rect 4430 6925 4436 6928
rect 4427 6916 4436 6925
rect 4120 6888 4436 6916
rect 4120 6876 4126 6888
rect 4427 6879 4436 6888
rect 4430 6876 4436 6879
rect 4488 6876 4494 6928
rect 6819 6919 6877 6925
rect 6819 6885 6831 6919
rect 6865 6916 6877 6919
rect 7098 6916 7104 6928
rect 6865 6888 7104 6916
rect 6865 6885 6877 6888
rect 6819 6879 6877 6885
rect 7098 6876 7104 6888
rect 7156 6876 7162 6928
rect 8772 6925 8800 6956
rect 9582 6944 9588 6996
rect 9640 6984 9646 6996
rect 9953 6987 10011 6993
rect 9953 6984 9965 6987
rect 9640 6956 9965 6984
rect 9640 6944 9646 6956
rect 9953 6953 9965 6956
rect 9999 6953 10011 6987
rect 11146 6984 11152 6996
rect 11107 6956 11152 6984
rect 9953 6947 10011 6953
rect 11146 6944 11152 6956
rect 11204 6944 11210 6996
rect 11790 6984 11796 6996
rect 11751 6956 11796 6984
rect 11790 6944 11796 6956
rect 11848 6944 11854 6996
rect 12434 6984 12440 6996
rect 12395 6956 12440 6984
rect 12434 6944 12440 6956
rect 12492 6944 12498 6996
rect 12710 6944 12716 6996
rect 12768 6984 12774 6996
rect 13722 6984 13728 6996
rect 12768 6956 13728 6984
rect 12768 6944 12774 6956
rect 13722 6944 13728 6956
rect 13780 6984 13786 6996
rect 15565 6987 15623 6993
rect 13780 6956 13952 6984
rect 13780 6944 13786 6956
rect 8757 6919 8815 6925
rect 8757 6885 8769 6919
rect 8803 6916 8815 6919
rect 8846 6916 8852 6928
rect 8803 6888 8852 6916
rect 8803 6885 8815 6888
rect 8757 6879 8815 6885
rect 8846 6876 8852 6888
rect 8904 6876 8910 6928
rect 10873 6919 10931 6925
rect 10873 6885 10885 6919
rect 10919 6916 10931 6919
rect 11882 6916 11888 6928
rect 10919 6888 11888 6916
rect 10919 6885 10931 6888
rect 10873 6879 10931 6885
rect 11882 6876 11888 6888
rect 11940 6876 11946 6928
rect 12989 6919 13047 6925
rect 12989 6885 13001 6919
rect 13035 6916 13047 6919
rect 13354 6916 13360 6928
rect 13035 6888 13360 6916
rect 13035 6885 13047 6888
rect 12989 6879 13047 6885
rect 13354 6876 13360 6888
rect 13412 6876 13418 6928
rect 2406 6848 2412 6860
rect 2367 6820 2412 6848
rect 2406 6808 2412 6820
rect 2464 6808 2470 6860
rect 2498 6808 2504 6860
rect 2556 6848 2562 6860
rect 2869 6851 2927 6857
rect 2869 6848 2881 6851
rect 2556 6820 2881 6848
rect 2556 6808 2562 6820
rect 2869 6817 2881 6820
rect 2915 6817 2927 6851
rect 8202 6848 8208 6860
rect 8163 6820 8208 6848
rect 2869 6811 2927 6817
rect 8202 6808 8208 6820
rect 8260 6808 8266 6860
rect 8386 6848 8392 6860
rect 8347 6820 8392 6848
rect 8386 6808 8392 6820
rect 8444 6808 8450 6860
rect 10134 6848 10140 6860
rect 10095 6820 10140 6848
rect 10134 6808 10140 6820
rect 10192 6808 10198 6860
rect 10413 6851 10471 6857
rect 10413 6817 10425 6851
rect 10459 6848 10471 6851
rect 10778 6848 10784 6860
rect 10459 6820 10784 6848
rect 10459 6817 10471 6820
rect 10413 6811 10471 6817
rect 10778 6808 10784 6820
rect 10836 6808 10842 6860
rect 3145 6783 3203 6789
rect 3145 6749 3157 6783
rect 3191 6780 3203 6783
rect 4065 6783 4123 6789
rect 4065 6780 4077 6783
rect 3191 6752 4077 6780
rect 3191 6749 3203 6752
rect 3145 6743 3203 6749
rect 4065 6749 4077 6752
rect 4111 6780 4123 6783
rect 5718 6780 5724 6792
rect 4111 6752 5724 6780
rect 4111 6749 4123 6752
rect 4065 6743 4123 6749
rect 5718 6740 5724 6752
rect 5776 6740 5782 6792
rect 6086 6740 6092 6792
rect 6144 6780 6150 6792
rect 6457 6783 6515 6789
rect 6457 6780 6469 6783
rect 6144 6752 6469 6780
rect 6144 6740 6150 6752
rect 6457 6749 6469 6752
rect 6503 6749 6515 6783
rect 6457 6743 6515 6749
rect 12158 6740 12164 6792
rect 12216 6780 12222 6792
rect 12897 6783 12955 6789
rect 12897 6780 12909 6783
rect 12216 6752 12909 6780
rect 12216 6740 12222 6752
rect 12897 6749 12909 6752
rect 12943 6749 12955 6783
rect 12897 6743 12955 6749
rect 13541 6783 13599 6789
rect 13541 6749 13553 6783
rect 13587 6780 13599 6783
rect 13630 6780 13636 6792
rect 13587 6752 13636 6780
rect 13587 6749 13599 6752
rect 13541 6743 13599 6749
rect 13630 6740 13636 6752
rect 13688 6780 13694 6792
rect 13814 6780 13820 6792
rect 13688 6752 13820 6780
rect 13688 6740 13694 6752
rect 13814 6740 13820 6752
rect 13872 6740 13878 6792
rect 5442 6672 5448 6724
rect 5500 6712 5506 6724
rect 10229 6715 10287 6721
rect 10229 6712 10241 6715
rect 5500 6684 10241 6712
rect 5500 6672 5506 6684
rect 10229 6681 10241 6684
rect 10275 6712 10287 6715
rect 10410 6712 10416 6724
rect 10275 6684 10416 6712
rect 10275 6681 10287 6684
rect 10229 6675 10287 6681
rect 10410 6672 10416 6684
rect 10468 6672 10474 6724
rect 13924 6721 13952 6956
rect 15565 6953 15577 6987
rect 15611 6984 15623 6987
rect 16482 6984 16488 6996
rect 15611 6956 16488 6984
rect 15611 6953 15623 6956
rect 15565 6947 15623 6953
rect 16482 6944 16488 6956
rect 16540 6944 16546 6996
rect 21085 6987 21143 6993
rect 21085 6953 21097 6987
rect 21131 6984 21143 6987
rect 21358 6984 21364 6996
rect 21131 6956 21364 6984
rect 21131 6953 21143 6956
rect 21085 6947 21143 6953
rect 21358 6944 21364 6956
rect 21416 6944 21422 6996
rect 16298 6876 16304 6928
rect 16356 6916 16362 6928
rect 16577 6919 16635 6925
rect 16577 6916 16589 6919
rect 16356 6888 16589 6916
rect 16356 6876 16362 6888
rect 16577 6885 16589 6888
rect 16623 6916 16635 6919
rect 17402 6916 17408 6928
rect 16623 6888 17408 6916
rect 16623 6885 16635 6888
rect 16577 6879 16635 6885
rect 17402 6876 17408 6888
rect 17460 6916 17466 6928
rect 18506 6916 18512 6928
rect 17460 6888 18512 6916
rect 17460 6876 17466 6888
rect 18506 6876 18512 6888
rect 18564 6916 18570 6928
rect 18601 6919 18659 6925
rect 18601 6916 18613 6919
rect 18564 6888 18613 6916
rect 18564 6876 18570 6888
rect 18601 6885 18613 6888
rect 18647 6885 18659 6919
rect 18601 6879 18659 6885
rect 15724 6851 15782 6857
rect 15724 6817 15736 6851
rect 15770 6848 15782 6851
rect 15930 6848 15936 6860
rect 15770 6820 15936 6848
rect 15770 6817 15782 6820
rect 15724 6811 15782 6817
rect 15930 6808 15936 6820
rect 15988 6808 15994 6860
rect 16736 6851 16794 6857
rect 16736 6817 16748 6851
rect 16782 6848 16794 6851
rect 17126 6848 17132 6860
rect 16782 6820 17132 6848
rect 16782 6817 16794 6820
rect 16736 6811 16794 6817
rect 17126 6808 17132 6820
rect 17184 6808 17190 6860
rect 20438 6808 20444 6860
rect 20496 6848 20502 6860
rect 20901 6851 20959 6857
rect 20901 6848 20913 6851
rect 20496 6820 20913 6848
rect 20496 6808 20502 6820
rect 20901 6817 20913 6820
rect 20947 6817 20959 6851
rect 20901 6811 20959 6817
rect 18509 6783 18567 6789
rect 18509 6749 18521 6783
rect 18555 6780 18567 6783
rect 18598 6780 18604 6792
rect 18555 6752 18604 6780
rect 18555 6749 18567 6752
rect 18509 6743 18567 6749
rect 18598 6740 18604 6752
rect 18656 6740 18662 6792
rect 18690 6740 18696 6792
rect 18748 6780 18754 6792
rect 18785 6783 18843 6789
rect 18785 6780 18797 6783
rect 18748 6752 18797 6780
rect 18748 6740 18754 6752
rect 18785 6749 18797 6752
rect 18831 6749 18843 6783
rect 18785 6743 18843 6749
rect 13909 6715 13967 6721
rect 13909 6681 13921 6715
rect 13955 6712 13967 6715
rect 18325 6715 18383 6721
rect 13955 6684 16252 6712
rect 13955 6681 13967 6684
rect 13909 6675 13967 6681
rect 2958 6604 2964 6656
rect 3016 6644 3022 6656
rect 3421 6647 3479 6653
rect 3421 6644 3433 6647
rect 3016 6616 3433 6644
rect 3016 6604 3022 6616
rect 3421 6613 3433 6616
rect 3467 6613 3479 6647
rect 7374 6644 7380 6656
rect 7335 6616 7380 6644
rect 3421 6607 3479 6613
rect 7374 6604 7380 6616
rect 7432 6604 7438 6656
rect 9306 6644 9312 6656
rect 9267 6616 9312 6644
rect 9306 6604 9312 6616
rect 9364 6604 9370 6656
rect 14550 6644 14556 6656
rect 14511 6616 14556 6644
rect 14550 6604 14556 6616
rect 14608 6604 14614 6656
rect 15795 6647 15853 6653
rect 15795 6613 15807 6647
rect 15841 6644 15853 6647
rect 16022 6644 16028 6656
rect 15841 6616 16028 6644
rect 15841 6613 15853 6616
rect 15795 6607 15853 6613
rect 16022 6604 16028 6616
rect 16080 6604 16086 6656
rect 16224 6653 16252 6684
rect 18325 6681 18337 6715
rect 18371 6712 18383 6715
rect 18708 6712 18736 6740
rect 18371 6684 18736 6712
rect 18371 6681 18383 6684
rect 18325 6675 18383 6681
rect 16209 6647 16267 6653
rect 16209 6613 16221 6647
rect 16255 6644 16267 6647
rect 16482 6644 16488 6656
rect 16255 6616 16488 6644
rect 16255 6613 16267 6616
rect 16209 6607 16267 6613
rect 16482 6604 16488 6616
rect 16540 6604 16546 6656
rect 16666 6604 16672 6656
rect 16724 6644 16730 6656
rect 16807 6647 16865 6653
rect 16807 6644 16819 6647
rect 16724 6616 16819 6644
rect 16724 6604 16730 6616
rect 16807 6613 16819 6616
rect 16853 6613 16865 6647
rect 16807 6607 16865 6613
rect 19334 6604 19340 6656
rect 19392 6644 19398 6656
rect 19429 6647 19487 6653
rect 19429 6644 19441 6647
rect 19392 6616 19441 6644
rect 19392 6604 19398 6616
rect 19429 6613 19441 6616
rect 19475 6613 19487 6647
rect 19429 6607 19487 6613
rect 1104 6554 22816 6576
rect 1104 6502 4982 6554
rect 5034 6502 5046 6554
rect 5098 6502 5110 6554
rect 5162 6502 5174 6554
rect 5226 6502 12982 6554
rect 13034 6502 13046 6554
rect 13098 6502 13110 6554
rect 13162 6502 13174 6554
rect 13226 6502 20982 6554
rect 21034 6502 21046 6554
rect 21098 6502 21110 6554
rect 21162 6502 21174 6554
rect 21226 6502 22816 6554
rect 1104 6480 22816 6502
rect 4614 6440 4620 6452
rect 4575 6412 4620 6440
rect 4614 6400 4620 6412
rect 4672 6400 4678 6452
rect 5718 6440 5724 6452
rect 5679 6412 5724 6440
rect 5718 6400 5724 6412
rect 5776 6400 5782 6452
rect 6549 6443 6607 6449
rect 6549 6409 6561 6443
rect 6595 6440 6607 6443
rect 7098 6440 7104 6452
rect 6595 6412 7104 6440
rect 6595 6409 6607 6412
rect 6549 6403 6607 6409
rect 7098 6400 7104 6412
rect 7156 6400 7162 6452
rect 7374 6440 7380 6452
rect 7335 6412 7380 6440
rect 7374 6400 7380 6412
rect 7432 6400 7438 6452
rect 8202 6400 8208 6452
rect 8260 6440 8266 6452
rect 8573 6443 8631 6449
rect 8573 6440 8585 6443
rect 8260 6412 8585 6440
rect 8260 6400 8266 6412
rect 8573 6409 8585 6412
rect 8619 6440 8631 6443
rect 9950 6440 9956 6452
rect 8619 6412 9956 6440
rect 8619 6409 8631 6412
rect 8573 6403 8631 6409
rect 9950 6400 9956 6412
rect 10008 6400 10014 6452
rect 10410 6440 10416 6452
rect 10371 6412 10416 6440
rect 10410 6400 10416 6412
rect 10468 6400 10474 6452
rect 11330 6400 11336 6452
rect 11388 6440 11394 6452
rect 12158 6440 12164 6452
rect 11388 6412 12164 6440
rect 11388 6400 11394 6412
rect 12158 6400 12164 6412
rect 12216 6400 12222 6452
rect 13354 6400 13360 6452
rect 13412 6440 13418 6452
rect 14461 6443 14519 6449
rect 14461 6440 14473 6443
rect 13412 6412 14473 6440
rect 13412 6400 13418 6412
rect 14461 6409 14473 6412
rect 14507 6409 14519 6443
rect 14461 6403 14519 6409
rect 16758 6400 16764 6452
rect 16816 6440 16822 6452
rect 17126 6440 17132 6452
rect 16816 6412 17132 6440
rect 16816 6400 16822 6412
rect 17126 6400 17132 6412
rect 17184 6400 17190 6452
rect 18598 6400 18604 6452
rect 18656 6440 18662 6452
rect 18877 6443 18935 6449
rect 18877 6440 18889 6443
rect 18656 6412 18889 6440
rect 18656 6400 18662 6412
rect 18877 6409 18889 6412
rect 18923 6409 18935 6443
rect 18877 6403 18935 6409
rect 20622 6400 20628 6452
rect 20680 6440 20686 6452
rect 21453 6443 21511 6449
rect 21453 6440 21465 6443
rect 20680 6412 21465 6440
rect 20680 6400 20686 6412
rect 21453 6409 21465 6412
rect 21499 6409 21511 6443
rect 21453 6403 21511 6409
rect 658 6332 664 6384
rect 716 6372 722 6384
rect 9217 6375 9275 6381
rect 9217 6372 9229 6375
rect 716 6344 9229 6372
rect 716 6332 722 6344
rect 9217 6341 9229 6344
rect 9263 6372 9275 6375
rect 9306 6372 9312 6384
rect 9263 6344 9312 6372
rect 9263 6341 9275 6344
rect 9217 6335 9275 6341
rect 9306 6332 9312 6344
rect 9364 6372 9370 6384
rect 12575 6375 12633 6381
rect 9364 6344 9536 6372
rect 9364 6332 9370 6344
rect 1535 6307 1593 6313
rect 1535 6273 1547 6307
rect 1581 6304 1593 6307
rect 2958 6304 2964 6316
rect 1581 6276 2964 6304
rect 1581 6273 1593 6276
rect 1535 6267 1593 6273
rect 2958 6264 2964 6276
rect 3016 6264 3022 6316
rect 3605 6307 3663 6313
rect 3605 6273 3617 6307
rect 3651 6304 3663 6307
rect 7561 6307 7619 6313
rect 3651 6276 5488 6304
rect 3651 6273 3663 6276
rect 3605 6267 3663 6273
rect 1448 6239 1506 6245
rect 1448 6205 1460 6239
rect 1494 6236 1506 6239
rect 1854 6236 1860 6248
rect 1494 6208 1860 6236
rect 1494 6205 1506 6208
rect 1448 6199 1506 6205
rect 1854 6196 1860 6208
rect 1912 6196 1918 6248
rect 3050 6128 3056 6180
rect 3108 6168 3114 6180
rect 3108 6140 3153 6168
rect 3108 6128 3114 6140
rect 3234 6128 3240 6180
rect 3292 6168 3298 6180
rect 4798 6168 4804 6180
rect 3292 6140 4804 6168
rect 3292 6128 3298 6140
rect 4798 6128 4804 6140
rect 4856 6128 4862 6180
rect 5460 6177 5488 6276
rect 7561 6273 7573 6307
rect 7607 6304 7619 6307
rect 7650 6304 7656 6316
rect 7607 6276 7656 6304
rect 7607 6273 7619 6276
rect 7561 6267 7619 6273
rect 7650 6264 7656 6276
rect 7708 6264 7714 6316
rect 8386 6264 8392 6316
rect 8444 6304 8450 6316
rect 8941 6307 8999 6313
rect 8941 6304 8953 6307
rect 8444 6276 8953 6304
rect 8444 6264 8450 6276
rect 8941 6273 8953 6276
rect 8987 6304 8999 6307
rect 9401 6307 9459 6313
rect 9401 6304 9413 6307
rect 8987 6276 9413 6304
rect 8987 6273 8999 6276
rect 8941 6267 8999 6273
rect 9401 6273 9413 6276
rect 9447 6273 9459 6307
rect 9401 6267 9459 6273
rect 9508 6245 9536 6344
rect 12575 6341 12587 6375
rect 12621 6372 12633 6375
rect 14550 6372 14556 6384
rect 12621 6344 14556 6372
rect 12621 6341 12633 6344
rect 12575 6335 12633 6341
rect 14550 6332 14556 6344
rect 14608 6332 14614 6384
rect 10042 6264 10048 6316
rect 10100 6304 10106 6316
rect 12989 6307 13047 6313
rect 12989 6304 13001 6307
rect 10100 6276 11652 6304
rect 10100 6264 10106 6276
rect 9493 6239 9551 6245
rect 9493 6205 9505 6239
rect 9539 6205 9551 6239
rect 11000 6239 11058 6245
rect 11000 6236 11012 6239
rect 9493 6199 9551 6205
rect 10704 6208 11012 6236
rect 4893 6171 4951 6177
rect 4893 6137 4905 6171
rect 4939 6137 4951 6171
rect 4893 6131 4951 6137
rect 5445 6171 5503 6177
rect 5445 6137 5457 6171
rect 5491 6168 5503 6171
rect 6730 6168 6736 6180
rect 5491 6140 6736 6168
rect 5491 6137 5503 6140
rect 5445 6131 5503 6137
rect 2498 6100 2504 6112
rect 2459 6072 2504 6100
rect 2498 6060 2504 6072
rect 2556 6060 2562 6112
rect 4062 6100 4068 6112
rect 4023 6072 4068 6100
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 4614 6060 4620 6112
rect 4672 6100 4678 6112
rect 4908 6100 4936 6131
rect 6730 6128 6736 6140
rect 6788 6128 6794 6180
rect 7653 6171 7711 6177
rect 7653 6137 7665 6171
rect 7699 6137 7711 6171
rect 7653 6131 7711 6137
rect 8205 6171 8263 6177
rect 8205 6137 8217 6171
rect 8251 6168 8263 6171
rect 8386 6168 8392 6180
rect 8251 6140 8392 6168
rect 8251 6137 8263 6140
rect 8205 6131 8263 6137
rect 6086 6100 6092 6112
rect 4672 6072 4936 6100
rect 6047 6072 6092 6100
rect 4672 6060 4678 6072
rect 6086 6060 6092 6072
rect 6144 6060 6150 6112
rect 7374 6060 7380 6112
rect 7432 6100 7438 6112
rect 7668 6100 7696 6131
rect 8386 6128 8392 6140
rect 8444 6128 8450 6180
rect 8754 6128 8760 6180
rect 8812 6168 8818 6180
rect 10704 6168 10732 6208
rect 11000 6205 11012 6208
rect 11046 6236 11058 6239
rect 11425 6239 11483 6245
rect 11425 6236 11437 6239
rect 11046 6208 11437 6236
rect 11046 6205 11058 6208
rect 11000 6199 11058 6205
rect 11425 6205 11437 6208
rect 11471 6205 11483 6239
rect 11425 6199 11483 6205
rect 8812 6140 10732 6168
rect 8812 6128 8818 6140
rect 9508 6112 9536 6140
rect 10778 6128 10784 6180
rect 10836 6168 10842 6180
rect 10873 6171 10931 6177
rect 10873 6168 10885 6171
rect 10836 6140 10885 6168
rect 10836 6128 10842 6140
rect 10873 6137 10885 6140
rect 10919 6168 10931 6171
rect 11514 6168 11520 6180
rect 10919 6140 11520 6168
rect 10919 6137 10931 6140
rect 10873 6131 10931 6137
rect 11514 6128 11520 6140
rect 11572 6128 11578 6180
rect 11624 6168 11652 6276
rect 12519 6276 13001 6304
rect 12519 6245 12547 6276
rect 12989 6273 13001 6276
rect 13035 6304 13047 6307
rect 15286 6304 15292 6316
rect 13035 6276 15292 6304
rect 13035 6273 13047 6276
rect 12989 6267 13047 6273
rect 15286 6264 15292 6276
rect 15344 6264 15350 6316
rect 17972 6276 18368 6304
rect 12504 6239 12562 6245
rect 12504 6205 12516 6239
rect 12550 6205 12562 6239
rect 13262 6236 13268 6248
rect 13223 6208 13268 6236
rect 12504 6199 12562 6205
rect 13262 6196 13268 6208
rect 13320 6236 13326 6248
rect 13449 6239 13507 6245
rect 13449 6236 13461 6239
rect 13320 6208 13461 6236
rect 13320 6196 13326 6208
rect 13449 6205 13461 6208
rect 13495 6205 13507 6239
rect 13449 6199 13507 6205
rect 13722 6196 13728 6248
rect 13780 6236 13786 6248
rect 13909 6239 13967 6245
rect 13909 6236 13921 6239
rect 13780 6208 13921 6236
rect 13780 6196 13786 6208
rect 13909 6205 13921 6208
rect 13955 6205 13967 6239
rect 13909 6199 13967 6205
rect 14826 6196 14832 6248
rect 14884 6236 14890 6248
rect 15048 6239 15106 6245
rect 15048 6236 15060 6239
rect 14884 6208 15060 6236
rect 14884 6196 14890 6208
rect 15048 6205 15060 6208
rect 15094 6236 15106 6239
rect 15473 6239 15531 6245
rect 15473 6236 15485 6239
rect 15094 6208 15485 6236
rect 15094 6205 15106 6208
rect 15048 6199 15106 6205
rect 15473 6205 15485 6208
rect 15519 6205 15531 6239
rect 16114 6236 16120 6248
rect 16075 6208 16120 6236
rect 15473 6199 15531 6205
rect 16114 6196 16120 6208
rect 16172 6196 16178 6248
rect 16482 6196 16488 6248
rect 16540 6236 16546 6248
rect 17972 6245 18000 6276
rect 18340 6248 18368 6276
rect 19242 6264 19248 6316
rect 19300 6304 19306 6316
rect 19429 6307 19487 6313
rect 19429 6304 19441 6307
rect 19300 6276 19441 6304
rect 19300 6264 19306 6276
rect 19429 6273 19441 6276
rect 19475 6273 19487 6307
rect 19429 6267 19487 6273
rect 16577 6239 16635 6245
rect 16577 6236 16589 6239
rect 16540 6208 16589 6236
rect 16540 6196 16546 6208
rect 16577 6205 16589 6208
rect 16623 6205 16635 6239
rect 16577 6199 16635 6205
rect 17957 6239 18015 6245
rect 17957 6205 17969 6239
rect 18003 6205 18015 6239
rect 17957 6199 18015 6205
rect 18322 6196 18328 6248
rect 18380 6236 18386 6248
rect 20640 6245 20668 6400
rect 18509 6239 18567 6245
rect 18509 6236 18521 6239
rect 18380 6208 18521 6236
rect 18380 6196 18386 6208
rect 18509 6205 18521 6208
rect 18555 6205 18567 6239
rect 20640 6239 20718 6245
rect 20640 6208 20672 6239
rect 18509 6199 18567 6205
rect 20660 6205 20672 6208
rect 20706 6205 20718 6239
rect 20660 6199 20718 6205
rect 13280 6168 13308 6196
rect 14182 6168 14188 6180
rect 11624 6140 13308 6168
rect 14143 6140 14188 6168
rect 14182 6128 14188 6140
rect 14240 6128 14246 6180
rect 16850 6168 16856 6180
rect 16811 6140 16856 6168
rect 16850 6128 16856 6140
rect 16908 6128 16914 6180
rect 19153 6171 19211 6177
rect 19153 6137 19165 6171
rect 19199 6137 19211 6171
rect 19153 6131 19211 6137
rect 19245 6171 19303 6177
rect 19245 6137 19257 6171
rect 19291 6168 19303 6171
rect 19334 6168 19340 6180
rect 19291 6140 19340 6168
rect 19291 6137 19303 6140
rect 19245 6131 19303 6137
rect 7432 6072 7696 6100
rect 7432 6060 7438 6072
rect 9490 6060 9496 6112
rect 9548 6060 9554 6112
rect 11103 6103 11161 6109
rect 11103 6069 11115 6103
rect 11149 6100 11161 6103
rect 11238 6100 11244 6112
rect 11149 6072 11244 6100
rect 11149 6069 11161 6072
rect 11103 6063 11161 6069
rect 11238 6060 11244 6072
rect 11296 6060 11302 6112
rect 13814 6060 13820 6112
rect 13872 6100 13878 6112
rect 14458 6100 14464 6112
rect 13872 6072 14464 6100
rect 13872 6060 13878 6072
rect 14458 6060 14464 6072
rect 14516 6060 14522 6112
rect 15102 6060 15108 6112
rect 15160 6100 15166 6112
rect 15289 6103 15347 6109
rect 15289 6100 15301 6103
rect 15160 6072 15301 6100
rect 15160 6060 15166 6072
rect 15289 6069 15301 6072
rect 15335 6069 15347 6103
rect 15930 6100 15936 6112
rect 15891 6072 15936 6100
rect 15289 6063 15347 6069
rect 15930 6060 15936 6072
rect 15988 6060 15994 6112
rect 18187 6103 18245 6109
rect 18187 6069 18199 6103
rect 18233 6100 18245 6103
rect 18414 6100 18420 6112
rect 18233 6072 18420 6100
rect 18233 6069 18245 6072
rect 18187 6063 18245 6069
rect 18414 6060 18420 6072
rect 18472 6060 18478 6112
rect 19168 6100 19196 6131
rect 19334 6128 19340 6140
rect 19392 6128 19398 6180
rect 20438 6128 20444 6180
rect 20496 6168 20502 6180
rect 21085 6171 21143 6177
rect 21085 6168 21097 6171
rect 20496 6140 21097 6168
rect 20496 6128 20502 6140
rect 21085 6137 21097 6140
rect 21131 6137 21143 6171
rect 21085 6131 21143 6137
rect 20165 6103 20223 6109
rect 20165 6100 20177 6103
rect 19168 6072 20177 6100
rect 20165 6069 20177 6072
rect 20211 6100 20223 6103
rect 20763 6103 20821 6109
rect 20763 6100 20775 6103
rect 20211 6072 20775 6100
rect 20211 6069 20223 6072
rect 20165 6063 20223 6069
rect 20763 6069 20775 6072
rect 20809 6069 20821 6103
rect 20763 6063 20821 6069
rect 1104 6010 22816 6032
rect 1104 5958 8982 6010
rect 9034 5958 9046 6010
rect 9098 5958 9110 6010
rect 9162 5958 9174 6010
rect 9226 5958 16982 6010
rect 17034 5958 17046 6010
rect 17098 5958 17110 6010
rect 17162 5958 17174 6010
rect 17226 5958 22816 6010
rect 1104 5936 22816 5958
rect 3050 5856 3056 5908
rect 3108 5896 3114 5908
rect 3421 5899 3479 5905
rect 3421 5896 3433 5899
rect 3108 5868 3433 5896
rect 3108 5856 3114 5868
rect 3421 5865 3433 5868
rect 3467 5896 3479 5899
rect 3510 5896 3516 5908
rect 3467 5868 3516 5896
rect 3467 5865 3479 5868
rect 3421 5859 3479 5865
rect 3510 5856 3516 5868
rect 3568 5856 3574 5908
rect 4154 5856 4160 5908
rect 4212 5896 4218 5908
rect 4212 5868 4257 5896
rect 4212 5856 4218 5868
rect 4798 5856 4804 5908
rect 4856 5896 4862 5908
rect 5537 5899 5595 5905
rect 5537 5896 5549 5899
rect 4856 5868 5549 5896
rect 4856 5856 4862 5868
rect 5537 5865 5549 5868
rect 5583 5865 5595 5899
rect 6086 5896 6092 5908
rect 6047 5868 6092 5896
rect 5537 5859 5595 5865
rect 6086 5856 6092 5868
rect 6144 5856 6150 5908
rect 7650 5896 7656 5908
rect 7611 5868 7656 5896
rect 7650 5856 7656 5868
rect 7708 5856 7714 5908
rect 10134 5856 10140 5908
rect 10192 5896 10198 5908
rect 10781 5899 10839 5905
rect 10781 5896 10793 5899
rect 10192 5868 10793 5896
rect 10192 5856 10198 5868
rect 10781 5865 10793 5868
rect 10827 5865 10839 5899
rect 14182 5896 14188 5908
rect 14143 5868 14188 5896
rect 10781 5859 10839 5865
rect 14182 5856 14188 5868
rect 14240 5856 14246 5908
rect 16022 5856 16028 5908
rect 16080 5896 16086 5908
rect 16669 5899 16727 5905
rect 16669 5896 16681 5899
rect 16080 5868 16681 5896
rect 16080 5856 16086 5868
rect 16669 5865 16681 5868
rect 16715 5865 16727 5899
rect 18506 5896 18512 5908
rect 18467 5868 18512 5896
rect 16669 5859 16727 5865
rect 18506 5856 18512 5868
rect 18564 5856 18570 5908
rect 19334 5856 19340 5908
rect 19392 5856 19398 5908
rect 19426 5856 19432 5908
rect 19484 5896 19490 5908
rect 21039 5899 21097 5905
rect 21039 5896 21051 5899
rect 19484 5868 21051 5896
rect 19484 5856 19490 5868
rect 21039 5865 21051 5868
rect 21085 5865 21097 5899
rect 21039 5859 21097 5865
rect 2498 5788 2504 5840
rect 2556 5828 2562 5840
rect 4246 5828 4252 5840
rect 2556 5800 4252 5828
rect 2556 5788 2562 5800
rect 4246 5788 4252 5800
rect 4304 5828 4310 5840
rect 5261 5831 5319 5837
rect 4304 5800 4660 5828
rect 4304 5788 4310 5800
rect 2866 5720 2872 5772
rect 2924 5760 2930 5772
rect 2996 5763 3054 5769
rect 2996 5760 3008 5763
rect 2924 5732 3008 5760
rect 2924 5720 2930 5732
rect 2996 5729 3008 5732
rect 3042 5729 3054 5763
rect 2996 5723 3054 5729
rect 3099 5763 3157 5769
rect 3099 5729 3111 5763
rect 3145 5760 3157 5763
rect 3234 5760 3240 5772
rect 3145 5732 3240 5760
rect 3145 5729 3157 5732
rect 3099 5723 3157 5729
rect 3234 5720 3240 5732
rect 3292 5720 3298 5772
rect 4341 5763 4399 5769
rect 4341 5729 4353 5763
rect 4387 5760 4399 5763
rect 4430 5760 4436 5772
rect 4387 5732 4436 5760
rect 4387 5729 4399 5732
rect 4341 5723 4399 5729
rect 4430 5720 4436 5732
rect 4488 5720 4494 5772
rect 4632 5769 4660 5800
rect 5261 5797 5273 5831
rect 5307 5828 5319 5831
rect 8202 5828 8208 5840
rect 5307 5800 6224 5828
rect 8163 5800 8208 5828
rect 5307 5797 5319 5800
rect 5261 5791 5319 5797
rect 4617 5763 4675 5769
rect 4617 5729 4629 5763
rect 4663 5760 4675 5763
rect 5276 5760 5304 5791
rect 6196 5772 6224 5800
rect 8202 5788 8208 5800
rect 8260 5788 8266 5840
rect 13081 5831 13139 5837
rect 10336 5800 11928 5828
rect 4663 5732 5304 5760
rect 6089 5763 6147 5769
rect 4663 5729 4675 5732
rect 4617 5723 4675 5729
rect 6089 5729 6101 5763
rect 6135 5729 6147 5763
rect 6089 5723 6147 5729
rect 6104 5692 6132 5723
rect 6178 5720 6184 5772
rect 6236 5760 6242 5772
rect 6273 5763 6331 5769
rect 6273 5760 6285 5763
rect 6236 5732 6285 5760
rect 6236 5720 6242 5732
rect 6273 5729 6285 5732
rect 6319 5729 6331 5763
rect 10042 5760 10048 5772
rect 10003 5732 10048 5760
rect 6273 5723 6331 5729
rect 10042 5720 10048 5732
rect 10100 5720 10106 5772
rect 10134 5720 10140 5772
rect 10192 5760 10198 5772
rect 10336 5769 10364 5800
rect 11900 5772 11928 5800
rect 13081 5797 13093 5831
rect 13127 5828 13139 5831
rect 13354 5828 13360 5840
rect 13127 5800 13360 5828
rect 13127 5797 13139 5800
rect 13081 5791 13139 5797
rect 13354 5788 13360 5800
rect 13412 5788 13418 5840
rect 15470 5828 15476 5840
rect 15431 5800 15476 5828
rect 15470 5788 15476 5800
rect 15528 5788 15534 5840
rect 17215 5831 17273 5837
rect 17215 5797 17227 5831
rect 17261 5828 17273 5831
rect 17402 5828 17408 5840
rect 17261 5800 17408 5828
rect 17261 5797 17273 5800
rect 17215 5791 17273 5797
rect 17402 5788 17408 5800
rect 17460 5788 17466 5840
rect 18877 5831 18935 5837
rect 18877 5828 18889 5831
rect 17788 5800 18889 5828
rect 10321 5763 10379 5769
rect 10321 5760 10333 5763
rect 10192 5732 10333 5760
rect 10192 5720 10198 5732
rect 10321 5729 10333 5732
rect 10367 5729 10379 5763
rect 11333 5763 11391 5769
rect 11333 5760 11345 5763
rect 10321 5723 10379 5729
rect 11164 5732 11345 5760
rect 6638 5692 6644 5704
rect 6104 5664 6644 5692
rect 6638 5652 6644 5664
rect 6696 5652 6702 5704
rect 6730 5652 6736 5704
rect 6788 5692 6794 5704
rect 8110 5692 8116 5704
rect 6788 5664 8116 5692
rect 6788 5652 6794 5664
rect 8110 5652 8116 5664
rect 8168 5652 8174 5704
rect 8386 5692 8392 5704
rect 8347 5664 8392 5692
rect 8386 5652 8392 5664
rect 8444 5652 8450 5704
rect 10410 5692 10416 5704
rect 10371 5664 10416 5692
rect 10410 5652 10416 5664
rect 10468 5652 10474 5704
rect 5442 5584 5448 5636
rect 5500 5624 5506 5636
rect 10870 5624 10876 5636
rect 5500 5596 10876 5624
rect 5500 5584 5506 5596
rect 10870 5584 10876 5596
rect 10928 5584 10934 5636
rect 11164 5624 11192 5732
rect 11333 5729 11345 5732
rect 11379 5729 11391 5763
rect 11882 5760 11888 5772
rect 11843 5732 11888 5760
rect 11333 5723 11391 5729
rect 11882 5720 11888 5732
rect 11940 5720 11946 5772
rect 16850 5760 16856 5772
rect 16811 5732 16856 5760
rect 16850 5720 16856 5732
rect 16908 5720 16914 5772
rect 12066 5692 12072 5704
rect 12027 5664 12072 5692
rect 12066 5652 12072 5664
rect 12124 5652 12130 5704
rect 12802 5652 12808 5704
rect 12860 5692 12866 5704
rect 12989 5695 13047 5701
rect 12989 5692 13001 5695
rect 12860 5664 13001 5692
rect 12860 5652 12866 5664
rect 12989 5661 13001 5664
rect 13035 5661 13047 5695
rect 13262 5692 13268 5704
rect 13223 5664 13268 5692
rect 12989 5655 13047 5661
rect 13262 5652 13268 5664
rect 13320 5652 13326 5704
rect 15102 5652 15108 5704
rect 15160 5692 15166 5704
rect 15381 5695 15439 5701
rect 15381 5692 15393 5695
rect 15160 5664 15393 5692
rect 15160 5652 15166 5664
rect 15381 5661 15393 5664
rect 15427 5661 15439 5695
rect 15381 5655 15439 5661
rect 16025 5695 16083 5701
rect 16025 5661 16037 5695
rect 16071 5692 16083 5695
rect 16574 5692 16580 5704
rect 16071 5664 16580 5692
rect 16071 5661 16083 5664
rect 16025 5655 16083 5661
rect 16574 5652 16580 5664
rect 16632 5652 16638 5704
rect 12342 5624 12348 5636
rect 11164 5596 12348 5624
rect 2406 5516 2412 5568
rect 2464 5556 2470 5568
rect 2501 5559 2559 5565
rect 2501 5556 2513 5559
rect 2464 5528 2513 5556
rect 2464 5516 2470 5528
rect 2501 5525 2513 5528
rect 2547 5556 2559 5559
rect 3970 5556 3976 5568
rect 2547 5528 3976 5556
rect 2547 5525 2559 5528
rect 2501 5519 2559 5525
rect 3970 5516 3976 5528
rect 4028 5516 4034 5568
rect 7282 5556 7288 5568
rect 7243 5528 7288 5556
rect 7282 5516 7288 5528
rect 7340 5516 7346 5568
rect 7466 5516 7472 5568
rect 7524 5556 7530 5568
rect 11164 5565 11192 5596
rect 12342 5584 12348 5596
rect 12400 5624 12406 5636
rect 16114 5624 16120 5636
rect 12400 5596 16120 5624
rect 12400 5584 12406 5596
rect 16114 5584 16120 5596
rect 16172 5624 16178 5636
rect 16301 5627 16359 5633
rect 16301 5624 16313 5627
rect 16172 5596 16313 5624
rect 16172 5584 16178 5596
rect 16301 5593 16313 5596
rect 16347 5593 16359 5627
rect 16301 5587 16359 5593
rect 11149 5559 11207 5565
rect 11149 5556 11161 5559
rect 7524 5528 11161 5556
rect 7524 5516 7530 5528
rect 11149 5525 11161 5528
rect 11195 5525 11207 5559
rect 11149 5519 11207 5525
rect 16390 5516 16396 5568
rect 16448 5556 16454 5568
rect 17788 5565 17816 5800
rect 18877 5797 18889 5800
rect 18923 5828 18935 5831
rect 19352 5828 19380 5856
rect 18923 5800 19380 5828
rect 18923 5797 18935 5800
rect 18877 5791 18935 5797
rect 20968 5763 21026 5769
rect 20968 5729 20980 5763
rect 21014 5760 21026 5763
rect 21542 5760 21548 5772
rect 21014 5732 21548 5760
rect 21014 5729 21026 5732
rect 20968 5723 21026 5729
rect 21542 5720 21548 5732
rect 21600 5720 21606 5772
rect 18506 5652 18512 5704
rect 18564 5692 18570 5704
rect 18785 5695 18843 5701
rect 18785 5692 18797 5695
rect 18564 5664 18797 5692
rect 18564 5652 18570 5664
rect 18785 5661 18797 5664
rect 18831 5692 18843 5695
rect 19610 5692 19616 5704
rect 18831 5664 19616 5692
rect 18831 5661 18843 5664
rect 18785 5655 18843 5661
rect 19610 5652 19616 5664
rect 19668 5652 19674 5704
rect 19334 5624 19340 5636
rect 19295 5596 19340 5624
rect 19334 5584 19340 5596
rect 19392 5584 19398 5636
rect 17773 5559 17831 5565
rect 17773 5556 17785 5559
rect 16448 5528 17785 5556
rect 16448 5516 16454 5528
rect 17773 5525 17785 5528
rect 17819 5525 17831 5559
rect 17773 5519 17831 5525
rect 1104 5466 22816 5488
rect 1104 5414 4982 5466
rect 5034 5414 5046 5466
rect 5098 5414 5110 5466
rect 5162 5414 5174 5466
rect 5226 5414 12982 5466
rect 13034 5414 13046 5466
rect 13098 5414 13110 5466
rect 13162 5414 13174 5466
rect 13226 5414 20982 5466
rect 21034 5414 21046 5466
rect 21098 5414 21110 5466
rect 21162 5414 21174 5466
rect 21226 5414 22816 5466
rect 1104 5392 22816 5414
rect 3510 5352 3516 5364
rect 3471 5324 3516 5352
rect 3510 5312 3516 5324
rect 3568 5312 3574 5364
rect 4246 5352 4252 5364
rect 4207 5324 4252 5352
rect 4246 5312 4252 5324
rect 4304 5312 4310 5364
rect 6178 5352 6184 5364
rect 6139 5324 6184 5352
rect 6178 5312 6184 5324
rect 6236 5312 6242 5364
rect 7098 5352 7104 5364
rect 7059 5324 7104 5352
rect 7098 5312 7104 5324
rect 7156 5312 7162 5364
rect 8202 5312 8208 5364
rect 8260 5352 8266 5364
rect 8481 5355 8539 5361
rect 8481 5352 8493 5355
rect 8260 5324 8493 5352
rect 8260 5312 8266 5324
rect 8481 5321 8493 5324
rect 8527 5321 8539 5355
rect 8481 5315 8539 5321
rect 9861 5355 9919 5361
rect 9861 5321 9873 5355
rect 9907 5352 9919 5355
rect 10042 5352 10048 5364
rect 9907 5324 10048 5352
rect 9907 5321 9919 5324
rect 9861 5315 9919 5321
rect 10042 5312 10048 5324
rect 10100 5312 10106 5364
rect 11701 5355 11759 5361
rect 11701 5321 11713 5355
rect 11747 5352 11759 5355
rect 11882 5352 11888 5364
rect 11747 5324 11888 5352
rect 11747 5321 11759 5324
rect 11701 5315 11759 5321
rect 11882 5312 11888 5324
rect 11940 5312 11946 5364
rect 12253 5355 12311 5361
rect 12253 5321 12265 5355
rect 12299 5352 12311 5355
rect 12526 5352 12532 5364
rect 12299 5324 12532 5352
rect 12299 5321 12311 5324
rect 12253 5315 12311 5321
rect 12526 5312 12532 5324
rect 12584 5312 12590 5364
rect 13354 5352 13360 5364
rect 13315 5324 13360 5352
rect 13354 5312 13360 5324
rect 13412 5352 13418 5364
rect 13633 5355 13691 5361
rect 13633 5352 13645 5355
rect 13412 5324 13645 5352
rect 13412 5312 13418 5324
rect 13633 5321 13645 5324
rect 13679 5321 13691 5355
rect 18506 5352 18512 5364
rect 18467 5324 18512 5352
rect 13633 5315 13691 5321
rect 18506 5312 18512 5324
rect 18564 5312 18570 5364
rect 19426 5312 19432 5364
rect 19484 5352 19490 5364
rect 19613 5355 19671 5361
rect 19613 5352 19625 5355
rect 19484 5324 19625 5352
rect 19484 5312 19490 5324
rect 19613 5321 19625 5324
rect 19659 5321 19671 5355
rect 19613 5315 19671 5321
rect 2866 5244 2872 5296
rect 2924 5284 2930 5296
rect 3789 5287 3847 5293
rect 3789 5284 3801 5287
rect 2924 5256 3801 5284
rect 2924 5244 2930 5256
rect 3789 5253 3801 5256
rect 3835 5284 3847 5287
rect 7558 5284 7564 5296
rect 3835 5256 7564 5284
rect 3835 5253 3847 5256
rect 3789 5247 3847 5253
rect 7558 5244 7564 5256
rect 7616 5244 7622 5296
rect 12544 5284 12572 5312
rect 14001 5287 14059 5293
rect 14001 5284 14013 5287
rect 12544 5256 14013 5284
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5216 2191 5219
rect 2593 5219 2651 5225
rect 2593 5216 2605 5219
rect 2179 5188 2605 5216
rect 2179 5185 2191 5188
rect 2133 5179 2191 5185
rect 2593 5185 2605 5188
rect 2639 5216 2651 5219
rect 4154 5216 4160 5228
rect 2639 5188 4160 5216
rect 2639 5185 2651 5188
rect 2593 5179 2651 5185
rect 4154 5176 4160 5188
rect 4212 5176 4218 5228
rect 5905 5219 5963 5225
rect 5905 5185 5917 5219
rect 5951 5216 5963 5219
rect 7282 5216 7288 5228
rect 5951 5188 7288 5216
rect 5951 5185 5963 5188
rect 5905 5179 5963 5185
rect 7282 5176 7288 5188
rect 7340 5176 7346 5228
rect 10410 5216 10416 5228
rect 7662 5188 9674 5216
rect 10371 5188 10416 5216
rect 5077 5151 5135 5157
rect 5077 5117 5089 5151
rect 5123 5148 5135 5151
rect 5445 5151 5503 5157
rect 5445 5148 5457 5151
rect 5123 5120 5457 5148
rect 5123 5117 5135 5120
rect 5077 5111 5135 5117
rect 5445 5117 5457 5120
rect 5491 5148 5503 5151
rect 5534 5148 5540 5160
rect 5491 5120 5540 5148
rect 5491 5117 5503 5120
rect 5445 5111 5503 5117
rect 5534 5108 5540 5120
rect 5592 5108 5598 5160
rect 5721 5151 5779 5157
rect 5721 5117 5733 5151
rect 5767 5148 5779 5151
rect 5810 5148 5816 5160
rect 5767 5120 5816 5148
rect 5767 5117 5779 5120
rect 5721 5111 5779 5117
rect 5810 5108 5816 5120
rect 5868 5148 5874 5160
rect 6178 5148 6184 5160
rect 5868 5120 6184 5148
rect 5868 5108 5874 5120
rect 6178 5108 6184 5120
rect 6236 5108 6242 5160
rect 7098 5108 7104 5160
rect 7156 5148 7162 5160
rect 7662 5148 7690 5188
rect 7156 5120 7690 5148
rect 7156 5108 7162 5120
rect 7662 5092 7690 5120
rect 7742 5108 7748 5160
rect 7800 5148 7806 5160
rect 8205 5151 8263 5157
rect 8205 5148 8217 5151
rect 7800 5120 8217 5148
rect 7800 5108 7806 5120
rect 8205 5117 8217 5120
rect 8251 5148 8263 5151
rect 8570 5148 8576 5160
rect 8251 5120 8576 5148
rect 8251 5117 8263 5120
rect 8205 5111 8263 5117
rect 8570 5108 8576 5120
rect 8628 5108 8634 5160
rect 2914 5083 2972 5089
rect 2914 5080 2926 5083
rect 2424 5052 2926 5080
rect 1486 4972 1492 5024
rect 1544 5012 1550 5024
rect 2424 5021 2452 5052
rect 2914 5049 2926 5052
rect 2960 5080 2972 5083
rect 4062 5080 4068 5092
rect 2960 5052 4068 5080
rect 2960 5049 2972 5052
rect 2914 5043 2972 5049
rect 4062 5040 4068 5052
rect 4120 5040 4126 5092
rect 7466 5080 7472 5092
rect 4540 5052 7472 5080
rect 2409 5015 2467 5021
rect 2409 5012 2421 5015
rect 1544 4984 2421 5012
rect 1544 4972 1550 4984
rect 2409 4981 2421 4984
rect 2455 4981 2467 5015
rect 2409 4975 2467 4981
rect 4430 4972 4436 5024
rect 4488 5012 4494 5024
rect 4540 5021 4568 5052
rect 7466 5040 7472 5052
rect 7524 5040 7530 5092
rect 7650 5089 7656 5092
rect 7647 5080 7656 5089
rect 7563 5052 7656 5080
rect 7647 5043 7656 5052
rect 7650 5040 7656 5043
rect 7708 5040 7714 5092
rect 8294 5040 8300 5092
rect 8352 5080 8358 5092
rect 9033 5083 9091 5089
rect 9033 5080 9045 5083
rect 8352 5052 9045 5080
rect 8352 5040 8358 5052
rect 9033 5049 9045 5052
rect 9079 5049 9091 5083
rect 9646 5080 9674 5188
rect 10410 5176 10416 5188
rect 10468 5176 10474 5228
rect 12066 5176 12072 5228
rect 12124 5216 12130 5228
rect 12434 5216 12440 5228
rect 12124 5188 12440 5216
rect 12124 5176 12130 5188
rect 12434 5176 12440 5188
rect 12492 5176 12498 5228
rect 10321 5083 10379 5089
rect 10321 5080 10333 5083
rect 9646 5052 10333 5080
rect 9033 5043 9091 5049
rect 10321 5049 10333 5052
rect 10367 5080 10379 5083
rect 10502 5080 10508 5092
rect 10367 5052 10508 5080
rect 10367 5049 10379 5052
rect 10321 5043 10379 5049
rect 10502 5040 10508 5052
rect 10560 5080 10566 5092
rect 12773 5089 12801 5256
rect 14001 5253 14013 5256
rect 14047 5253 14059 5287
rect 19242 5284 19248 5296
rect 19203 5256 19248 5284
rect 14001 5247 14059 5253
rect 10775 5083 10833 5089
rect 10775 5080 10787 5083
rect 10560 5052 10787 5080
rect 10560 5040 10566 5052
rect 10775 5049 10787 5052
rect 10821 5080 10833 5083
rect 12758 5083 12816 5089
rect 12758 5080 12770 5083
rect 10821 5052 12770 5080
rect 10821 5049 10833 5052
rect 10775 5043 10833 5049
rect 12758 5049 12770 5052
rect 12804 5049 12816 5083
rect 14016 5080 14044 5247
rect 19242 5244 19248 5256
rect 19300 5244 19306 5296
rect 14182 5216 14188 5228
rect 14143 5188 14188 5216
rect 14182 5176 14188 5188
rect 14240 5176 14246 5228
rect 16022 5176 16028 5228
rect 16080 5216 16086 5228
rect 16301 5219 16359 5225
rect 16301 5216 16313 5219
rect 16080 5188 16313 5216
rect 16080 5176 16086 5188
rect 16301 5185 16313 5188
rect 16347 5185 16359 5219
rect 16574 5216 16580 5228
rect 16535 5188 16580 5216
rect 16301 5179 16359 5185
rect 16574 5176 16580 5188
rect 16632 5176 16638 5228
rect 18414 5176 18420 5228
rect 18472 5216 18478 5228
rect 18693 5219 18751 5225
rect 18693 5216 18705 5219
rect 18472 5188 18705 5216
rect 18472 5176 18478 5188
rect 18693 5185 18705 5188
rect 18739 5216 18751 5219
rect 19981 5219 20039 5225
rect 19981 5216 19993 5219
rect 18739 5188 19993 5216
rect 18739 5185 18751 5188
rect 18693 5179 18751 5185
rect 19981 5185 19993 5188
rect 20027 5185 20039 5219
rect 20438 5216 20444 5228
rect 19981 5179 20039 5185
rect 20247 5188 20444 5216
rect 20247 5157 20275 5188
rect 20438 5176 20444 5188
rect 20496 5216 20502 5228
rect 20622 5216 20628 5228
rect 20496 5188 20628 5216
rect 20496 5176 20502 5188
rect 20622 5176 20628 5188
rect 20680 5176 20686 5228
rect 20216 5151 20275 5157
rect 20216 5117 20228 5151
rect 20262 5120 20275 5151
rect 20262 5117 20274 5120
rect 20216 5111 20274 5117
rect 20530 5108 20536 5160
rect 20588 5148 20594 5160
rect 21212 5151 21270 5157
rect 21212 5148 21224 5151
rect 20588 5120 21224 5148
rect 20588 5108 20594 5120
rect 21212 5117 21224 5120
rect 21258 5148 21270 5151
rect 21637 5151 21695 5157
rect 21637 5148 21649 5151
rect 21258 5120 21649 5148
rect 21258 5117 21270 5120
rect 21212 5111 21270 5117
rect 21637 5117 21649 5120
rect 21683 5117 21695 5151
rect 21637 5111 21695 5117
rect 14506 5083 14564 5089
rect 14506 5080 14518 5083
rect 14016 5052 14518 5080
rect 12758 5043 12816 5049
rect 14506 5049 14518 5052
rect 14552 5049 14564 5083
rect 14506 5043 14564 5049
rect 16117 5083 16175 5089
rect 16117 5049 16129 5083
rect 16163 5080 16175 5083
rect 16390 5080 16396 5092
rect 16163 5052 16396 5080
rect 16163 5049 16175 5052
rect 16117 5043 16175 5049
rect 16390 5040 16396 5052
rect 16448 5040 16454 5092
rect 17865 5083 17923 5089
rect 17865 5080 17877 5083
rect 17144 5052 17877 5080
rect 4525 5015 4583 5021
rect 4525 5012 4537 5015
rect 4488 4984 4537 5012
rect 4488 4972 4494 4984
rect 4525 4981 4537 4984
rect 4571 4981 4583 5015
rect 6638 5012 6644 5024
rect 6599 4984 6644 5012
rect 4525 4975 4583 4981
rect 6638 4972 6644 4984
rect 6696 4972 6702 5024
rect 8846 5012 8852 5024
rect 8807 4984 8852 5012
rect 8846 4972 8852 4984
rect 8904 4972 8910 5024
rect 11330 5012 11336 5024
rect 11291 4984 11336 5012
rect 11330 4972 11336 4984
rect 11388 4972 11394 5024
rect 15105 5015 15163 5021
rect 15105 4981 15117 5015
rect 15151 5012 15163 5015
rect 15470 5012 15476 5024
rect 15151 4984 15476 5012
rect 15151 4981 15163 4984
rect 15105 4975 15163 4981
rect 15470 4972 15476 4984
rect 15528 5012 15534 5024
rect 17144 5012 17172 5052
rect 17865 5049 17877 5052
rect 17911 5080 17923 5083
rect 18782 5080 18788 5092
rect 17911 5052 18788 5080
rect 17911 5049 17923 5052
rect 17865 5043 17923 5049
rect 18782 5040 18788 5052
rect 18840 5040 18846 5092
rect 19886 5040 19892 5092
rect 19944 5080 19950 5092
rect 20303 5083 20361 5089
rect 20303 5080 20315 5083
rect 19944 5052 20315 5080
rect 19944 5040 19950 5052
rect 20303 5049 20315 5052
rect 20349 5049 20361 5083
rect 20303 5043 20361 5049
rect 20714 5040 20720 5092
rect 20772 5080 20778 5092
rect 21315 5083 21373 5089
rect 21315 5080 21327 5083
rect 20772 5052 21327 5080
rect 20772 5040 20778 5052
rect 21315 5049 21327 5052
rect 21361 5049 21373 5083
rect 21315 5043 21373 5049
rect 15528 4984 17172 5012
rect 17313 5015 17371 5021
rect 15528 4972 15534 4984
rect 17313 4981 17325 5015
rect 17359 5012 17371 5015
rect 17402 5012 17408 5024
rect 17359 4984 17408 5012
rect 17359 4981 17371 4984
rect 17313 4975 17371 4981
rect 17402 4972 17408 4984
rect 17460 4972 17466 5024
rect 21085 5015 21143 5021
rect 21085 4981 21097 5015
rect 21131 5012 21143 5015
rect 21542 5012 21548 5024
rect 21131 4984 21548 5012
rect 21131 4981 21143 4984
rect 21085 4975 21143 4981
rect 21542 4972 21548 4984
rect 21600 4972 21606 5024
rect 1104 4922 22816 4944
rect 1104 4870 8982 4922
rect 9034 4870 9046 4922
rect 9098 4870 9110 4922
rect 9162 4870 9174 4922
rect 9226 4870 16982 4922
rect 17034 4870 17046 4922
rect 17098 4870 17110 4922
rect 17162 4870 17174 4922
rect 17226 4870 22816 4922
rect 1104 4848 22816 4870
rect 3418 4808 3424 4820
rect 3379 4780 3424 4808
rect 3418 4768 3424 4780
rect 3476 4808 3482 4820
rect 4798 4808 4804 4820
rect 3476 4780 4804 4808
rect 3476 4768 3482 4780
rect 4798 4768 4804 4780
rect 4856 4768 4862 4820
rect 7650 4768 7656 4820
rect 7708 4808 7714 4820
rect 7745 4811 7803 4817
rect 7745 4808 7757 4811
rect 7708 4780 7757 4808
rect 7708 4768 7714 4780
rect 7745 4777 7757 4780
rect 7791 4777 7803 4811
rect 7745 4771 7803 4777
rect 8202 4768 8208 4820
rect 8260 4808 8266 4820
rect 8297 4811 8355 4817
rect 8297 4808 8309 4811
rect 8260 4780 8309 4808
rect 8260 4768 8266 4780
rect 8297 4777 8309 4780
rect 8343 4777 8355 4811
rect 8570 4808 8576 4820
rect 8531 4780 8576 4808
rect 8297 4771 8355 4777
rect 8570 4768 8576 4780
rect 8628 4768 8634 4820
rect 10410 4768 10416 4820
rect 10468 4808 10474 4820
rect 10689 4811 10747 4817
rect 10689 4808 10701 4811
rect 10468 4780 10701 4808
rect 10468 4768 10474 4780
rect 10689 4777 10701 4780
rect 10735 4777 10747 4811
rect 12434 4808 12440 4820
rect 12395 4780 12440 4808
rect 10689 4771 10747 4777
rect 12434 4768 12440 4780
rect 12492 4768 12498 4820
rect 12802 4768 12808 4820
rect 12860 4808 12866 4820
rect 12897 4811 12955 4817
rect 12897 4808 12909 4811
rect 12860 4780 12909 4808
rect 12860 4768 12866 4780
rect 12897 4777 12909 4780
rect 12943 4808 12955 4811
rect 13219 4811 13277 4817
rect 13219 4808 13231 4811
rect 12943 4780 13231 4808
rect 12943 4777 12955 4780
rect 12897 4771 12955 4777
rect 13219 4777 13231 4780
rect 13265 4777 13277 4811
rect 15102 4808 15108 4820
rect 15063 4780 15108 4808
rect 13219 4771 13277 4777
rect 15102 4768 15108 4780
rect 15160 4768 15166 4820
rect 15378 4808 15384 4820
rect 15339 4780 15384 4808
rect 15378 4768 15384 4780
rect 15436 4768 15442 4820
rect 16761 4811 16819 4817
rect 16761 4777 16773 4811
rect 16807 4808 16819 4811
rect 16850 4808 16856 4820
rect 16807 4780 16856 4808
rect 16807 4777 16819 4780
rect 16761 4771 16819 4777
rect 16850 4768 16856 4780
rect 16908 4768 16914 4820
rect 3145 4743 3203 4749
rect 3145 4709 3157 4743
rect 3191 4740 3203 4743
rect 4430 4740 4436 4752
rect 3191 4712 4436 4740
rect 3191 4709 3203 4712
rect 3145 4703 3203 4709
rect 4430 4700 4436 4712
rect 4488 4700 4494 4752
rect 11330 4700 11336 4752
rect 11388 4740 11394 4752
rect 11425 4743 11483 4749
rect 11425 4740 11437 4743
rect 11388 4712 11437 4740
rect 11388 4700 11394 4712
rect 11425 4709 11437 4712
rect 11471 4709 11483 4743
rect 13446 4740 13452 4752
rect 11425 4703 11483 4709
rect 13163 4712 13452 4740
rect 2314 4632 2320 4684
rect 2372 4672 2378 4684
rect 2409 4675 2467 4681
rect 2409 4672 2421 4675
rect 2372 4644 2421 4672
rect 2372 4632 2378 4644
rect 2409 4641 2421 4644
rect 2455 4641 2467 4675
rect 2682 4672 2688 4684
rect 2643 4644 2688 4672
rect 2409 4635 2467 4641
rect 2682 4632 2688 4644
rect 2740 4672 2746 4684
rect 4338 4672 4344 4684
rect 2740 4644 4154 4672
rect 4299 4644 4344 4672
rect 2740 4632 2746 4644
rect 4126 4604 4154 4644
rect 4338 4632 4344 4644
rect 4396 4632 4402 4684
rect 6086 4672 6092 4684
rect 6047 4644 6092 4672
rect 6086 4632 6092 4644
rect 6144 4632 6150 4684
rect 6178 4632 6184 4684
rect 6236 4672 6242 4684
rect 6273 4675 6331 4681
rect 6273 4672 6285 4675
rect 6236 4644 6285 4672
rect 6236 4632 6242 4644
rect 6273 4641 6285 4644
rect 6319 4672 6331 4675
rect 6362 4672 6368 4684
rect 6319 4644 6368 4672
rect 6319 4641 6331 4644
rect 6273 4635 6331 4641
rect 6362 4632 6368 4644
rect 6420 4632 6426 4684
rect 9766 4672 9772 4684
rect 9727 4644 9772 4672
rect 9766 4632 9772 4644
rect 9824 4632 9830 4684
rect 10134 4672 10140 4684
rect 10095 4644 10140 4672
rect 10134 4632 10140 4644
rect 10192 4632 10198 4684
rect 13163 4681 13191 4712
rect 13446 4700 13452 4712
rect 13504 4740 13510 4752
rect 15654 4740 15660 4752
rect 13504 4712 15660 4740
rect 13504 4700 13510 4712
rect 15654 4700 15660 4712
rect 15712 4700 15718 4752
rect 16482 4740 16488 4752
rect 15856 4712 16488 4740
rect 13148 4675 13206 4681
rect 13148 4641 13160 4675
rect 13194 4641 13206 4675
rect 14090 4672 14096 4684
rect 14051 4644 14096 4672
rect 13148 4635 13206 4641
rect 14090 4632 14096 4644
rect 14148 4632 14154 4684
rect 15470 4672 15476 4684
rect 15431 4644 15476 4672
rect 15470 4632 15476 4644
rect 15528 4632 15534 4684
rect 15562 4632 15568 4684
rect 15620 4672 15626 4684
rect 15856 4681 15884 4712
rect 16482 4700 16488 4712
rect 16540 4740 16546 4752
rect 18782 4740 18788 4752
rect 16540 4712 17356 4740
rect 18743 4712 18788 4740
rect 16540 4700 16546 4712
rect 17328 4684 17356 4712
rect 18782 4700 18788 4712
rect 18840 4700 18846 4752
rect 19334 4740 19340 4752
rect 19295 4712 19340 4740
rect 19334 4700 19340 4712
rect 19392 4700 19398 4752
rect 15841 4675 15899 4681
rect 15841 4672 15853 4675
rect 15620 4644 15853 4672
rect 15620 4632 15626 4644
rect 15841 4641 15853 4644
rect 15887 4641 15899 4675
rect 17034 4672 17040 4684
rect 16995 4644 17040 4672
rect 15841 4635 15899 4641
rect 17034 4632 17040 4644
rect 17092 4632 17098 4684
rect 17310 4672 17316 4684
rect 17271 4644 17316 4672
rect 17310 4632 17316 4644
rect 17368 4632 17374 4684
rect 20806 4632 20812 4684
rect 20864 4672 20870 4684
rect 20936 4675 20994 4681
rect 20936 4672 20948 4675
rect 20864 4644 20948 4672
rect 20864 4632 20870 4644
rect 20936 4641 20948 4644
rect 20982 4641 20994 4675
rect 20936 4635 20994 4641
rect 4246 4604 4252 4616
rect 4126 4576 4252 4604
rect 4246 4564 4252 4576
rect 4304 4564 4310 4616
rect 6546 4604 6552 4616
rect 6507 4576 6552 4604
rect 6546 4564 6552 4576
rect 6604 4604 6610 4616
rect 7377 4607 7435 4613
rect 7377 4604 7389 4607
rect 6604 4576 7389 4604
rect 6604 4564 6610 4576
rect 7377 4573 7389 4576
rect 7423 4573 7435 4607
rect 7377 4567 7435 4573
rect 10042 4564 10048 4616
rect 10100 4604 10106 4616
rect 10229 4607 10287 4613
rect 10229 4604 10241 4607
rect 10100 4576 10241 4604
rect 10100 4564 10106 4576
rect 10229 4573 10241 4576
rect 10275 4573 10287 4607
rect 10229 4567 10287 4573
rect 11333 4607 11391 4613
rect 11333 4573 11345 4607
rect 11379 4573 11391 4607
rect 11333 4567 11391 4573
rect 11977 4607 12035 4613
rect 11977 4573 11989 4607
rect 12023 4604 12035 4607
rect 13262 4604 13268 4616
rect 12023 4576 13268 4604
rect 12023 4573 12035 4576
rect 11977 4567 12035 4573
rect 2498 4536 2504 4548
rect 2459 4508 2504 4536
rect 2498 4496 2504 4508
rect 2556 4496 2562 4548
rect 6178 4496 6184 4548
rect 6236 4536 6242 4548
rect 8754 4536 8760 4548
rect 6236 4508 8760 4536
rect 6236 4496 6242 4508
rect 8754 4496 8760 4508
rect 8812 4496 8818 4548
rect 8846 4496 8852 4548
rect 8904 4536 8910 4548
rect 9122 4536 9128 4548
rect 8904 4508 9128 4536
rect 8904 4496 8910 4508
rect 9122 4496 9128 4508
rect 9180 4536 9186 4548
rect 10134 4536 10140 4548
rect 9180 4508 10140 4536
rect 9180 4496 9186 4508
rect 10134 4496 10140 4508
rect 10192 4496 10198 4548
rect 11238 4496 11244 4548
rect 11296 4536 11302 4548
rect 11348 4536 11376 4567
rect 13262 4564 13268 4576
rect 13320 4564 13326 4616
rect 17586 4604 17592 4616
rect 17547 4576 17592 4604
rect 17586 4564 17592 4576
rect 17644 4564 17650 4616
rect 18509 4607 18567 4613
rect 18509 4573 18521 4607
rect 18555 4604 18567 4607
rect 18693 4607 18751 4613
rect 18693 4604 18705 4607
rect 18555 4576 18705 4604
rect 18555 4573 18567 4576
rect 18509 4567 18567 4573
rect 18693 4573 18705 4576
rect 18739 4604 18751 4607
rect 21039 4607 21097 4613
rect 21039 4604 21051 4607
rect 18739 4576 21051 4604
rect 18739 4573 18751 4576
rect 18693 4567 18751 4573
rect 21039 4573 21051 4576
rect 21085 4573 21097 4607
rect 21039 4567 21097 4573
rect 11296 4508 11376 4536
rect 14277 4539 14335 4545
rect 11296 4496 11302 4508
rect 14277 4505 14289 4539
rect 14323 4536 14335 4539
rect 17494 4536 17500 4548
rect 14323 4508 17500 4536
rect 14323 4505 14335 4508
rect 14277 4499 14335 4505
rect 17494 4496 17500 4508
rect 17552 4496 17558 4548
rect 1670 4468 1676 4480
rect 1631 4440 1676 4468
rect 1670 4428 1676 4440
rect 1728 4428 1734 4480
rect 3510 4428 3516 4480
rect 3568 4468 3574 4480
rect 4706 4468 4712 4480
rect 3568 4440 4712 4468
rect 3568 4428 3574 4440
rect 4706 4428 4712 4440
rect 4764 4428 4770 4480
rect 4798 4428 4804 4480
rect 4856 4468 4862 4480
rect 5261 4471 5319 4477
rect 5261 4468 5273 4471
rect 4856 4440 5273 4468
rect 4856 4428 4862 4440
rect 5261 4437 5273 4440
rect 5307 4437 5319 4471
rect 5261 4431 5319 4437
rect 7285 4471 7343 4477
rect 7285 4437 7297 4471
rect 7331 4468 7343 4471
rect 8110 4468 8116 4480
rect 7331 4440 8116 4468
rect 7331 4437 7343 4440
rect 7285 4431 7343 4437
rect 8110 4428 8116 4440
rect 8168 4468 8174 4480
rect 8938 4468 8944 4480
rect 8168 4440 8944 4468
rect 8168 4428 8174 4440
rect 8938 4428 8944 4440
rect 8996 4428 9002 4480
rect 9033 4471 9091 4477
rect 9033 4437 9045 4471
rect 9079 4468 9091 4471
rect 9214 4468 9220 4480
rect 9079 4440 9220 4468
rect 9079 4437 9091 4440
rect 9033 4431 9091 4437
rect 9214 4428 9220 4440
rect 9272 4428 9278 4480
rect 14550 4428 14556 4480
rect 14608 4468 14614 4480
rect 14645 4471 14703 4477
rect 14645 4468 14657 4471
rect 14608 4440 14657 4468
rect 14608 4428 14614 4440
rect 14645 4437 14657 4440
rect 14691 4437 14703 4471
rect 16298 4468 16304 4480
rect 16259 4440 16304 4468
rect 14645 4431 14703 4437
rect 16298 4428 16304 4440
rect 16356 4428 16362 4480
rect 1104 4378 22816 4400
rect 1104 4326 4982 4378
rect 5034 4326 5046 4378
rect 5098 4326 5110 4378
rect 5162 4326 5174 4378
rect 5226 4326 12982 4378
rect 13034 4326 13046 4378
rect 13098 4326 13110 4378
rect 13162 4326 13174 4378
rect 13226 4326 20982 4378
rect 21034 4326 21046 4378
rect 21098 4326 21110 4378
rect 21162 4326 21174 4378
rect 21226 4326 22816 4378
rect 1104 4304 22816 4326
rect 1578 4264 1584 4276
rect 1539 4236 1584 4264
rect 1578 4224 1584 4236
rect 1636 4224 1642 4276
rect 6546 4264 6552 4276
rect 4126 4236 5948 4264
rect 6507 4236 6552 4264
rect 4126 4196 4154 4236
rect 5810 4196 5816 4208
rect 2608 4168 4154 4196
rect 5771 4168 5816 4196
rect 2133 4131 2191 4137
rect 2133 4097 2145 4131
rect 2179 4128 2191 4131
rect 2498 4128 2504 4140
rect 2179 4100 2504 4128
rect 2179 4097 2191 4100
rect 2133 4091 2191 4097
rect 2498 4088 2504 4100
rect 2556 4088 2562 4140
rect 1397 4063 1455 4069
rect 1397 4029 1409 4063
rect 1443 4060 1455 4063
rect 1670 4060 1676 4072
rect 1443 4032 1676 4060
rect 1443 4029 1455 4032
rect 1397 4023 1455 4029
rect 1670 4020 1676 4032
rect 1728 4060 1734 4072
rect 2608 4060 2636 4168
rect 5810 4156 5816 4168
rect 5868 4156 5874 4208
rect 5920 4196 5948 4236
rect 6546 4224 6552 4236
rect 6604 4224 6610 4276
rect 9674 4264 9680 4276
rect 6748 4236 9680 4264
rect 6748 4196 6776 4236
rect 9674 4224 9680 4236
rect 9732 4224 9738 4276
rect 11241 4267 11299 4273
rect 11241 4233 11253 4267
rect 11287 4264 11299 4267
rect 11330 4264 11336 4276
rect 11287 4236 11336 4264
rect 11287 4233 11299 4236
rect 11241 4227 11299 4233
rect 11330 4224 11336 4236
rect 11388 4224 11394 4276
rect 13446 4264 13452 4276
rect 11440 4236 12296 4264
rect 13407 4236 13452 4264
rect 5920 4168 6776 4196
rect 7469 4199 7527 4205
rect 7469 4165 7481 4199
rect 7515 4196 7527 4199
rect 7558 4196 7564 4208
rect 7515 4168 7564 4196
rect 7515 4165 7527 4168
rect 7469 4159 7527 4165
rect 7558 4156 7564 4168
rect 7616 4156 7622 4208
rect 7650 4156 7656 4208
rect 7708 4196 7714 4208
rect 7745 4199 7803 4205
rect 7745 4196 7757 4199
rect 7708 4168 7757 4196
rect 7708 4156 7714 4168
rect 7745 4165 7757 4168
rect 7791 4165 7803 4199
rect 7745 4159 7803 4165
rect 9122 4156 9128 4208
rect 9180 4196 9186 4208
rect 9217 4199 9275 4205
rect 9217 4196 9229 4199
rect 9180 4168 9229 4196
rect 9180 4156 9186 4168
rect 9217 4165 9229 4168
rect 9263 4165 9275 4199
rect 9766 4196 9772 4208
rect 9679 4168 9772 4196
rect 9217 4159 9275 4165
rect 9766 4156 9772 4168
rect 9824 4196 9830 4208
rect 10873 4199 10931 4205
rect 10873 4196 10885 4199
rect 9824 4168 10885 4196
rect 9824 4156 9830 4168
rect 10873 4165 10885 4168
rect 10919 4196 10931 4199
rect 11440 4196 11468 4236
rect 10919 4168 11468 4196
rect 12268 4196 12296 4236
rect 13446 4224 13452 4236
rect 13504 4224 13510 4276
rect 14090 4264 14096 4276
rect 14051 4236 14096 4264
rect 14090 4224 14096 4236
rect 14148 4224 14154 4276
rect 15562 4264 15568 4276
rect 15523 4236 15568 4264
rect 15562 4224 15568 4236
rect 15620 4224 15626 4276
rect 17129 4267 17187 4273
rect 17129 4233 17141 4267
rect 17175 4264 17187 4267
rect 17310 4264 17316 4276
rect 17175 4236 17316 4264
rect 17175 4233 17187 4236
rect 17129 4227 17187 4233
rect 17310 4224 17316 4236
rect 17368 4264 17374 4276
rect 18690 4264 18696 4276
rect 17368 4236 18696 4264
rect 17368 4224 17374 4236
rect 18690 4224 18696 4236
rect 18748 4224 18754 4276
rect 18782 4224 18788 4276
rect 18840 4264 18846 4276
rect 19245 4267 19303 4273
rect 19245 4264 19257 4267
rect 18840 4236 19257 4264
rect 18840 4224 18846 4236
rect 19245 4233 19257 4236
rect 19291 4233 19303 4267
rect 19245 4227 19303 4233
rect 20162 4224 20168 4276
rect 20220 4264 20226 4276
rect 21499 4267 21557 4273
rect 21499 4264 21511 4267
rect 20220 4236 21511 4264
rect 20220 4224 20226 4236
rect 21499 4233 21511 4236
rect 21545 4233 21557 4267
rect 21499 4227 21557 4233
rect 15746 4196 15752 4208
rect 12268 4168 15752 4196
rect 10919 4165 10931 4168
rect 10873 4159 10931 4165
rect 15746 4156 15752 4168
rect 15804 4196 15810 4208
rect 16206 4196 16212 4208
rect 15804 4168 16212 4196
rect 15804 4156 15810 4168
rect 16206 4156 16212 4168
rect 16264 4156 16270 4208
rect 17034 4156 17040 4208
rect 17092 4196 17098 4208
rect 17405 4199 17463 4205
rect 17405 4196 17417 4199
rect 17092 4168 17417 4196
rect 17092 4156 17098 4168
rect 17405 4165 17417 4168
rect 17451 4165 17463 4199
rect 17405 4159 17463 4165
rect 19702 4156 19708 4208
rect 19760 4196 19766 4208
rect 20806 4196 20812 4208
rect 19760 4168 20812 4196
rect 19760 4156 19766 4168
rect 20806 4156 20812 4168
rect 20864 4196 20870 4208
rect 20901 4199 20959 4205
rect 20901 4196 20913 4199
rect 20864 4168 20913 4196
rect 20864 4156 20870 4168
rect 20901 4165 20913 4168
rect 20947 4165 20959 4199
rect 20901 4159 20959 4165
rect 3329 4131 3387 4137
rect 3329 4128 3341 4131
rect 1728 4032 2636 4060
rect 2884 4100 3341 4128
rect 1728 4020 1734 4032
rect 2498 3952 2504 4004
rect 2556 3992 2562 4004
rect 2884 3992 2912 4100
rect 3329 4097 3341 4100
rect 3375 4128 3387 4131
rect 3418 4128 3424 4140
rect 3375 4100 3424 4128
rect 3375 4097 3387 4100
rect 3329 4091 3387 4097
rect 3418 4088 3424 4100
rect 3476 4088 3482 4140
rect 3970 4128 3976 4140
rect 3931 4100 3976 4128
rect 3970 4088 3976 4100
rect 4028 4088 4034 4140
rect 4246 4088 4252 4140
rect 4304 4128 4310 4140
rect 8938 4128 8944 4140
rect 4304 4100 5120 4128
rect 8899 4100 8944 4128
rect 4304 4088 4310 4100
rect 3234 4060 3240 4072
rect 3195 4032 3240 4060
rect 3234 4020 3240 4032
rect 3292 4020 3298 4072
rect 3513 4063 3571 4069
rect 3513 4029 3525 4063
rect 3559 4060 3571 4063
rect 4798 4060 4804 4072
rect 3559 4032 4154 4060
rect 4759 4032 4804 4060
rect 3559 4029 3571 4032
rect 3513 4023 3571 4029
rect 2556 3964 2912 3992
rect 3145 3995 3203 4001
rect 2556 3952 2562 3964
rect 3145 3961 3157 3995
rect 3191 3992 3203 3995
rect 3528 3992 3556 4023
rect 3191 3964 3556 3992
rect 3191 3961 3203 3964
rect 3145 3955 3203 3961
rect 2314 3884 2320 3936
rect 2372 3924 2378 3936
rect 2409 3927 2467 3933
rect 2409 3924 2421 3927
rect 2372 3896 2421 3924
rect 2372 3884 2378 3896
rect 2409 3893 2421 3896
rect 2455 3893 2467 3927
rect 4126 3924 4154 4032
rect 4798 4020 4804 4032
rect 4856 4020 4862 4072
rect 4890 4020 4896 4072
rect 4948 4060 4954 4072
rect 5092 4069 5120 4100
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 9677 4131 9735 4137
rect 9677 4097 9689 4131
rect 9723 4128 9735 4131
rect 10134 4128 10140 4140
rect 9723 4100 10140 4128
rect 9723 4097 9735 4100
rect 9677 4091 9735 4097
rect 10134 4088 10140 4100
rect 10192 4128 10198 4140
rect 16758 4128 16764 4140
rect 10192 4100 10272 4128
rect 10192 4088 10198 4100
rect 5077 4063 5135 4069
rect 4948 4032 4993 4060
rect 4948 4020 4954 4032
rect 5077 4029 5089 4063
rect 5123 4060 5135 4063
rect 5258 4060 5264 4072
rect 5123 4032 5264 4060
rect 5123 4029 5135 4032
rect 5077 4023 5135 4029
rect 5258 4020 5264 4032
rect 5316 4020 5322 4072
rect 6825 4063 6883 4069
rect 6825 4029 6837 4063
rect 6871 4060 6883 4063
rect 7558 4060 7564 4072
rect 6871 4032 7564 4060
rect 6871 4029 6883 4032
rect 6825 4023 6883 4029
rect 7558 4020 7564 4032
rect 7616 4020 7622 4072
rect 10244 4069 10272 4100
rect 12268 4100 12940 4128
rect 16719 4100 16764 4128
rect 9953 4063 10011 4069
rect 9953 4029 9965 4063
rect 9999 4060 10011 4063
rect 10229 4063 10287 4069
rect 9999 4032 10180 4060
rect 9999 4029 10011 4032
rect 9953 4023 10011 4029
rect 4709 3995 4767 4001
rect 4709 3961 4721 3995
rect 4755 3992 4767 3995
rect 4908 3992 4936 4020
rect 10152 4004 10180 4032
rect 10229 4029 10241 4063
rect 10275 4029 10287 4063
rect 10229 4023 10287 4029
rect 10594 4020 10600 4072
rect 10652 4060 10658 4072
rect 11368 4063 11426 4069
rect 11368 4060 11380 4063
rect 10652 4032 11380 4060
rect 10652 4020 10658 4032
rect 11368 4029 11380 4032
rect 11414 4060 11426 4063
rect 11793 4063 11851 4069
rect 11793 4060 11805 4063
rect 11414 4032 11805 4060
rect 11414 4029 11426 4032
rect 11368 4023 11426 4029
rect 11793 4029 11805 4032
rect 11839 4029 11851 4063
rect 11793 4023 11851 4029
rect 11882 4020 11888 4072
rect 11940 4060 11946 4072
rect 12161 4063 12219 4069
rect 12161 4060 12173 4063
rect 11940 4032 12173 4060
rect 11940 4020 11946 4032
rect 12161 4029 12173 4032
rect 12207 4060 12219 4063
rect 12268 4060 12296 4100
rect 12434 4060 12440 4072
rect 12207 4032 12296 4060
rect 12395 4032 12440 4060
rect 12207 4029 12219 4032
rect 12161 4023 12219 4029
rect 12434 4020 12440 4032
rect 12492 4020 12498 4072
rect 12912 4069 12940 4100
rect 16758 4088 16764 4100
rect 16816 4088 16822 4140
rect 17586 4088 17592 4140
rect 17644 4128 17650 4140
rect 18046 4128 18052 4140
rect 17644 4100 18052 4128
rect 17644 4088 17650 4100
rect 18046 4088 18052 4100
rect 18104 4088 18110 4140
rect 18782 4088 18788 4140
rect 18840 4128 18846 4140
rect 19058 4128 19064 4140
rect 18840 4100 19064 4128
rect 18840 4088 18846 4100
rect 19058 4088 19064 4100
rect 19116 4128 19122 4140
rect 20165 4131 20223 4137
rect 20165 4128 20177 4131
rect 19116 4100 20177 4128
rect 19116 4088 19122 4100
rect 20165 4097 20177 4100
rect 20211 4097 20223 4131
rect 20165 4091 20223 4097
rect 12897 4063 12955 4069
rect 12897 4029 12909 4063
rect 12943 4029 12955 4063
rect 12897 4023 12955 4029
rect 4755 3964 4936 3992
rect 5537 3995 5595 4001
rect 4755 3961 4767 3964
rect 4709 3955 4767 3961
rect 5537 3961 5549 3995
rect 5583 3961 5595 3995
rect 5537 3955 5595 3961
rect 8297 3995 8355 4001
rect 8297 3961 8309 3995
rect 8343 3961 8355 3995
rect 8297 3955 8355 3961
rect 8389 3995 8447 4001
rect 8389 3961 8401 3995
rect 8435 3992 8447 3995
rect 8570 3992 8576 4004
rect 8435 3964 8576 3992
rect 8435 3961 8447 3964
rect 8389 3955 8447 3961
rect 4338 3924 4344 3936
rect 4126 3896 4344 3924
rect 2409 3887 2467 3893
rect 4338 3884 4344 3896
rect 4396 3884 4402 3936
rect 5552 3924 5580 3955
rect 6086 3924 6092 3936
rect 5552 3896 6092 3924
rect 6086 3884 6092 3896
rect 6144 3924 6150 3936
rect 6270 3924 6276 3936
rect 6144 3896 6276 3924
rect 6144 3884 6150 3896
rect 6270 3884 6276 3896
rect 6328 3884 6334 3936
rect 7009 3927 7067 3933
rect 7009 3893 7021 3927
rect 7055 3924 7067 3927
rect 7098 3924 7104 3936
rect 7055 3896 7104 3924
rect 7055 3893 7067 3896
rect 7009 3887 7067 3893
rect 7098 3884 7104 3896
rect 7156 3884 7162 3936
rect 8312 3924 8340 3955
rect 8570 3952 8576 3964
rect 8628 3952 8634 4004
rect 9214 3952 9220 4004
rect 9272 3952 9278 4004
rect 10134 3952 10140 4004
rect 10192 3992 10198 4004
rect 10962 3992 10968 4004
rect 10192 3964 10968 3992
rect 10192 3952 10198 3964
rect 10962 3952 10968 3964
rect 11020 3952 11026 4004
rect 12452 3992 12480 4020
rect 14550 3992 14556 4004
rect 12452 3964 12731 3992
rect 14511 3964 14556 3992
rect 9232 3924 9260 3952
rect 9858 3924 9864 3936
rect 8312 3896 9260 3924
rect 9819 3896 9864 3924
rect 9858 3884 9864 3896
rect 9916 3884 9922 3936
rect 11471 3927 11529 3933
rect 11471 3893 11483 3927
rect 11517 3924 11529 3927
rect 12342 3924 12348 3936
rect 11517 3896 12348 3924
rect 11517 3893 11529 3896
rect 11471 3887 11529 3893
rect 12342 3884 12348 3896
rect 12400 3884 12406 3936
rect 12526 3924 12532 3936
rect 12487 3896 12532 3924
rect 12526 3884 12532 3896
rect 12584 3884 12590 3936
rect 12703 3924 12731 3964
rect 14550 3952 14556 3964
rect 14608 3952 14614 4004
rect 14642 3952 14648 4004
rect 14700 3992 14706 4004
rect 15197 3995 15255 4001
rect 14700 3964 14745 3992
rect 14700 3952 14706 3964
rect 15197 3961 15209 3995
rect 15243 3992 15255 3995
rect 16114 3992 16120 4004
rect 15243 3964 16120 3992
rect 15243 3961 15255 3964
rect 15197 3955 15255 3961
rect 16114 3952 16120 3964
rect 16172 3952 16178 4004
rect 16209 3995 16267 4001
rect 16209 3961 16221 3995
rect 16255 3992 16267 3995
rect 16298 3992 16304 4004
rect 16255 3964 16304 3992
rect 16255 3961 16267 3964
rect 16209 3955 16267 3961
rect 16298 3952 16304 3964
rect 16356 3952 16362 4004
rect 16776 3992 16804 4088
rect 18598 4020 18604 4072
rect 18656 4060 18662 4072
rect 19334 4060 19340 4072
rect 18656 4032 19340 4060
rect 18656 4020 18662 4032
rect 19334 4020 19340 4032
rect 19392 4020 19398 4072
rect 21396 4063 21454 4069
rect 21396 4060 21408 4063
rect 21376 4029 21408 4060
rect 21442 4029 21454 4063
rect 21376 4023 21454 4029
rect 18874 3992 18880 4004
rect 16776 3964 18880 3992
rect 18874 3952 18880 3964
rect 18932 3952 18938 4004
rect 19886 3992 19892 4004
rect 19847 3964 19892 3992
rect 19886 3952 19892 3964
rect 19944 3952 19950 4004
rect 19981 3995 20039 4001
rect 19981 3961 19993 3995
rect 20027 3961 20039 3995
rect 19981 3955 20039 3961
rect 14274 3924 14280 3936
rect 12703 3896 14280 3924
rect 14274 3884 14280 3896
rect 14332 3924 14338 3936
rect 15470 3924 15476 3936
rect 14332 3896 15476 3924
rect 14332 3884 14338 3896
rect 15470 3884 15476 3896
rect 15528 3924 15534 3936
rect 15841 3927 15899 3933
rect 15841 3924 15853 3927
rect 15528 3896 15853 3924
rect 15528 3884 15534 3896
rect 15841 3893 15853 3896
rect 15887 3893 15899 3927
rect 15841 3887 15899 3893
rect 17310 3884 17316 3936
rect 17368 3924 17374 3936
rect 17865 3927 17923 3933
rect 17865 3924 17877 3927
rect 17368 3896 17877 3924
rect 17368 3884 17374 3896
rect 17865 3893 17877 3896
rect 17911 3924 17923 3927
rect 18417 3927 18475 3933
rect 18417 3924 18429 3927
rect 17911 3896 18429 3924
rect 17911 3893 17923 3896
rect 17865 3887 17923 3893
rect 18417 3893 18429 3896
rect 18463 3893 18475 3927
rect 18966 3924 18972 3936
rect 18927 3896 18972 3924
rect 18417 3887 18475 3893
rect 18966 3884 18972 3896
rect 19024 3884 19030 3936
rect 19150 3884 19156 3936
rect 19208 3924 19214 3936
rect 19613 3927 19671 3933
rect 19613 3924 19625 3927
rect 19208 3896 19625 3924
rect 19208 3884 19214 3896
rect 19613 3893 19625 3896
rect 19659 3924 19671 3927
rect 19996 3924 20024 3955
rect 21376 3936 21404 4023
rect 19659 3896 20024 3924
rect 19659 3893 19671 3896
rect 19613 3887 19671 3893
rect 21358 3884 21364 3936
rect 21416 3924 21422 3936
rect 21821 3927 21879 3933
rect 21821 3924 21833 3927
rect 21416 3896 21833 3924
rect 21416 3884 21422 3896
rect 21821 3893 21833 3896
rect 21867 3893 21879 3927
rect 21821 3887 21879 3893
rect 1104 3834 22816 3856
rect 1104 3782 8982 3834
rect 9034 3782 9046 3834
rect 9098 3782 9110 3834
rect 9162 3782 9174 3834
rect 9226 3782 16982 3834
rect 17034 3782 17046 3834
rect 17098 3782 17110 3834
rect 17162 3782 17174 3834
rect 17226 3782 22816 3834
rect 1104 3760 22816 3782
rect 2501 3723 2559 3729
rect 2501 3689 2513 3723
rect 2547 3720 2559 3723
rect 2682 3720 2688 3732
rect 2547 3692 2688 3720
rect 2547 3689 2559 3692
rect 2501 3683 2559 3689
rect 2682 3680 2688 3692
rect 2740 3680 2746 3732
rect 3418 3720 3424 3732
rect 3379 3692 3424 3720
rect 3418 3680 3424 3692
rect 3476 3680 3482 3732
rect 5258 3720 5264 3732
rect 5219 3692 5264 3720
rect 5258 3680 5264 3692
rect 5316 3680 5322 3732
rect 6454 3720 6460 3732
rect 6415 3692 6460 3720
rect 6454 3680 6460 3692
rect 6512 3680 6518 3732
rect 7742 3720 7748 3732
rect 7655 3692 7748 3720
rect 7742 3680 7748 3692
rect 7800 3720 7806 3732
rect 8294 3720 8300 3732
rect 7800 3692 8300 3720
rect 7800 3680 7806 3692
rect 8294 3680 8300 3692
rect 8352 3680 8358 3732
rect 9309 3723 9367 3729
rect 9309 3689 9321 3723
rect 9355 3720 9367 3723
rect 9398 3720 9404 3732
rect 9355 3692 9404 3720
rect 9355 3689 9367 3692
rect 9309 3683 9367 3689
rect 9398 3680 9404 3692
rect 9456 3680 9462 3732
rect 10134 3720 10140 3732
rect 10060 3692 10140 3720
rect 1670 3652 1676 3664
rect 1412 3624 1676 3652
rect 1412 3593 1440 3624
rect 1670 3612 1676 3624
rect 1728 3652 1734 3664
rect 6178 3652 6184 3664
rect 1728 3624 6184 3652
rect 1728 3612 1734 3624
rect 6178 3612 6184 3624
rect 6236 3612 6242 3664
rect 6638 3612 6644 3664
rect 6696 3652 6702 3664
rect 8665 3655 8723 3661
rect 6696 3624 7373 3652
rect 6696 3612 6702 3624
rect 1397 3587 1455 3593
rect 1397 3553 1409 3587
rect 1443 3553 1455 3587
rect 2958 3584 2964 3596
rect 2919 3556 2964 3584
rect 1397 3547 1455 3553
rect 2958 3544 2964 3556
rect 3016 3544 3022 3596
rect 3418 3544 3424 3596
rect 3476 3584 3482 3596
rect 4890 3584 4896 3596
rect 3476 3556 4896 3584
rect 3476 3544 3482 3556
rect 4890 3544 4896 3556
rect 4948 3584 4954 3596
rect 5718 3584 5724 3596
rect 4948 3556 5724 3584
rect 4948 3544 4954 3556
rect 5718 3544 5724 3556
rect 5776 3544 5782 3596
rect 6549 3587 6607 3593
rect 6549 3553 6561 3587
rect 6595 3584 6607 3587
rect 6730 3584 6736 3596
rect 6595 3556 6736 3584
rect 6595 3553 6607 3556
rect 6549 3547 6607 3553
rect 6730 3544 6736 3556
rect 6788 3544 6794 3596
rect 6825 3587 6883 3593
rect 6825 3553 6837 3587
rect 6871 3553 6883 3587
rect 6825 3547 6883 3553
rect 3099 3519 3157 3525
rect 3099 3485 3111 3519
rect 3145 3516 3157 3519
rect 3145 3488 6316 3516
rect 3145 3485 3157 3488
rect 3099 3479 3157 3485
rect 1578 3380 1584 3392
rect 1539 3352 1584 3380
rect 1578 3340 1584 3352
rect 1636 3340 1642 3392
rect 4706 3380 4712 3392
rect 4667 3352 4712 3380
rect 4706 3340 4712 3352
rect 4764 3340 4770 3392
rect 6288 3380 6316 3488
rect 6362 3408 6368 3460
rect 6420 3448 6426 3460
rect 6840 3448 6868 3547
rect 7345 3516 7373 3624
rect 8665 3621 8677 3655
rect 8711 3652 8723 3655
rect 9950 3652 9956 3664
rect 8711 3624 9956 3652
rect 8711 3621 8723 3624
rect 8665 3615 8723 3621
rect 9950 3612 9956 3624
rect 10008 3612 10014 3664
rect 7926 3584 7932 3596
rect 7887 3556 7932 3584
rect 7926 3544 7932 3556
rect 7984 3544 7990 3596
rect 8202 3584 8208 3596
rect 8163 3556 8208 3584
rect 8202 3544 8208 3556
rect 8260 3544 8266 3596
rect 9861 3587 9919 3593
rect 9861 3584 9873 3587
rect 8864 3556 9873 3584
rect 8864 3516 8892 3556
rect 9861 3553 9873 3556
rect 9907 3584 9919 3587
rect 10060 3584 10088 3692
rect 10134 3680 10140 3692
rect 10192 3680 10198 3732
rect 11238 3720 11244 3732
rect 11199 3692 11244 3720
rect 11238 3680 11244 3692
rect 11296 3680 11302 3732
rect 12434 3720 12440 3732
rect 12395 3692 12440 3720
rect 12434 3680 12440 3692
rect 12492 3680 12498 3732
rect 14553 3723 14611 3729
rect 14553 3689 14565 3723
rect 14599 3720 14611 3723
rect 14642 3720 14648 3732
rect 14599 3692 14648 3720
rect 14599 3689 14611 3692
rect 14553 3683 14611 3689
rect 14642 3680 14648 3692
rect 14700 3680 14706 3732
rect 16209 3723 16267 3729
rect 16209 3689 16221 3723
rect 16255 3720 16267 3723
rect 16298 3720 16304 3732
rect 16255 3692 16304 3720
rect 16255 3689 16267 3692
rect 16209 3683 16267 3689
rect 16298 3680 16304 3692
rect 16356 3680 16362 3732
rect 18046 3720 18052 3732
rect 18007 3692 18052 3720
rect 18046 3680 18052 3692
rect 18104 3680 18110 3732
rect 19886 3720 19892 3732
rect 19847 3692 19892 3720
rect 19886 3680 19892 3692
rect 19944 3680 19950 3732
rect 10318 3652 10324 3664
rect 10279 3624 10324 3652
rect 10318 3612 10324 3624
rect 10376 3612 10382 3664
rect 13081 3655 13139 3661
rect 13081 3621 13093 3655
rect 13127 3652 13139 3655
rect 13354 3652 13360 3664
rect 13127 3624 13360 3652
rect 13127 3621 13139 3624
rect 13081 3615 13139 3621
rect 13354 3612 13360 3624
rect 13412 3612 13418 3664
rect 15651 3655 15709 3661
rect 15651 3621 15663 3655
rect 15697 3652 15709 3655
rect 15746 3652 15752 3664
rect 15697 3624 15752 3652
rect 15697 3621 15709 3624
rect 15651 3615 15709 3621
rect 15746 3612 15752 3624
rect 15804 3612 15810 3664
rect 16114 3612 16120 3664
rect 16172 3652 16178 3664
rect 16485 3655 16543 3661
rect 16485 3652 16497 3655
rect 16172 3624 16497 3652
rect 16172 3612 16178 3624
rect 16485 3621 16497 3624
rect 16531 3652 16543 3655
rect 16574 3652 16580 3664
rect 16531 3624 16580 3652
rect 16531 3621 16543 3624
rect 16485 3615 16543 3621
rect 16574 3612 16580 3624
rect 16632 3612 16638 3664
rect 18414 3612 18420 3664
rect 18472 3652 18478 3664
rect 18693 3655 18751 3661
rect 18693 3652 18705 3655
rect 18472 3624 18705 3652
rect 18472 3612 18478 3624
rect 18693 3621 18705 3624
rect 18739 3652 18751 3655
rect 18966 3652 18972 3664
rect 18739 3624 18972 3652
rect 18739 3621 18751 3624
rect 18693 3615 18751 3621
rect 18966 3612 18972 3624
rect 19024 3612 19030 3664
rect 11790 3584 11796 3596
rect 9907 3556 10088 3584
rect 11751 3556 11796 3584
rect 9907 3553 9919 3556
rect 9861 3547 9919 3553
rect 11790 3544 11796 3556
rect 11848 3544 11854 3596
rect 15289 3587 15347 3593
rect 15289 3553 15301 3587
rect 15335 3584 15347 3587
rect 15378 3584 15384 3596
rect 15335 3556 15384 3584
rect 15335 3553 15347 3556
rect 15289 3547 15347 3553
rect 15378 3544 15384 3556
rect 15436 3544 15442 3596
rect 16666 3544 16672 3596
rect 16724 3584 16730 3596
rect 17037 3587 17095 3593
rect 17037 3584 17049 3587
rect 16724 3556 17049 3584
rect 16724 3544 16730 3556
rect 17037 3553 17049 3556
rect 17083 3584 17095 3587
rect 17589 3587 17647 3593
rect 17589 3584 17601 3587
rect 17083 3556 17601 3584
rect 17083 3553 17095 3556
rect 17037 3547 17095 3553
rect 17589 3553 17601 3556
rect 17635 3553 17647 3587
rect 17589 3547 17647 3553
rect 20968 3587 21026 3593
rect 20968 3553 20980 3587
rect 21014 3584 21026 3587
rect 21266 3584 21272 3596
rect 21014 3556 21272 3584
rect 21014 3553 21026 3556
rect 20968 3547 21026 3553
rect 21266 3544 21272 3556
rect 21324 3544 21330 3596
rect 10229 3519 10287 3525
rect 10229 3516 10241 3519
rect 7345 3488 8892 3516
rect 8956 3488 10241 3516
rect 8018 3448 8024 3460
rect 6420 3420 6868 3448
rect 7979 3420 8024 3448
rect 6420 3408 6426 3420
rect 8018 3408 8024 3420
rect 8076 3408 8082 3460
rect 8956 3380 8984 3488
rect 10229 3485 10241 3488
rect 10275 3516 10287 3519
rect 11330 3516 11336 3528
rect 10275 3488 11336 3516
rect 10275 3485 10287 3488
rect 10229 3479 10287 3485
rect 11330 3476 11336 3488
rect 11388 3476 11394 3528
rect 12989 3519 13047 3525
rect 12989 3485 13001 3519
rect 13035 3516 13047 3519
rect 13262 3516 13268 3528
rect 13035 3488 13268 3516
rect 13035 3485 13047 3488
rect 12989 3479 13047 3485
rect 13262 3476 13268 3488
rect 13320 3516 13326 3528
rect 13909 3519 13967 3525
rect 13909 3516 13921 3519
rect 13320 3488 13921 3516
rect 13320 3476 13326 3488
rect 13909 3485 13921 3488
rect 13955 3485 13967 3519
rect 13909 3479 13967 3485
rect 18601 3519 18659 3525
rect 18601 3485 18613 3519
rect 18647 3516 18659 3519
rect 18782 3516 18788 3528
rect 18647 3488 18788 3516
rect 18647 3485 18659 3488
rect 18601 3479 18659 3485
rect 18782 3476 18788 3488
rect 18840 3476 18846 3528
rect 18874 3476 18880 3528
rect 18932 3516 18938 3528
rect 18969 3519 19027 3525
rect 18969 3516 18981 3519
rect 18932 3488 18981 3516
rect 18932 3476 18938 3488
rect 18969 3485 18981 3488
rect 19015 3485 19027 3519
rect 18969 3479 19027 3485
rect 10781 3451 10839 3457
rect 10781 3417 10793 3451
rect 10827 3448 10839 3451
rect 13541 3451 13599 3457
rect 13541 3448 13553 3451
rect 10827 3420 13553 3448
rect 10827 3417 10839 3420
rect 10781 3411 10839 3417
rect 13541 3417 13553 3420
rect 13587 3448 13599 3451
rect 13630 3448 13636 3460
rect 13587 3420 13636 3448
rect 13587 3417 13599 3420
rect 13541 3411 13599 3417
rect 13630 3408 13636 3420
rect 13688 3408 13694 3460
rect 6288 3352 8984 3380
rect 11701 3383 11759 3389
rect 11701 3349 11713 3383
rect 11747 3380 11759 3383
rect 11790 3380 11796 3392
rect 11747 3352 11796 3380
rect 11747 3349 11759 3352
rect 11701 3343 11759 3349
rect 11790 3340 11796 3352
rect 11848 3340 11854 3392
rect 11974 3380 11980 3392
rect 11935 3352 11980 3380
rect 11974 3340 11980 3352
rect 12032 3340 12038 3392
rect 15470 3340 15476 3392
rect 15528 3380 15534 3392
rect 17221 3383 17279 3389
rect 17221 3380 17233 3383
rect 15528 3352 17233 3380
rect 15528 3340 15534 3352
rect 17221 3349 17233 3352
rect 17267 3349 17279 3383
rect 17221 3343 17279 3349
rect 17402 3340 17408 3392
rect 17460 3380 17466 3392
rect 21039 3383 21097 3389
rect 21039 3380 21051 3383
rect 17460 3352 21051 3380
rect 17460 3340 17466 3352
rect 21039 3349 21051 3352
rect 21085 3349 21097 3383
rect 21039 3343 21097 3349
rect 1104 3290 22816 3312
rect 1104 3238 4982 3290
rect 5034 3238 5046 3290
rect 5098 3238 5110 3290
rect 5162 3238 5174 3290
rect 5226 3238 12982 3290
rect 13034 3238 13046 3290
rect 13098 3238 13110 3290
rect 13162 3238 13174 3290
rect 13226 3238 20982 3290
rect 21034 3238 21046 3290
rect 21098 3238 21110 3290
rect 21162 3238 21174 3290
rect 21226 3238 22816 3290
rect 1104 3216 22816 3238
rect 1670 3176 1676 3188
rect 1631 3148 1676 3176
rect 1670 3136 1676 3148
rect 1728 3136 1734 3188
rect 3234 3176 3240 3188
rect 3195 3148 3240 3176
rect 3234 3136 3240 3148
rect 3292 3136 3298 3188
rect 6362 3176 6368 3188
rect 6323 3148 6368 3176
rect 6362 3136 6368 3148
rect 6420 3136 6426 3188
rect 10042 3176 10048 3188
rect 10003 3148 10048 3176
rect 10042 3136 10048 3148
rect 10100 3176 10106 3188
rect 13354 3176 13360 3188
rect 10100 3148 10640 3176
rect 13315 3148 13360 3176
rect 10100 3136 10106 3148
rect 4706 3108 4712 3120
rect 4667 3080 4712 3108
rect 4706 3068 4712 3080
rect 4764 3068 4770 3120
rect 5626 3108 5632 3120
rect 5276 3080 5632 3108
rect 5276 3040 5304 3080
rect 5626 3068 5632 3080
rect 5684 3108 5690 3120
rect 7926 3108 7932 3120
rect 5684 3080 7932 3108
rect 5684 3068 5690 3080
rect 7926 3068 7932 3080
rect 7984 3108 7990 3120
rect 8665 3111 8723 3117
rect 8665 3108 8677 3111
rect 7984 3080 8677 3108
rect 7984 3068 7990 3080
rect 8665 3077 8677 3080
rect 8711 3077 8723 3111
rect 10502 3108 10508 3120
rect 10463 3080 10508 3108
rect 8665 3071 8723 3077
rect 10502 3068 10508 3080
rect 10560 3068 10566 3120
rect 4632 3012 5304 3040
rect 5353 3043 5411 3049
rect 4632 2981 4660 3012
rect 5353 3009 5365 3043
rect 5399 3040 5411 3043
rect 6638 3040 6644 3052
rect 5399 3012 6644 3040
rect 5399 3009 5411 3012
rect 5353 3003 5411 3009
rect 6638 3000 6644 3012
rect 6696 3000 6702 3052
rect 6730 3000 6736 3052
rect 6788 3040 6794 3052
rect 7101 3043 7159 3049
rect 7101 3040 7113 3043
rect 6788 3012 7113 3040
rect 6788 3000 6794 3012
rect 7101 3009 7113 3012
rect 7147 3040 7159 3043
rect 7190 3040 7196 3052
rect 7147 3012 7196 3040
rect 7147 3009 7159 3012
rect 7101 3003 7159 3009
rect 7190 3000 7196 3012
rect 7248 3000 7254 3052
rect 7742 3040 7748 3052
rect 7703 3012 7748 3040
rect 7742 3000 7748 3012
rect 7800 3000 7806 3052
rect 8386 3040 8392 3052
rect 8347 3012 8392 3040
rect 8386 3000 8392 3012
rect 8444 3000 8450 3052
rect 2685 2975 2743 2981
rect 2685 2941 2697 2975
rect 2731 2972 2743 2975
rect 3053 2975 3111 2981
rect 3053 2972 3065 2975
rect 2731 2944 3065 2972
rect 2731 2941 2743 2944
rect 2685 2935 2743 2941
rect 3053 2941 3065 2944
rect 3099 2972 3111 2975
rect 4433 2975 4491 2981
rect 4433 2972 4445 2975
rect 3099 2944 4445 2972
rect 3099 2941 3111 2944
rect 3053 2935 3111 2941
rect 4433 2941 4445 2944
rect 4479 2972 4491 2975
rect 4617 2975 4675 2981
rect 4617 2972 4629 2975
rect 4479 2944 4629 2972
rect 4479 2941 4491 2944
rect 4433 2935 4491 2941
rect 4617 2941 4629 2944
rect 4663 2941 4675 2975
rect 4617 2935 4675 2941
rect 4890 2932 4896 2984
rect 4948 2972 4954 2984
rect 4948 2944 4993 2972
rect 4948 2932 4954 2944
rect 5166 2932 5172 2984
rect 5224 2972 5230 2984
rect 6748 2972 6776 3000
rect 5224 2944 6776 2972
rect 9217 2975 9275 2981
rect 5224 2932 5230 2944
rect 9217 2941 9229 2975
rect 9263 2972 9275 2975
rect 9398 2972 9404 2984
rect 9263 2944 9404 2972
rect 9263 2941 9275 2944
rect 9217 2935 9275 2941
rect 9398 2932 9404 2944
rect 9456 2932 9462 2984
rect 10520 2972 10548 3068
rect 10612 3049 10640 3148
rect 13354 3136 13360 3148
rect 13412 3136 13418 3188
rect 14642 3136 14648 3188
rect 14700 3176 14706 3188
rect 15102 3176 15108 3188
rect 14700 3148 15108 3176
rect 14700 3136 14706 3148
rect 15102 3136 15108 3148
rect 15160 3136 15166 3188
rect 15562 3136 15568 3188
rect 15620 3176 15626 3188
rect 15749 3179 15807 3185
rect 15749 3176 15761 3179
rect 15620 3148 15761 3176
rect 15620 3136 15626 3148
rect 15749 3145 15761 3148
rect 15795 3145 15807 3179
rect 18414 3176 18420 3188
rect 18375 3148 18420 3176
rect 15749 3139 15807 3145
rect 10597 3043 10655 3049
rect 10597 3009 10609 3043
rect 10643 3009 10655 3043
rect 10597 3003 10655 3009
rect 11885 3043 11943 3049
rect 11885 3009 11897 3043
rect 11931 3040 11943 3043
rect 12437 3043 12495 3049
rect 12437 3040 12449 3043
rect 11931 3012 12449 3040
rect 11931 3009 11943 3012
rect 11885 3003 11943 3009
rect 12437 3009 12449 3012
rect 12483 3040 12495 3043
rect 12526 3040 12532 3052
rect 12483 3012 12532 3040
rect 12483 3009 12495 3012
rect 12437 3003 12495 3009
rect 12526 3000 12532 3012
rect 12584 3000 12590 3052
rect 14001 3043 14059 3049
rect 14001 3040 14013 3043
rect 12636 3012 14013 3040
rect 12161 2975 12219 2981
rect 12161 2972 12173 2975
rect 10520 2944 12173 2972
rect 2501 2907 2559 2913
rect 2501 2873 2513 2907
rect 2547 2904 2559 2907
rect 2958 2904 2964 2916
rect 2547 2876 2964 2904
rect 2547 2873 2559 2876
rect 2501 2867 2559 2873
rect 2958 2864 2964 2876
rect 3016 2904 3022 2916
rect 5902 2904 5908 2916
rect 3016 2876 5908 2904
rect 3016 2864 3022 2876
rect 5902 2864 5908 2876
rect 5960 2864 5966 2916
rect 7742 2904 7748 2916
rect 7024 2876 7748 2904
rect 2314 2796 2320 2848
rect 2372 2836 2378 2848
rect 2685 2839 2743 2845
rect 2685 2836 2697 2839
rect 2372 2808 2697 2836
rect 2372 2796 2378 2808
rect 2685 2805 2697 2808
rect 2731 2836 2743 2839
rect 2777 2839 2835 2845
rect 2777 2836 2789 2839
rect 2731 2808 2789 2836
rect 2731 2805 2743 2808
rect 2685 2799 2743 2805
rect 2777 2805 2789 2808
rect 2823 2805 2835 2839
rect 2777 2799 2835 2805
rect 4157 2839 4215 2845
rect 4157 2805 4169 2839
rect 4203 2836 4215 2839
rect 4338 2836 4344 2848
rect 4203 2808 4344 2836
rect 4203 2805 4215 2808
rect 4157 2799 4215 2805
rect 4338 2796 4344 2808
rect 4396 2836 4402 2848
rect 4890 2836 4896 2848
rect 4396 2808 4896 2836
rect 4396 2796 4402 2808
rect 4890 2796 4896 2808
rect 4948 2796 4954 2848
rect 5718 2836 5724 2848
rect 5631 2808 5724 2836
rect 5718 2796 5724 2808
rect 5776 2836 5782 2848
rect 7024 2836 7052 2876
rect 7742 2864 7748 2876
rect 7800 2864 7806 2916
rect 10933 2913 10961 2944
rect 12161 2941 12173 2944
rect 12207 2972 12219 2975
rect 12636 2972 12664 3012
rect 14001 3009 14013 3012
rect 14047 3040 14059 3043
rect 15764 3040 15792 3139
rect 18414 3136 18420 3148
rect 18472 3136 18478 3188
rect 18690 3136 18696 3188
rect 18748 3176 18754 3188
rect 19889 3179 19947 3185
rect 19889 3176 19901 3179
rect 18748 3148 19901 3176
rect 18748 3136 18754 3148
rect 19889 3145 19901 3148
rect 19935 3145 19947 3179
rect 19889 3139 19947 3145
rect 18782 3068 18788 3120
rect 18840 3108 18846 3120
rect 19521 3111 19579 3117
rect 19521 3108 19533 3111
rect 18840 3080 19533 3108
rect 18840 3068 18846 3080
rect 19521 3077 19533 3080
rect 19567 3077 19579 3111
rect 19521 3071 19579 3077
rect 18874 3040 18880 3052
rect 14047 3012 14549 3040
rect 15764 3012 16436 3040
rect 18835 3012 18880 3040
rect 14047 3009 14059 3012
rect 14001 3003 14059 3009
rect 14185 2975 14243 2981
rect 12207 2944 12801 2972
rect 12207 2941 12219 2944
rect 12161 2935 12219 2941
rect 12773 2913 12801 2944
rect 14185 2941 14197 2975
rect 14231 2941 14243 2975
rect 14185 2935 14243 2941
rect 7837 2907 7895 2913
rect 7837 2873 7849 2907
rect 7883 2873 7895 2907
rect 9033 2907 9091 2913
rect 9033 2904 9045 2907
rect 7837 2867 7895 2873
rect 8588 2876 9045 2904
rect 5776 2808 7052 2836
rect 7561 2839 7619 2845
rect 5776 2796 5782 2808
rect 7561 2805 7573 2839
rect 7607 2836 7619 2839
rect 7650 2836 7656 2848
rect 7607 2808 7656 2836
rect 7607 2805 7619 2808
rect 7561 2799 7619 2805
rect 7650 2796 7656 2808
rect 7708 2796 7714 2848
rect 7852 2836 7880 2867
rect 7926 2836 7932 2848
rect 7839 2808 7932 2836
rect 7926 2796 7932 2808
rect 7984 2836 7990 2848
rect 8588 2836 8616 2876
rect 9033 2873 9045 2876
rect 9079 2873 9091 2907
rect 10918 2907 10976 2913
rect 10918 2904 10930 2907
rect 10896 2876 10930 2904
rect 9033 2867 9091 2873
rect 10918 2873 10930 2876
rect 10964 2873 10976 2907
rect 10918 2867 10976 2873
rect 12758 2907 12816 2913
rect 12758 2873 12770 2907
rect 12804 2873 12816 2907
rect 12758 2867 12816 2873
rect 13725 2907 13783 2913
rect 13725 2873 13737 2907
rect 13771 2904 13783 2907
rect 14200 2904 14228 2935
rect 14521 2913 14549 3012
rect 16206 2972 16212 2984
rect 16167 2944 16212 2972
rect 16206 2932 16212 2944
rect 16264 2932 16270 2984
rect 16408 2981 16436 3012
rect 18874 3000 18880 3012
rect 18932 3000 18938 3052
rect 19334 3000 19340 3052
rect 19392 3000 19398 3052
rect 19904 3040 19932 3139
rect 19904 3012 20576 3040
rect 16393 2975 16451 2981
rect 16393 2941 16405 2975
rect 16439 2941 16451 2975
rect 19352 2972 19380 3000
rect 20070 2972 20076 2984
rect 19352 2944 20076 2972
rect 16393 2935 16451 2941
rect 20070 2932 20076 2944
rect 20128 2932 20134 2984
rect 20548 2981 20576 3012
rect 20533 2975 20591 2981
rect 20533 2941 20545 2975
rect 20579 2941 20591 2975
rect 20533 2935 20591 2941
rect 13771 2876 14228 2904
rect 13771 2873 13783 2876
rect 13725 2867 13783 2873
rect 9398 2836 9404 2848
rect 7984 2808 8616 2836
rect 9359 2808 9404 2836
rect 7984 2796 7990 2808
rect 9398 2796 9404 2808
rect 9456 2796 9462 2848
rect 11517 2839 11575 2845
rect 11517 2805 11529 2839
rect 11563 2836 11575 2839
rect 12066 2836 12072 2848
rect 11563 2808 12072 2836
rect 11563 2805 11575 2808
rect 11517 2799 11575 2805
rect 12066 2796 12072 2808
rect 12124 2796 12130 2848
rect 14200 2836 14228 2876
rect 14506 2907 14564 2913
rect 14506 2873 14518 2907
rect 14552 2873 14564 2907
rect 14506 2867 14564 2873
rect 15473 2907 15531 2913
rect 15473 2873 15485 2907
rect 15519 2904 15531 2907
rect 15746 2904 15752 2916
rect 15519 2876 15752 2904
rect 15519 2873 15531 2876
rect 15473 2867 15531 2873
rect 15746 2864 15752 2876
rect 15804 2864 15810 2916
rect 16224 2904 16252 2932
rect 16945 2907 17003 2913
rect 16945 2904 16957 2907
rect 16224 2876 16957 2904
rect 16945 2873 16957 2876
rect 16991 2873 17003 2907
rect 16945 2867 17003 2873
rect 17497 2907 17555 2913
rect 17497 2873 17509 2907
rect 17543 2904 17555 2907
rect 18598 2904 18604 2916
rect 17543 2876 18604 2904
rect 17543 2873 17555 2876
rect 17497 2867 17555 2873
rect 18598 2864 18604 2876
rect 18656 2864 18662 2916
rect 18693 2907 18751 2913
rect 18693 2873 18705 2907
rect 18739 2873 18751 2907
rect 18693 2867 18751 2873
rect 16025 2839 16083 2845
rect 16025 2836 16037 2839
rect 14200 2808 16037 2836
rect 16025 2805 16037 2808
rect 16071 2805 16083 2839
rect 17862 2836 17868 2848
rect 17775 2808 17868 2836
rect 16025 2799 16083 2805
rect 17862 2796 17868 2808
rect 17920 2836 17926 2848
rect 18708 2836 18736 2867
rect 19058 2864 19064 2916
rect 19116 2904 19122 2916
rect 20714 2904 20720 2916
rect 19116 2876 20720 2904
rect 19116 2864 19122 2876
rect 20714 2864 20720 2876
rect 20772 2864 20778 2916
rect 20162 2836 20168 2848
rect 17920 2808 18736 2836
rect 20123 2808 20168 2836
rect 17920 2796 17926 2808
rect 20162 2796 20168 2808
rect 20220 2796 20226 2848
rect 21177 2839 21235 2845
rect 21177 2805 21189 2839
rect 21223 2836 21235 2839
rect 21266 2836 21272 2848
rect 21223 2808 21272 2836
rect 21223 2805 21235 2808
rect 21177 2799 21235 2805
rect 21266 2796 21272 2808
rect 21324 2836 21330 2848
rect 22462 2836 22468 2848
rect 21324 2808 22468 2836
rect 21324 2796 21330 2808
rect 22462 2796 22468 2808
rect 22520 2796 22526 2848
rect 1104 2746 22816 2768
rect 1104 2694 8982 2746
rect 9034 2694 9046 2746
rect 9098 2694 9110 2746
rect 9162 2694 9174 2746
rect 9226 2694 16982 2746
rect 17034 2694 17046 2746
rect 17098 2694 17110 2746
rect 17162 2694 17174 2746
rect 17226 2694 22816 2746
rect 1104 2672 22816 2694
rect 3510 2632 3516 2644
rect 3471 2604 3516 2632
rect 3510 2592 3516 2604
rect 3568 2592 3574 2644
rect 4341 2635 4399 2641
rect 4341 2601 4353 2635
rect 4387 2632 4399 2635
rect 4890 2632 4896 2644
rect 4387 2604 4896 2632
rect 4387 2601 4399 2604
rect 4341 2595 4399 2601
rect 4890 2592 4896 2604
rect 4948 2592 4954 2644
rect 6365 2635 6423 2641
rect 6365 2601 6377 2635
rect 6411 2632 6423 2635
rect 6454 2632 6460 2644
rect 6411 2604 6460 2632
rect 6411 2601 6423 2604
rect 6365 2595 6423 2601
rect 6454 2592 6460 2604
rect 6512 2632 6518 2644
rect 7926 2632 7932 2644
rect 6512 2604 7052 2632
rect 7887 2604 7932 2632
rect 6512 2592 6518 2604
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2465 1455 2499
rect 1397 2459 1455 2465
rect 2869 2499 2927 2505
rect 2869 2465 2881 2499
rect 2915 2496 2927 2499
rect 3528 2496 3556 2592
rect 4798 2564 4804 2576
rect 4448 2536 4804 2564
rect 4448 2505 4476 2536
rect 4798 2524 4804 2536
rect 4856 2564 4862 2576
rect 5813 2567 5871 2573
rect 5813 2564 5825 2567
rect 4856 2536 5825 2564
rect 4856 2524 4862 2536
rect 5813 2533 5825 2536
rect 5859 2533 5871 2567
rect 5813 2527 5871 2533
rect 6641 2567 6699 2573
rect 6641 2533 6653 2567
rect 6687 2533 6699 2567
rect 6641 2527 6699 2533
rect 2915 2468 3556 2496
rect 4433 2499 4491 2505
rect 2915 2465 2927 2468
rect 2869 2459 2927 2465
rect 4433 2465 4445 2499
rect 4479 2465 4491 2499
rect 4433 2459 4491 2465
rect 4709 2499 4767 2505
rect 4709 2465 4721 2499
rect 4755 2496 4767 2499
rect 4890 2496 4896 2508
rect 4755 2468 4896 2496
rect 4755 2465 4767 2468
rect 4709 2459 4767 2465
rect 1412 2428 1440 2459
rect 4890 2456 4896 2468
rect 4948 2456 4954 2508
rect 5166 2496 5172 2508
rect 5127 2468 5172 2496
rect 5166 2456 5172 2468
rect 5224 2456 5230 2508
rect 2038 2428 2044 2440
rect 1412 2400 2044 2428
rect 2038 2388 2044 2400
rect 2096 2388 2102 2440
rect 3881 2431 3939 2437
rect 3881 2397 3893 2431
rect 3927 2428 3939 2431
rect 5445 2431 5503 2437
rect 5445 2428 5457 2431
rect 3927 2400 4568 2428
rect 3927 2397 3939 2400
rect 3881 2391 3939 2397
rect 4540 2369 4568 2400
rect 5000 2400 5457 2428
rect 3053 2363 3111 2369
rect 3053 2329 3065 2363
rect 3099 2360 3111 2363
rect 4525 2363 4583 2369
rect 3099 2332 4476 2360
rect 3099 2329 3111 2332
rect 3053 2323 3111 2329
rect 106 2252 112 2304
rect 164 2292 170 2304
rect 1581 2295 1639 2301
rect 1581 2292 1593 2295
rect 164 2264 1593 2292
rect 164 2252 170 2264
rect 1581 2261 1593 2264
rect 1627 2261 1639 2295
rect 4448 2292 4476 2332
rect 4525 2329 4537 2363
rect 4571 2360 4583 2363
rect 4706 2360 4712 2372
rect 4571 2332 4712 2360
rect 4571 2329 4583 2332
rect 4525 2323 4583 2329
rect 4706 2320 4712 2332
rect 4764 2360 4770 2372
rect 5000 2360 5028 2400
rect 5445 2397 5457 2400
rect 5491 2397 5503 2431
rect 6656 2428 6684 2527
rect 7024 2505 7052 2604
rect 7926 2592 7932 2604
rect 7984 2592 7990 2644
rect 10318 2592 10324 2644
rect 10376 2632 10382 2644
rect 10689 2635 10747 2641
rect 10689 2632 10701 2635
rect 10376 2604 10701 2632
rect 10376 2592 10382 2604
rect 10689 2601 10701 2604
rect 10735 2632 10747 2635
rect 10965 2635 11023 2641
rect 10965 2632 10977 2635
rect 10735 2604 10977 2632
rect 10735 2601 10747 2604
rect 10689 2595 10747 2601
rect 10965 2601 10977 2604
rect 11011 2601 11023 2635
rect 11330 2632 11336 2644
rect 11291 2604 11336 2632
rect 10965 2595 11023 2601
rect 11330 2592 11336 2604
rect 11388 2592 11394 2644
rect 11655 2635 11713 2641
rect 11655 2601 11667 2635
rect 11701 2632 11713 2635
rect 11790 2632 11796 2644
rect 11701 2604 11796 2632
rect 11701 2601 11713 2604
rect 11655 2595 11713 2601
rect 11790 2592 11796 2604
rect 11848 2592 11854 2644
rect 12066 2592 12072 2644
rect 12124 2632 12130 2644
rect 12345 2635 12403 2641
rect 12345 2632 12357 2635
rect 12124 2604 12357 2632
rect 12124 2592 12130 2604
rect 12345 2601 12357 2604
rect 12391 2601 12403 2635
rect 12345 2595 12403 2601
rect 7330 2567 7388 2573
rect 7330 2533 7342 2567
rect 7376 2564 7388 2567
rect 9493 2567 9551 2573
rect 9493 2564 9505 2567
rect 7376 2536 9505 2564
rect 7376 2533 7388 2536
rect 7330 2527 7388 2533
rect 9493 2533 9505 2536
rect 9539 2564 9551 2567
rect 10131 2567 10189 2573
rect 10131 2564 10143 2567
rect 9539 2536 10143 2564
rect 9539 2533 9551 2536
rect 9493 2527 9551 2533
rect 10131 2533 10143 2536
rect 10177 2564 10189 2567
rect 10502 2564 10508 2576
rect 10177 2536 10508 2564
rect 10177 2533 10189 2536
rect 10131 2527 10189 2533
rect 7009 2499 7067 2505
rect 7009 2465 7021 2499
rect 7055 2465 7067 2499
rect 7009 2459 7067 2465
rect 7345 2428 7373 2527
rect 10502 2524 10508 2536
rect 10560 2524 10566 2576
rect 12360 2564 12388 2595
rect 13354 2592 13360 2644
rect 13412 2632 13418 2644
rect 13633 2635 13691 2641
rect 13633 2632 13645 2635
rect 13412 2604 13645 2632
rect 13412 2592 13418 2604
rect 13633 2601 13645 2604
rect 13679 2601 13691 2635
rect 13633 2595 13691 2601
rect 15289 2635 15347 2641
rect 15289 2601 15301 2635
rect 15335 2632 15347 2635
rect 15378 2632 15384 2644
rect 15335 2604 15384 2632
rect 15335 2601 15347 2604
rect 15289 2595 15347 2601
rect 15378 2592 15384 2604
rect 15436 2592 15442 2644
rect 17405 2635 17463 2641
rect 17405 2601 17417 2635
rect 17451 2632 17463 2635
rect 17862 2632 17868 2644
rect 17451 2604 17868 2632
rect 17451 2601 17463 2604
rect 17405 2595 17463 2601
rect 17862 2592 17868 2604
rect 17920 2592 17926 2644
rect 20162 2632 20168 2644
rect 18064 2604 20168 2632
rect 12805 2567 12863 2573
rect 12805 2564 12817 2567
rect 12360 2536 12817 2564
rect 12805 2533 12817 2536
rect 12851 2533 12863 2567
rect 12805 2527 12863 2533
rect 13722 2524 13728 2576
rect 13780 2564 13786 2576
rect 13780 2536 14504 2564
rect 13780 2524 13786 2536
rect 7650 2456 7656 2508
rect 7708 2496 7714 2508
rect 8202 2496 8208 2508
rect 7708 2468 8208 2496
rect 7708 2456 7714 2468
rect 8202 2456 8208 2468
rect 8260 2456 8266 2508
rect 9217 2499 9275 2505
rect 9217 2465 9229 2499
rect 9263 2496 9275 2499
rect 9769 2499 9827 2505
rect 9769 2496 9781 2499
rect 9263 2468 9781 2496
rect 9263 2465 9275 2468
rect 9217 2459 9275 2465
rect 9769 2465 9781 2468
rect 9815 2496 9827 2499
rect 9858 2496 9864 2508
rect 9815 2468 9864 2496
rect 9815 2465 9827 2468
rect 9769 2459 9827 2465
rect 9858 2456 9864 2468
rect 9916 2456 9922 2508
rect 11552 2499 11610 2505
rect 11552 2465 11564 2499
rect 11598 2496 11610 2499
rect 11977 2499 12035 2505
rect 11977 2496 11989 2499
rect 11598 2468 11989 2496
rect 11598 2465 11610 2468
rect 11552 2459 11610 2465
rect 11977 2465 11989 2468
rect 12023 2465 12035 2499
rect 11977 2459 12035 2465
rect 14185 2499 14243 2505
rect 14185 2465 14197 2499
rect 14231 2465 14243 2499
rect 14476 2496 14504 2536
rect 14550 2524 14556 2576
rect 14608 2564 14614 2576
rect 15611 2567 15669 2573
rect 15611 2564 15623 2567
rect 14608 2536 15623 2564
rect 14608 2524 14614 2536
rect 15611 2533 15623 2536
rect 15657 2533 15669 2567
rect 15611 2527 15669 2533
rect 15746 2524 15752 2576
rect 15804 2564 15810 2576
rect 16393 2567 16451 2573
rect 16393 2564 16405 2567
rect 15804 2536 16405 2564
rect 15804 2524 15810 2536
rect 16393 2533 16405 2536
rect 16439 2564 16451 2567
rect 16847 2567 16905 2573
rect 16847 2564 16859 2567
rect 16439 2536 16859 2564
rect 16439 2533 16451 2536
rect 16393 2527 16451 2533
rect 16847 2533 16859 2536
rect 16893 2564 16905 2567
rect 17310 2564 17316 2576
rect 16893 2536 17316 2564
rect 16893 2533 16905 2536
rect 16847 2527 16905 2533
rect 17310 2524 17316 2536
rect 17368 2524 17374 2576
rect 17773 2567 17831 2573
rect 17773 2533 17785 2567
rect 17819 2564 17831 2567
rect 18064 2564 18092 2604
rect 20162 2592 20168 2604
rect 20220 2592 20226 2644
rect 17819 2536 18092 2564
rect 18141 2567 18199 2573
rect 17819 2533 17831 2536
rect 17773 2527 17831 2533
rect 18141 2533 18153 2567
rect 18187 2564 18199 2567
rect 19058 2564 19064 2576
rect 18187 2536 19064 2564
rect 18187 2533 18199 2536
rect 18141 2527 18199 2533
rect 15286 2496 15292 2508
rect 14476 2468 15292 2496
rect 14185 2459 14243 2465
rect 6656 2400 7373 2428
rect 5445 2391 5503 2397
rect 8386 2388 8392 2440
rect 8444 2428 8450 2440
rect 11567 2428 11595 2459
rect 8444 2400 11595 2428
rect 8444 2388 8450 2400
rect 12342 2388 12348 2440
rect 12400 2428 12406 2440
rect 12713 2431 12771 2437
rect 12713 2428 12725 2431
rect 12400 2400 12725 2428
rect 12400 2388 12406 2400
rect 12713 2397 12725 2400
rect 12759 2428 12771 2431
rect 14001 2431 14059 2437
rect 14001 2428 14013 2431
rect 12759 2400 14013 2428
rect 12759 2397 12771 2400
rect 12713 2391 12771 2397
rect 14001 2397 14013 2400
rect 14047 2397 14059 2431
rect 14200 2428 14228 2459
rect 15286 2456 15292 2468
rect 15344 2496 15350 2508
rect 15508 2499 15566 2505
rect 15508 2496 15520 2499
rect 15344 2468 15520 2496
rect 15344 2456 15350 2468
rect 15508 2465 15520 2468
rect 15554 2496 15566 2499
rect 15933 2499 15991 2505
rect 15933 2496 15945 2499
rect 15554 2468 15945 2496
rect 15554 2465 15566 2468
rect 15508 2459 15566 2465
rect 15933 2465 15945 2468
rect 15979 2465 15991 2499
rect 15933 2459 15991 2465
rect 16485 2499 16543 2505
rect 16485 2465 16497 2499
rect 16531 2496 16543 2499
rect 17788 2496 17816 2527
rect 19058 2524 19064 2536
rect 19116 2524 19122 2576
rect 19150 2524 19156 2576
rect 19208 2564 19214 2576
rect 20070 2564 20076 2576
rect 19208 2536 19253 2564
rect 20031 2536 20076 2564
rect 19208 2524 19214 2536
rect 20070 2524 20076 2536
rect 20128 2524 20134 2576
rect 16531 2468 17816 2496
rect 16531 2465 16543 2468
rect 16485 2459 16543 2465
rect 20438 2456 20444 2508
rect 20496 2496 20502 2508
rect 21177 2499 21235 2505
rect 21177 2496 21189 2499
rect 20496 2468 21189 2496
rect 20496 2456 20502 2468
rect 21177 2465 21189 2468
rect 21223 2496 21235 2499
rect 21729 2499 21787 2505
rect 21729 2496 21741 2499
rect 21223 2468 21741 2496
rect 21223 2465 21235 2468
rect 21177 2459 21235 2465
rect 21729 2465 21741 2468
rect 21775 2465 21787 2499
rect 21729 2459 21787 2465
rect 14274 2428 14280 2440
rect 14187 2400 14280 2428
rect 14001 2391 14059 2397
rect 14274 2388 14280 2400
rect 14332 2428 14338 2440
rect 14332 2400 14872 2428
rect 14332 2388 14338 2400
rect 7558 2360 7564 2372
rect 4764 2332 5028 2360
rect 5368 2332 7564 2360
rect 4764 2320 4770 2332
rect 5368 2292 5396 2332
rect 7558 2320 7564 2332
rect 7616 2320 7622 2372
rect 13262 2360 13268 2372
rect 13223 2332 13268 2360
rect 13262 2320 13268 2332
rect 13320 2320 13326 2372
rect 14844 2369 14872 2400
rect 15102 2388 15108 2440
rect 15160 2428 15166 2440
rect 18785 2431 18843 2437
rect 18785 2428 18797 2431
rect 15160 2400 18797 2428
rect 15160 2388 15166 2400
rect 18785 2397 18797 2400
rect 18831 2428 18843 2431
rect 19058 2428 19064 2440
rect 18831 2400 19064 2428
rect 18831 2397 18843 2400
rect 18785 2391 18843 2397
rect 19058 2388 19064 2400
rect 19116 2388 19122 2440
rect 19337 2431 19395 2437
rect 19337 2428 19349 2431
rect 19168 2400 19349 2428
rect 14369 2363 14427 2369
rect 14369 2360 14381 2363
rect 13786 2332 14381 2360
rect 4448 2264 5396 2292
rect 1581 2255 1639 2261
rect 8018 2252 8024 2304
rect 8076 2292 8082 2304
rect 8297 2295 8355 2301
rect 8297 2292 8309 2295
rect 8076 2264 8309 2292
rect 8076 2252 8082 2264
rect 8297 2261 8309 2264
rect 8343 2292 8355 2295
rect 12434 2292 12440 2304
rect 8343 2264 12440 2292
rect 8343 2261 8355 2264
rect 8297 2255 8355 2261
rect 12434 2252 12440 2264
rect 12492 2252 12498 2304
rect 12710 2252 12716 2304
rect 12768 2292 12774 2304
rect 13786 2292 13814 2332
rect 14369 2329 14381 2332
rect 14415 2329 14427 2363
rect 14369 2323 14427 2329
rect 14829 2363 14887 2369
rect 14829 2329 14841 2363
rect 14875 2360 14887 2363
rect 18230 2360 18236 2372
rect 14875 2332 18236 2360
rect 14875 2329 14887 2332
rect 14829 2323 14887 2329
rect 18230 2320 18236 2332
rect 18288 2320 18294 2372
rect 18598 2320 18604 2372
rect 18656 2360 18662 2372
rect 19168 2360 19196 2400
rect 19337 2397 19349 2400
rect 19383 2397 19395 2431
rect 19337 2391 19395 2397
rect 21361 2363 21419 2369
rect 21361 2360 21373 2363
rect 18656 2332 19196 2360
rect 19996 2332 21373 2360
rect 18656 2320 18662 2332
rect 12768 2264 13814 2292
rect 12768 2252 12774 2264
rect 18874 2252 18880 2304
rect 18932 2292 18938 2304
rect 19996 2292 20024 2332
rect 21361 2329 21373 2332
rect 21407 2329 21419 2363
rect 21361 2323 21419 2329
rect 18932 2264 20024 2292
rect 18932 2252 18938 2264
rect 1104 2202 22816 2224
rect 1104 2150 4982 2202
rect 5034 2150 5046 2202
rect 5098 2150 5110 2202
rect 5162 2150 5174 2202
rect 5226 2150 12982 2202
rect 13034 2150 13046 2202
rect 13098 2150 13110 2202
rect 13162 2150 13174 2202
rect 13226 2150 20982 2202
rect 21034 2150 21046 2202
rect 21098 2150 21110 2202
rect 21162 2150 21174 2202
rect 21226 2150 22816 2202
rect 1104 2128 22816 2150
rect 11974 1708 11980 1760
rect 12032 1748 12038 1760
rect 17034 1748 17040 1760
rect 12032 1720 17040 1748
rect 12032 1708 12038 1720
rect 17034 1708 17040 1720
rect 17092 1708 17098 1760
rect 13814 76 13820 128
rect 13872 116 13878 128
rect 14458 116 14464 128
rect 13872 88 14464 116
rect 13872 76 13878 88
rect 14458 76 14464 88
rect 14516 76 14522 128
<< via1 >>
rect 22100 23536 22152 23588
rect 23296 23536 23348 23588
rect 4982 21734 5034 21786
rect 5046 21734 5098 21786
rect 5110 21734 5162 21786
rect 5174 21734 5226 21786
rect 12982 21734 13034 21786
rect 13046 21734 13098 21786
rect 13110 21734 13162 21786
rect 13174 21734 13226 21786
rect 20982 21734 21034 21786
rect 21046 21734 21098 21786
rect 21110 21734 21162 21786
rect 21174 21734 21226 21786
rect 8982 21190 9034 21242
rect 9046 21190 9098 21242
rect 9110 21190 9162 21242
rect 9174 21190 9226 21242
rect 16982 21190 17034 21242
rect 17046 21190 17098 21242
rect 17110 21190 17162 21242
rect 17174 21190 17226 21242
rect 572 21088 624 21140
rect 6460 21088 6512 21140
rect 11428 21088 11480 21140
rect 11060 20952 11112 21004
rect 15016 20952 15068 21004
rect 8668 20791 8720 20800
rect 8668 20757 8677 20791
rect 8677 20757 8711 20791
rect 8711 20757 8720 20791
rect 8668 20748 8720 20757
rect 13728 20748 13780 20800
rect 4982 20646 5034 20698
rect 5046 20646 5098 20698
rect 5110 20646 5162 20698
rect 5174 20646 5226 20698
rect 12982 20646 13034 20698
rect 13046 20646 13098 20698
rect 13110 20646 13162 20698
rect 13174 20646 13226 20698
rect 20982 20646 21034 20698
rect 21046 20646 21098 20698
rect 21110 20646 21162 20698
rect 21174 20646 21226 20698
rect 4344 20544 4396 20596
rect 1860 20383 1912 20392
rect 1860 20349 1869 20383
rect 1869 20349 1903 20383
rect 1903 20349 1912 20383
rect 1860 20340 1912 20349
rect 2228 20340 2280 20392
rect 3700 20340 3752 20392
rect 8392 20544 8444 20596
rect 10140 20544 10192 20596
rect 14096 20587 14148 20596
rect 14096 20553 14105 20587
rect 14105 20553 14139 20587
rect 14139 20553 14148 20587
rect 14096 20544 14148 20553
rect 15016 20544 15068 20596
rect 8668 20451 8720 20460
rect 8668 20417 8677 20451
rect 8677 20417 8711 20451
rect 8711 20417 8720 20451
rect 8668 20408 8720 20417
rect 6460 20272 6512 20324
rect 2504 20204 2556 20256
rect 2780 20204 2832 20256
rect 3700 20204 3752 20256
rect 7380 20204 7432 20256
rect 7840 20204 7892 20256
rect 8760 20315 8812 20324
rect 8760 20281 8769 20315
rect 8769 20281 8803 20315
rect 8803 20281 8812 20315
rect 8760 20272 8812 20281
rect 9312 20315 9364 20324
rect 9312 20281 9321 20315
rect 9321 20281 9355 20315
rect 9355 20281 9364 20315
rect 9312 20272 9364 20281
rect 14096 20340 14148 20392
rect 16396 20544 16448 20596
rect 19064 20544 19116 20596
rect 21456 20587 21508 20596
rect 21456 20553 21465 20587
rect 21465 20553 21499 20587
rect 21499 20553 21508 20587
rect 21456 20544 21508 20553
rect 21456 20340 21508 20392
rect 11060 20247 11112 20256
rect 11060 20213 11069 20247
rect 11069 20213 11103 20247
rect 11103 20213 11112 20247
rect 11060 20204 11112 20213
rect 13820 20204 13872 20256
rect 15384 20204 15436 20256
rect 18604 20204 18656 20256
rect 18696 20204 18748 20256
rect 8982 20102 9034 20154
rect 9046 20102 9098 20154
rect 9110 20102 9162 20154
rect 9174 20102 9226 20154
rect 16982 20102 17034 20154
rect 17046 20102 17098 20154
rect 17110 20102 17162 20154
rect 17174 20102 17226 20154
rect 1584 20043 1636 20052
rect 1584 20009 1593 20043
rect 1593 20009 1627 20043
rect 1627 20009 1636 20043
rect 1584 20000 1636 20009
rect 8668 20000 8720 20052
rect 13544 20000 13596 20052
rect 112 19932 164 19984
rect 8760 19932 8812 19984
rect 9772 19932 9824 19984
rect 15476 19975 15528 19984
rect 15476 19941 15485 19975
rect 15485 19941 15519 19975
rect 15519 19941 15528 19975
rect 15476 19932 15528 19941
rect 2136 19907 2188 19916
rect 2136 19873 2154 19907
rect 2154 19873 2188 19907
rect 2136 19864 2188 19873
rect 3056 19864 3108 19916
rect 7380 19907 7432 19916
rect 7380 19873 7389 19907
rect 7389 19873 7423 19907
rect 7423 19873 7432 19907
rect 7380 19864 7432 19873
rect 8484 19907 8536 19916
rect 8484 19873 8528 19907
rect 8528 19873 8536 19907
rect 8484 19864 8536 19873
rect 12716 19864 12768 19916
rect 16948 19907 17000 19916
rect 16948 19873 16966 19907
rect 16966 19873 17000 19907
rect 16948 19864 17000 19873
rect 17684 19864 17736 19916
rect 21180 19864 21232 19916
rect 9956 19839 10008 19848
rect 9956 19805 9965 19839
rect 9965 19805 9999 19839
rect 9999 19805 10008 19839
rect 9956 19796 10008 19805
rect 10140 19796 10192 19848
rect 10416 19796 10468 19848
rect 13728 19796 13780 19848
rect 14280 19839 14332 19848
rect 14280 19805 14289 19839
rect 14289 19805 14323 19839
rect 14323 19805 14332 19839
rect 14280 19796 14332 19805
rect 15384 19839 15436 19848
rect 15384 19805 15393 19839
rect 15393 19805 15427 19839
rect 15427 19805 15436 19839
rect 15384 19796 15436 19805
rect 2044 19660 2096 19712
rect 6828 19703 6880 19712
rect 6828 19669 6837 19703
rect 6837 19669 6871 19703
rect 6871 19669 6880 19703
rect 6828 19660 6880 19669
rect 8852 19660 8904 19712
rect 13360 19660 13412 19712
rect 16856 19660 16908 19712
rect 17408 19660 17460 19712
rect 4982 19558 5034 19610
rect 5046 19558 5098 19610
rect 5110 19558 5162 19610
rect 5174 19558 5226 19610
rect 12982 19558 13034 19610
rect 13046 19558 13098 19610
rect 13110 19558 13162 19610
rect 13174 19558 13226 19610
rect 20982 19558 21034 19610
rect 21046 19558 21098 19610
rect 21110 19558 21162 19610
rect 21174 19558 21226 19610
rect 2136 19499 2188 19508
rect 2136 19465 2145 19499
rect 2145 19465 2179 19499
rect 2179 19465 2188 19499
rect 2136 19456 2188 19465
rect 7380 19456 7432 19508
rect 8484 19499 8536 19508
rect 8484 19465 8493 19499
rect 8493 19465 8527 19499
rect 8527 19465 8536 19499
rect 8484 19456 8536 19465
rect 9772 19499 9824 19508
rect 9772 19465 9781 19499
rect 9781 19465 9815 19499
rect 9815 19465 9824 19499
rect 9772 19456 9824 19465
rect 15384 19456 15436 19508
rect 16948 19499 17000 19508
rect 16948 19465 16957 19499
rect 16957 19465 16991 19499
rect 16991 19465 17000 19499
rect 16948 19456 17000 19465
rect 7012 19388 7064 19440
rect 1584 19320 1636 19372
rect 6920 19320 6972 19372
rect 8852 19363 8904 19372
rect 8852 19329 8861 19363
rect 8861 19329 8895 19363
rect 8895 19329 8904 19363
rect 8852 19320 8904 19329
rect 10140 19320 10192 19372
rect 10416 19363 10468 19372
rect 10416 19329 10425 19363
rect 10425 19329 10459 19363
rect 10459 19329 10468 19363
rect 10416 19320 10468 19329
rect 14096 19388 14148 19440
rect 12072 19320 12124 19372
rect 14372 19363 14424 19372
rect 14372 19329 14381 19363
rect 14381 19329 14415 19363
rect 14415 19329 14424 19363
rect 14372 19320 14424 19329
rect 12716 19252 12768 19304
rect 13728 19252 13780 19304
rect 20720 19456 20772 19508
rect 21272 19456 21324 19508
rect 21732 19456 21784 19508
rect 22468 19456 22520 19508
rect 5264 19184 5316 19236
rect 6828 19116 6880 19168
rect 7012 19227 7064 19236
rect 7012 19193 7021 19227
rect 7021 19193 7055 19227
rect 7055 19193 7064 19227
rect 7012 19184 7064 19193
rect 8852 19184 8904 19236
rect 10508 19227 10560 19236
rect 10508 19193 10517 19227
rect 10517 19193 10551 19227
rect 10551 19193 10560 19227
rect 10508 19184 10560 19193
rect 14096 19227 14148 19236
rect 14096 19193 14105 19227
rect 14105 19193 14139 19227
rect 14139 19193 14148 19227
rect 14096 19184 14148 19193
rect 14188 19227 14240 19236
rect 14188 19193 14197 19227
rect 14197 19193 14231 19227
rect 14231 19193 14240 19227
rect 14188 19184 14240 19193
rect 15476 19184 15528 19236
rect 7380 19116 7432 19168
rect 12808 19116 12860 19168
rect 13452 19116 13504 19168
rect 13636 19116 13688 19168
rect 15384 19116 15436 19168
rect 18144 19116 18196 19168
rect 18972 19116 19024 19168
rect 20812 19116 20864 19168
rect 8982 19014 9034 19066
rect 9046 19014 9098 19066
rect 9110 19014 9162 19066
rect 9174 19014 9226 19066
rect 16982 19014 17034 19066
rect 17046 19014 17098 19066
rect 17110 19014 17162 19066
rect 17174 19014 17226 19066
rect 204 18912 256 18964
rect 14096 18912 14148 18964
rect 16304 18955 16356 18964
rect 16304 18921 16313 18955
rect 16313 18921 16347 18955
rect 16347 18921 16356 18955
rect 16304 18912 16356 18921
rect 16856 18912 16908 18964
rect 18144 18955 18196 18964
rect 5264 18887 5316 18896
rect 5264 18853 5273 18887
rect 5273 18853 5307 18887
rect 5307 18853 5316 18887
rect 5264 18844 5316 18853
rect 5448 18844 5500 18896
rect 6644 18844 6696 18896
rect 10508 18844 10560 18896
rect 12808 18844 12860 18896
rect 13452 18844 13504 18896
rect 13728 18844 13780 18896
rect 14372 18844 14424 18896
rect 15844 18844 15896 18896
rect 18144 18921 18153 18955
rect 18153 18921 18187 18955
rect 18187 18921 18196 18955
rect 18144 18912 18196 18921
rect 17040 18887 17092 18896
rect 17040 18853 17049 18887
rect 17049 18853 17083 18887
rect 17083 18853 17092 18887
rect 17040 18844 17092 18853
rect 1952 18776 2004 18828
rect 7564 18776 7616 18828
rect 8300 18819 8352 18828
rect 8300 18785 8344 18819
rect 8344 18785 8352 18819
rect 9956 18819 10008 18828
rect 8300 18776 8352 18785
rect 9956 18785 9965 18819
rect 9965 18785 9999 18819
rect 9999 18785 10008 18819
rect 9956 18776 10008 18785
rect 2504 18751 2556 18760
rect 2504 18717 2513 18751
rect 2513 18717 2547 18751
rect 2547 18717 2556 18751
rect 2504 18708 2556 18717
rect 6828 18751 6880 18760
rect 6828 18717 6837 18751
rect 6837 18717 6871 18751
rect 6871 18717 6880 18751
rect 6828 18708 6880 18717
rect 10876 18751 10928 18760
rect 6920 18640 6972 18692
rect 10876 18717 10885 18751
rect 10885 18717 10919 18751
rect 10919 18717 10928 18751
rect 10876 18708 10928 18717
rect 10692 18640 10744 18692
rect 13360 18708 13412 18760
rect 15476 18708 15528 18760
rect 15568 18708 15620 18760
rect 16672 18708 16724 18760
rect 17224 18751 17276 18760
rect 17224 18717 17233 18751
rect 17233 18717 17267 18751
rect 17267 18717 17276 18751
rect 17224 18708 17276 18717
rect 8576 18572 8628 18624
rect 8852 18615 8904 18624
rect 8852 18581 8861 18615
rect 8861 18581 8895 18615
rect 8895 18581 8904 18615
rect 8852 18572 8904 18581
rect 10508 18572 10560 18624
rect 14188 18572 14240 18624
rect 14740 18572 14792 18624
rect 4982 18470 5034 18522
rect 5046 18470 5098 18522
rect 5110 18470 5162 18522
rect 5174 18470 5226 18522
rect 12982 18470 13034 18522
rect 13046 18470 13098 18522
rect 13110 18470 13162 18522
rect 13174 18470 13226 18522
rect 20982 18470 21034 18522
rect 21046 18470 21098 18522
rect 21110 18470 21162 18522
rect 21174 18470 21226 18522
rect 1952 18411 2004 18420
rect 1952 18377 1961 18411
rect 1961 18377 1995 18411
rect 1995 18377 2004 18411
rect 1952 18368 2004 18377
rect 5356 18368 5408 18420
rect 6644 18411 6696 18420
rect 6644 18377 6653 18411
rect 6653 18377 6687 18411
rect 6687 18377 6696 18411
rect 6644 18368 6696 18377
rect 8300 18411 8352 18420
rect 8300 18377 8309 18411
rect 8309 18377 8343 18411
rect 8343 18377 8352 18411
rect 8300 18368 8352 18377
rect 16856 18368 16908 18420
rect 5448 18300 5500 18352
rect 9312 18343 9364 18352
rect 9312 18309 9321 18343
rect 9321 18309 9355 18343
rect 9355 18309 9364 18343
rect 9312 18300 9364 18309
rect 10876 18300 10928 18352
rect 6920 18275 6972 18284
rect 6920 18241 6929 18275
rect 6929 18241 6963 18275
rect 6963 18241 6972 18275
rect 6920 18232 6972 18241
rect 8576 18232 8628 18284
rect 2320 18164 2372 18216
rect 10968 18232 11020 18284
rect 10692 18164 10744 18216
rect 12072 18232 12124 18284
rect 12532 18275 12584 18284
rect 12532 18241 12541 18275
rect 12541 18241 12575 18275
rect 12575 18241 12584 18275
rect 12532 18232 12584 18241
rect 15568 18300 15620 18352
rect 15936 18300 15988 18352
rect 17040 18343 17092 18352
rect 17040 18309 17049 18343
rect 17049 18309 17083 18343
rect 17083 18309 17092 18343
rect 17040 18300 17092 18309
rect 18236 18300 18288 18352
rect 15384 18232 15436 18284
rect 16304 18232 16356 18284
rect 17224 18232 17276 18284
rect 18144 18275 18196 18284
rect 18144 18241 18153 18275
rect 18153 18241 18187 18275
rect 18187 18241 18196 18275
rect 18144 18232 18196 18241
rect 112 18028 164 18080
rect 2780 18028 2832 18080
rect 4528 18071 4580 18080
rect 4528 18037 4537 18071
rect 4537 18037 4571 18071
rect 4571 18037 4580 18071
rect 4528 18028 4580 18037
rect 6276 18071 6328 18080
rect 6276 18037 6285 18071
rect 6285 18037 6319 18071
rect 6319 18037 6328 18071
rect 6276 18028 6328 18037
rect 7656 18096 7708 18148
rect 8852 18139 8904 18148
rect 8852 18105 8861 18139
rect 8861 18105 8895 18139
rect 8895 18105 8904 18139
rect 8852 18096 8904 18105
rect 9864 18096 9916 18148
rect 10508 18028 10560 18080
rect 10784 18028 10836 18080
rect 10968 18139 11020 18148
rect 10968 18105 10977 18139
rect 10977 18105 11011 18139
rect 11011 18105 11020 18139
rect 10968 18096 11020 18105
rect 11152 18096 11204 18148
rect 11244 18096 11296 18148
rect 14556 18139 14608 18148
rect 12164 18071 12216 18080
rect 12164 18037 12173 18071
rect 12173 18037 12207 18071
rect 12207 18037 12216 18071
rect 14556 18105 14565 18139
rect 14565 18105 14599 18139
rect 14599 18105 14608 18139
rect 14556 18096 14608 18105
rect 13452 18071 13504 18080
rect 12164 18028 12216 18037
rect 13452 18037 13461 18071
rect 13461 18037 13495 18071
rect 13495 18037 13504 18071
rect 13452 18028 13504 18037
rect 15844 18071 15896 18080
rect 15844 18037 15853 18071
rect 15853 18037 15887 18071
rect 15887 18037 15896 18071
rect 15844 18028 15896 18037
rect 17592 18028 17644 18080
rect 8982 17926 9034 17978
rect 9046 17926 9098 17978
rect 9110 17926 9162 17978
rect 9174 17926 9226 17978
rect 16982 17926 17034 17978
rect 17046 17926 17098 17978
rect 17110 17926 17162 17978
rect 17174 17926 17226 17978
rect 6276 17824 6328 17876
rect 6920 17824 6972 17876
rect 8576 17824 8628 17876
rect 10968 17824 11020 17876
rect 11152 17824 11204 17876
rect 12532 17867 12584 17876
rect 12532 17833 12541 17867
rect 12541 17833 12575 17867
rect 12575 17833 12584 17867
rect 12532 17824 12584 17833
rect 12808 17824 12860 17876
rect 15476 17867 15528 17876
rect 15476 17833 15485 17867
rect 15485 17833 15519 17867
rect 15519 17833 15528 17867
rect 15476 17824 15528 17833
rect 5632 17756 5684 17808
rect 6828 17756 6880 17808
rect 15936 17756 15988 17808
rect 17592 17756 17644 17808
rect 2228 17731 2280 17740
rect 2228 17697 2237 17731
rect 2237 17697 2271 17731
rect 2271 17697 2280 17731
rect 2228 17688 2280 17697
rect 4712 17688 4764 17740
rect 8024 17731 8076 17740
rect 8024 17697 8033 17731
rect 8033 17697 8067 17731
rect 8067 17697 8076 17731
rect 8024 17688 8076 17697
rect 8484 17731 8536 17740
rect 8484 17697 8493 17731
rect 8493 17697 8527 17731
rect 8527 17697 8536 17731
rect 8484 17688 8536 17697
rect 12716 17688 12768 17740
rect 13544 17731 13596 17740
rect 13544 17697 13553 17731
rect 13553 17697 13587 17731
rect 13587 17697 13596 17731
rect 13544 17688 13596 17697
rect 4620 17663 4672 17672
rect 4620 17629 4629 17663
rect 4629 17629 4663 17663
rect 4663 17629 4672 17663
rect 4620 17620 4672 17629
rect 6092 17620 6144 17672
rect 8576 17663 8628 17672
rect 8576 17629 8585 17663
rect 8585 17629 8619 17663
rect 8619 17629 8628 17663
rect 8576 17620 8628 17629
rect 10692 17663 10744 17672
rect 10692 17629 10701 17663
rect 10701 17629 10735 17663
rect 10735 17629 10744 17663
rect 10692 17620 10744 17629
rect 13912 17620 13964 17672
rect 15200 17620 15252 17672
rect 17316 17663 17368 17672
rect 17316 17629 17325 17663
rect 17325 17629 17359 17663
rect 17359 17629 17368 17663
rect 17316 17620 17368 17629
rect 11612 17552 11664 17604
rect 17868 17595 17920 17604
rect 17868 17561 17877 17595
rect 17877 17561 17911 17595
rect 17911 17561 17920 17595
rect 17868 17552 17920 17561
rect 1952 17527 2004 17536
rect 1952 17493 1961 17527
rect 1961 17493 1995 17527
rect 1995 17493 2004 17527
rect 1952 17484 2004 17493
rect 7104 17484 7156 17536
rect 10600 17484 10652 17536
rect 18328 17527 18380 17536
rect 18328 17493 18337 17527
rect 18337 17493 18371 17527
rect 18371 17493 18380 17527
rect 18328 17484 18380 17493
rect 4982 17382 5034 17434
rect 5046 17382 5098 17434
rect 5110 17382 5162 17434
rect 5174 17382 5226 17434
rect 12982 17382 13034 17434
rect 13046 17382 13098 17434
rect 13110 17382 13162 17434
rect 13174 17382 13226 17434
rect 20982 17382 21034 17434
rect 21046 17382 21098 17434
rect 21110 17382 21162 17434
rect 21174 17382 21226 17434
rect 2504 17280 2556 17332
rect 7012 17280 7064 17332
rect 8484 17280 8536 17332
rect 9772 17280 9824 17332
rect 12164 17280 12216 17332
rect 13544 17280 13596 17332
rect 14556 17280 14608 17332
rect 15936 17280 15988 17332
rect 17316 17323 17368 17332
rect 17316 17289 17325 17323
rect 17325 17289 17359 17323
rect 17359 17289 17368 17323
rect 17316 17280 17368 17289
rect 21272 17280 21324 17332
rect 8024 17212 8076 17264
rect 12716 17255 12768 17264
rect 12716 17221 12725 17255
rect 12725 17221 12759 17255
rect 12759 17221 12768 17255
rect 12716 17212 12768 17221
rect 2320 17187 2372 17196
rect 2320 17153 2329 17187
rect 2329 17153 2363 17187
rect 2363 17153 2372 17187
rect 2320 17144 2372 17153
rect 8576 17187 8628 17196
rect 8576 17153 8585 17187
rect 8585 17153 8619 17187
rect 8619 17153 8628 17187
rect 8576 17144 8628 17153
rect 10692 17144 10744 17196
rect 13912 17187 13964 17196
rect 13912 17153 13921 17187
rect 13921 17153 13955 17187
rect 13955 17153 13964 17187
rect 13912 17144 13964 17153
rect 18236 17187 18288 17196
rect 18236 17153 18245 17187
rect 18245 17153 18279 17187
rect 18279 17153 18288 17187
rect 18236 17144 18288 17153
rect 18696 17187 18748 17196
rect 18696 17153 18705 17187
rect 18705 17153 18739 17187
rect 18739 17153 18748 17187
rect 18696 17144 18748 17153
rect 2872 17076 2924 17128
rect 4252 17119 4304 17128
rect 4252 17085 4261 17119
rect 4261 17085 4295 17119
rect 4295 17085 4304 17119
rect 4252 17076 4304 17085
rect 4712 17076 4764 17128
rect 6552 17119 6604 17128
rect 6552 17085 6561 17119
rect 6561 17085 6595 17119
rect 6595 17085 6604 17119
rect 6552 17076 6604 17085
rect 7104 17119 7156 17128
rect 7104 17085 7113 17119
rect 7113 17085 7147 17119
rect 7147 17085 7156 17119
rect 7104 17076 7156 17085
rect 7196 17076 7248 17128
rect 10600 17076 10652 17128
rect 20812 17076 20864 17128
rect 1952 17008 2004 17060
rect 5632 17051 5684 17060
rect 5632 17017 5641 17051
rect 5641 17017 5675 17051
rect 5675 17017 5684 17051
rect 5632 17008 5684 17017
rect 6092 17051 6144 17060
rect 6092 17017 6101 17051
rect 6101 17017 6135 17051
rect 6135 17017 6144 17051
rect 6092 17008 6144 17017
rect 2964 16983 3016 16992
rect 2964 16949 2973 16983
rect 2973 16949 3007 16983
rect 3007 16949 3016 16983
rect 2964 16940 3016 16949
rect 3516 16940 3568 16992
rect 4344 16940 4396 16992
rect 8392 16983 8444 16992
rect 8392 16949 8401 16983
rect 8401 16949 8435 16983
rect 8435 16949 8444 16983
rect 8392 16940 8444 16949
rect 13544 17008 13596 17060
rect 13820 17008 13872 17060
rect 16120 17051 16172 17060
rect 16120 17017 16129 17051
rect 16129 17017 16163 17051
rect 16163 17017 16172 17051
rect 16120 17008 16172 17017
rect 10968 16940 11020 16992
rect 13912 16940 13964 16992
rect 15200 16983 15252 16992
rect 15200 16949 15209 16983
rect 15209 16949 15243 16983
rect 15243 16949 15252 16983
rect 15200 16940 15252 16949
rect 15844 16983 15896 16992
rect 15844 16949 15853 16983
rect 15853 16949 15887 16983
rect 15887 16949 15896 16983
rect 17868 17008 17920 17060
rect 18328 17051 18380 17060
rect 18328 17017 18337 17051
rect 18337 17017 18371 17051
rect 18371 17017 18380 17051
rect 18328 17008 18380 17017
rect 17592 16983 17644 16992
rect 15844 16940 15896 16949
rect 17592 16949 17601 16983
rect 17601 16949 17635 16983
rect 17635 16949 17644 16983
rect 17592 16940 17644 16949
rect 8982 16838 9034 16890
rect 9046 16838 9098 16890
rect 9110 16838 9162 16890
rect 9174 16838 9226 16890
rect 16982 16838 17034 16890
rect 17046 16838 17098 16890
rect 17110 16838 17162 16890
rect 17174 16838 17226 16890
rect 1952 16736 2004 16788
rect 4252 16736 4304 16788
rect 5448 16736 5500 16788
rect 6736 16736 6788 16788
rect 8576 16779 8628 16788
rect 8576 16745 8585 16779
rect 8585 16745 8619 16779
rect 8619 16745 8628 16779
rect 8576 16736 8628 16745
rect 11704 16779 11756 16788
rect 11704 16745 11713 16779
rect 11713 16745 11747 16779
rect 11747 16745 11756 16779
rect 11704 16736 11756 16745
rect 16120 16779 16172 16788
rect 16120 16745 16129 16779
rect 16129 16745 16163 16779
rect 16163 16745 16172 16779
rect 16120 16736 16172 16745
rect 18328 16736 18380 16788
rect 2228 16668 2280 16720
rect 2964 16668 3016 16720
rect 6552 16668 6604 16720
rect 7196 16668 7248 16720
rect 8392 16668 8444 16720
rect 10692 16668 10744 16720
rect 4160 16643 4212 16652
rect 4160 16609 4169 16643
rect 4169 16609 4203 16643
rect 4203 16609 4212 16643
rect 4160 16600 4212 16609
rect 4712 16600 4764 16652
rect 6092 16600 6144 16652
rect 7104 16600 7156 16652
rect 10324 16643 10376 16652
rect 10324 16609 10333 16643
rect 10333 16609 10367 16643
rect 10367 16609 10376 16643
rect 10324 16600 10376 16609
rect 10416 16600 10468 16652
rect 11612 16643 11664 16652
rect 11612 16609 11621 16643
rect 11621 16609 11655 16643
rect 11655 16609 11664 16643
rect 11612 16600 11664 16609
rect 11980 16600 12032 16652
rect 15200 16668 15252 16720
rect 17408 16668 17460 16720
rect 13268 16643 13320 16652
rect 13268 16609 13277 16643
rect 13277 16609 13311 16643
rect 13311 16609 13320 16643
rect 13268 16600 13320 16609
rect 13820 16643 13872 16652
rect 13820 16609 13829 16643
rect 13829 16609 13863 16643
rect 13863 16609 13872 16643
rect 13820 16600 13872 16609
rect 15384 16600 15436 16652
rect 2320 16575 2372 16584
rect 2320 16541 2329 16575
rect 2329 16541 2363 16575
rect 2363 16541 2372 16575
rect 2320 16532 2372 16541
rect 7564 16532 7616 16584
rect 14004 16575 14056 16584
rect 14004 16541 14013 16575
rect 14013 16541 14047 16575
rect 14047 16541 14056 16575
rect 14004 16532 14056 16541
rect 18236 16600 18288 16652
rect 17316 16575 17368 16584
rect 17316 16541 17325 16575
rect 17325 16541 17359 16575
rect 17359 16541 17368 16575
rect 17316 16532 17368 16541
rect 2412 16464 2464 16516
rect 4160 16464 4212 16516
rect 8024 16464 8076 16516
rect 10876 16464 10928 16516
rect 11060 16464 11112 16516
rect 16120 16464 16172 16516
rect 3884 16439 3936 16448
rect 3884 16405 3893 16439
rect 3893 16405 3927 16439
rect 3927 16405 3936 16439
rect 3884 16396 3936 16405
rect 6276 16396 6328 16448
rect 9312 16396 9364 16448
rect 4982 16294 5034 16346
rect 5046 16294 5098 16346
rect 5110 16294 5162 16346
rect 5174 16294 5226 16346
rect 12982 16294 13034 16346
rect 13046 16294 13098 16346
rect 13110 16294 13162 16346
rect 13174 16294 13226 16346
rect 20982 16294 21034 16346
rect 21046 16294 21098 16346
rect 21110 16294 21162 16346
rect 21174 16294 21226 16346
rect 112 16192 164 16244
rect 5356 16235 5408 16244
rect 3884 16167 3936 16176
rect 3884 16133 3893 16167
rect 3893 16133 3927 16167
rect 3927 16133 3936 16167
rect 3884 16124 3936 16133
rect 5356 16201 5365 16235
rect 5365 16201 5399 16235
rect 5399 16201 5408 16235
rect 5356 16192 5408 16201
rect 6644 16192 6696 16244
rect 9128 16192 9180 16244
rect 9772 16192 9824 16244
rect 10324 16192 10376 16244
rect 6092 16124 6144 16176
rect 8484 16124 8536 16176
rect 9404 16124 9456 16176
rect 10416 16124 10468 16176
rect 15844 16192 15896 16244
rect 16120 16235 16172 16244
rect 16120 16201 16129 16235
rect 16129 16201 16163 16235
rect 16163 16201 16172 16235
rect 16120 16192 16172 16201
rect 20812 16192 20864 16244
rect 18696 16167 18748 16176
rect 2044 16099 2096 16108
rect 2044 16065 2053 16099
rect 2053 16065 2087 16099
rect 2087 16065 2096 16099
rect 2044 16056 2096 16065
rect 2412 16099 2464 16108
rect 2412 16065 2421 16099
rect 2421 16065 2455 16099
rect 2455 16065 2464 16099
rect 2412 16056 2464 16065
rect 4160 16056 4212 16108
rect 4620 16056 4672 16108
rect 4344 15988 4396 16040
rect 8760 16056 8812 16108
rect 9312 16056 9364 16108
rect 1860 15895 1912 15904
rect 1860 15861 1869 15895
rect 1869 15861 1903 15895
rect 1903 15861 1912 15895
rect 3884 15920 3936 15972
rect 4620 15920 4672 15972
rect 7196 15988 7248 16040
rect 8392 15988 8444 16040
rect 10784 16031 10836 16040
rect 10784 15997 10793 16031
rect 10793 15997 10827 16031
rect 10827 15997 10836 16031
rect 10784 15988 10836 15997
rect 11612 15988 11664 16040
rect 13268 16056 13320 16108
rect 14004 16056 14056 16108
rect 7564 15963 7616 15972
rect 7564 15929 7573 15963
rect 7573 15929 7607 15963
rect 7607 15929 7616 15963
rect 7564 15920 7616 15929
rect 9128 15963 9180 15972
rect 9128 15929 9137 15963
rect 9137 15929 9171 15963
rect 9171 15929 9180 15963
rect 9128 15920 9180 15929
rect 9956 15920 10008 15972
rect 12256 15920 12308 15972
rect 15384 16031 15436 16040
rect 15384 15997 15393 16031
rect 15393 15997 15427 16031
rect 15427 15997 15436 16031
rect 15384 15988 15436 15997
rect 16120 15988 16172 16040
rect 18696 16133 18705 16167
rect 18705 16133 18739 16167
rect 18739 16133 18748 16167
rect 18696 16124 18748 16133
rect 17316 16056 17368 16108
rect 17868 16056 17920 16108
rect 16580 15988 16632 16040
rect 18236 15963 18288 15972
rect 18236 15929 18245 15963
rect 18245 15929 18279 15963
rect 18279 15929 18288 15963
rect 18236 15920 18288 15929
rect 1860 15852 1912 15861
rect 2596 15852 2648 15904
rect 2964 15895 3016 15904
rect 2964 15861 2973 15895
rect 2973 15861 3007 15895
rect 3007 15861 3016 15895
rect 2964 15852 3016 15861
rect 4436 15852 4488 15904
rect 6092 15895 6144 15904
rect 6092 15861 6101 15895
rect 6101 15861 6135 15895
rect 6135 15861 6144 15895
rect 6092 15852 6144 15861
rect 10600 15895 10652 15904
rect 10600 15861 10609 15895
rect 10609 15861 10643 15895
rect 10643 15861 10652 15895
rect 10600 15852 10652 15861
rect 12532 15895 12584 15904
rect 12532 15861 12541 15895
rect 12541 15861 12575 15895
rect 12575 15861 12584 15895
rect 12532 15852 12584 15861
rect 13268 15852 13320 15904
rect 13912 15852 13964 15904
rect 14464 15895 14516 15904
rect 14464 15861 14473 15895
rect 14473 15861 14507 15895
rect 14507 15861 14516 15895
rect 14464 15852 14516 15861
rect 15752 15895 15804 15904
rect 15752 15861 15761 15895
rect 15761 15861 15795 15895
rect 15795 15861 15804 15895
rect 15752 15852 15804 15861
rect 17316 15895 17368 15904
rect 17316 15861 17325 15895
rect 17325 15861 17359 15895
rect 17359 15861 17368 15895
rect 17316 15852 17368 15861
rect 17960 15852 18012 15904
rect 8982 15750 9034 15802
rect 9046 15750 9098 15802
rect 9110 15750 9162 15802
rect 9174 15750 9226 15802
rect 16982 15750 17034 15802
rect 17046 15750 17098 15802
rect 17110 15750 17162 15802
rect 17174 15750 17226 15802
rect 1860 15648 1912 15700
rect 2044 15648 2096 15700
rect 5356 15648 5408 15700
rect 3516 15580 3568 15632
rect 4252 15580 4304 15632
rect 4344 15623 4396 15632
rect 4344 15589 4353 15623
rect 4353 15589 4387 15623
rect 4387 15589 4396 15623
rect 4344 15580 4396 15589
rect 6276 15580 6328 15632
rect 7564 15648 7616 15700
rect 10416 15691 10468 15700
rect 10416 15657 10425 15691
rect 10425 15657 10459 15691
rect 10459 15657 10468 15691
rect 10416 15648 10468 15657
rect 11612 15691 11664 15700
rect 11612 15657 11621 15691
rect 11621 15657 11655 15691
rect 11655 15657 11664 15691
rect 11612 15648 11664 15657
rect 11980 15691 12032 15700
rect 11980 15657 11989 15691
rect 11989 15657 12023 15691
rect 12023 15657 12032 15691
rect 11980 15648 12032 15657
rect 14004 15648 14056 15700
rect 16580 15691 16632 15700
rect 16580 15657 16589 15691
rect 16589 15657 16623 15691
rect 16623 15657 16632 15691
rect 16580 15648 16632 15657
rect 18236 15648 18288 15700
rect 21456 15648 21508 15700
rect 7012 15580 7064 15632
rect 10324 15580 10376 15632
rect 14464 15580 14516 15632
rect 16856 15580 16908 15632
rect 17316 15580 17368 15632
rect 2504 15512 2556 15564
rect 8300 15512 8352 15564
rect 11704 15512 11756 15564
rect 12532 15512 12584 15564
rect 4252 15487 4304 15496
rect 4252 15453 4261 15487
rect 4261 15453 4295 15487
rect 4295 15453 4304 15487
rect 4252 15444 4304 15453
rect 7380 15487 7432 15496
rect 7380 15453 7389 15487
rect 7389 15453 7423 15487
rect 7423 15453 7432 15487
rect 7380 15444 7432 15453
rect 10784 15444 10836 15496
rect 15108 15512 15160 15564
rect 15752 15512 15804 15564
rect 20812 15512 20864 15564
rect 17500 15444 17552 15496
rect 4804 15419 4856 15428
rect 4804 15385 4813 15419
rect 4813 15385 4847 15419
rect 4847 15385 4856 15419
rect 4804 15376 4856 15385
rect 6092 15376 6144 15428
rect 10692 15376 10744 15428
rect 7932 15308 7984 15360
rect 8760 15351 8812 15360
rect 8760 15317 8769 15351
rect 8769 15317 8803 15351
rect 8803 15317 8812 15351
rect 8760 15308 8812 15317
rect 10508 15308 10560 15360
rect 12440 15308 12492 15360
rect 13452 15308 13504 15360
rect 13820 15308 13872 15360
rect 4982 15206 5034 15258
rect 5046 15206 5098 15258
rect 5110 15206 5162 15258
rect 5174 15206 5226 15258
rect 12982 15206 13034 15258
rect 13046 15206 13098 15258
rect 13110 15206 13162 15258
rect 13174 15206 13226 15258
rect 20982 15206 21034 15258
rect 21046 15206 21098 15258
rect 21110 15206 21162 15258
rect 21174 15206 21226 15258
rect 4344 15104 4396 15156
rect 4528 15104 4580 15156
rect 6276 15147 6328 15156
rect 2412 15079 2464 15088
rect 2412 15045 2421 15079
rect 2421 15045 2455 15079
rect 2455 15045 2464 15079
rect 2412 15036 2464 15045
rect 6276 15113 6285 15147
rect 6285 15113 6319 15147
rect 6319 15113 6328 15147
rect 6276 15104 6328 15113
rect 7012 15104 7064 15156
rect 11704 15104 11756 15156
rect 13636 15104 13688 15156
rect 14464 15104 14516 15156
rect 15108 15147 15160 15156
rect 15108 15113 15117 15147
rect 15117 15113 15151 15147
rect 15151 15113 15160 15147
rect 15108 15104 15160 15113
rect 17500 15147 17552 15156
rect 17500 15113 17509 15147
rect 17509 15113 17543 15147
rect 17543 15113 17552 15147
rect 17500 15104 17552 15113
rect 21272 15104 21324 15156
rect 4804 15036 4856 15088
rect 7380 15036 7432 15088
rect 7932 14968 7984 15020
rect 8760 14968 8812 15020
rect 13268 15036 13320 15088
rect 13820 15036 13872 15088
rect 15752 15036 15804 15088
rect 16212 15036 16264 15088
rect 11428 14968 11480 15020
rect 11980 14968 12032 15020
rect 9404 14900 9456 14952
rect 5356 14832 5408 14884
rect 7288 14875 7340 14884
rect 7288 14841 7297 14875
rect 7297 14841 7331 14875
rect 7331 14841 7340 14875
rect 7288 14832 7340 14841
rect 8300 14875 8352 14884
rect 8300 14841 8309 14875
rect 8309 14841 8343 14875
rect 8343 14841 8352 14875
rect 8300 14832 8352 14841
rect 8852 14832 8904 14884
rect 10508 14875 10560 14884
rect 10508 14841 10517 14875
rect 10517 14841 10551 14875
rect 10551 14841 10560 14875
rect 10508 14832 10560 14841
rect 10600 14832 10652 14884
rect 13452 14900 13504 14952
rect 15568 14943 15620 14952
rect 15568 14909 15577 14943
rect 15577 14909 15611 14943
rect 15611 14909 15620 14943
rect 15568 14900 15620 14909
rect 13636 14832 13688 14884
rect 16488 14832 16540 14884
rect 19340 14832 19392 14884
rect 20812 14832 20864 14884
rect 2504 14764 2556 14816
rect 3792 14807 3844 14816
rect 3792 14773 3801 14807
rect 3801 14773 3835 14807
rect 3835 14773 3844 14807
rect 3792 14764 3844 14773
rect 8760 14807 8812 14816
rect 8760 14773 8769 14807
rect 8769 14773 8803 14807
rect 8803 14773 8812 14807
rect 8760 14764 8812 14773
rect 10416 14764 10468 14816
rect 12716 14764 12768 14816
rect 12808 14764 12860 14816
rect 14740 14764 14792 14816
rect 16856 14764 16908 14816
rect 8982 14662 9034 14714
rect 9046 14662 9098 14714
rect 9110 14662 9162 14714
rect 9174 14662 9226 14714
rect 16982 14662 17034 14714
rect 17046 14662 17098 14714
rect 17110 14662 17162 14714
rect 17174 14662 17226 14714
rect 1952 14560 2004 14612
rect 2596 14603 2648 14612
rect 2596 14569 2605 14603
rect 2605 14569 2639 14603
rect 2639 14569 2648 14603
rect 2596 14560 2648 14569
rect 4252 14560 4304 14612
rect 7288 14560 7340 14612
rect 7932 14603 7984 14612
rect 7932 14569 7941 14603
rect 7941 14569 7975 14603
rect 7975 14569 7984 14603
rect 7932 14560 7984 14569
rect 9312 14560 9364 14612
rect 12532 14603 12584 14612
rect 12532 14569 12541 14603
rect 12541 14569 12575 14603
rect 12575 14569 12584 14603
rect 12532 14560 12584 14569
rect 15568 14560 15620 14612
rect 4804 14492 4856 14544
rect 5356 14492 5408 14544
rect 6736 14492 6788 14544
rect 9404 14492 9456 14544
rect 9864 14535 9916 14544
rect 9864 14501 9873 14535
rect 9873 14501 9907 14535
rect 9907 14501 9916 14535
rect 9864 14492 9916 14501
rect 10784 14535 10836 14544
rect 10784 14501 10793 14535
rect 10793 14501 10827 14535
rect 10827 14501 10836 14535
rect 10784 14492 10836 14501
rect 12440 14492 12492 14544
rect 15752 14492 15804 14544
rect 16856 14492 16908 14544
rect 3240 14356 3292 14408
rect 3884 14356 3936 14408
rect 6368 14424 6420 14476
rect 10692 14424 10744 14476
rect 11796 14424 11848 14476
rect 14096 14424 14148 14476
rect 15568 14424 15620 14476
rect 6828 14399 6880 14408
rect 6828 14365 6837 14399
rect 6837 14365 6871 14399
rect 6871 14365 6880 14399
rect 6828 14356 6880 14365
rect 8116 14399 8168 14408
rect 8116 14365 8125 14399
rect 8125 14365 8159 14399
rect 8159 14365 8168 14399
rect 8116 14356 8168 14365
rect 9772 14399 9824 14408
rect 7380 14288 7432 14340
rect 9772 14365 9781 14399
rect 9781 14365 9815 14399
rect 9815 14365 9824 14399
rect 9772 14356 9824 14365
rect 9956 14356 10008 14408
rect 10600 14356 10652 14408
rect 12164 14356 12216 14408
rect 12716 14399 12768 14408
rect 12716 14365 12725 14399
rect 12725 14365 12759 14399
rect 12759 14365 12768 14399
rect 12716 14356 12768 14365
rect 13544 14356 13596 14408
rect 14924 14356 14976 14408
rect 16488 14356 16540 14408
rect 4252 14263 4304 14272
rect 4252 14229 4261 14263
rect 4261 14229 4295 14263
rect 4295 14229 4304 14263
rect 4252 14220 4304 14229
rect 6276 14263 6328 14272
rect 6276 14229 6285 14263
rect 6285 14229 6319 14263
rect 6319 14229 6328 14263
rect 6276 14220 6328 14229
rect 6368 14220 6420 14272
rect 7656 14220 7708 14272
rect 13452 14220 13504 14272
rect 14648 14263 14700 14272
rect 14648 14229 14657 14263
rect 14657 14229 14691 14263
rect 14691 14229 14700 14263
rect 14648 14220 14700 14229
rect 16580 14220 16632 14272
rect 17592 14220 17644 14272
rect 4982 14118 5034 14170
rect 5046 14118 5098 14170
rect 5110 14118 5162 14170
rect 5174 14118 5226 14170
rect 12982 14118 13034 14170
rect 13046 14118 13098 14170
rect 13110 14118 13162 14170
rect 13174 14118 13226 14170
rect 20982 14118 21034 14170
rect 21046 14118 21098 14170
rect 21110 14118 21162 14170
rect 21174 14118 21226 14170
rect 2504 14059 2556 14068
rect 2504 14025 2513 14059
rect 2513 14025 2547 14059
rect 2547 14025 2556 14059
rect 2504 14016 2556 14025
rect 5356 14016 5408 14068
rect 6736 14016 6788 14068
rect 8116 14016 8168 14068
rect 8484 14016 8536 14068
rect 9864 14059 9916 14068
rect 9864 14025 9873 14059
rect 9873 14025 9907 14059
rect 9907 14025 9916 14059
rect 9864 14016 9916 14025
rect 11796 14059 11848 14068
rect 11796 14025 11805 14059
rect 11805 14025 11839 14059
rect 11839 14025 11848 14059
rect 11796 14016 11848 14025
rect 12256 14059 12308 14068
rect 12256 14025 12265 14059
rect 12265 14025 12299 14059
rect 12299 14025 12308 14059
rect 12256 14016 12308 14025
rect 6184 13948 6236 14000
rect 9404 13948 9456 14000
rect 4252 13923 4304 13932
rect 4252 13889 4261 13923
rect 4261 13889 4295 13923
rect 4295 13889 4304 13923
rect 4252 13880 4304 13889
rect 7380 13880 7432 13932
rect 7656 13923 7708 13932
rect 7656 13889 7665 13923
rect 7665 13889 7699 13923
rect 7699 13889 7708 13923
rect 7656 13880 7708 13889
rect 8760 13880 8812 13932
rect 10784 13880 10836 13932
rect 16856 13948 16908 14000
rect 13452 13923 13504 13932
rect 2044 13812 2096 13864
rect 1952 13787 2004 13796
rect 1952 13753 1968 13787
rect 1968 13753 2004 13787
rect 4436 13812 4488 13864
rect 1952 13744 2004 13753
rect 3240 13787 3292 13796
rect 3240 13753 3249 13787
rect 3249 13753 3283 13787
rect 3283 13753 3292 13787
rect 3240 13744 3292 13753
rect 10968 13812 11020 13864
rect 7288 13744 7340 13796
rect 4804 13676 4856 13728
rect 5632 13676 5684 13728
rect 6828 13676 6880 13728
rect 12624 13812 12676 13864
rect 13452 13889 13461 13923
rect 13461 13889 13495 13923
rect 13495 13889 13504 13923
rect 13452 13880 13504 13889
rect 14648 13923 14700 13932
rect 14648 13889 14657 13923
rect 14657 13889 14691 13923
rect 14691 13889 14700 13923
rect 14648 13880 14700 13889
rect 14924 13923 14976 13932
rect 14924 13889 14933 13923
rect 14933 13889 14967 13923
rect 14967 13889 14976 13923
rect 14924 13880 14976 13889
rect 16580 13880 16632 13932
rect 16672 13880 16724 13932
rect 11520 13787 11572 13796
rect 11520 13753 11529 13787
rect 11529 13753 11563 13787
rect 11563 13753 11572 13787
rect 11520 13744 11572 13753
rect 18328 13812 18380 13864
rect 10416 13676 10468 13728
rect 14096 13744 14148 13796
rect 14740 13787 14792 13796
rect 14740 13753 14749 13787
rect 14749 13753 14783 13787
rect 14783 13753 14792 13787
rect 14740 13744 14792 13753
rect 15936 13676 15988 13728
rect 16580 13787 16632 13796
rect 16580 13753 16589 13787
rect 16589 13753 16623 13787
rect 16623 13753 16632 13787
rect 16580 13744 16632 13753
rect 17500 13719 17552 13728
rect 17500 13685 17509 13719
rect 17509 13685 17543 13719
rect 17543 13685 17552 13719
rect 17500 13676 17552 13685
rect 8982 13574 9034 13626
rect 9046 13574 9098 13626
rect 9110 13574 9162 13626
rect 9174 13574 9226 13626
rect 16982 13574 17034 13626
rect 17046 13574 17098 13626
rect 17110 13574 17162 13626
rect 17174 13574 17226 13626
rect 112 13472 164 13524
rect 2780 13472 2832 13524
rect 4252 13515 4304 13524
rect 4252 13481 4261 13515
rect 4261 13481 4295 13515
rect 4295 13481 4304 13515
rect 4252 13472 4304 13481
rect 5632 13515 5684 13524
rect 5632 13481 5641 13515
rect 5641 13481 5675 13515
rect 5675 13481 5684 13515
rect 5632 13472 5684 13481
rect 6644 13472 6696 13524
rect 7288 13515 7340 13524
rect 7288 13481 7297 13515
rect 7297 13481 7331 13515
rect 7331 13481 7340 13515
rect 7288 13472 7340 13481
rect 7380 13472 7432 13524
rect 8116 13472 8168 13524
rect 8760 13472 8812 13524
rect 12164 13515 12216 13524
rect 12164 13481 12173 13515
rect 12173 13481 12207 13515
rect 12207 13481 12216 13515
rect 12164 13472 12216 13481
rect 12440 13515 12492 13524
rect 12440 13481 12449 13515
rect 12449 13481 12483 13515
rect 12483 13481 12492 13515
rect 12440 13472 12492 13481
rect 10692 13447 10744 13456
rect 10692 13413 10701 13447
rect 10701 13413 10735 13447
rect 10735 13413 10744 13447
rect 10692 13404 10744 13413
rect 11244 13447 11296 13456
rect 11244 13413 11253 13447
rect 11253 13413 11287 13447
rect 11287 13413 11296 13447
rect 11244 13404 11296 13413
rect 12716 13404 12768 13456
rect 13636 13472 13688 13524
rect 14740 13472 14792 13524
rect 16488 13515 16540 13524
rect 16488 13481 16497 13515
rect 16497 13481 16531 13515
rect 16531 13481 16540 13515
rect 16488 13472 16540 13481
rect 21088 13515 21140 13524
rect 16856 13404 16908 13456
rect 21088 13481 21097 13515
rect 21097 13481 21131 13515
rect 21131 13481 21140 13515
rect 21088 13472 21140 13481
rect 18880 13404 18932 13456
rect 1676 13336 1728 13388
rect 3148 13336 3200 13388
rect 3700 13336 3752 13388
rect 4712 13379 4764 13388
rect 4712 13345 4721 13379
rect 4721 13345 4755 13379
rect 4755 13345 4764 13379
rect 4712 13336 4764 13345
rect 8208 13336 8260 13388
rect 11520 13336 11572 13388
rect 13636 13336 13688 13388
rect 15200 13379 15252 13388
rect 15200 13345 15209 13379
rect 15209 13345 15243 13379
rect 15243 13345 15252 13379
rect 15200 13336 15252 13345
rect 20812 13336 20864 13388
rect 6368 13311 6420 13320
rect 6368 13277 6377 13311
rect 6377 13277 6411 13311
rect 6411 13277 6420 13311
rect 6368 13268 6420 13277
rect 10600 13311 10652 13320
rect 10600 13277 10609 13311
rect 10609 13277 10643 13311
rect 10643 13277 10652 13311
rect 10600 13268 10652 13277
rect 16672 13311 16724 13320
rect 16672 13277 16681 13311
rect 16681 13277 16715 13311
rect 16715 13277 16724 13311
rect 16672 13268 16724 13277
rect 18512 13311 18564 13320
rect 18512 13277 18521 13311
rect 18521 13277 18555 13311
rect 18555 13277 18564 13311
rect 18512 13268 18564 13277
rect 18696 13268 18748 13320
rect 10784 13200 10836 13252
rect 15752 13200 15804 13252
rect 1952 13175 2004 13184
rect 1952 13141 1961 13175
rect 1961 13141 1995 13175
rect 1995 13141 2004 13175
rect 1952 13132 2004 13141
rect 2044 13132 2096 13184
rect 2320 13175 2372 13184
rect 2320 13141 2329 13175
rect 2329 13141 2363 13175
rect 2363 13141 2372 13175
rect 2320 13132 2372 13141
rect 5356 13132 5408 13184
rect 9864 13175 9916 13184
rect 9864 13141 9873 13175
rect 9873 13141 9907 13175
rect 9907 13141 9916 13175
rect 9864 13132 9916 13141
rect 14004 13132 14056 13184
rect 14280 13175 14332 13184
rect 14280 13141 14289 13175
rect 14289 13141 14323 13175
rect 14323 13141 14332 13175
rect 14280 13132 14332 13141
rect 14740 13132 14792 13184
rect 15568 13132 15620 13184
rect 15844 13175 15896 13184
rect 15844 13141 15853 13175
rect 15853 13141 15887 13175
rect 15887 13141 15896 13175
rect 15844 13132 15896 13141
rect 4982 13030 5034 13082
rect 5046 13030 5098 13082
rect 5110 13030 5162 13082
rect 5174 13030 5226 13082
rect 12982 13030 13034 13082
rect 13046 13030 13098 13082
rect 13110 13030 13162 13082
rect 13174 13030 13226 13082
rect 20982 13030 21034 13082
rect 21046 13030 21098 13082
rect 21110 13030 21162 13082
rect 21174 13030 21226 13082
rect 6276 12928 6328 12980
rect 9864 12928 9916 12980
rect 10600 12928 10652 12980
rect 11428 12928 11480 12980
rect 13636 12971 13688 12980
rect 13636 12937 13645 12971
rect 13645 12937 13679 12971
rect 13679 12937 13688 12971
rect 13636 12928 13688 12937
rect 14004 12971 14056 12980
rect 14004 12937 14013 12971
rect 14013 12937 14047 12971
rect 14047 12937 14056 12971
rect 14004 12928 14056 12937
rect 17500 12928 17552 12980
rect 18880 12971 18932 12980
rect 18880 12937 18889 12971
rect 18889 12937 18923 12971
rect 18923 12937 18932 12971
rect 18880 12928 18932 12937
rect 4436 12860 4488 12912
rect 6644 12860 6696 12912
rect 8852 12860 8904 12912
rect 2596 12724 2648 12776
rect 3792 12724 3844 12776
rect 4160 12767 4212 12776
rect 4160 12733 4204 12767
rect 4204 12733 4212 12767
rect 4160 12724 4212 12733
rect 5356 12767 5408 12776
rect 5356 12733 5365 12767
rect 5365 12733 5399 12767
rect 5399 12733 5408 12767
rect 5356 12724 5408 12733
rect 4712 12656 4764 12708
rect 6368 12724 6420 12776
rect 6644 12724 6696 12776
rect 8208 12767 8260 12776
rect 8208 12733 8217 12767
rect 8217 12733 8251 12767
rect 8251 12733 8260 12767
rect 8208 12724 8260 12733
rect 9128 12767 9180 12776
rect 9128 12733 9137 12767
rect 9137 12733 9171 12767
rect 9171 12733 9180 12767
rect 9128 12724 9180 12733
rect 9588 12767 9640 12776
rect 9588 12733 9597 12767
rect 9597 12733 9631 12767
rect 9631 12733 9640 12767
rect 9588 12724 9640 12733
rect 6828 12699 6880 12708
rect 2504 12631 2556 12640
rect 2504 12597 2513 12631
rect 2513 12597 2547 12631
rect 2547 12597 2556 12631
rect 2504 12588 2556 12597
rect 3148 12631 3200 12640
rect 3148 12597 3157 12631
rect 3157 12597 3191 12631
rect 3191 12597 3200 12631
rect 3148 12588 3200 12597
rect 3700 12631 3752 12640
rect 3700 12597 3709 12631
rect 3709 12597 3743 12631
rect 3743 12597 3752 12631
rect 3700 12588 3752 12597
rect 6828 12665 6837 12699
rect 6837 12665 6871 12699
rect 6871 12665 6880 12699
rect 6828 12656 6880 12665
rect 9312 12656 9364 12708
rect 10324 12724 10376 12776
rect 18512 12860 18564 12912
rect 20812 12860 20864 12912
rect 12808 12792 12860 12844
rect 14556 12835 14608 12844
rect 14556 12801 14565 12835
rect 14565 12801 14599 12835
rect 14599 12801 14608 12835
rect 14556 12792 14608 12801
rect 16672 12792 16724 12844
rect 11796 12724 11848 12776
rect 15384 12724 15436 12776
rect 15752 12767 15804 12776
rect 15752 12733 15761 12767
rect 15761 12733 15795 12767
rect 15795 12733 15804 12767
rect 15752 12724 15804 12733
rect 15844 12724 15896 12776
rect 14280 12699 14332 12708
rect 14280 12665 14289 12699
rect 14289 12665 14323 12699
rect 14323 12665 14332 12699
rect 14280 12656 14332 12665
rect 18696 12724 18748 12776
rect 20720 12724 20772 12776
rect 9680 12588 9732 12640
rect 9864 12631 9916 12640
rect 9864 12597 9873 12631
rect 9873 12597 9907 12631
rect 9907 12597 9916 12631
rect 9864 12588 9916 12597
rect 10692 12631 10744 12640
rect 10692 12597 10701 12631
rect 10701 12597 10735 12631
rect 10735 12597 10744 12631
rect 10692 12588 10744 12597
rect 12716 12588 12768 12640
rect 13360 12631 13412 12640
rect 13360 12597 13369 12631
rect 13369 12597 13403 12631
rect 13403 12597 13412 12631
rect 13360 12588 13412 12597
rect 14004 12588 14056 12640
rect 14464 12588 14516 12640
rect 15200 12588 15252 12640
rect 16856 12631 16908 12640
rect 16856 12597 16865 12631
rect 16865 12597 16899 12631
rect 16899 12597 16908 12631
rect 16856 12588 16908 12597
rect 19892 12588 19944 12640
rect 8982 12486 9034 12538
rect 9046 12486 9098 12538
rect 9110 12486 9162 12538
rect 9174 12486 9226 12538
rect 16982 12486 17034 12538
rect 17046 12486 17098 12538
rect 17110 12486 17162 12538
rect 17174 12486 17226 12538
rect 6368 12427 6420 12436
rect 6368 12393 6377 12427
rect 6377 12393 6411 12427
rect 6411 12393 6420 12427
rect 6368 12384 6420 12393
rect 7748 12384 7800 12436
rect 8668 12384 8720 12436
rect 9588 12384 9640 12436
rect 10416 12427 10468 12436
rect 10416 12393 10425 12427
rect 10425 12393 10459 12427
rect 10459 12393 10468 12427
rect 10416 12384 10468 12393
rect 10692 12384 10744 12436
rect 12716 12384 12768 12436
rect 14740 12427 14792 12436
rect 14740 12393 14749 12427
rect 14749 12393 14783 12427
rect 14783 12393 14792 12427
rect 14740 12384 14792 12393
rect 2504 12359 2556 12368
rect 2504 12325 2513 12359
rect 2513 12325 2547 12359
rect 2547 12325 2556 12359
rect 2504 12316 2556 12325
rect 5356 12316 5408 12368
rect 13360 12316 13412 12368
rect 14004 12359 14056 12368
rect 14004 12325 14013 12359
rect 14013 12325 14047 12359
rect 14047 12325 14056 12359
rect 14004 12316 14056 12325
rect 14556 12316 14608 12368
rect 15476 12359 15528 12368
rect 15476 12325 15485 12359
rect 15485 12325 15519 12359
rect 15519 12325 15528 12359
rect 15476 12316 15528 12325
rect 8024 12291 8076 12300
rect 8024 12257 8033 12291
rect 8033 12257 8067 12291
rect 8067 12257 8076 12291
rect 8024 12248 8076 12257
rect 9864 12248 9916 12300
rect 19892 12248 19944 12300
rect 20812 12248 20864 12300
rect 5632 12180 5684 12232
rect 7748 12223 7800 12232
rect 7748 12189 7757 12223
rect 7757 12189 7791 12223
rect 7791 12189 7800 12223
rect 7748 12180 7800 12189
rect 13728 12180 13780 12232
rect 14556 12180 14608 12232
rect 3056 12112 3108 12164
rect 4344 12112 4396 12164
rect 5448 12155 5500 12164
rect 5448 12121 5457 12155
rect 5457 12121 5491 12155
rect 5491 12121 5500 12155
rect 5448 12112 5500 12121
rect 14280 12112 14332 12164
rect 1676 12087 1728 12096
rect 1676 12053 1685 12087
rect 1685 12053 1719 12087
rect 1719 12053 1728 12087
rect 1676 12044 1728 12053
rect 2136 12087 2188 12096
rect 2136 12053 2145 12087
rect 2145 12053 2179 12087
rect 2179 12053 2188 12087
rect 2136 12044 2188 12053
rect 6644 12044 6696 12096
rect 7196 12087 7248 12096
rect 7196 12053 7205 12087
rect 7205 12053 7239 12087
rect 7239 12053 7248 12087
rect 7196 12044 7248 12053
rect 12808 12087 12860 12096
rect 12808 12053 12817 12087
rect 12817 12053 12851 12087
rect 12851 12053 12860 12087
rect 12808 12044 12860 12053
rect 23572 12044 23624 12096
rect 4982 11942 5034 11994
rect 5046 11942 5098 11994
rect 5110 11942 5162 11994
rect 5174 11942 5226 11994
rect 12982 11942 13034 11994
rect 13046 11942 13098 11994
rect 13110 11942 13162 11994
rect 13174 11942 13226 11994
rect 20982 11942 21034 11994
rect 21046 11942 21098 11994
rect 21110 11942 21162 11994
rect 21174 11942 21226 11994
rect 2136 11840 2188 11892
rect 2504 11840 2556 11892
rect 5632 11883 5684 11892
rect 5632 11849 5641 11883
rect 5641 11849 5675 11883
rect 5675 11849 5684 11883
rect 5632 11840 5684 11849
rect 6828 11840 6880 11892
rect 7196 11840 7248 11892
rect 9864 11840 9916 11892
rect 3056 11815 3108 11824
rect 3056 11781 3065 11815
rect 3065 11781 3099 11815
rect 3099 11781 3108 11815
rect 3056 11772 3108 11781
rect 3148 11772 3200 11824
rect 8392 11772 8444 11824
rect 4344 11747 4396 11756
rect 4344 11713 4353 11747
rect 4353 11713 4387 11747
rect 4387 11713 4396 11747
rect 4344 11704 4396 11713
rect 5448 11704 5500 11756
rect 7196 11704 7248 11756
rect 7380 11747 7432 11756
rect 7380 11713 7389 11747
rect 7389 11713 7423 11747
rect 7423 11713 7432 11747
rect 7380 11704 7432 11713
rect 8668 11747 8720 11756
rect 8668 11713 8677 11747
rect 8677 11713 8711 11747
rect 8711 11713 8720 11747
rect 8668 11704 8720 11713
rect 11244 11840 11296 11892
rect 12256 11883 12308 11892
rect 12256 11849 12265 11883
rect 12265 11849 12299 11883
rect 12299 11849 12308 11883
rect 12256 11840 12308 11849
rect 13360 11840 13412 11892
rect 13728 11840 13780 11892
rect 14556 11883 14608 11892
rect 14556 11849 14565 11883
rect 14565 11849 14599 11883
rect 14599 11849 14608 11883
rect 14556 11840 14608 11849
rect 15660 11883 15712 11892
rect 15660 11849 15669 11883
rect 15669 11849 15703 11883
rect 15703 11849 15712 11883
rect 15660 11840 15712 11849
rect 20812 11840 20864 11892
rect 2504 11611 2556 11620
rect 2504 11577 2513 11611
rect 2513 11577 2547 11611
rect 2547 11577 2556 11611
rect 2504 11568 2556 11577
rect 2596 11611 2648 11620
rect 2596 11577 2605 11611
rect 2605 11577 2639 11611
rect 2639 11577 2648 11611
rect 2596 11568 2648 11577
rect 4804 11568 4856 11620
rect 2044 11500 2096 11552
rect 2872 11500 2924 11552
rect 5356 11543 5408 11552
rect 5356 11509 5365 11543
rect 5365 11509 5399 11543
rect 5399 11509 5408 11543
rect 5356 11500 5408 11509
rect 6828 11500 6880 11552
rect 8024 11543 8076 11552
rect 8024 11509 8033 11543
rect 8033 11509 8067 11543
rect 8067 11509 8076 11543
rect 8024 11500 8076 11509
rect 9588 11568 9640 11620
rect 12808 11704 12860 11756
rect 16212 11679 16264 11688
rect 9404 11500 9456 11552
rect 10416 11500 10468 11552
rect 11704 11500 11756 11552
rect 16212 11645 16221 11679
rect 16221 11645 16255 11679
rect 16255 11645 16264 11679
rect 16212 11636 16264 11645
rect 14740 11611 14792 11620
rect 14740 11577 14749 11611
rect 14749 11577 14783 11611
rect 14783 11577 14792 11611
rect 14740 11568 14792 11577
rect 15476 11568 15528 11620
rect 14280 11500 14332 11552
rect 15384 11500 15436 11552
rect 16488 11543 16540 11552
rect 16488 11509 16497 11543
rect 16497 11509 16531 11543
rect 16531 11509 16540 11543
rect 16488 11500 16540 11509
rect 8982 11398 9034 11450
rect 9046 11398 9098 11450
rect 9110 11398 9162 11450
rect 9174 11398 9226 11450
rect 16982 11398 17034 11450
rect 17046 11398 17098 11450
rect 17110 11398 17162 11450
rect 17174 11398 17226 11450
rect 2136 11339 2188 11348
rect 2136 11305 2145 11339
rect 2145 11305 2179 11339
rect 2179 11305 2188 11339
rect 2136 11296 2188 11305
rect 2504 11296 2556 11348
rect 4436 11339 4488 11348
rect 4436 11305 4445 11339
rect 4445 11305 4479 11339
rect 4479 11305 4488 11339
rect 4436 11296 4488 11305
rect 4804 11296 4856 11348
rect 5632 11296 5684 11348
rect 13360 11296 13412 11348
rect 6644 11228 6696 11280
rect 10784 11228 10836 11280
rect 11704 11228 11756 11280
rect 12716 11228 12768 11280
rect 14004 11271 14056 11280
rect 14004 11237 14013 11271
rect 14013 11237 14047 11271
rect 14047 11237 14056 11271
rect 14004 11228 14056 11237
rect 14832 11228 14884 11280
rect 15476 11271 15528 11280
rect 15476 11237 15485 11271
rect 15485 11237 15519 11271
rect 15519 11237 15528 11271
rect 15476 11228 15528 11237
rect 18696 11271 18748 11280
rect 18696 11237 18705 11271
rect 18705 11237 18739 11271
rect 18739 11237 18748 11271
rect 18696 11228 18748 11237
rect 2596 11160 2648 11212
rect 9956 11203 10008 11212
rect 9956 11169 9965 11203
rect 9965 11169 9999 11203
rect 9999 11169 10008 11203
rect 9956 11160 10008 11169
rect 3332 11092 3384 11144
rect 4068 11135 4120 11144
rect 4068 11101 4077 11135
rect 4077 11101 4111 11135
rect 4111 11101 4120 11135
rect 4068 11092 4120 11101
rect 7380 11135 7432 11144
rect 6276 11024 6328 11076
rect 7380 11101 7389 11135
rect 7389 11101 7423 11135
rect 7423 11101 7432 11135
rect 7380 11092 7432 11101
rect 7932 11092 7984 11144
rect 20812 11160 20864 11212
rect 22100 11160 22152 11212
rect 10692 11092 10744 11144
rect 11612 11092 11664 11144
rect 15384 11135 15436 11144
rect 9772 11024 9824 11076
rect 10416 11024 10468 11076
rect 13544 11024 13596 11076
rect 15384 11101 15393 11135
rect 15393 11101 15427 11135
rect 15427 11101 15436 11135
rect 15384 11092 15436 11101
rect 18788 11092 18840 11144
rect 19156 11067 19208 11076
rect 19156 11033 19165 11067
rect 19165 11033 19199 11067
rect 19199 11033 19208 11067
rect 19156 11024 19208 11033
rect 11796 10956 11848 11008
rect 15200 10956 15252 11008
rect 16396 10956 16448 11008
rect 17316 10956 17368 11008
rect 19248 10956 19300 11008
rect 4982 10854 5034 10906
rect 5046 10854 5098 10906
rect 5110 10854 5162 10906
rect 5174 10854 5226 10906
rect 12982 10854 13034 10906
rect 13046 10854 13098 10906
rect 13110 10854 13162 10906
rect 13174 10854 13226 10906
rect 20982 10854 21034 10906
rect 21046 10854 21098 10906
rect 21110 10854 21162 10906
rect 21174 10854 21226 10906
rect 1584 10795 1636 10804
rect 1584 10761 1593 10795
rect 1593 10761 1627 10795
rect 1627 10761 1636 10795
rect 1584 10752 1636 10761
rect 2136 10752 2188 10804
rect 2504 10752 2556 10804
rect 4068 10752 4120 10804
rect 5448 10752 5500 10804
rect 6276 10795 6328 10804
rect 6276 10761 6285 10795
rect 6285 10761 6319 10795
rect 6319 10761 6328 10795
rect 6276 10752 6328 10761
rect 7748 10795 7800 10804
rect 7748 10761 7757 10795
rect 7757 10761 7791 10795
rect 7791 10761 7800 10795
rect 7748 10752 7800 10761
rect 9956 10752 10008 10804
rect 11244 10752 11296 10804
rect 11704 10752 11756 10804
rect 13360 10795 13412 10804
rect 13360 10761 13369 10795
rect 13369 10761 13403 10795
rect 13403 10761 13412 10795
rect 13360 10752 13412 10761
rect 14832 10795 14884 10804
rect 14832 10761 14841 10795
rect 14841 10761 14875 10795
rect 14875 10761 14884 10795
rect 14832 10752 14884 10761
rect 16212 10795 16264 10804
rect 16212 10761 16221 10795
rect 16221 10761 16255 10795
rect 16255 10761 16264 10795
rect 16212 10752 16264 10761
rect 20812 10752 20864 10804
rect 13544 10684 13596 10736
rect 13820 10684 13872 10736
rect 17960 10684 18012 10736
rect 18604 10684 18656 10736
rect 18880 10684 18932 10736
rect 5356 10616 5408 10668
rect 7932 10659 7984 10668
rect 7932 10625 7941 10659
rect 7941 10625 7975 10659
rect 7975 10625 7984 10659
rect 7932 10616 7984 10625
rect 8392 10659 8444 10668
rect 8392 10625 8401 10659
rect 8401 10625 8435 10659
rect 8435 10625 8444 10659
rect 8392 10616 8444 10625
rect 9496 10659 9548 10668
rect 9496 10625 9505 10659
rect 9505 10625 9539 10659
rect 9539 10625 9548 10659
rect 9496 10616 9548 10625
rect 9772 10659 9824 10668
rect 9772 10625 9781 10659
rect 9781 10625 9815 10659
rect 9815 10625 9824 10659
rect 9772 10616 9824 10625
rect 14004 10616 14056 10668
rect 18696 10616 18748 10668
rect 2228 10548 2280 10600
rect 3608 10548 3660 10600
rect 4804 10591 4856 10600
rect 4804 10557 4813 10591
rect 4813 10557 4847 10591
rect 4847 10557 4856 10591
rect 4804 10548 4856 10557
rect 12532 10591 12584 10600
rect 12532 10557 12550 10591
rect 12550 10557 12584 10591
rect 4712 10480 4764 10532
rect 12532 10548 12584 10557
rect 13912 10591 13964 10600
rect 13912 10557 13921 10591
rect 13921 10557 13955 10591
rect 13955 10557 13964 10591
rect 13912 10548 13964 10557
rect 16212 10548 16264 10600
rect 16764 10548 16816 10600
rect 17316 10548 17368 10600
rect 7564 10480 7616 10532
rect 7748 10480 7800 10532
rect 2044 10455 2096 10464
rect 2044 10421 2053 10455
rect 2053 10421 2087 10455
rect 2087 10421 2096 10455
rect 2044 10412 2096 10421
rect 3332 10455 3384 10464
rect 3332 10421 3341 10455
rect 3341 10421 3375 10455
rect 3375 10421 3384 10455
rect 3332 10412 3384 10421
rect 5448 10455 5500 10464
rect 5448 10421 5457 10455
rect 5457 10421 5491 10455
rect 5491 10421 5500 10455
rect 5448 10412 5500 10421
rect 6644 10455 6696 10464
rect 6644 10421 6653 10455
rect 6653 10421 6687 10455
rect 6687 10421 6696 10455
rect 6644 10412 6696 10421
rect 14004 10480 14056 10532
rect 16856 10480 16908 10532
rect 17776 10480 17828 10532
rect 18604 10523 18656 10532
rect 18604 10489 18613 10523
rect 18613 10489 18647 10523
rect 18647 10489 18656 10523
rect 18604 10480 18656 10489
rect 10416 10455 10468 10464
rect 10416 10421 10425 10455
rect 10425 10421 10459 10455
rect 10459 10421 10468 10455
rect 10416 10412 10468 10421
rect 10692 10412 10744 10464
rect 11612 10412 11664 10464
rect 12256 10412 12308 10464
rect 15384 10412 15436 10464
rect 15752 10455 15804 10464
rect 15752 10421 15761 10455
rect 15761 10421 15795 10455
rect 15795 10421 15804 10455
rect 15752 10412 15804 10421
rect 17408 10412 17460 10464
rect 18788 10480 18840 10532
rect 18880 10412 18932 10464
rect 19892 10455 19944 10464
rect 19892 10421 19901 10455
rect 19901 10421 19935 10455
rect 19935 10421 19944 10455
rect 19892 10412 19944 10421
rect 8982 10310 9034 10362
rect 9046 10310 9098 10362
rect 9110 10310 9162 10362
rect 9174 10310 9226 10362
rect 16982 10310 17034 10362
rect 17046 10310 17098 10362
rect 17110 10310 17162 10362
rect 17174 10310 17226 10362
rect 1676 10208 1728 10260
rect 3884 10208 3936 10260
rect 4252 10251 4304 10260
rect 4252 10217 4261 10251
rect 4261 10217 4295 10251
rect 4295 10217 4304 10251
rect 4252 10208 4304 10217
rect 4436 10208 4488 10260
rect 3976 10140 4028 10192
rect 6644 10208 6696 10260
rect 9496 10251 9548 10260
rect 9496 10217 9505 10251
rect 9505 10217 9539 10251
rect 9539 10217 9548 10251
rect 9496 10208 9548 10217
rect 12532 10251 12584 10260
rect 12532 10217 12541 10251
rect 12541 10217 12575 10251
rect 12575 10217 12584 10251
rect 12532 10208 12584 10217
rect 4068 10072 4120 10124
rect 4160 10072 4212 10124
rect 4804 10115 4856 10124
rect 4804 10081 4813 10115
rect 4813 10081 4847 10115
rect 4847 10081 4856 10115
rect 4804 10072 4856 10081
rect 7104 10140 7156 10192
rect 11612 10183 11664 10192
rect 11612 10149 11621 10183
rect 11621 10149 11655 10183
rect 11655 10149 11664 10183
rect 11612 10140 11664 10149
rect 5540 10115 5592 10124
rect 5540 10081 5549 10115
rect 5549 10081 5583 10115
rect 5583 10081 5592 10115
rect 5540 10072 5592 10081
rect 6092 10115 6144 10124
rect 6092 10081 6101 10115
rect 6101 10081 6135 10115
rect 6135 10081 6144 10115
rect 6092 10072 6144 10081
rect 10968 10115 11020 10124
rect 10968 10081 10977 10115
rect 10977 10081 11011 10115
rect 11011 10081 11020 10115
rect 10968 10072 11020 10081
rect 11336 10072 11388 10124
rect 12164 10072 12216 10124
rect 12348 10072 12400 10124
rect 15660 10208 15712 10260
rect 16856 10251 16908 10260
rect 16856 10217 16865 10251
rect 16865 10217 16899 10251
rect 16899 10217 16908 10251
rect 16856 10208 16908 10217
rect 18696 10208 18748 10260
rect 16120 10140 16172 10192
rect 13912 10115 13964 10124
rect 7380 10004 7432 10056
rect 12808 10004 12860 10056
rect 13912 10081 13921 10115
rect 13921 10081 13955 10115
rect 13955 10081 13964 10115
rect 13912 10072 13964 10081
rect 15844 10072 15896 10124
rect 16488 10115 16540 10124
rect 16488 10081 16497 10115
rect 16497 10081 16531 10115
rect 16531 10081 16540 10115
rect 16488 10072 16540 10081
rect 18328 10140 18380 10192
rect 20720 10072 20772 10124
rect 13544 10004 13596 10056
rect 17776 10004 17828 10056
rect 1584 9979 1636 9988
rect 1584 9945 1593 9979
rect 1593 9945 1627 9979
rect 1627 9945 1636 9979
rect 1584 9936 1636 9945
rect 2412 9936 2464 9988
rect 3976 9936 4028 9988
rect 10784 9936 10836 9988
rect 15752 9936 15804 9988
rect 20168 9936 20220 9988
rect 21088 9979 21140 9988
rect 21088 9945 21097 9979
rect 21097 9945 21131 9979
rect 21131 9945 21140 9979
rect 21088 9936 21140 9945
rect 2504 9868 2556 9920
rect 2596 9868 2648 9920
rect 3792 9868 3844 9920
rect 8116 9868 8168 9920
rect 10600 9911 10652 9920
rect 10600 9877 10609 9911
rect 10609 9877 10643 9911
rect 10643 9877 10652 9911
rect 10600 9868 10652 9877
rect 14556 9868 14608 9920
rect 15844 9911 15896 9920
rect 15844 9877 15853 9911
rect 15853 9877 15887 9911
rect 15887 9877 15896 9911
rect 15844 9868 15896 9877
rect 17408 9911 17460 9920
rect 17408 9877 17417 9911
rect 17417 9877 17451 9911
rect 17451 9877 17460 9911
rect 17408 9868 17460 9877
rect 4982 9766 5034 9818
rect 5046 9766 5098 9818
rect 5110 9766 5162 9818
rect 5174 9766 5226 9818
rect 12982 9766 13034 9818
rect 13046 9766 13098 9818
rect 13110 9766 13162 9818
rect 13174 9766 13226 9818
rect 20982 9766 21034 9818
rect 21046 9766 21098 9818
rect 21110 9766 21162 9818
rect 21174 9766 21226 9818
rect 6092 9664 6144 9716
rect 7104 9707 7156 9716
rect 7104 9673 7113 9707
rect 7113 9673 7147 9707
rect 7147 9673 7156 9707
rect 7104 9664 7156 9673
rect 7380 9707 7432 9716
rect 7380 9673 7389 9707
rect 7389 9673 7423 9707
rect 7423 9673 7432 9707
rect 7380 9664 7432 9673
rect 10600 9664 10652 9716
rect 11336 9707 11388 9716
rect 11336 9673 11345 9707
rect 11345 9673 11379 9707
rect 11379 9673 11388 9707
rect 11336 9664 11388 9673
rect 14004 9664 14056 9716
rect 16488 9664 16540 9716
rect 17776 9707 17828 9716
rect 17776 9673 17785 9707
rect 17785 9673 17819 9707
rect 17819 9673 17828 9707
rect 17776 9664 17828 9673
rect 5448 9596 5500 9648
rect 1952 9460 2004 9512
rect 2596 9528 2648 9580
rect 2412 9503 2464 9512
rect 2412 9469 2421 9503
rect 2421 9469 2455 9503
rect 2455 9469 2464 9503
rect 2412 9460 2464 9469
rect 2504 9460 2556 9512
rect 3148 9503 3200 9512
rect 3148 9469 3157 9503
rect 3157 9469 3191 9503
rect 3191 9469 3200 9503
rect 3148 9460 3200 9469
rect 3792 9460 3844 9512
rect 9772 9528 9824 9580
rect 10416 9528 10468 9580
rect 10784 9528 10836 9580
rect 11520 9528 11572 9580
rect 1768 9367 1820 9376
rect 1768 9333 1777 9367
rect 1777 9333 1811 9367
rect 1811 9333 1820 9367
rect 1768 9324 1820 9333
rect 2320 9324 2372 9376
rect 4068 9367 4120 9376
rect 4068 9333 4077 9367
rect 4077 9333 4111 9367
rect 4111 9333 4120 9367
rect 5264 9460 5316 9512
rect 6092 9460 6144 9512
rect 8116 9435 8168 9444
rect 8116 9401 8125 9435
rect 8125 9401 8159 9435
rect 8159 9401 8168 9435
rect 8116 9392 8168 9401
rect 4068 9324 4120 9333
rect 5540 9324 5592 9376
rect 6000 9367 6052 9376
rect 6000 9333 6009 9367
rect 6009 9333 6043 9367
rect 6043 9333 6052 9367
rect 6000 9324 6052 9333
rect 8024 9324 8076 9376
rect 8392 9392 8444 9444
rect 9680 9367 9732 9376
rect 9680 9333 9689 9367
rect 9689 9333 9723 9367
rect 9723 9333 9732 9367
rect 9680 9324 9732 9333
rect 10416 9324 10468 9376
rect 10968 9324 11020 9376
rect 15844 9596 15896 9648
rect 19064 9596 19116 9648
rect 17316 9528 17368 9580
rect 19248 9528 19300 9580
rect 12348 9324 12400 9376
rect 12992 9324 13044 9376
rect 13544 9460 13596 9512
rect 15568 9460 15620 9512
rect 13268 9324 13320 9376
rect 14004 9367 14056 9376
rect 14004 9333 14013 9367
rect 14013 9333 14047 9367
rect 14047 9333 14056 9367
rect 14004 9324 14056 9333
rect 14648 9324 14700 9376
rect 18052 9392 18104 9444
rect 19892 9392 19944 9444
rect 16212 9324 16264 9376
rect 16856 9324 16908 9376
rect 18328 9367 18380 9376
rect 18328 9333 18337 9367
rect 18337 9333 18371 9367
rect 18371 9333 18380 9367
rect 18328 9324 18380 9333
rect 20720 9324 20772 9376
rect 8982 9222 9034 9274
rect 9046 9222 9098 9274
rect 9110 9222 9162 9274
rect 9174 9222 9226 9274
rect 16982 9222 17034 9274
rect 17046 9222 17098 9274
rect 17110 9222 17162 9274
rect 17174 9222 17226 9274
rect 3792 9120 3844 9172
rect 3240 9052 3292 9104
rect 1952 9027 2004 9036
rect 1952 8993 1961 9027
rect 1961 8993 1995 9027
rect 1995 8993 2004 9027
rect 1952 8984 2004 8993
rect 2320 9027 2372 9036
rect 2320 8993 2329 9027
rect 2329 8993 2363 9027
rect 2363 8993 2372 9027
rect 2320 8984 2372 8993
rect 2504 9027 2556 9036
rect 2504 8993 2513 9027
rect 2513 8993 2547 9027
rect 2547 8993 2556 9027
rect 2504 8984 2556 8993
rect 2964 9027 3016 9036
rect 2964 8993 2973 9027
rect 2973 8993 3007 9027
rect 3007 8993 3016 9027
rect 5264 9120 5316 9172
rect 8392 9163 8444 9172
rect 8392 9129 8401 9163
rect 8401 9129 8435 9163
rect 8435 9129 8444 9163
rect 8392 9120 8444 9129
rect 10324 9163 10376 9172
rect 10324 9129 10333 9163
rect 10333 9129 10367 9163
rect 10367 9129 10376 9163
rect 10324 9120 10376 9129
rect 12808 9120 12860 9172
rect 12992 9120 13044 9172
rect 14924 9120 14976 9172
rect 15660 9163 15712 9172
rect 15660 9129 15669 9163
rect 15669 9129 15703 9163
rect 15703 9129 15712 9163
rect 15660 9120 15712 9129
rect 16212 9163 16264 9172
rect 16212 9129 16221 9163
rect 16221 9129 16255 9163
rect 16255 9129 16264 9163
rect 16212 9120 16264 9129
rect 19248 9120 19300 9172
rect 4804 9095 4856 9104
rect 4804 9061 4813 9095
rect 4813 9061 4847 9095
rect 4847 9061 4856 9095
rect 4804 9052 4856 9061
rect 5908 9052 5960 9104
rect 7104 9052 7156 9104
rect 9312 9052 9364 9104
rect 18052 9095 18104 9104
rect 18052 9061 18061 9095
rect 18061 9061 18095 9095
rect 18095 9061 18104 9095
rect 18052 9052 18104 9061
rect 20812 9052 20864 9104
rect 2964 8984 3016 8993
rect 6000 9027 6052 9036
rect 3976 8916 4028 8968
rect 4344 8916 4396 8968
rect 6000 8993 6009 9027
rect 6009 8993 6043 9027
rect 6043 8993 6052 9027
rect 6000 8984 6052 8993
rect 6368 9027 6420 9036
rect 6368 8993 6377 9027
rect 6377 8993 6411 9027
rect 6411 8993 6420 9027
rect 6368 8984 6420 8993
rect 9680 9027 9732 9036
rect 9680 8993 9689 9027
rect 9689 8993 9723 9027
rect 9723 8993 9732 9027
rect 9680 8984 9732 8993
rect 9864 9027 9916 9036
rect 9864 8993 9870 9027
rect 9870 8993 9916 9027
rect 9864 8984 9916 8993
rect 10600 8984 10652 9036
rect 11244 9027 11296 9036
rect 11244 8993 11253 9027
rect 11253 8993 11287 9027
rect 11287 8993 11296 9027
rect 11244 8984 11296 8993
rect 11520 9027 11572 9036
rect 11520 8993 11529 9027
rect 11529 8993 11563 9027
rect 11563 8993 11572 9027
rect 11520 8984 11572 8993
rect 13912 9027 13964 9036
rect 13912 8993 13921 9027
rect 13921 8993 13955 9027
rect 13955 8993 13964 9027
rect 13912 8984 13964 8993
rect 14280 8984 14332 9036
rect 21272 8984 21324 9036
rect 6460 8916 6512 8968
rect 7472 8959 7524 8968
rect 7472 8925 7481 8959
rect 7481 8925 7515 8959
rect 7515 8925 7524 8959
rect 7472 8916 7524 8925
rect 10692 8916 10744 8968
rect 15016 8916 15068 8968
rect 17960 8959 18012 8968
rect 17960 8925 17969 8959
rect 17969 8925 18003 8959
rect 18003 8925 18012 8959
rect 17960 8916 18012 8925
rect 18604 8959 18656 8968
rect 18604 8925 18613 8959
rect 18613 8925 18647 8959
rect 18647 8925 18656 8959
rect 18604 8916 18656 8925
rect 10784 8848 10836 8900
rect 9588 8780 9640 8832
rect 10416 8780 10468 8832
rect 4982 8678 5034 8730
rect 5046 8678 5098 8730
rect 5110 8678 5162 8730
rect 5174 8678 5226 8730
rect 12982 8678 13034 8730
rect 13046 8678 13098 8730
rect 13110 8678 13162 8730
rect 13174 8678 13226 8730
rect 20982 8678 21034 8730
rect 21046 8678 21098 8730
rect 21110 8678 21162 8730
rect 21174 8678 21226 8730
rect 3976 8619 4028 8628
rect 3976 8585 3985 8619
rect 3985 8585 4019 8619
rect 4019 8585 4028 8619
rect 3976 8576 4028 8585
rect 4344 8576 4396 8628
rect 6460 8619 6512 8628
rect 1768 8483 1820 8492
rect 1768 8449 1777 8483
rect 1777 8449 1811 8483
rect 1811 8449 1820 8483
rect 1768 8440 1820 8449
rect 3148 8440 3200 8492
rect 3332 8483 3384 8492
rect 3332 8449 3341 8483
rect 3341 8449 3375 8483
rect 3375 8449 3384 8483
rect 3332 8440 3384 8449
rect 6460 8585 6469 8619
rect 6469 8585 6503 8619
rect 6503 8585 6512 8619
rect 14648 8619 14700 8628
rect 6460 8576 6512 8585
rect 4804 8551 4856 8560
rect 4804 8517 4813 8551
rect 4813 8517 4847 8551
rect 4847 8517 4856 8551
rect 4804 8508 4856 8517
rect 6736 8508 6788 8560
rect 14648 8585 14657 8619
rect 14657 8585 14691 8619
rect 14691 8585 14700 8619
rect 14648 8576 14700 8585
rect 18052 8576 18104 8628
rect 10784 8551 10836 8560
rect 10784 8517 10793 8551
rect 10793 8517 10827 8551
rect 10827 8517 10836 8551
rect 10784 8508 10836 8517
rect 17960 8508 18012 8560
rect 1952 8415 2004 8424
rect 1952 8381 1961 8415
rect 1961 8381 1995 8415
rect 1995 8381 2004 8415
rect 1952 8372 2004 8381
rect 2136 8372 2188 8424
rect 2504 8372 2556 8424
rect 5632 8440 5684 8492
rect 6368 8440 6420 8492
rect 7104 8483 7156 8492
rect 7104 8449 7113 8483
rect 7113 8449 7147 8483
rect 7147 8449 7156 8483
rect 7104 8440 7156 8449
rect 5356 8304 5408 8356
rect 7288 8372 7340 8424
rect 9588 8440 9640 8492
rect 8208 8415 8260 8424
rect 8208 8381 8217 8415
rect 8217 8381 8251 8415
rect 8251 8381 8260 8415
rect 8208 8372 8260 8381
rect 9312 8372 9364 8424
rect 9772 8440 9824 8492
rect 13544 8483 13596 8492
rect 8484 8304 8536 8356
rect 8852 8304 8904 8356
rect 5540 8236 5592 8288
rect 8208 8236 8260 8288
rect 10416 8279 10468 8288
rect 10416 8245 10425 8279
rect 10425 8245 10459 8279
rect 10459 8245 10468 8279
rect 10416 8236 10468 8245
rect 10692 8236 10744 8288
rect 11520 8236 11572 8288
rect 13268 8372 13320 8424
rect 13544 8449 13553 8483
rect 13553 8449 13587 8483
rect 13587 8449 13596 8483
rect 13544 8440 13596 8449
rect 14924 8483 14976 8492
rect 14924 8449 14933 8483
rect 14933 8449 14967 8483
rect 14967 8449 14976 8483
rect 14924 8440 14976 8449
rect 15660 8440 15712 8492
rect 17500 8440 17552 8492
rect 18604 8440 18656 8492
rect 13452 8372 13504 8424
rect 14648 8304 14700 8356
rect 15568 8347 15620 8356
rect 15568 8313 15577 8347
rect 15577 8313 15611 8347
rect 15611 8313 15620 8347
rect 15568 8304 15620 8313
rect 16764 8372 16816 8424
rect 18052 8415 18104 8424
rect 18052 8381 18061 8415
rect 18061 8381 18095 8415
rect 18095 8381 18104 8415
rect 18052 8372 18104 8381
rect 18328 8304 18380 8356
rect 13912 8279 13964 8288
rect 13912 8245 13921 8279
rect 13921 8245 13955 8279
rect 13955 8245 13964 8279
rect 13912 8236 13964 8245
rect 14280 8279 14332 8288
rect 14280 8245 14289 8279
rect 14289 8245 14323 8279
rect 14323 8245 14332 8279
rect 14280 8236 14332 8245
rect 16212 8279 16264 8288
rect 16212 8245 16221 8279
rect 16221 8245 16255 8279
rect 16255 8245 16264 8279
rect 16212 8236 16264 8245
rect 17500 8236 17552 8288
rect 18972 8279 19024 8288
rect 18972 8245 18981 8279
rect 18981 8245 19015 8279
rect 19015 8245 19024 8279
rect 18972 8236 19024 8245
rect 19524 8236 19576 8288
rect 19800 8236 19852 8288
rect 19984 8347 20036 8356
rect 19984 8313 19993 8347
rect 19993 8313 20027 8347
rect 20027 8313 20036 8347
rect 19984 8304 20036 8313
rect 21272 8236 21324 8288
rect 23204 8236 23256 8288
rect 8982 8134 9034 8186
rect 9046 8134 9098 8186
rect 9110 8134 9162 8186
rect 9174 8134 9226 8186
rect 16982 8134 17034 8186
rect 17046 8134 17098 8186
rect 17110 8134 17162 8186
rect 17174 8134 17226 8186
rect 2320 8075 2372 8084
rect 2320 8041 2329 8075
rect 2329 8041 2363 8075
rect 2363 8041 2372 8075
rect 2320 8032 2372 8041
rect 2964 8032 3016 8084
rect 3424 8032 3476 8084
rect 3792 8032 3844 8084
rect 4252 8032 4304 8084
rect 7288 8032 7340 8084
rect 7472 8075 7524 8084
rect 7472 8041 7481 8075
rect 7481 8041 7515 8075
rect 7515 8041 7524 8075
rect 7472 8032 7524 8041
rect 5540 8007 5592 8016
rect 5540 7973 5549 8007
rect 5549 7973 5583 8007
rect 5583 7973 5592 8007
rect 5540 7964 5592 7973
rect 9588 8032 9640 8084
rect 9864 8075 9916 8084
rect 9864 8041 9873 8075
rect 9873 8041 9907 8075
rect 9907 8041 9916 8075
rect 9864 8032 9916 8041
rect 11244 8032 11296 8084
rect 14004 8032 14056 8084
rect 15016 8075 15068 8084
rect 15016 8041 15025 8075
rect 15025 8041 15059 8075
rect 15059 8041 15068 8075
rect 15016 8032 15068 8041
rect 15384 8075 15436 8084
rect 15384 8041 15393 8075
rect 15393 8041 15427 8075
rect 15427 8041 15436 8075
rect 15384 8032 15436 8041
rect 1952 7896 2004 7948
rect 2136 7939 2188 7948
rect 2136 7905 2145 7939
rect 2145 7905 2179 7939
rect 2179 7905 2188 7939
rect 2136 7896 2188 7905
rect 8484 7939 8536 7948
rect 8484 7905 8493 7939
rect 8493 7905 8527 7939
rect 8527 7905 8536 7939
rect 8484 7896 8536 7905
rect 8852 7896 8904 7948
rect 9680 7896 9732 7948
rect 10232 7939 10284 7948
rect 10232 7905 10241 7939
rect 10241 7905 10275 7939
rect 10275 7905 10284 7939
rect 10232 7896 10284 7905
rect 11060 7964 11112 8016
rect 16212 7964 16264 8016
rect 5908 7871 5960 7880
rect 5908 7837 5917 7871
rect 5917 7837 5951 7871
rect 5951 7837 5960 7871
rect 5908 7828 5960 7837
rect 5448 7760 5500 7812
rect 10784 7896 10836 7948
rect 11152 7896 11204 7948
rect 11796 7939 11848 7948
rect 11796 7905 11805 7939
rect 11805 7905 11839 7939
rect 11839 7905 11848 7939
rect 11796 7896 11848 7905
rect 11888 7896 11940 7948
rect 13912 7896 13964 7948
rect 12440 7871 12492 7880
rect 12440 7837 12449 7871
rect 12449 7837 12483 7871
rect 12483 7837 12492 7871
rect 12440 7828 12492 7837
rect 13452 7871 13504 7880
rect 13452 7837 13461 7871
rect 13461 7837 13495 7871
rect 13495 7837 13504 7871
rect 13452 7828 13504 7837
rect 15936 7896 15988 7948
rect 15660 7828 15712 7880
rect 16764 8032 16816 8084
rect 18052 8075 18104 8084
rect 18052 8041 18061 8075
rect 18061 8041 18095 8075
rect 18095 8041 18104 8075
rect 18052 8032 18104 8041
rect 19524 8032 19576 8084
rect 19984 8032 20036 8084
rect 17868 7964 17920 8016
rect 18972 7964 19024 8016
rect 19156 8007 19208 8016
rect 19156 7973 19165 8007
rect 19165 7973 19199 8007
rect 19199 7973 19208 8007
rect 19156 7964 19208 7973
rect 16856 7939 16908 7948
rect 16856 7905 16865 7939
rect 16865 7905 16899 7939
rect 16899 7905 16908 7939
rect 16856 7896 16908 7905
rect 18512 7871 18564 7880
rect 18512 7837 18521 7871
rect 18521 7837 18555 7871
rect 18555 7837 18564 7871
rect 18512 7828 18564 7837
rect 18604 7828 18656 7880
rect 1952 7735 2004 7744
rect 1952 7701 1961 7735
rect 1961 7701 1995 7735
rect 1995 7701 2004 7735
rect 1952 7692 2004 7701
rect 5356 7692 5408 7744
rect 6184 7735 6236 7744
rect 6184 7701 6193 7735
rect 6193 7701 6227 7735
rect 6227 7701 6236 7735
rect 6184 7692 6236 7701
rect 8208 7692 8260 7744
rect 10784 7760 10836 7812
rect 12716 7760 12768 7812
rect 14372 7735 14424 7744
rect 14372 7701 14381 7735
rect 14381 7701 14415 7735
rect 14415 7701 14424 7735
rect 14372 7692 14424 7701
rect 16488 7692 16540 7744
rect 19432 7735 19484 7744
rect 19432 7701 19441 7735
rect 19441 7701 19475 7735
rect 19475 7701 19484 7735
rect 19432 7692 19484 7701
rect 19800 7735 19852 7744
rect 19800 7701 19809 7735
rect 19809 7701 19843 7735
rect 19843 7701 19852 7735
rect 19800 7692 19852 7701
rect 4982 7590 5034 7642
rect 5046 7590 5098 7642
rect 5110 7590 5162 7642
rect 5174 7590 5226 7642
rect 12982 7590 13034 7642
rect 13046 7590 13098 7642
rect 13110 7590 13162 7642
rect 13174 7590 13226 7642
rect 20982 7590 21034 7642
rect 21046 7590 21098 7642
rect 21110 7590 21162 7642
rect 21174 7590 21226 7642
rect 1584 7531 1636 7540
rect 1584 7497 1593 7531
rect 1593 7497 1627 7531
rect 1627 7497 1636 7531
rect 1584 7488 1636 7497
rect 2504 7531 2556 7540
rect 2504 7497 2513 7531
rect 2513 7497 2547 7531
rect 2547 7497 2556 7531
rect 2504 7488 2556 7497
rect 2688 7488 2740 7540
rect 1492 7352 1544 7404
rect 4068 7488 4120 7540
rect 3884 7420 3936 7472
rect 5356 7488 5408 7540
rect 6736 7488 6788 7540
rect 7748 7488 7800 7540
rect 8484 7488 8536 7540
rect 9312 7488 9364 7540
rect 10140 7488 10192 7540
rect 10232 7488 10284 7540
rect 11888 7531 11940 7540
rect 11888 7497 11897 7531
rect 11897 7497 11931 7531
rect 11931 7497 11940 7531
rect 11888 7488 11940 7497
rect 13452 7488 13504 7540
rect 15384 7488 15436 7540
rect 15660 7531 15712 7540
rect 15660 7497 15669 7531
rect 15669 7497 15703 7531
rect 15703 7497 15712 7531
rect 15660 7488 15712 7497
rect 17868 7531 17920 7540
rect 5908 7420 5960 7472
rect 8208 7420 8260 7472
rect 7656 7352 7708 7404
rect 12440 7395 12492 7404
rect 12440 7361 12449 7395
rect 12449 7361 12483 7395
rect 12483 7361 12492 7395
rect 12440 7352 12492 7361
rect 5448 7284 5500 7336
rect 6736 7284 6788 7336
rect 9588 7327 9640 7336
rect 9588 7293 9597 7327
rect 9597 7293 9631 7327
rect 9631 7293 9640 7327
rect 9588 7284 9640 7293
rect 9956 7327 10008 7336
rect 9956 7293 9965 7327
rect 9965 7293 9999 7327
rect 9999 7293 10008 7327
rect 9956 7284 10008 7293
rect 1952 7148 2004 7200
rect 2596 7148 2648 7200
rect 7748 7259 7800 7268
rect 7748 7225 7757 7259
rect 7757 7225 7791 7259
rect 7791 7225 7800 7259
rect 7748 7216 7800 7225
rect 9312 7216 9364 7268
rect 12532 7216 12584 7268
rect 14004 7420 14056 7472
rect 14372 7463 14424 7472
rect 14372 7429 14381 7463
rect 14381 7429 14415 7463
rect 14415 7429 14424 7463
rect 14372 7420 14424 7429
rect 14740 7420 14792 7472
rect 15568 7420 15620 7472
rect 17868 7497 17877 7531
rect 17877 7497 17911 7531
rect 17911 7497 17920 7531
rect 17868 7488 17920 7497
rect 19800 7488 19852 7540
rect 19524 7420 19576 7472
rect 15936 7395 15988 7404
rect 15936 7361 15945 7395
rect 15945 7361 15979 7395
rect 15979 7361 15988 7395
rect 15936 7352 15988 7361
rect 16488 7352 16540 7404
rect 18236 7284 18288 7336
rect 19248 7352 19300 7404
rect 19892 7395 19944 7404
rect 19892 7361 19901 7395
rect 19901 7361 19935 7395
rect 19935 7361 19944 7395
rect 19892 7352 19944 7361
rect 4620 7148 4672 7200
rect 4988 7148 5040 7200
rect 10784 7191 10836 7200
rect 10784 7157 10793 7191
rect 10793 7157 10827 7191
rect 10827 7157 10836 7191
rect 10784 7148 10836 7157
rect 11336 7191 11388 7200
rect 11336 7157 11345 7191
rect 11345 7157 11379 7191
rect 11379 7157 11388 7191
rect 11336 7148 11388 7157
rect 13360 7191 13412 7200
rect 13360 7157 13369 7191
rect 13369 7157 13403 7191
rect 13403 7157 13412 7191
rect 13360 7148 13412 7157
rect 14556 7148 14608 7200
rect 14740 7259 14792 7268
rect 14740 7225 14749 7259
rect 14749 7225 14783 7259
rect 14783 7225 14792 7259
rect 14740 7216 14792 7225
rect 16304 7259 16356 7268
rect 16304 7225 16313 7259
rect 16313 7225 16347 7259
rect 16347 7225 16356 7259
rect 16304 7216 16356 7225
rect 19432 7259 19484 7268
rect 19432 7225 19441 7259
rect 19441 7225 19475 7259
rect 19475 7225 19484 7259
rect 19432 7216 19484 7225
rect 19524 7259 19576 7268
rect 19524 7225 19533 7259
rect 19533 7225 19567 7259
rect 19567 7225 19576 7259
rect 19524 7216 19576 7225
rect 16028 7148 16080 7200
rect 16856 7148 16908 7200
rect 19616 7148 19668 7200
rect 8982 7046 9034 7098
rect 9046 7046 9098 7098
rect 9110 7046 9162 7098
rect 9174 7046 9226 7098
rect 16982 7046 17034 7098
rect 17046 7046 17098 7098
rect 17110 7046 17162 7098
rect 17174 7046 17226 7098
rect 1492 6944 1544 6996
rect 4988 6987 5040 6996
rect 4988 6953 4997 6987
rect 4997 6953 5031 6987
rect 5031 6953 5040 6987
rect 4988 6944 5040 6953
rect 5540 6944 5592 6996
rect 4068 6876 4120 6928
rect 4436 6919 4488 6928
rect 4436 6885 4439 6919
rect 4439 6885 4473 6919
rect 4473 6885 4488 6919
rect 4436 6876 4488 6885
rect 7104 6876 7156 6928
rect 9588 6944 9640 6996
rect 11152 6987 11204 6996
rect 11152 6953 11161 6987
rect 11161 6953 11195 6987
rect 11195 6953 11204 6987
rect 11152 6944 11204 6953
rect 11796 6987 11848 6996
rect 11796 6953 11805 6987
rect 11805 6953 11839 6987
rect 11839 6953 11848 6987
rect 11796 6944 11848 6953
rect 12440 6987 12492 6996
rect 12440 6953 12449 6987
rect 12449 6953 12483 6987
rect 12483 6953 12492 6987
rect 12440 6944 12492 6953
rect 12716 6944 12768 6996
rect 13728 6944 13780 6996
rect 8852 6876 8904 6928
rect 11888 6876 11940 6928
rect 13360 6876 13412 6928
rect 2412 6851 2464 6860
rect 2412 6817 2421 6851
rect 2421 6817 2455 6851
rect 2455 6817 2464 6851
rect 2412 6808 2464 6817
rect 2504 6808 2556 6860
rect 8208 6851 8260 6860
rect 8208 6817 8217 6851
rect 8217 6817 8251 6851
rect 8251 6817 8260 6851
rect 8208 6808 8260 6817
rect 8392 6851 8444 6860
rect 8392 6817 8401 6851
rect 8401 6817 8435 6851
rect 8435 6817 8444 6851
rect 8392 6808 8444 6817
rect 10140 6851 10192 6860
rect 10140 6817 10149 6851
rect 10149 6817 10183 6851
rect 10183 6817 10192 6851
rect 10140 6808 10192 6817
rect 10784 6808 10836 6860
rect 5724 6740 5776 6792
rect 6092 6740 6144 6792
rect 12164 6740 12216 6792
rect 13636 6740 13688 6792
rect 13820 6740 13872 6792
rect 5448 6672 5500 6724
rect 10416 6672 10468 6724
rect 16488 6944 16540 6996
rect 21364 6944 21416 6996
rect 16304 6876 16356 6928
rect 17408 6876 17460 6928
rect 18512 6876 18564 6928
rect 15936 6808 15988 6860
rect 17132 6808 17184 6860
rect 20444 6808 20496 6860
rect 18604 6740 18656 6792
rect 18696 6740 18748 6792
rect 2964 6604 3016 6656
rect 7380 6647 7432 6656
rect 7380 6613 7389 6647
rect 7389 6613 7423 6647
rect 7423 6613 7432 6647
rect 7380 6604 7432 6613
rect 9312 6647 9364 6656
rect 9312 6613 9321 6647
rect 9321 6613 9355 6647
rect 9355 6613 9364 6647
rect 9312 6604 9364 6613
rect 14556 6647 14608 6656
rect 14556 6613 14565 6647
rect 14565 6613 14599 6647
rect 14599 6613 14608 6647
rect 14556 6604 14608 6613
rect 16028 6604 16080 6656
rect 16488 6604 16540 6656
rect 16672 6604 16724 6656
rect 19340 6604 19392 6656
rect 4982 6502 5034 6554
rect 5046 6502 5098 6554
rect 5110 6502 5162 6554
rect 5174 6502 5226 6554
rect 12982 6502 13034 6554
rect 13046 6502 13098 6554
rect 13110 6502 13162 6554
rect 13174 6502 13226 6554
rect 20982 6502 21034 6554
rect 21046 6502 21098 6554
rect 21110 6502 21162 6554
rect 21174 6502 21226 6554
rect 4620 6443 4672 6452
rect 4620 6409 4629 6443
rect 4629 6409 4663 6443
rect 4663 6409 4672 6443
rect 4620 6400 4672 6409
rect 5724 6443 5776 6452
rect 5724 6409 5733 6443
rect 5733 6409 5767 6443
rect 5767 6409 5776 6443
rect 5724 6400 5776 6409
rect 7104 6400 7156 6452
rect 7380 6443 7432 6452
rect 7380 6409 7389 6443
rect 7389 6409 7423 6443
rect 7423 6409 7432 6443
rect 7380 6400 7432 6409
rect 8208 6400 8260 6452
rect 9956 6400 10008 6452
rect 10416 6443 10468 6452
rect 10416 6409 10425 6443
rect 10425 6409 10459 6443
rect 10459 6409 10468 6443
rect 10416 6400 10468 6409
rect 11336 6400 11388 6452
rect 12164 6443 12216 6452
rect 12164 6409 12173 6443
rect 12173 6409 12207 6443
rect 12207 6409 12216 6443
rect 12164 6400 12216 6409
rect 13360 6400 13412 6452
rect 16764 6400 16816 6452
rect 17132 6443 17184 6452
rect 17132 6409 17141 6443
rect 17141 6409 17175 6443
rect 17175 6409 17184 6443
rect 17132 6400 17184 6409
rect 18604 6400 18656 6452
rect 20628 6400 20680 6452
rect 664 6332 716 6384
rect 9312 6332 9364 6384
rect 2964 6307 3016 6316
rect 2964 6273 2973 6307
rect 2973 6273 3007 6307
rect 3007 6273 3016 6307
rect 2964 6264 3016 6273
rect 1860 6239 1912 6248
rect 1860 6205 1869 6239
rect 1869 6205 1903 6239
rect 1903 6205 1912 6239
rect 1860 6196 1912 6205
rect 3056 6171 3108 6180
rect 3056 6137 3065 6171
rect 3065 6137 3099 6171
rect 3099 6137 3108 6171
rect 3056 6128 3108 6137
rect 3240 6128 3292 6180
rect 4804 6171 4856 6180
rect 4804 6137 4813 6171
rect 4813 6137 4847 6171
rect 4847 6137 4856 6171
rect 4804 6128 4856 6137
rect 7656 6264 7708 6316
rect 8392 6264 8444 6316
rect 14556 6332 14608 6384
rect 10048 6264 10100 6316
rect 2504 6103 2556 6112
rect 2504 6069 2513 6103
rect 2513 6069 2547 6103
rect 2547 6069 2556 6103
rect 2504 6060 2556 6069
rect 4068 6103 4120 6112
rect 4068 6069 4077 6103
rect 4077 6069 4111 6103
rect 4111 6069 4120 6103
rect 4068 6060 4120 6069
rect 4620 6060 4672 6112
rect 6736 6128 6788 6180
rect 6092 6103 6144 6112
rect 6092 6069 6101 6103
rect 6101 6069 6135 6103
rect 6135 6069 6144 6103
rect 6092 6060 6144 6069
rect 7380 6060 7432 6112
rect 8392 6128 8444 6180
rect 8760 6128 8812 6180
rect 10784 6128 10836 6180
rect 11520 6128 11572 6180
rect 15292 6264 15344 6316
rect 13268 6239 13320 6248
rect 13268 6205 13277 6239
rect 13277 6205 13311 6239
rect 13311 6205 13320 6239
rect 13268 6196 13320 6205
rect 13728 6196 13780 6248
rect 14832 6196 14884 6248
rect 16120 6239 16172 6248
rect 16120 6205 16129 6239
rect 16129 6205 16163 6239
rect 16163 6205 16172 6239
rect 16120 6196 16172 6205
rect 16488 6196 16540 6248
rect 19248 6264 19300 6316
rect 18328 6196 18380 6248
rect 14188 6171 14240 6180
rect 14188 6137 14197 6171
rect 14197 6137 14231 6171
rect 14231 6137 14240 6171
rect 14188 6128 14240 6137
rect 16856 6171 16908 6180
rect 16856 6137 16865 6171
rect 16865 6137 16899 6171
rect 16899 6137 16908 6171
rect 16856 6128 16908 6137
rect 9496 6060 9548 6112
rect 11244 6060 11296 6112
rect 13820 6060 13872 6112
rect 14464 6060 14516 6112
rect 15108 6060 15160 6112
rect 15936 6103 15988 6112
rect 15936 6069 15945 6103
rect 15945 6069 15979 6103
rect 15979 6069 15988 6103
rect 15936 6060 15988 6069
rect 18420 6060 18472 6112
rect 19340 6128 19392 6180
rect 20444 6128 20496 6180
rect 8982 5958 9034 6010
rect 9046 5958 9098 6010
rect 9110 5958 9162 6010
rect 9174 5958 9226 6010
rect 16982 5958 17034 6010
rect 17046 5958 17098 6010
rect 17110 5958 17162 6010
rect 17174 5958 17226 6010
rect 3056 5856 3108 5908
rect 3516 5856 3568 5908
rect 4160 5899 4212 5908
rect 4160 5865 4169 5899
rect 4169 5865 4203 5899
rect 4203 5865 4212 5899
rect 4160 5856 4212 5865
rect 4804 5856 4856 5908
rect 6092 5899 6144 5908
rect 6092 5865 6101 5899
rect 6101 5865 6135 5899
rect 6135 5865 6144 5899
rect 6092 5856 6144 5865
rect 7656 5899 7708 5908
rect 7656 5865 7665 5899
rect 7665 5865 7699 5899
rect 7699 5865 7708 5899
rect 7656 5856 7708 5865
rect 10140 5856 10192 5908
rect 14188 5899 14240 5908
rect 14188 5865 14197 5899
rect 14197 5865 14231 5899
rect 14231 5865 14240 5899
rect 14188 5856 14240 5865
rect 16028 5856 16080 5908
rect 18512 5899 18564 5908
rect 18512 5865 18521 5899
rect 18521 5865 18555 5899
rect 18555 5865 18564 5899
rect 18512 5856 18564 5865
rect 19340 5856 19392 5908
rect 19432 5856 19484 5908
rect 2504 5788 2556 5840
rect 4252 5788 4304 5840
rect 2872 5720 2924 5772
rect 3240 5720 3292 5772
rect 4436 5720 4488 5772
rect 8208 5831 8260 5840
rect 8208 5797 8217 5831
rect 8217 5797 8251 5831
rect 8251 5797 8260 5831
rect 8208 5788 8260 5797
rect 6184 5720 6236 5772
rect 10048 5763 10100 5772
rect 10048 5729 10057 5763
rect 10057 5729 10091 5763
rect 10091 5729 10100 5763
rect 10048 5720 10100 5729
rect 10140 5720 10192 5772
rect 13360 5788 13412 5840
rect 15476 5831 15528 5840
rect 15476 5797 15485 5831
rect 15485 5797 15519 5831
rect 15519 5797 15528 5831
rect 15476 5788 15528 5797
rect 17408 5788 17460 5840
rect 6644 5652 6696 5704
rect 6736 5652 6788 5704
rect 8116 5695 8168 5704
rect 8116 5661 8125 5695
rect 8125 5661 8159 5695
rect 8159 5661 8168 5695
rect 8116 5652 8168 5661
rect 8392 5695 8444 5704
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 10416 5695 10468 5704
rect 10416 5661 10425 5695
rect 10425 5661 10459 5695
rect 10459 5661 10468 5695
rect 10416 5652 10468 5661
rect 5448 5584 5500 5636
rect 10876 5584 10928 5636
rect 11888 5763 11940 5772
rect 11888 5729 11897 5763
rect 11897 5729 11931 5763
rect 11931 5729 11940 5763
rect 11888 5720 11940 5729
rect 16856 5763 16908 5772
rect 16856 5729 16865 5763
rect 16865 5729 16899 5763
rect 16899 5729 16908 5763
rect 16856 5720 16908 5729
rect 12072 5695 12124 5704
rect 12072 5661 12081 5695
rect 12081 5661 12115 5695
rect 12115 5661 12124 5695
rect 12072 5652 12124 5661
rect 12808 5652 12860 5704
rect 13268 5695 13320 5704
rect 13268 5661 13277 5695
rect 13277 5661 13311 5695
rect 13311 5661 13320 5695
rect 13268 5652 13320 5661
rect 15108 5652 15160 5704
rect 16580 5652 16632 5704
rect 2412 5516 2464 5568
rect 3976 5516 4028 5568
rect 7288 5559 7340 5568
rect 7288 5525 7297 5559
rect 7297 5525 7331 5559
rect 7331 5525 7340 5559
rect 7288 5516 7340 5525
rect 7472 5516 7524 5568
rect 12348 5584 12400 5636
rect 16120 5584 16172 5636
rect 16396 5516 16448 5568
rect 21548 5720 21600 5772
rect 18512 5652 18564 5704
rect 19616 5652 19668 5704
rect 19340 5627 19392 5636
rect 19340 5593 19349 5627
rect 19349 5593 19383 5627
rect 19383 5593 19392 5627
rect 19340 5584 19392 5593
rect 4982 5414 5034 5466
rect 5046 5414 5098 5466
rect 5110 5414 5162 5466
rect 5174 5414 5226 5466
rect 12982 5414 13034 5466
rect 13046 5414 13098 5466
rect 13110 5414 13162 5466
rect 13174 5414 13226 5466
rect 20982 5414 21034 5466
rect 21046 5414 21098 5466
rect 21110 5414 21162 5466
rect 21174 5414 21226 5466
rect 3516 5355 3568 5364
rect 3516 5321 3525 5355
rect 3525 5321 3559 5355
rect 3559 5321 3568 5355
rect 3516 5312 3568 5321
rect 4252 5355 4304 5364
rect 4252 5321 4261 5355
rect 4261 5321 4295 5355
rect 4295 5321 4304 5355
rect 4252 5312 4304 5321
rect 6184 5355 6236 5364
rect 6184 5321 6193 5355
rect 6193 5321 6227 5355
rect 6227 5321 6236 5355
rect 6184 5312 6236 5321
rect 7104 5355 7156 5364
rect 7104 5321 7113 5355
rect 7113 5321 7147 5355
rect 7147 5321 7156 5355
rect 7104 5312 7156 5321
rect 8208 5312 8260 5364
rect 10048 5312 10100 5364
rect 11888 5312 11940 5364
rect 12532 5312 12584 5364
rect 13360 5355 13412 5364
rect 13360 5321 13369 5355
rect 13369 5321 13403 5355
rect 13403 5321 13412 5355
rect 13360 5312 13412 5321
rect 18512 5355 18564 5364
rect 18512 5321 18521 5355
rect 18521 5321 18555 5355
rect 18555 5321 18564 5355
rect 18512 5312 18564 5321
rect 19432 5312 19484 5364
rect 2872 5244 2924 5296
rect 7564 5244 7616 5296
rect 4160 5176 4212 5228
rect 7288 5219 7340 5228
rect 7288 5185 7297 5219
rect 7297 5185 7331 5219
rect 7331 5185 7340 5219
rect 7288 5176 7340 5185
rect 10416 5219 10468 5228
rect 5540 5108 5592 5160
rect 5816 5108 5868 5160
rect 6184 5108 6236 5160
rect 7104 5108 7156 5160
rect 7748 5108 7800 5160
rect 8576 5108 8628 5160
rect 1492 4972 1544 5024
rect 4068 5040 4120 5092
rect 4436 4972 4488 5024
rect 7472 5040 7524 5092
rect 7656 5083 7708 5092
rect 7656 5049 7659 5083
rect 7659 5049 7693 5083
rect 7693 5049 7708 5083
rect 7656 5040 7708 5049
rect 8300 5040 8352 5092
rect 10416 5185 10425 5219
rect 10425 5185 10459 5219
rect 10459 5185 10468 5219
rect 10416 5176 10468 5185
rect 12072 5176 12124 5228
rect 12440 5219 12492 5228
rect 12440 5185 12449 5219
rect 12449 5185 12483 5219
rect 12483 5185 12492 5219
rect 12440 5176 12492 5185
rect 10508 5040 10560 5092
rect 19248 5287 19300 5296
rect 19248 5253 19257 5287
rect 19257 5253 19291 5287
rect 19291 5253 19300 5287
rect 19248 5244 19300 5253
rect 14188 5219 14240 5228
rect 14188 5185 14197 5219
rect 14197 5185 14231 5219
rect 14231 5185 14240 5219
rect 14188 5176 14240 5185
rect 16028 5176 16080 5228
rect 16580 5219 16632 5228
rect 16580 5185 16589 5219
rect 16589 5185 16623 5219
rect 16623 5185 16632 5219
rect 16580 5176 16632 5185
rect 18420 5176 18472 5228
rect 20444 5176 20496 5228
rect 20628 5219 20680 5228
rect 20628 5185 20637 5219
rect 20637 5185 20671 5219
rect 20671 5185 20680 5219
rect 20628 5176 20680 5185
rect 20536 5108 20588 5160
rect 16396 5083 16448 5092
rect 16396 5049 16405 5083
rect 16405 5049 16439 5083
rect 16439 5049 16448 5083
rect 16396 5040 16448 5049
rect 6644 5015 6696 5024
rect 6644 4981 6653 5015
rect 6653 4981 6687 5015
rect 6687 4981 6696 5015
rect 6644 4972 6696 4981
rect 8852 5015 8904 5024
rect 8852 4981 8861 5015
rect 8861 4981 8895 5015
rect 8895 4981 8904 5015
rect 8852 4972 8904 4981
rect 11336 5015 11388 5024
rect 11336 4981 11345 5015
rect 11345 4981 11379 5015
rect 11379 4981 11388 5015
rect 11336 4972 11388 4981
rect 15476 5015 15528 5024
rect 15476 4981 15485 5015
rect 15485 4981 15519 5015
rect 15519 4981 15528 5015
rect 18788 5083 18840 5092
rect 18788 5049 18797 5083
rect 18797 5049 18831 5083
rect 18831 5049 18840 5083
rect 18788 5040 18840 5049
rect 19892 5040 19944 5092
rect 20720 5040 20772 5092
rect 15476 4972 15528 4981
rect 17408 4972 17460 5024
rect 21548 4972 21600 5024
rect 8982 4870 9034 4922
rect 9046 4870 9098 4922
rect 9110 4870 9162 4922
rect 9174 4870 9226 4922
rect 16982 4870 17034 4922
rect 17046 4870 17098 4922
rect 17110 4870 17162 4922
rect 17174 4870 17226 4922
rect 3424 4811 3476 4820
rect 3424 4777 3433 4811
rect 3433 4777 3467 4811
rect 3467 4777 3476 4811
rect 3424 4768 3476 4777
rect 4804 4768 4856 4820
rect 7656 4768 7708 4820
rect 8208 4768 8260 4820
rect 8576 4811 8628 4820
rect 8576 4777 8585 4811
rect 8585 4777 8619 4811
rect 8619 4777 8628 4811
rect 8576 4768 8628 4777
rect 10416 4768 10468 4820
rect 12440 4811 12492 4820
rect 12440 4777 12449 4811
rect 12449 4777 12483 4811
rect 12483 4777 12492 4811
rect 12440 4768 12492 4777
rect 12808 4768 12860 4820
rect 15108 4811 15160 4820
rect 15108 4777 15117 4811
rect 15117 4777 15151 4811
rect 15151 4777 15160 4811
rect 15108 4768 15160 4777
rect 15384 4811 15436 4820
rect 15384 4777 15393 4811
rect 15393 4777 15427 4811
rect 15427 4777 15436 4811
rect 15384 4768 15436 4777
rect 16856 4768 16908 4820
rect 4436 4700 4488 4752
rect 11336 4700 11388 4752
rect 2320 4632 2372 4684
rect 2688 4675 2740 4684
rect 2688 4641 2697 4675
rect 2697 4641 2731 4675
rect 2731 4641 2740 4675
rect 4344 4675 4396 4684
rect 2688 4632 2740 4641
rect 4344 4641 4353 4675
rect 4353 4641 4387 4675
rect 4387 4641 4396 4675
rect 4344 4632 4396 4641
rect 6092 4675 6144 4684
rect 6092 4641 6101 4675
rect 6101 4641 6135 4675
rect 6135 4641 6144 4675
rect 6092 4632 6144 4641
rect 6184 4632 6236 4684
rect 6368 4632 6420 4684
rect 9772 4675 9824 4684
rect 9772 4641 9781 4675
rect 9781 4641 9815 4675
rect 9815 4641 9824 4675
rect 9772 4632 9824 4641
rect 10140 4675 10192 4684
rect 10140 4641 10149 4675
rect 10149 4641 10183 4675
rect 10183 4641 10192 4675
rect 10140 4632 10192 4641
rect 13452 4700 13504 4752
rect 15660 4700 15712 4752
rect 14096 4675 14148 4684
rect 14096 4641 14105 4675
rect 14105 4641 14139 4675
rect 14139 4641 14148 4675
rect 14096 4632 14148 4641
rect 15476 4675 15528 4684
rect 15476 4641 15485 4675
rect 15485 4641 15519 4675
rect 15519 4641 15528 4675
rect 15476 4632 15528 4641
rect 15568 4632 15620 4684
rect 16488 4700 16540 4752
rect 18788 4743 18840 4752
rect 18788 4709 18797 4743
rect 18797 4709 18831 4743
rect 18831 4709 18840 4743
rect 18788 4700 18840 4709
rect 19340 4743 19392 4752
rect 19340 4709 19349 4743
rect 19349 4709 19383 4743
rect 19383 4709 19392 4743
rect 19340 4700 19392 4709
rect 17040 4675 17092 4684
rect 17040 4641 17049 4675
rect 17049 4641 17083 4675
rect 17083 4641 17092 4675
rect 17040 4632 17092 4641
rect 17316 4675 17368 4684
rect 17316 4641 17325 4675
rect 17325 4641 17359 4675
rect 17359 4641 17368 4675
rect 17316 4632 17368 4641
rect 20812 4632 20864 4684
rect 4252 4607 4304 4616
rect 4252 4573 4261 4607
rect 4261 4573 4295 4607
rect 4295 4573 4304 4607
rect 4252 4564 4304 4573
rect 6552 4607 6604 4616
rect 6552 4573 6561 4607
rect 6561 4573 6595 4607
rect 6595 4573 6604 4607
rect 6552 4564 6604 4573
rect 10048 4564 10100 4616
rect 2504 4539 2556 4548
rect 2504 4505 2513 4539
rect 2513 4505 2547 4539
rect 2547 4505 2556 4539
rect 2504 4496 2556 4505
rect 6184 4496 6236 4548
rect 8760 4496 8812 4548
rect 8852 4496 8904 4548
rect 9128 4496 9180 4548
rect 10140 4496 10192 4548
rect 11244 4496 11296 4548
rect 13268 4564 13320 4616
rect 17592 4607 17644 4616
rect 17592 4573 17601 4607
rect 17601 4573 17635 4607
rect 17635 4573 17644 4607
rect 17592 4564 17644 4573
rect 17500 4496 17552 4548
rect 1676 4471 1728 4480
rect 1676 4437 1685 4471
rect 1685 4437 1719 4471
rect 1719 4437 1728 4471
rect 1676 4428 1728 4437
rect 3516 4428 3568 4480
rect 4712 4428 4764 4480
rect 4804 4428 4856 4480
rect 8116 4428 8168 4480
rect 8944 4428 8996 4480
rect 9220 4428 9272 4480
rect 14556 4428 14608 4480
rect 16304 4471 16356 4480
rect 16304 4437 16313 4471
rect 16313 4437 16347 4471
rect 16347 4437 16356 4471
rect 16304 4428 16356 4437
rect 4982 4326 5034 4378
rect 5046 4326 5098 4378
rect 5110 4326 5162 4378
rect 5174 4326 5226 4378
rect 12982 4326 13034 4378
rect 13046 4326 13098 4378
rect 13110 4326 13162 4378
rect 13174 4326 13226 4378
rect 20982 4326 21034 4378
rect 21046 4326 21098 4378
rect 21110 4326 21162 4378
rect 21174 4326 21226 4378
rect 1584 4267 1636 4276
rect 1584 4233 1593 4267
rect 1593 4233 1627 4267
rect 1627 4233 1636 4267
rect 1584 4224 1636 4233
rect 6552 4267 6604 4276
rect 5816 4199 5868 4208
rect 2504 4088 2556 4140
rect 1676 4020 1728 4072
rect 5816 4165 5825 4199
rect 5825 4165 5859 4199
rect 5859 4165 5868 4199
rect 5816 4156 5868 4165
rect 6552 4233 6561 4267
rect 6561 4233 6595 4267
rect 6595 4233 6604 4267
rect 6552 4224 6604 4233
rect 9680 4224 9732 4276
rect 11336 4224 11388 4276
rect 13452 4267 13504 4276
rect 7564 4156 7616 4208
rect 7656 4156 7708 4208
rect 9128 4156 9180 4208
rect 9772 4156 9824 4208
rect 13452 4233 13461 4267
rect 13461 4233 13495 4267
rect 13495 4233 13504 4267
rect 13452 4224 13504 4233
rect 14096 4267 14148 4276
rect 14096 4233 14105 4267
rect 14105 4233 14139 4267
rect 14139 4233 14148 4267
rect 14096 4224 14148 4233
rect 15568 4267 15620 4276
rect 15568 4233 15577 4267
rect 15577 4233 15611 4267
rect 15611 4233 15620 4267
rect 15568 4224 15620 4233
rect 17316 4224 17368 4276
rect 18696 4224 18748 4276
rect 18788 4224 18840 4276
rect 20168 4224 20220 4276
rect 15752 4156 15804 4208
rect 16212 4156 16264 4208
rect 17040 4156 17092 4208
rect 19708 4156 19760 4208
rect 20812 4156 20864 4208
rect 2504 3952 2556 4004
rect 3424 4088 3476 4140
rect 3976 4131 4028 4140
rect 3976 4097 3985 4131
rect 3985 4097 4019 4131
rect 4019 4097 4028 4131
rect 3976 4088 4028 4097
rect 4252 4088 4304 4140
rect 8944 4131 8996 4140
rect 3240 4063 3292 4072
rect 3240 4029 3249 4063
rect 3249 4029 3283 4063
rect 3283 4029 3292 4063
rect 3240 4020 3292 4029
rect 4804 4063 4856 4072
rect 2320 3884 2372 3936
rect 4804 4029 4813 4063
rect 4813 4029 4847 4063
rect 4847 4029 4856 4063
rect 4804 4020 4856 4029
rect 4896 4063 4948 4072
rect 4896 4029 4905 4063
rect 4905 4029 4939 4063
rect 4939 4029 4948 4063
rect 8944 4097 8953 4131
rect 8953 4097 8987 4131
rect 8987 4097 8996 4131
rect 8944 4088 8996 4097
rect 10140 4088 10192 4140
rect 16764 4131 16816 4140
rect 4896 4020 4948 4029
rect 5264 4020 5316 4072
rect 7564 4020 7616 4072
rect 10600 4020 10652 4072
rect 11888 4020 11940 4072
rect 12440 4063 12492 4072
rect 12440 4029 12449 4063
rect 12449 4029 12483 4063
rect 12483 4029 12492 4063
rect 12440 4020 12492 4029
rect 16764 4097 16773 4131
rect 16773 4097 16807 4131
rect 16807 4097 16816 4131
rect 16764 4088 16816 4097
rect 17592 4088 17644 4140
rect 18052 4131 18104 4140
rect 18052 4097 18061 4131
rect 18061 4097 18095 4131
rect 18095 4097 18104 4131
rect 18052 4088 18104 4097
rect 18788 4088 18840 4140
rect 19064 4088 19116 4140
rect 4344 3927 4396 3936
rect 4344 3893 4353 3927
rect 4353 3893 4387 3927
rect 4387 3893 4396 3927
rect 4344 3884 4396 3893
rect 6092 3884 6144 3936
rect 6276 3927 6328 3936
rect 6276 3893 6285 3927
rect 6285 3893 6319 3927
rect 6319 3893 6328 3927
rect 6276 3884 6328 3893
rect 7104 3884 7156 3936
rect 8576 3952 8628 4004
rect 9220 3952 9272 4004
rect 10140 3952 10192 4004
rect 10968 3952 11020 4004
rect 14556 3995 14608 4004
rect 9864 3927 9916 3936
rect 9864 3893 9873 3927
rect 9873 3893 9907 3927
rect 9907 3893 9916 3927
rect 9864 3884 9916 3893
rect 12348 3884 12400 3936
rect 12532 3927 12584 3936
rect 12532 3893 12541 3927
rect 12541 3893 12575 3927
rect 12575 3893 12584 3927
rect 12532 3884 12584 3893
rect 14556 3961 14565 3995
rect 14565 3961 14599 3995
rect 14599 3961 14608 3995
rect 14556 3952 14608 3961
rect 14648 3995 14700 4004
rect 14648 3961 14657 3995
rect 14657 3961 14691 3995
rect 14691 3961 14700 3995
rect 14648 3952 14700 3961
rect 16120 3995 16172 4004
rect 16120 3961 16129 3995
rect 16129 3961 16163 3995
rect 16163 3961 16172 3995
rect 16120 3952 16172 3961
rect 16304 3952 16356 4004
rect 18604 4020 18656 4072
rect 19340 4020 19392 4072
rect 18880 3952 18932 4004
rect 19892 3995 19944 4004
rect 19892 3961 19901 3995
rect 19901 3961 19935 3995
rect 19935 3961 19944 3995
rect 19892 3952 19944 3961
rect 14280 3884 14332 3936
rect 15476 3884 15528 3936
rect 17316 3884 17368 3936
rect 18972 3927 19024 3936
rect 18972 3893 18981 3927
rect 18981 3893 19015 3927
rect 19015 3893 19024 3927
rect 18972 3884 19024 3893
rect 19156 3884 19208 3936
rect 21364 3884 21416 3936
rect 8982 3782 9034 3834
rect 9046 3782 9098 3834
rect 9110 3782 9162 3834
rect 9174 3782 9226 3834
rect 16982 3782 17034 3834
rect 17046 3782 17098 3834
rect 17110 3782 17162 3834
rect 17174 3782 17226 3834
rect 2688 3680 2740 3732
rect 3424 3723 3476 3732
rect 3424 3689 3433 3723
rect 3433 3689 3467 3723
rect 3467 3689 3476 3723
rect 3424 3680 3476 3689
rect 5264 3723 5316 3732
rect 5264 3689 5273 3723
rect 5273 3689 5307 3723
rect 5307 3689 5316 3723
rect 5264 3680 5316 3689
rect 6460 3723 6512 3732
rect 6460 3689 6469 3723
rect 6469 3689 6503 3723
rect 6503 3689 6512 3723
rect 6460 3680 6512 3689
rect 7748 3723 7800 3732
rect 7748 3689 7757 3723
rect 7757 3689 7791 3723
rect 7791 3689 7800 3723
rect 7748 3680 7800 3689
rect 8300 3680 8352 3732
rect 9404 3680 9456 3732
rect 1676 3612 1728 3664
rect 6184 3612 6236 3664
rect 6644 3612 6696 3664
rect 2964 3587 3016 3596
rect 2964 3553 2973 3587
rect 2973 3553 3007 3587
rect 3007 3553 3016 3587
rect 2964 3544 3016 3553
rect 3424 3544 3476 3596
rect 4896 3587 4948 3596
rect 4896 3553 4905 3587
rect 4905 3553 4939 3587
rect 4939 3553 4948 3587
rect 4896 3544 4948 3553
rect 5724 3544 5776 3596
rect 6736 3544 6788 3596
rect 1584 3383 1636 3392
rect 1584 3349 1593 3383
rect 1593 3349 1627 3383
rect 1627 3349 1636 3383
rect 1584 3340 1636 3349
rect 4712 3383 4764 3392
rect 4712 3349 4721 3383
rect 4721 3349 4755 3383
rect 4755 3349 4764 3383
rect 4712 3340 4764 3349
rect 6368 3408 6420 3460
rect 9956 3612 10008 3664
rect 7932 3587 7984 3596
rect 7932 3553 7941 3587
rect 7941 3553 7975 3587
rect 7975 3553 7984 3587
rect 7932 3544 7984 3553
rect 8208 3587 8260 3596
rect 8208 3553 8217 3587
rect 8217 3553 8251 3587
rect 8251 3553 8260 3587
rect 8208 3544 8260 3553
rect 10140 3680 10192 3732
rect 11244 3723 11296 3732
rect 11244 3689 11253 3723
rect 11253 3689 11287 3723
rect 11287 3689 11296 3723
rect 11244 3680 11296 3689
rect 12440 3723 12492 3732
rect 12440 3689 12449 3723
rect 12449 3689 12483 3723
rect 12483 3689 12492 3723
rect 12440 3680 12492 3689
rect 14648 3680 14700 3732
rect 16304 3680 16356 3732
rect 18052 3723 18104 3732
rect 18052 3689 18061 3723
rect 18061 3689 18095 3723
rect 18095 3689 18104 3723
rect 18052 3680 18104 3689
rect 19892 3723 19944 3732
rect 19892 3689 19901 3723
rect 19901 3689 19935 3723
rect 19935 3689 19944 3723
rect 19892 3680 19944 3689
rect 10324 3655 10376 3664
rect 10324 3621 10333 3655
rect 10333 3621 10367 3655
rect 10367 3621 10376 3655
rect 10324 3612 10376 3621
rect 13360 3612 13412 3664
rect 15752 3612 15804 3664
rect 16120 3612 16172 3664
rect 16580 3612 16632 3664
rect 18420 3612 18472 3664
rect 18972 3612 19024 3664
rect 11796 3587 11848 3596
rect 11796 3553 11805 3587
rect 11805 3553 11839 3587
rect 11839 3553 11848 3587
rect 11796 3544 11848 3553
rect 15384 3544 15436 3596
rect 16672 3544 16724 3596
rect 21272 3544 21324 3596
rect 8024 3451 8076 3460
rect 8024 3417 8033 3451
rect 8033 3417 8067 3451
rect 8067 3417 8076 3451
rect 8024 3408 8076 3417
rect 11336 3476 11388 3528
rect 13268 3476 13320 3528
rect 18788 3476 18840 3528
rect 18880 3476 18932 3528
rect 13636 3408 13688 3460
rect 11796 3340 11848 3392
rect 11980 3383 12032 3392
rect 11980 3349 11989 3383
rect 11989 3349 12023 3383
rect 12023 3349 12032 3383
rect 11980 3340 12032 3349
rect 15476 3340 15528 3392
rect 17408 3340 17460 3392
rect 4982 3238 5034 3290
rect 5046 3238 5098 3290
rect 5110 3238 5162 3290
rect 5174 3238 5226 3290
rect 12982 3238 13034 3290
rect 13046 3238 13098 3290
rect 13110 3238 13162 3290
rect 13174 3238 13226 3290
rect 20982 3238 21034 3290
rect 21046 3238 21098 3290
rect 21110 3238 21162 3290
rect 21174 3238 21226 3290
rect 1676 3179 1728 3188
rect 1676 3145 1685 3179
rect 1685 3145 1719 3179
rect 1719 3145 1728 3179
rect 1676 3136 1728 3145
rect 3240 3179 3292 3188
rect 3240 3145 3249 3179
rect 3249 3145 3283 3179
rect 3283 3145 3292 3179
rect 3240 3136 3292 3145
rect 6368 3179 6420 3188
rect 6368 3145 6377 3179
rect 6377 3145 6411 3179
rect 6411 3145 6420 3179
rect 6368 3136 6420 3145
rect 10048 3179 10100 3188
rect 10048 3145 10057 3179
rect 10057 3145 10091 3179
rect 10091 3145 10100 3179
rect 13360 3179 13412 3188
rect 10048 3136 10100 3145
rect 4712 3111 4764 3120
rect 4712 3077 4721 3111
rect 4721 3077 4755 3111
rect 4755 3077 4764 3111
rect 4712 3068 4764 3077
rect 5632 3068 5684 3120
rect 7932 3068 7984 3120
rect 10508 3111 10560 3120
rect 10508 3077 10517 3111
rect 10517 3077 10551 3111
rect 10551 3077 10560 3111
rect 10508 3068 10560 3077
rect 6644 3000 6696 3052
rect 6736 3000 6788 3052
rect 7196 3000 7248 3052
rect 7748 3043 7800 3052
rect 7748 3009 7757 3043
rect 7757 3009 7791 3043
rect 7791 3009 7800 3043
rect 7748 3000 7800 3009
rect 8392 3043 8444 3052
rect 8392 3009 8401 3043
rect 8401 3009 8435 3043
rect 8435 3009 8444 3043
rect 8392 3000 8444 3009
rect 4896 2975 4948 2984
rect 4896 2941 4905 2975
rect 4905 2941 4939 2975
rect 4939 2941 4948 2975
rect 4896 2932 4948 2941
rect 5172 2932 5224 2984
rect 9404 2932 9456 2984
rect 13360 3145 13369 3179
rect 13369 3145 13403 3179
rect 13403 3145 13412 3179
rect 13360 3136 13412 3145
rect 14648 3136 14700 3188
rect 15108 3179 15160 3188
rect 15108 3145 15117 3179
rect 15117 3145 15151 3179
rect 15151 3145 15160 3179
rect 15108 3136 15160 3145
rect 15568 3136 15620 3188
rect 18420 3179 18472 3188
rect 12532 3000 12584 3052
rect 2964 2864 3016 2916
rect 5908 2864 5960 2916
rect 2320 2796 2372 2848
rect 4344 2796 4396 2848
rect 4896 2796 4948 2848
rect 5724 2839 5776 2848
rect 5724 2805 5733 2839
rect 5733 2805 5767 2839
rect 5767 2805 5776 2839
rect 7748 2864 7800 2916
rect 18420 3145 18429 3179
rect 18429 3145 18463 3179
rect 18463 3145 18472 3179
rect 18420 3136 18472 3145
rect 18696 3136 18748 3188
rect 18788 3068 18840 3120
rect 18880 3043 18932 3052
rect 5724 2796 5776 2805
rect 7656 2796 7708 2848
rect 7932 2796 7984 2848
rect 16212 2975 16264 2984
rect 16212 2941 16221 2975
rect 16221 2941 16255 2975
rect 16255 2941 16264 2975
rect 16212 2932 16264 2941
rect 18880 3009 18889 3043
rect 18889 3009 18923 3043
rect 18923 3009 18932 3043
rect 18880 3000 18932 3009
rect 19340 3000 19392 3052
rect 20076 2975 20128 2984
rect 20076 2941 20085 2975
rect 20085 2941 20119 2975
rect 20119 2941 20128 2975
rect 20076 2932 20128 2941
rect 9404 2839 9456 2848
rect 9404 2805 9413 2839
rect 9413 2805 9447 2839
rect 9447 2805 9456 2839
rect 9404 2796 9456 2805
rect 12072 2796 12124 2848
rect 15752 2864 15804 2916
rect 18604 2907 18656 2916
rect 18604 2873 18613 2907
rect 18613 2873 18647 2907
rect 18647 2873 18656 2907
rect 18604 2864 18656 2873
rect 17868 2839 17920 2848
rect 17868 2805 17877 2839
rect 17877 2805 17911 2839
rect 17911 2805 17920 2839
rect 19064 2864 19116 2916
rect 20720 2864 20772 2916
rect 20168 2839 20220 2848
rect 17868 2796 17920 2805
rect 20168 2805 20177 2839
rect 20177 2805 20211 2839
rect 20211 2805 20220 2839
rect 20168 2796 20220 2805
rect 21272 2796 21324 2848
rect 22468 2796 22520 2848
rect 8982 2694 9034 2746
rect 9046 2694 9098 2746
rect 9110 2694 9162 2746
rect 9174 2694 9226 2746
rect 16982 2694 17034 2746
rect 17046 2694 17098 2746
rect 17110 2694 17162 2746
rect 17174 2694 17226 2746
rect 3516 2635 3568 2644
rect 3516 2601 3525 2635
rect 3525 2601 3559 2635
rect 3559 2601 3568 2635
rect 3516 2592 3568 2601
rect 4896 2592 4948 2644
rect 6460 2592 6512 2644
rect 7932 2635 7984 2644
rect 4804 2524 4856 2576
rect 4896 2456 4948 2508
rect 5172 2499 5224 2508
rect 5172 2465 5181 2499
rect 5181 2465 5215 2499
rect 5215 2465 5224 2499
rect 5172 2456 5224 2465
rect 2044 2431 2096 2440
rect 2044 2397 2053 2431
rect 2053 2397 2087 2431
rect 2087 2397 2096 2431
rect 2044 2388 2096 2397
rect 112 2252 164 2304
rect 4712 2320 4764 2372
rect 7932 2601 7941 2635
rect 7941 2601 7975 2635
rect 7975 2601 7984 2635
rect 7932 2592 7984 2601
rect 10324 2592 10376 2644
rect 11336 2635 11388 2644
rect 11336 2601 11345 2635
rect 11345 2601 11379 2635
rect 11379 2601 11388 2635
rect 11336 2592 11388 2601
rect 11796 2592 11848 2644
rect 12072 2592 12124 2644
rect 10508 2524 10560 2576
rect 13360 2592 13412 2644
rect 15384 2592 15436 2644
rect 17868 2592 17920 2644
rect 13728 2524 13780 2576
rect 7656 2456 7708 2508
rect 8208 2456 8260 2508
rect 9864 2456 9916 2508
rect 14556 2524 14608 2576
rect 15752 2524 15804 2576
rect 17316 2524 17368 2576
rect 20168 2592 20220 2644
rect 19064 2567 19116 2576
rect 8392 2388 8444 2440
rect 12348 2388 12400 2440
rect 15292 2456 15344 2508
rect 19064 2533 19073 2567
rect 19073 2533 19107 2567
rect 19107 2533 19116 2567
rect 19064 2524 19116 2533
rect 19156 2567 19208 2576
rect 19156 2533 19165 2567
rect 19165 2533 19199 2567
rect 19199 2533 19208 2567
rect 20076 2567 20128 2576
rect 19156 2524 19208 2533
rect 20076 2533 20085 2567
rect 20085 2533 20119 2567
rect 20119 2533 20128 2567
rect 20076 2524 20128 2533
rect 20444 2456 20496 2508
rect 14280 2388 14332 2440
rect 7564 2320 7616 2372
rect 13268 2363 13320 2372
rect 13268 2329 13277 2363
rect 13277 2329 13311 2363
rect 13311 2329 13320 2363
rect 13268 2320 13320 2329
rect 15108 2388 15160 2440
rect 19064 2388 19116 2440
rect 8024 2252 8076 2304
rect 12440 2252 12492 2304
rect 12716 2252 12768 2304
rect 18236 2320 18288 2372
rect 18604 2320 18656 2372
rect 18880 2252 18932 2304
rect 4982 2150 5034 2202
rect 5046 2150 5098 2202
rect 5110 2150 5162 2202
rect 5174 2150 5226 2202
rect 12982 2150 13034 2202
rect 13046 2150 13098 2202
rect 13110 2150 13162 2202
rect 13174 2150 13226 2202
rect 20982 2150 21034 2202
rect 21046 2150 21098 2202
rect 21110 2150 21162 2202
rect 21174 2150 21226 2202
rect 11980 1708 12032 1760
rect 17040 1708 17092 1760
rect 13820 76 13872 128
rect 14464 76 14516 128
<< metal2 >>
rect 662 23610 718 24000
rect 584 23582 718 23610
rect 584 21146 612 23582
rect 662 23520 718 23582
rect 1950 23610 2006 24000
rect 3330 23610 3386 24000
rect 4618 23610 4674 24000
rect 1950 23582 2268 23610
rect 1950 23520 2006 23582
rect 1582 22672 1638 22681
rect 1582 22607 1638 22616
rect 572 21140 624 21146
rect 572 21082 624 21088
rect 110 20360 166 20369
rect 110 20295 166 20304
rect 124 19990 152 20295
rect 1596 20058 1624 22607
rect 1858 21312 1914 21321
rect 1858 21247 1914 21256
rect 1872 20398 1900 21247
rect 2240 20398 2268 23582
rect 3068 23582 3386 23610
rect 1860 20392 1912 20398
rect 1860 20334 1912 20340
rect 2228 20392 2280 20398
rect 2228 20334 2280 20340
rect 2504 20256 2556 20262
rect 2780 20256 2832 20262
rect 2504 20198 2556 20204
rect 2700 20216 2780 20244
rect 1584 20052 1636 20058
rect 1584 19994 1636 20000
rect 112 19984 164 19990
rect 112 19926 164 19932
rect 1596 19378 1624 19994
rect 2136 19916 2188 19922
rect 2136 19858 2188 19864
rect 2044 19712 2096 19718
rect 2044 19654 2096 19660
rect 1584 19372 1636 19378
rect 1584 19314 1636 19320
rect 110 19000 166 19009
rect 166 18970 244 18986
rect 166 18964 256 18970
rect 166 18958 204 18964
rect 110 18935 166 18944
rect 204 18906 256 18912
rect 1952 18828 2004 18834
rect 1952 18770 2004 18776
rect 1964 18426 1992 18770
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 112 18080 164 18086
rect 112 18022 164 18028
rect 124 17649 152 18022
rect 110 17640 166 17649
rect 110 17575 166 17584
rect 1952 17536 2004 17542
rect 1952 17478 2004 17484
rect 1964 17066 1992 17478
rect 1952 17060 2004 17066
rect 1952 17002 2004 17008
rect 1964 16794 1992 17002
rect 1952 16788 2004 16794
rect 1952 16730 2004 16736
rect 112 16244 164 16250
rect 112 16186 164 16192
rect 124 16153 152 16186
rect 110 16144 166 16153
rect 2056 16114 2084 19654
rect 2148 19514 2176 19858
rect 2136 19508 2188 19514
rect 2136 19450 2188 19456
rect 2516 19281 2544 20198
rect 2502 19272 2558 19281
rect 2502 19207 2558 19216
rect 2504 18760 2556 18766
rect 2504 18702 2556 18708
rect 2320 18216 2372 18222
rect 2320 18158 2372 18164
rect 2228 17740 2280 17746
rect 2228 17682 2280 17688
rect 2240 16726 2268 17682
rect 2332 17202 2360 18158
rect 2516 17338 2544 18702
rect 2504 17332 2556 17338
rect 2504 17274 2556 17280
rect 2320 17196 2372 17202
rect 2320 17138 2372 17144
rect 2228 16720 2280 16726
rect 2228 16662 2280 16668
rect 2332 16590 2360 17138
rect 2320 16584 2372 16590
rect 2320 16526 2372 16532
rect 2412 16516 2464 16522
rect 2412 16458 2464 16464
rect 2424 16114 2452 16458
rect 110 16079 166 16088
rect 2044 16108 2096 16114
rect 2044 16050 2096 16056
rect 2412 16108 2464 16114
rect 2412 16050 2464 16056
rect 1860 15904 1912 15910
rect 1860 15846 1912 15852
rect 1872 15706 1900 15846
rect 2056 15706 2084 16050
rect 1860 15700 1912 15706
rect 1860 15642 1912 15648
rect 2044 15700 2096 15706
rect 2044 15642 2096 15648
rect 2424 15094 2452 16050
rect 2596 15904 2648 15910
rect 2596 15846 2648 15852
rect 2504 15564 2556 15570
rect 2504 15506 2556 15512
rect 2412 15088 2464 15094
rect 2412 15030 2464 15036
rect 2516 14822 2544 15506
rect 2504 14816 2556 14822
rect 2504 14758 2556 14764
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 1964 13802 1992 14554
rect 2516 14074 2544 14758
rect 2608 14618 2636 15846
rect 2596 14612 2648 14618
rect 2596 14554 2648 14560
rect 2504 14068 2556 14074
rect 2504 14010 2556 14016
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 1952 13796 2004 13802
rect 1952 13738 2004 13744
rect 112 13524 164 13530
rect 112 13466 164 13472
rect 124 13433 152 13466
rect 110 13424 166 13433
rect 110 13359 166 13368
rect 1676 13388 1728 13394
rect 1676 13330 1728 13336
rect 1688 12102 1716 13330
rect 1964 13190 1992 13738
rect 2056 13190 2084 13806
rect 1952 13184 2004 13190
rect 1952 13126 2004 13132
rect 2044 13184 2096 13190
rect 2044 13126 2096 13132
rect 2320 13184 2372 13190
rect 2320 13126 2372 13132
rect 1676 12096 1728 12102
rect 1676 12038 1728 12044
rect 1582 11384 1638 11393
rect 1582 11319 1638 11328
rect 1596 10810 1624 11319
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 1582 10296 1638 10305
rect 1688 10266 1716 12038
rect 1964 11778 1992 13126
rect 2136 12096 2188 12102
rect 2136 12038 2188 12044
rect 2148 11898 2176 12038
rect 2136 11892 2188 11898
rect 2136 11834 2188 11840
rect 1964 11750 2176 11778
rect 2044 11552 2096 11558
rect 2044 11494 2096 11500
rect 2056 10470 2084 11494
rect 2148 11354 2176 11750
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 2148 10810 2176 11290
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 2228 10600 2280 10606
rect 2228 10542 2280 10548
rect 2044 10464 2096 10470
rect 2044 10406 2096 10412
rect 1582 10231 1638 10240
rect 1676 10260 1728 10266
rect 1596 9994 1624 10231
rect 1676 10202 1728 10208
rect 1584 9988 1636 9994
rect 1584 9930 1636 9936
rect 1952 9512 2004 9518
rect 1952 9454 2004 9460
rect 1768 9376 1820 9382
rect 1768 9318 1820 9324
rect 1582 8664 1638 8673
rect 1582 8599 1638 8608
rect 1596 7546 1624 8599
rect 1780 8498 1808 9318
rect 1964 9042 1992 9454
rect 1952 9036 2004 9042
rect 1952 8978 2004 8984
rect 1768 8492 1820 8498
rect 1768 8434 1820 8440
rect 1964 8430 1992 8978
rect 1952 8424 2004 8430
rect 1952 8366 2004 8372
rect 1952 7948 2004 7954
rect 1952 7890 2004 7896
rect 1964 7750 1992 7890
rect 1952 7744 2004 7750
rect 1952 7686 2004 7692
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 1492 7404 1544 7410
rect 1492 7346 1544 7352
rect 1504 7313 1532 7346
rect 1490 7304 1546 7313
rect 1490 7239 1546 7248
rect 1504 7002 1532 7239
rect 1964 7206 1992 7686
rect 1952 7200 2004 7206
rect 1858 7168 1914 7177
rect 1952 7142 2004 7148
rect 1858 7103 1914 7112
rect 1492 6996 1544 7002
rect 1492 6938 1544 6944
rect 664 6384 716 6390
rect 664 6326 716 6332
rect 112 2304 164 2310
rect 112 2246 164 2252
rect 124 2145 152 2246
rect 110 2136 166 2145
rect 110 2071 166 2080
rect 386 82 442 480
rect 676 82 704 6326
rect 1872 6254 1900 7103
rect 1860 6248 1912 6254
rect 1860 6190 1912 6196
rect 1492 5024 1544 5030
rect 1492 4966 1544 4972
rect 386 54 704 82
rect 1214 82 1270 480
rect 1504 82 1532 4966
rect 1676 4480 1728 4486
rect 1582 4448 1638 4457
rect 1676 4422 1728 4428
rect 1582 4383 1638 4392
rect 1596 4282 1624 4383
rect 1584 4276 1636 4282
rect 1584 4218 1636 4224
rect 1688 4078 1716 4422
rect 2056 4154 2084 10406
rect 2136 8424 2188 8430
rect 2136 8366 2188 8372
rect 2148 7954 2176 8366
rect 2136 7948 2188 7954
rect 2136 7890 2188 7896
rect 2240 6905 2268 10542
rect 2332 9382 2360 13126
rect 2596 12776 2648 12782
rect 2596 12718 2648 12724
rect 2504 12640 2556 12646
rect 2504 12582 2556 12588
rect 2516 12374 2544 12582
rect 2504 12368 2556 12374
rect 2504 12310 2556 12316
rect 2516 11898 2544 12310
rect 2504 11892 2556 11898
rect 2504 11834 2556 11840
rect 2608 11626 2636 12718
rect 2504 11620 2556 11626
rect 2504 11562 2556 11568
rect 2596 11620 2648 11626
rect 2596 11562 2648 11568
rect 2516 11354 2544 11562
rect 2504 11348 2556 11354
rect 2504 11290 2556 11296
rect 2516 10810 2544 11290
rect 2608 11218 2636 11562
rect 2596 11212 2648 11218
rect 2596 11154 2648 11160
rect 2504 10804 2556 10810
rect 2504 10746 2556 10752
rect 2412 9988 2464 9994
rect 2412 9930 2464 9936
rect 2424 9518 2452 9930
rect 2504 9920 2556 9926
rect 2504 9862 2556 9868
rect 2596 9920 2648 9926
rect 2596 9862 2648 9868
rect 2516 9518 2544 9862
rect 2608 9586 2636 9862
rect 2596 9580 2648 9586
rect 2596 9522 2648 9528
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 2504 9512 2556 9518
rect 2504 9454 2556 9460
rect 2320 9376 2372 9382
rect 2320 9318 2372 9324
rect 2320 9036 2372 9042
rect 2424 9024 2452 9454
rect 2516 9042 2544 9454
rect 2372 8996 2452 9024
rect 2504 9036 2556 9042
rect 2320 8978 2372 8984
rect 2504 8978 2556 8984
rect 2332 8090 2360 8978
rect 2516 8430 2544 8978
rect 2504 8424 2556 8430
rect 2504 8366 2556 8372
rect 2320 8084 2372 8090
rect 2320 8026 2372 8032
rect 2516 7546 2544 8366
rect 2700 7546 2728 20216
rect 2780 20198 2832 20204
rect 3068 19922 3096 23582
rect 3330 23520 3386 23582
rect 4356 23582 4674 23610
rect 4356 20602 4384 23582
rect 4618 23520 4674 23582
rect 5998 23610 6054 24000
rect 7286 23610 7342 24000
rect 8666 23610 8722 24000
rect 5998 23582 6224 23610
rect 5998 23520 6054 23582
rect 4956 21788 5252 21808
rect 5012 21786 5036 21788
rect 5092 21786 5116 21788
rect 5172 21786 5196 21788
rect 5034 21734 5036 21786
rect 5098 21734 5110 21786
rect 5172 21734 5174 21786
rect 5012 21732 5036 21734
rect 5092 21732 5116 21734
rect 5172 21732 5196 21734
rect 4956 21712 5252 21732
rect 4956 20700 5252 20720
rect 5012 20698 5036 20700
rect 5092 20698 5116 20700
rect 5172 20698 5196 20700
rect 5034 20646 5036 20698
rect 5098 20646 5110 20698
rect 5172 20646 5174 20698
rect 5012 20644 5036 20646
rect 5092 20644 5116 20646
rect 5172 20644 5196 20646
rect 4956 20624 5252 20644
rect 4344 20596 4396 20602
rect 4344 20538 4396 20544
rect 3700 20392 3752 20398
rect 3700 20334 3752 20340
rect 3712 20262 3740 20334
rect 3700 20256 3752 20262
rect 3700 20198 3752 20204
rect 3056 19916 3108 19922
rect 3056 19858 3108 19864
rect 2780 18080 2832 18086
rect 2780 18022 2832 18028
rect 2792 13530 2820 18022
rect 2872 17128 2924 17134
rect 2872 17070 2924 17076
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2884 11558 2912 17070
rect 2964 16992 3016 16998
rect 2964 16934 3016 16940
rect 3516 16992 3568 16998
rect 3516 16934 3568 16940
rect 2976 16726 3004 16934
rect 2964 16720 3016 16726
rect 2964 16662 3016 16668
rect 2976 15910 3004 16662
rect 2964 15904 3016 15910
rect 2964 15846 3016 15852
rect 3528 15638 3556 16934
rect 3516 15632 3568 15638
rect 3516 15574 3568 15580
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 3252 13802 3280 14350
rect 3422 14240 3478 14249
rect 3422 14175 3478 14184
rect 3240 13796 3292 13802
rect 3240 13738 3292 13744
rect 3148 13388 3200 13394
rect 3148 13330 3200 13336
rect 3160 12646 3188 13330
rect 3148 12640 3200 12646
rect 3148 12582 3200 12588
rect 3056 12164 3108 12170
rect 3056 12106 3108 12112
rect 3068 11830 3096 12106
rect 3160 11830 3188 12582
rect 3056 11824 3108 11830
rect 3056 11766 3108 11772
rect 3148 11824 3200 11830
rect 3148 11766 3200 11772
rect 2872 11552 2924 11558
rect 2872 11494 2924 11500
rect 3148 9512 3200 9518
rect 3148 9454 3200 9460
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 2976 8090 3004 8978
rect 3160 8498 3188 9454
rect 3252 9110 3280 13738
rect 3332 11144 3384 11150
rect 3332 11086 3384 11092
rect 3344 10470 3372 11086
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 3240 9104 3292 9110
rect 3240 9046 3292 9052
rect 3344 8498 3372 10406
rect 3436 8537 3464 14175
rect 3712 13814 3740 20198
rect 4956 19612 5252 19632
rect 5012 19610 5036 19612
rect 5092 19610 5116 19612
rect 5172 19610 5196 19612
rect 5034 19558 5036 19610
rect 5098 19558 5110 19610
rect 5172 19558 5174 19610
rect 5012 19556 5036 19558
rect 5092 19556 5116 19558
rect 5172 19556 5196 19558
rect 4956 19536 5252 19556
rect 5264 19236 5316 19242
rect 5264 19178 5316 19184
rect 5276 18902 5304 19178
rect 5264 18896 5316 18902
rect 5448 18896 5500 18902
rect 5316 18856 5396 18884
rect 5264 18838 5316 18844
rect 4956 18524 5252 18544
rect 5012 18522 5036 18524
rect 5092 18522 5116 18524
rect 5172 18522 5196 18524
rect 5034 18470 5036 18522
rect 5098 18470 5110 18522
rect 5172 18470 5174 18522
rect 5012 18468 5036 18470
rect 5092 18468 5116 18470
rect 5172 18468 5196 18470
rect 4956 18448 5252 18468
rect 5368 18426 5396 18856
rect 5448 18838 5500 18844
rect 5356 18420 5408 18426
rect 5356 18362 5408 18368
rect 5460 18358 5488 18838
rect 5448 18352 5500 18358
rect 5448 18294 5500 18300
rect 4528 18080 4580 18086
rect 4528 18022 4580 18028
rect 4252 17128 4304 17134
rect 4252 17070 4304 17076
rect 4264 16794 4292 17070
rect 4344 16992 4396 16998
rect 4344 16934 4396 16940
rect 4252 16788 4304 16794
rect 4252 16730 4304 16736
rect 4160 16652 4212 16658
rect 4160 16594 4212 16600
rect 4172 16522 4200 16594
rect 4160 16516 4212 16522
rect 4160 16458 4212 16464
rect 3884 16448 3936 16454
rect 3884 16390 3936 16396
rect 3896 16182 3924 16390
rect 3884 16176 3936 16182
rect 3884 16118 3936 16124
rect 3896 15978 3924 16118
rect 4172 16114 4200 16458
rect 4160 16108 4212 16114
rect 4160 16050 4212 16056
rect 4356 16046 4384 16934
rect 4344 16040 4396 16046
rect 4396 16000 4476 16028
rect 4344 15982 4396 15988
rect 3884 15972 3936 15978
rect 3884 15914 3936 15920
rect 4448 15910 4476 16000
rect 4436 15904 4488 15910
rect 4436 15846 4488 15852
rect 4252 15632 4304 15638
rect 4252 15574 4304 15580
rect 4344 15632 4396 15638
rect 4344 15574 4396 15580
rect 4264 15502 4292 15574
rect 4252 15496 4304 15502
rect 4252 15438 4304 15444
rect 3792 14816 3844 14822
rect 3792 14758 3844 14764
rect 3620 13786 3740 13814
rect 3620 10606 3648 13786
rect 3700 13388 3752 13394
rect 3700 13330 3752 13336
rect 3712 12646 3740 13330
rect 3804 12782 3832 14758
rect 4264 14618 4292 15438
rect 4356 15162 4384 15574
rect 4344 15156 4396 15162
rect 4344 15098 4396 15104
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 3884 14408 3936 14414
rect 3884 14350 3936 14356
rect 3792 12776 3844 12782
rect 3792 12718 3844 12724
rect 3700 12640 3752 12646
rect 3700 12582 3752 12588
rect 3712 11801 3740 12582
rect 3698 11792 3754 11801
rect 3698 11727 3754 11736
rect 3608 10600 3660 10606
rect 3608 10542 3660 10548
rect 3896 10266 3924 14350
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 4264 13938 4292 14214
rect 4252 13932 4304 13938
rect 4252 13874 4304 13880
rect 4264 13530 4292 13874
rect 4448 13870 4476 15846
rect 4540 15162 4568 18022
rect 4712 17740 4764 17746
rect 4712 17682 4764 17688
rect 4620 17672 4672 17678
rect 4620 17614 4672 17620
rect 4632 16114 4660 17614
rect 4724 17134 4752 17682
rect 4956 17436 5252 17456
rect 5012 17434 5036 17436
rect 5092 17434 5116 17436
rect 5172 17434 5196 17436
rect 5034 17382 5036 17434
rect 5098 17382 5110 17434
rect 5172 17382 5174 17434
rect 5012 17380 5036 17382
rect 5092 17380 5116 17382
rect 5172 17380 5196 17382
rect 4956 17360 5252 17380
rect 4712 17128 4764 17134
rect 4712 17070 4764 17076
rect 4724 16658 4752 17070
rect 5460 16794 5488 18294
rect 5632 17808 5684 17814
rect 5632 17750 5684 17756
rect 5644 17066 5672 17750
rect 6092 17672 6144 17678
rect 6092 17614 6144 17620
rect 6104 17066 6132 17614
rect 5632 17060 5684 17066
rect 5632 17002 5684 17008
rect 6092 17060 6144 17066
rect 6092 17002 6144 17008
rect 5448 16788 5500 16794
rect 5448 16730 5500 16736
rect 4712 16652 4764 16658
rect 4712 16594 4764 16600
rect 6092 16652 6144 16658
rect 6092 16594 6144 16600
rect 4620 16108 4672 16114
rect 4620 16050 4672 16056
rect 4620 15972 4672 15978
rect 4724 15960 4752 16594
rect 4956 16348 5252 16368
rect 5012 16346 5036 16348
rect 5092 16346 5116 16348
rect 5172 16346 5196 16348
rect 5034 16294 5036 16346
rect 5098 16294 5110 16346
rect 5172 16294 5174 16346
rect 5012 16292 5036 16294
rect 5092 16292 5116 16294
rect 5172 16292 5196 16294
rect 4956 16272 5252 16292
rect 5356 16244 5408 16250
rect 5356 16186 5408 16192
rect 4672 15932 4752 15960
rect 4620 15914 4672 15920
rect 4528 15156 4580 15162
rect 4528 15098 4580 15104
rect 4436 13864 4488 13870
rect 4436 13806 4488 13812
rect 4252 13524 4304 13530
rect 4252 13466 4304 13472
rect 4448 12918 4476 13806
rect 4724 13394 4752 15932
rect 5368 15706 5396 16186
rect 6104 16182 6132 16594
rect 6092 16176 6144 16182
rect 6092 16118 6144 16124
rect 6104 15910 6132 16118
rect 6092 15904 6144 15910
rect 6092 15846 6144 15852
rect 5356 15700 5408 15706
rect 5356 15642 5408 15648
rect 4804 15428 4856 15434
rect 4804 15370 4856 15376
rect 4816 15094 4844 15370
rect 4956 15260 5252 15280
rect 5012 15258 5036 15260
rect 5092 15258 5116 15260
rect 5172 15258 5196 15260
rect 5034 15206 5036 15258
rect 5098 15206 5110 15258
rect 5172 15206 5174 15258
rect 5012 15204 5036 15206
rect 5092 15204 5116 15206
rect 5172 15204 5196 15206
rect 4956 15184 5252 15204
rect 4804 15088 4856 15094
rect 4804 15030 4856 15036
rect 4816 14550 4844 15030
rect 5368 14890 5396 15642
rect 6104 15434 6132 15846
rect 6092 15428 6144 15434
rect 6092 15370 6144 15376
rect 5356 14884 5408 14890
rect 5356 14826 5408 14832
rect 4804 14544 4856 14550
rect 4804 14486 4856 14492
rect 5356 14544 5408 14550
rect 5356 14486 5408 14492
rect 4816 13734 4844 14486
rect 4956 14172 5252 14192
rect 5012 14170 5036 14172
rect 5092 14170 5116 14172
rect 5172 14170 5196 14172
rect 5034 14118 5036 14170
rect 5098 14118 5110 14170
rect 5172 14118 5174 14170
rect 5012 14116 5036 14118
rect 5092 14116 5116 14118
rect 5172 14116 5196 14118
rect 4956 14096 5252 14116
rect 5368 14074 5396 14486
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 6196 14006 6224 23582
rect 7286 23582 7604 23610
rect 7286 23520 7342 23582
rect 6460 21140 6512 21146
rect 6460 21082 6512 21088
rect 6472 20330 6500 21082
rect 6460 20324 6512 20330
rect 6460 20266 6512 20272
rect 6276 18080 6328 18086
rect 6276 18022 6328 18028
rect 6288 17882 6316 18022
rect 6276 17876 6328 17882
rect 6276 17818 6328 17824
rect 6276 16448 6328 16454
rect 6276 16390 6328 16396
rect 6288 15638 6316 16390
rect 6276 15632 6328 15638
rect 6276 15574 6328 15580
rect 6288 15162 6316 15574
rect 6276 15156 6328 15162
rect 6276 15098 6328 15104
rect 6368 14476 6420 14482
rect 6368 14418 6420 14424
rect 6380 14278 6408 14418
rect 6276 14272 6328 14278
rect 6276 14214 6328 14220
rect 6368 14272 6420 14278
rect 6368 14214 6420 14220
rect 6184 14000 6236 14006
rect 6184 13942 6236 13948
rect 4804 13728 4856 13734
rect 4804 13670 4856 13676
rect 5632 13728 5684 13734
rect 5632 13670 5684 13676
rect 5644 13530 5672 13670
rect 5632 13524 5684 13530
rect 5632 13466 5684 13472
rect 4712 13388 4764 13394
rect 4712 13330 4764 13336
rect 4436 12912 4488 12918
rect 4436 12854 4488 12860
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 4080 10810 4108 11086
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 3884 10260 3936 10266
rect 3884 10202 3936 10208
rect 3976 10192 4028 10198
rect 3976 10134 4028 10140
rect 3988 9994 4016 10134
rect 4172 10130 4200 12718
rect 4724 12714 4752 13330
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 4956 13084 5252 13104
rect 5012 13082 5036 13084
rect 5092 13082 5116 13084
rect 5172 13082 5196 13084
rect 5034 13030 5036 13082
rect 5098 13030 5110 13082
rect 5172 13030 5174 13082
rect 5012 13028 5036 13030
rect 5092 13028 5116 13030
rect 5172 13028 5196 13030
rect 4956 13008 5252 13028
rect 5368 12782 5396 13126
rect 6288 12986 6316 14214
rect 6472 13814 6500 20266
rect 7380 20256 7432 20262
rect 7380 20198 7432 20204
rect 7392 19922 7420 20198
rect 7380 19916 7432 19922
rect 7380 19858 7432 19864
rect 6828 19712 6880 19718
rect 6828 19654 6880 19660
rect 6840 19174 6868 19654
rect 7392 19514 7420 19858
rect 7380 19508 7432 19514
rect 7380 19450 7432 19456
rect 7012 19440 7064 19446
rect 7012 19382 7064 19388
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 6644 18896 6696 18902
rect 6644 18838 6696 18844
rect 6826 18864 6882 18873
rect 6656 18426 6684 18838
rect 6826 18799 6882 18808
rect 6840 18766 6868 18799
rect 6828 18760 6880 18766
rect 6828 18702 6880 18708
rect 6644 18420 6696 18426
rect 6644 18362 6696 18368
rect 6552 17128 6604 17134
rect 6552 17070 6604 17076
rect 6564 16726 6592 17070
rect 6552 16720 6604 16726
rect 6552 16662 6604 16668
rect 6656 16250 6684 18362
rect 6840 17814 6868 18702
rect 6932 18698 6960 19314
rect 7024 19242 7052 19382
rect 7012 19236 7064 19242
rect 7012 19178 7064 19184
rect 6920 18692 6972 18698
rect 6920 18634 6972 18640
rect 6932 18290 6960 18634
rect 6920 18284 6972 18290
rect 6920 18226 6972 18232
rect 6932 17882 6960 18226
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6828 17808 6880 17814
rect 6828 17750 6880 17756
rect 7024 17338 7052 19178
rect 7380 19168 7432 19174
rect 7380 19110 7432 19116
rect 7392 18329 7420 19110
rect 7576 18834 7604 23582
rect 8404 23582 8722 23610
rect 8404 20602 8432 23582
rect 8666 23520 8722 23582
rect 9954 23610 10010 24000
rect 11334 23610 11390 24000
rect 12622 23610 12678 24000
rect 14002 23610 14058 24000
rect 15290 23610 15346 24000
rect 16670 23610 16726 24000
rect 17958 23610 18014 24000
rect 19338 23610 19394 24000
rect 9954 23582 10180 23610
rect 9954 23520 10010 23582
rect 8956 21244 9252 21264
rect 9012 21242 9036 21244
rect 9092 21242 9116 21244
rect 9172 21242 9196 21244
rect 9034 21190 9036 21242
rect 9098 21190 9110 21242
rect 9172 21190 9174 21242
rect 9012 21188 9036 21190
rect 9092 21188 9116 21190
rect 9172 21188 9196 21190
rect 8956 21168 9252 21188
rect 8668 20800 8720 20806
rect 8668 20742 8720 20748
rect 8392 20596 8444 20602
rect 8392 20538 8444 20544
rect 8680 20466 8708 20742
rect 10152 20602 10180 23582
rect 11334 23582 11468 23610
rect 11334 23520 11390 23582
rect 11440 21146 11468 23582
rect 12622 23582 12756 23610
rect 12622 23520 12678 23582
rect 11428 21140 11480 21146
rect 11428 21082 11480 21088
rect 11060 21004 11112 21010
rect 11060 20946 11112 20952
rect 10140 20596 10192 20602
rect 10140 20538 10192 20544
rect 8668 20460 8720 20466
rect 8668 20402 8720 20408
rect 7840 20256 7892 20262
rect 7840 20198 7892 20204
rect 7564 18828 7616 18834
rect 7484 18788 7564 18816
rect 7378 18320 7434 18329
rect 7378 18255 7434 18264
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 7012 17332 7064 17338
rect 7012 17274 7064 17280
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 6644 16244 6696 16250
rect 6644 16186 6696 16192
rect 6748 14550 6776 16730
rect 7024 15638 7052 17274
rect 7116 17134 7144 17478
rect 7104 17128 7156 17134
rect 7104 17070 7156 17076
rect 7196 17128 7248 17134
rect 7196 17070 7248 17076
rect 7116 16658 7144 17070
rect 7208 16726 7236 17070
rect 7196 16720 7248 16726
rect 7196 16662 7248 16668
rect 7104 16652 7156 16658
rect 7104 16594 7156 16600
rect 7208 16046 7236 16662
rect 7196 16040 7248 16046
rect 7196 15982 7248 15988
rect 7012 15632 7064 15638
rect 7012 15574 7064 15580
rect 7024 15162 7052 15574
rect 7380 15496 7432 15502
rect 7380 15438 7432 15444
rect 7012 15156 7064 15162
rect 7012 15098 7064 15104
rect 7392 15094 7420 15438
rect 7380 15088 7432 15094
rect 7380 15030 7432 15036
rect 7288 14884 7340 14890
rect 7288 14826 7340 14832
rect 7300 14618 7328 14826
rect 7288 14612 7340 14618
rect 7288 14554 7340 14560
rect 6736 14544 6788 14550
rect 6736 14486 6788 14492
rect 6748 14074 6776 14486
rect 6828 14408 6880 14414
rect 6828 14350 6880 14356
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 6472 13786 6776 13814
rect 6644 13524 6696 13530
rect 6644 13466 6696 13472
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 6276 12980 6328 12986
rect 6276 12922 6328 12928
rect 6380 12782 6408 13262
rect 6656 12918 6684 13466
rect 6644 12912 6696 12918
rect 6644 12854 6696 12860
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 6368 12776 6420 12782
rect 6368 12718 6420 12724
rect 6644 12776 6696 12782
rect 6644 12718 6696 12724
rect 4712 12708 4764 12714
rect 4712 12650 4764 12656
rect 6380 12442 6408 12718
rect 6368 12436 6420 12442
rect 6368 12378 6420 12384
rect 5356 12368 5408 12374
rect 5356 12310 5408 12316
rect 4344 12164 4396 12170
rect 4344 12106 4396 12112
rect 4356 11762 4384 12106
rect 4956 11996 5252 12016
rect 5012 11994 5036 11996
rect 5092 11994 5116 11996
rect 5172 11994 5196 11996
rect 5034 11942 5036 11994
rect 5098 11942 5110 11994
rect 5172 11942 5174 11994
rect 5012 11940 5036 11942
rect 5092 11940 5116 11942
rect 5172 11940 5196 11942
rect 4956 11920 5252 11940
rect 4344 11756 4396 11762
rect 4344 11698 4396 11704
rect 4804 11620 4856 11626
rect 4804 11562 4856 11568
rect 4816 11354 4844 11562
rect 5368 11558 5396 12310
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 5448 12164 5500 12170
rect 5448 12106 5500 12112
rect 5460 11762 5488 12106
rect 5644 11898 5672 12174
rect 6656 12102 6684 12718
rect 6644 12096 6696 12102
rect 6644 12038 6696 12044
rect 5632 11892 5684 11898
rect 5632 11834 5684 11840
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5460 11665 5488 11698
rect 5446 11656 5502 11665
rect 5446 11591 5502 11600
rect 5356 11552 5408 11558
rect 5356 11494 5408 11500
rect 4436 11348 4488 11354
rect 4436 11290 4488 11296
rect 4804 11348 4856 11354
rect 4804 11290 4856 11296
rect 4448 10266 4476 11290
rect 4816 10606 4844 11290
rect 4956 10908 5252 10928
rect 5012 10906 5036 10908
rect 5092 10906 5116 10908
rect 5172 10906 5196 10908
rect 5034 10854 5036 10906
rect 5098 10854 5110 10906
rect 5172 10854 5174 10906
rect 5012 10852 5036 10854
rect 5092 10852 5116 10854
rect 5172 10852 5196 10854
rect 4956 10832 5252 10852
rect 5368 10674 5396 11494
rect 5644 11354 5672 11834
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 6656 11286 6684 12038
rect 6644 11280 6696 11286
rect 6644 11222 6696 11228
rect 6276 11076 6328 11082
rect 6276 11018 6328 11024
rect 6288 10810 6316 11018
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4712 10532 4764 10538
rect 4712 10474 4764 10480
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 4436 10260 4488 10266
rect 4436 10202 4488 10208
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 4160 10124 4212 10130
rect 4160 10066 4212 10072
rect 3976 9988 4028 9994
rect 3976 9930 4028 9936
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3804 9518 3832 9862
rect 4080 9625 4108 10066
rect 4066 9616 4122 9625
rect 4066 9551 4122 9560
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 3804 9178 3832 9454
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 3792 9172 3844 9178
rect 3792 9114 3844 9120
rect 3422 8528 3478 8537
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 3332 8492 3384 8498
rect 3422 8463 3478 8472
rect 3332 8434 3384 8440
rect 3804 8090 3832 9114
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 3988 8634 4016 8910
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3792 8084 3844 8090
rect 3792 8026 3844 8032
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 2688 7540 2740 7546
rect 2688 7482 2740 7488
rect 2596 7200 2648 7206
rect 2596 7142 2648 7148
rect 2226 6896 2282 6905
rect 2226 6831 2282 6840
rect 2412 6860 2464 6866
rect 2412 6802 2464 6808
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 2424 5574 2452 6802
rect 2516 6118 2544 6802
rect 2504 6112 2556 6118
rect 2504 6054 2556 6060
rect 2516 5846 2544 6054
rect 2504 5840 2556 5846
rect 2504 5782 2556 5788
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2320 4684 2372 4690
rect 2320 4626 2372 4632
rect 1964 4126 2084 4154
rect 1676 4072 1728 4078
rect 1676 4014 1728 4020
rect 1676 3664 1728 3670
rect 1676 3606 1728 3612
rect 1584 3392 1636 3398
rect 1584 3334 1636 3340
rect 1596 3233 1624 3334
rect 1582 3224 1638 3233
rect 1688 3194 1716 3606
rect 1582 3159 1638 3168
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 1964 1329 1992 4126
rect 2332 3942 2360 4626
rect 2504 4548 2556 4554
rect 2504 4490 2556 4496
rect 2516 4146 2544 4490
rect 2504 4140 2556 4146
rect 2504 4082 2556 4088
rect 2516 4010 2544 4082
rect 2504 4004 2556 4010
rect 2504 3946 2556 3952
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 2332 2854 2360 3878
rect 2320 2848 2372 2854
rect 2320 2790 2372 2796
rect 2042 2544 2098 2553
rect 2042 2479 2098 2488
rect 2056 2446 2084 2479
rect 2044 2440 2096 2446
rect 2044 2382 2096 2388
rect 1950 1320 2006 1329
rect 1950 1255 2006 1264
rect 1214 54 1532 82
rect 2042 82 2098 480
rect 2332 82 2360 2790
rect 2042 54 2360 82
rect 2608 82 2636 7142
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2976 6322 3004 6598
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 3056 6180 3108 6186
rect 3056 6122 3108 6128
rect 3240 6180 3292 6186
rect 3240 6122 3292 6128
rect 3068 5914 3096 6122
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 3252 5778 3280 6122
rect 2872 5772 2924 5778
rect 2872 5714 2924 5720
rect 3240 5772 3292 5778
rect 3240 5714 3292 5720
rect 2884 5302 2912 5714
rect 2872 5296 2924 5302
rect 2872 5238 2924 5244
rect 3436 4826 3464 8026
rect 4080 7546 4108 9318
rect 4264 8090 4292 10202
rect 4344 8968 4396 8974
rect 4344 8910 4396 8916
rect 4356 8634 4384 8910
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 3884 7472 3936 7478
rect 3884 7414 3936 7420
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3528 5370 3556 5850
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 3424 4820 3476 4826
rect 3252 4780 3424 4808
rect 2688 4684 2740 4690
rect 2688 4626 2740 4632
rect 2700 3738 2728 4626
rect 3252 4078 3280 4780
rect 3424 4762 3476 4768
rect 3516 4480 3568 4486
rect 3516 4422 3568 4428
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 3240 4072 3292 4078
rect 3240 4014 3292 4020
rect 2688 3732 2740 3738
rect 2688 3674 2740 3680
rect 2964 3596 3016 3602
rect 2964 3538 3016 3544
rect 2976 2922 3004 3538
rect 3252 3194 3280 4014
rect 3436 3738 3464 4082
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3436 3602 3464 3674
rect 3424 3596 3476 3602
rect 3424 3538 3476 3544
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 2964 2916 3016 2922
rect 2964 2858 3016 2864
rect 3528 2650 3556 4422
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 2870 82 2926 480
rect 2608 54 2926 82
rect 386 0 442 54
rect 1214 0 1270 54
rect 2042 0 2098 54
rect 2870 0 2926 54
rect 3698 82 3754 480
rect 3896 82 3924 7414
rect 4448 6934 4476 10202
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4068 6928 4120 6934
rect 4068 6870 4120 6876
rect 4436 6928 4488 6934
rect 4436 6870 4488 6876
rect 4080 6118 4108 6870
rect 4632 6458 4660 7142
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 4632 6118 4660 6394
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 3988 4146 4016 5510
rect 4080 5098 4108 6054
rect 4160 5908 4212 5914
rect 4160 5850 4212 5856
rect 4172 5234 4200 5850
rect 4252 5840 4304 5846
rect 4252 5782 4304 5788
rect 4264 5370 4292 5782
rect 4436 5772 4488 5778
rect 4436 5714 4488 5720
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 4068 5092 4120 5098
rect 4068 5034 4120 5040
rect 4448 5030 4476 5714
rect 4436 5024 4488 5030
rect 4436 4966 4488 4972
rect 4448 4758 4476 4966
rect 4436 4752 4488 4758
rect 4436 4694 4488 4700
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4264 4146 4292 4558
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 3988 4049 4016 4082
rect 3974 4040 4030 4049
rect 3974 3975 4030 3984
rect 4356 3942 4384 4626
rect 4724 4486 4752 10474
rect 5460 10470 5488 10746
rect 6656 10470 6684 11222
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 6644 10464 6696 10470
rect 6644 10406 6696 10412
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 4816 9110 4844 10066
rect 4956 9820 5252 9840
rect 5012 9818 5036 9820
rect 5092 9818 5116 9820
rect 5172 9818 5196 9820
rect 5034 9766 5036 9818
rect 5098 9766 5110 9818
rect 5172 9766 5174 9818
rect 5012 9764 5036 9766
rect 5092 9764 5116 9766
rect 5172 9764 5196 9766
rect 4956 9744 5252 9764
rect 5460 9654 5488 10406
rect 6656 10266 6684 10406
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 6092 10124 6144 10130
rect 6092 10066 6144 10072
rect 5448 9648 5500 9654
rect 5448 9590 5500 9596
rect 5264 9512 5316 9518
rect 5264 9454 5316 9460
rect 5276 9178 5304 9454
rect 5552 9382 5580 10066
rect 6104 9722 6132 10066
rect 6092 9716 6144 9722
rect 6092 9658 6144 9664
rect 5814 9616 5870 9625
rect 5814 9551 5870 9560
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5264 9172 5316 9178
rect 5264 9114 5316 9120
rect 4804 9104 4856 9110
rect 4804 9046 4856 9052
rect 4816 8566 4844 9046
rect 4956 8732 5252 8752
rect 5012 8730 5036 8732
rect 5092 8730 5116 8732
rect 5172 8730 5196 8732
rect 5034 8678 5036 8730
rect 5098 8678 5110 8730
rect 5172 8678 5174 8730
rect 5012 8676 5036 8678
rect 5092 8676 5116 8678
rect 5172 8676 5196 8678
rect 4956 8656 5252 8676
rect 4804 8560 4856 8566
rect 4804 8502 4856 8508
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5356 8356 5408 8362
rect 5356 8298 5408 8304
rect 5368 7750 5396 8298
rect 5540 8288 5592 8294
rect 5540 8230 5592 8236
rect 5552 8022 5580 8230
rect 5540 8016 5592 8022
rect 5540 7958 5592 7964
rect 5448 7812 5500 7818
rect 5448 7754 5500 7760
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 4956 7644 5252 7664
rect 5012 7642 5036 7644
rect 5092 7642 5116 7644
rect 5172 7642 5196 7644
rect 5034 7590 5036 7642
rect 5098 7590 5110 7642
rect 5172 7590 5174 7642
rect 5012 7588 5036 7590
rect 5092 7588 5116 7590
rect 5172 7588 5196 7590
rect 4956 7568 5252 7588
rect 5368 7546 5396 7686
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5460 7342 5488 7754
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 5000 7002 5028 7142
rect 4988 6996 5040 7002
rect 4988 6938 5040 6944
rect 5460 6730 5488 7278
rect 5552 7002 5580 7958
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5448 6724 5500 6730
rect 5448 6666 5500 6672
rect 4956 6556 5252 6576
rect 5012 6554 5036 6556
rect 5092 6554 5116 6556
rect 5172 6554 5196 6556
rect 5034 6502 5036 6554
rect 5098 6502 5110 6554
rect 5172 6502 5174 6554
rect 5012 6500 5036 6502
rect 5092 6500 5116 6502
rect 5172 6500 5196 6502
rect 4956 6480 5252 6500
rect 4804 6180 4856 6186
rect 4804 6122 4856 6128
rect 4816 5914 4844 6122
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 5448 5636 5500 5642
rect 5448 5578 5500 5584
rect 4956 5468 5252 5488
rect 5012 5466 5036 5468
rect 5092 5466 5116 5468
rect 5172 5466 5196 5468
rect 5034 5414 5036 5466
rect 5098 5414 5110 5466
rect 5172 5414 5174 5466
rect 5012 5412 5036 5414
rect 5092 5412 5116 5414
rect 5172 5412 5196 5414
rect 4956 5392 5252 5412
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 4816 4486 4844 4762
rect 4712 4480 4764 4486
rect 4712 4422 4764 4428
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4816 4078 4844 4422
rect 4956 4380 5252 4400
rect 5012 4378 5036 4380
rect 5092 4378 5116 4380
rect 5172 4378 5196 4380
rect 5034 4326 5036 4378
rect 5098 4326 5110 4378
rect 5172 4326 5174 4378
rect 5012 4324 5036 4326
rect 5092 4324 5116 4326
rect 5172 4324 5196 4326
rect 4956 4304 5252 4324
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 4896 4072 4948 4078
rect 4896 4014 4948 4020
rect 5264 4072 5316 4078
rect 5264 4014 5316 4020
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 4356 2854 4384 3878
rect 4712 3392 4764 3398
rect 4712 3334 4764 3340
rect 4724 3126 4752 3334
rect 4712 3120 4764 3126
rect 4712 3062 4764 3068
rect 4344 2848 4396 2854
rect 4344 2790 4396 2796
rect 4434 2544 4490 2553
rect 4434 2479 4490 2488
rect 3698 54 3924 82
rect 4448 82 4476 2479
rect 4724 2378 4752 3062
rect 4816 2582 4844 4014
rect 4908 3602 4936 4014
rect 5276 3738 5304 4014
rect 5264 3732 5316 3738
rect 5264 3674 5316 3680
rect 4896 3596 4948 3602
rect 4896 3538 4948 3544
rect 4956 3292 5252 3312
rect 5012 3290 5036 3292
rect 5092 3290 5116 3292
rect 5172 3290 5196 3292
rect 5034 3238 5036 3290
rect 5098 3238 5110 3290
rect 5172 3238 5174 3290
rect 5012 3236 5036 3238
rect 5092 3236 5116 3238
rect 5172 3236 5196 3238
rect 4956 3216 5252 3236
rect 4896 2984 4948 2990
rect 4896 2926 4948 2932
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 4908 2854 4936 2926
rect 4896 2848 4948 2854
rect 4894 2816 4896 2825
rect 4948 2816 4950 2825
rect 4894 2751 4950 2760
rect 4908 2650 4936 2751
rect 4896 2644 4948 2650
rect 4896 2586 4948 2592
rect 4804 2576 4856 2582
rect 4804 2518 4856 2524
rect 4908 2514 4936 2586
rect 5184 2514 5212 2926
rect 4896 2508 4948 2514
rect 4896 2450 4948 2456
rect 5172 2508 5224 2514
rect 5172 2450 5224 2456
rect 4712 2372 4764 2378
rect 4712 2314 4764 2320
rect 4956 2204 5252 2224
rect 5012 2202 5036 2204
rect 5092 2202 5116 2204
rect 5172 2202 5196 2204
rect 5034 2150 5036 2202
rect 5098 2150 5110 2202
rect 5172 2150 5174 2202
rect 5012 2148 5036 2150
rect 5092 2148 5116 2150
rect 5172 2148 5196 2150
rect 4956 2128 5252 2148
rect 4526 82 4582 480
rect 4448 54 4582 82
rect 3698 0 3754 54
rect 4526 0 4582 54
rect 5354 82 5410 480
rect 5460 82 5488 5578
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 5552 4321 5580 5102
rect 5538 4312 5594 4321
rect 5538 4247 5594 4256
rect 5644 3126 5672 8434
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5736 6458 5764 6734
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 5828 5681 5856 9551
rect 6104 9518 6132 9658
rect 6092 9512 6144 9518
rect 6092 9454 6144 9460
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 5908 9104 5960 9110
rect 5908 9046 5960 9052
rect 5920 7886 5948 9046
rect 6012 9042 6040 9318
rect 6000 9036 6052 9042
rect 6000 8978 6052 8984
rect 6368 9036 6420 9042
rect 6368 8978 6420 8984
rect 6380 8498 6408 8978
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 6472 8634 6500 8910
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 6748 8566 6776 13786
rect 6840 13734 6868 14350
rect 7392 14346 7420 15030
rect 7380 14340 7432 14346
rect 7380 14282 7432 14288
rect 7392 13938 7420 14282
rect 7380 13932 7432 13938
rect 7380 13874 7432 13880
rect 7288 13796 7340 13802
rect 7288 13738 7340 13744
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 7300 13530 7328 13738
rect 7392 13530 7420 13874
rect 7484 13814 7512 18788
rect 7564 18770 7616 18776
rect 7656 18148 7708 18154
rect 7656 18090 7708 18096
rect 7564 16584 7616 16590
rect 7564 16526 7616 16532
rect 7576 15978 7604 16526
rect 7564 15972 7616 15978
rect 7564 15914 7616 15920
rect 7576 15706 7604 15914
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7668 14278 7696 18090
rect 7656 14272 7708 14278
rect 7656 14214 7708 14220
rect 7668 13938 7696 14214
rect 7656 13932 7708 13938
rect 7656 13874 7708 13880
rect 7852 13814 7880 20198
rect 8680 20058 8708 20402
rect 8760 20324 8812 20330
rect 8760 20266 8812 20272
rect 9312 20324 9364 20330
rect 9312 20266 9364 20272
rect 8668 20052 8720 20058
rect 8668 19994 8720 20000
rect 8772 19990 8800 20266
rect 8956 20156 9252 20176
rect 9012 20154 9036 20156
rect 9092 20154 9116 20156
rect 9172 20154 9196 20156
rect 9034 20102 9036 20154
rect 9098 20102 9110 20154
rect 9172 20102 9174 20154
rect 9012 20100 9036 20102
rect 9092 20100 9116 20102
rect 9172 20100 9196 20102
rect 8956 20080 9252 20100
rect 8760 19984 8812 19990
rect 8760 19926 8812 19932
rect 8484 19916 8536 19922
rect 8484 19858 8536 19864
rect 8496 19514 8524 19858
rect 8852 19712 8904 19718
rect 8852 19654 8904 19660
rect 8484 19508 8536 19514
rect 8484 19450 8536 19456
rect 8864 19378 8892 19654
rect 8852 19372 8904 19378
rect 8852 19314 8904 19320
rect 8852 19236 8904 19242
rect 8852 19178 8904 19184
rect 8300 18828 8352 18834
rect 8300 18770 8352 18776
rect 8312 18426 8340 18770
rect 8864 18630 8892 19178
rect 8956 19068 9252 19088
rect 9012 19066 9036 19068
rect 9092 19066 9116 19068
rect 9172 19066 9196 19068
rect 9034 19014 9036 19066
rect 9098 19014 9110 19066
rect 9172 19014 9174 19066
rect 9012 19012 9036 19014
rect 9092 19012 9116 19014
rect 9172 19012 9196 19014
rect 8956 18992 9252 19012
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 8852 18624 8904 18630
rect 8852 18566 8904 18572
rect 8300 18420 8352 18426
rect 8300 18362 8352 18368
rect 8588 18290 8616 18566
rect 8576 18284 8628 18290
rect 8576 18226 8628 18232
rect 8588 17882 8616 18226
rect 8864 18154 8892 18566
rect 9324 18358 9352 20266
rect 11072 20262 11100 20946
rect 11060 20256 11112 20262
rect 11060 20198 11112 20204
rect 9772 19984 9824 19990
rect 9772 19926 9824 19932
rect 9784 19514 9812 19926
rect 9956 19848 10008 19854
rect 9956 19790 10008 19796
rect 10140 19848 10192 19854
rect 10140 19790 10192 19796
rect 10416 19848 10468 19854
rect 10416 19790 10468 19796
rect 9772 19508 9824 19514
rect 9772 19450 9824 19456
rect 9312 18352 9364 18358
rect 9312 18294 9364 18300
rect 8852 18148 8904 18154
rect 8852 18090 8904 18096
rect 8956 17980 9252 18000
rect 9012 17978 9036 17980
rect 9092 17978 9116 17980
rect 9172 17978 9196 17980
rect 9034 17926 9036 17978
rect 9098 17926 9110 17978
rect 9172 17926 9174 17978
rect 9012 17924 9036 17926
rect 9092 17924 9116 17926
rect 9172 17924 9196 17926
rect 8956 17904 9252 17924
rect 8576 17876 8628 17882
rect 8576 17818 8628 17824
rect 8024 17740 8076 17746
rect 8024 17682 8076 17688
rect 8484 17740 8536 17746
rect 8484 17682 8536 17688
rect 8036 17270 8064 17682
rect 8496 17338 8524 17682
rect 8576 17672 8628 17678
rect 8576 17614 8628 17620
rect 8484 17332 8536 17338
rect 8484 17274 8536 17280
rect 8024 17264 8076 17270
rect 8024 17206 8076 17212
rect 8036 16522 8064 17206
rect 8392 16992 8444 16998
rect 8392 16934 8444 16940
rect 8404 16726 8432 16934
rect 8392 16720 8444 16726
rect 8392 16662 8444 16668
rect 8024 16516 8076 16522
rect 8024 16458 8076 16464
rect 8404 16046 8432 16662
rect 8496 16182 8524 17274
rect 8588 17202 8616 17614
rect 9784 17338 9812 19450
rect 9968 18834 9996 19790
rect 10152 19378 10180 19790
rect 10428 19378 10456 19790
rect 10140 19372 10192 19378
rect 10140 19314 10192 19320
rect 10416 19372 10468 19378
rect 10416 19314 10468 19320
rect 10508 19236 10560 19242
rect 10508 19178 10560 19184
rect 10520 18902 10548 19178
rect 10508 18896 10560 18902
rect 10508 18838 10560 18844
rect 9956 18828 10008 18834
rect 9956 18770 10008 18776
rect 9968 18737 9996 18770
rect 9954 18728 10010 18737
rect 9954 18663 10010 18672
rect 10520 18630 10548 18838
rect 10876 18760 10928 18766
rect 10876 18702 10928 18708
rect 10692 18692 10744 18698
rect 10692 18634 10744 18640
rect 10508 18624 10560 18630
rect 10508 18566 10560 18572
rect 9864 18148 9916 18154
rect 9864 18090 9916 18096
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 8576 17196 8628 17202
rect 8576 17138 8628 17144
rect 8588 16794 8616 17138
rect 8956 16892 9252 16912
rect 9012 16890 9036 16892
rect 9092 16890 9116 16892
rect 9172 16890 9196 16892
rect 9034 16838 9036 16890
rect 9098 16838 9110 16890
rect 9172 16838 9174 16890
rect 9012 16836 9036 16838
rect 9092 16836 9116 16838
rect 9172 16836 9196 16838
rect 8956 16816 9252 16836
rect 8576 16788 8628 16794
rect 8576 16730 8628 16736
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 9128 16244 9180 16250
rect 9128 16186 9180 16192
rect 8484 16176 8536 16182
rect 8484 16118 8536 16124
rect 8760 16108 8812 16114
rect 8760 16050 8812 16056
rect 8392 16040 8444 16046
rect 8392 15982 8444 15988
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 7932 15360 7984 15366
rect 7932 15302 7984 15308
rect 7944 15026 7972 15302
rect 7932 15020 7984 15026
rect 7932 14962 7984 14968
rect 7944 14618 7972 14962
rect 8312 14890 8340 15506
rect 8300 14884 8352 14890
rect 8300 14826 8352 14832
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 8116 14408 8168 14414
rect 8116 14350 8168 14356
rect 8128 14074 8156 14350
rect 8116 14068 8168 14074
rect 8404 14056 8432 15982
rect 8772 15366 8800 16050
rect 9140 15978 9168 16186
rect 9324 16114 9352 16390
rect 9784 16250 9812 17274
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9404 16176 9456 16182
rect 9404 16118 9456 16124
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 9128 15972 9180 15978
rect 9128 15914 9180 15920
rect 8956 15804 9252 15824
rect 9012 15802 9036 15804
rect 9092 15802 9116 15804
rect 9172 15802 9196 15804
rect 9034 15750 9036 15802
rect 9098 15750 9110 15802
rect 9172 15750 9174 15802
rect 9012 15748 9036 15750
rect 9092 15748 9116 15750
rect 9172 15748 9196 15750
rect 8956 15728 9252 15748
rect 8760 15360 8812 15366
rect 8760 15302 8812 15308
rect 8772 15026 8800 15302
rect 8760 15020 8812 15026
rect 8760 14962 8812 14968
rect 8852 14884 8904 14890
rect 8852 14826 8904 14832
rect 8760 14816 8812 14822
rect 8760 14758 8812 14764
rect 8484 14068 8536 14074
rect 8404 14028 8484 14056
rect 8116 14010 8168 14016
rect 8484 14010 8536 14016
rect 7484 13786 7604 13814
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 6828 12708 6880 12714
rect 6828 12650 6880 12656
rect 6840 11898 6868 12650
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7208 11898 7236 12038
rect 6828 11892 6880 11898
rect 6828 11834 6880 11840
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 6840 11558 6868 11834
rect 7208 11762 7236 11834
rect 7196 11756 7248 11762
rect 7196 11698 7248 11704
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 7392 11150 7420 11698
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7576 10538 7604 13786
rect 7760 13786 7880 13814
rect 7760 12442 7788 13786
rect 8128 13530 8156 14010
rect 8772 13938 8800 14758
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 8772 13530 8800 13874
rect 8116 13524 8168 13530
rect 8116 13466 8168 13472
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 8208 13388 8260 13394
rect 8208 13330 8260 13336
rect 8220 12782 8248 13330
rect 8864 12918 8892 14826
rect 8956 14716 9252 14736
rect 9012 14714 9036 14716
rect 9092 14714 9116 14716
rect 9172 14714 9196 14716
rect 9034 14662 9036 14714
rect 9098 14662 9110 14714
rect 9172 14662 9174 14714
rect 9012 14660 9036 14662
rect 9092 14660 9116 14662
rect 9172 14660 9196 14662
rect 8956 14640 9252 14660
rect 9324 14618 9352 16050
rect 9416 14958 9444 16118
rect 9404 14952 9456 14958
rect 9404 14894 9456 14900
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 9416 14550 9444 14894
rect 9876 14550 9904 18090
rect 10520 18086 10548 18566
rect 10704 18222 10732 18634
rect 10888 18358 10916 18702
rect 10876 18352 10928 18358
rect 10876 18294 10928 18300
rect 10692 18216 10744 18222
rect 10888 18193 10916 18294
rect 10968 18284 11020 18290
rect 10968 18226 11020 18232
rect 10692 18158 10744 18164
rect 10874 18184 10930 18193
rect 10508 18080 10560 18086
rect 10704 18068 10732 18158
rect 10980 18154 11008 18226
rect 10874 18119 10930 18128
rect 10968 18148 11020 18154
rect 10968 18090 11020 18096
rect 10784 18080 10836 18086
rect 10704 18040 10784 18068
rect 10508 18022 10560 18028
rect 10784 18022 10836 18028
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 10416 16652 10468 16658
rect 10416 16594 10468 16600
rect 10336 16250 10364 16594
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 9956 15972 10008 15978
rect 9956 15914 10008 15920
rect 9404 14544 9456 14550
rect 9324 14492 9404 14498
rect 9324 14486 9456 14492
rect 9864 14544 9916 14550
rect 9864 14486 9916 14492
rect 9324 14470 9444 14486
rect 8956 13628 9252 13648
rect 9012 13626 9036 13628
rect 9092 13626 9116 13628
rect 9172 13626 9196 13628
rect 9034 13574 9036 13626
rect 9098 13574 9110 13626
rect 9172 13574 9174 13626
rect 9012 13572 9036 13574
rect 9092 13572 9116 13574
rect 9172 13572 9196 13574
rect 8956 13552 9252 13572
rect 8852 12912 8904 12918
rect 8852 12854 8904 12860
rect 9126 12880 9182 12889
rect 9126 12815 9182 12824
rect 9140 12782 9168 12815
rect 8208 12776 8260 12782
rect 8208 12718 8260 12724
rect 9128 12776 9180 12782
rect 9128 12718 9180 12724
rect 9324 12714 9352 14470
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 9404 14000 9456 14006
rect 9404 13942 9456 13948
rect 9416 13705 9444 13942
rect 9402 13696 9458 13705
rect 9402 13631 9458 13640
rect 9312 12708 9364 12714
rect 9312 12650 9364 12656
rect 8956 12540 9252 12560
rect 9012 12538 9036 12540
rect 9092 12538 9116 12540
rect 9172 12538 9196 12540
rect 9034 12486 9036 12538
rect 9098 12486 9110 12538
rect 9172 12486 9174 12538
rect 9012 12484 9036 12486
rect 9092 12484 9116 12486
rect 9172 12484 9196 12486
rect 8956 12464 9252 12484
rect 7748 12436 7800 12442
rect 7748 12378 7800 12384
rect 8668 12436 8720 12442
rect 8668 12378 8720 12384
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 7760 10810 7788 12174
rect 8036 11558 8064 12242
rect 8392 11824 8444 11830
rect 8392 11766 8444 11772
rect 8024 11552 8076 11558
rect 8024 11494 8076 11500
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 7760 10538 7788 10746
rect 7944 10674 7972 11086
rect 7932 10668 7984 10674
rect 7932 10610 7984 10616
rect 7564 10532 7616 10538
rect 7564 10474 7616 10480
rect 7748 10532 7800 10538
rect 7748 10474 7800 10480
rect 7104 10192 7156 10198
rect 7104 10134 7156 10140
rect 7116 9722 7144 10134
rect 7380 10056 7432 10062
rect 7380 9998 7432 10004
rect 7392 9722 7420 9998
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 7380 9716 7432 9722
rect 7380 9658 7432 9664
rect 7116 9110 7144 9658
rect 8036 9382 8064 11494
rect 8404 10674 8432 11766
rect 8680 11762 8708 12378
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 9416 11642 9444 13631
rect 9784 13172 9812 14350
rect 9876 14074 9904 14486
rect 9968 14414 9996 15914
rect 10336 15638 10364 16186
rect 10428 16182 10456 16594
rect 10416 16176 10468 16182
rect 10416 16118 10468 16124
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 10324 15632 10376 15638
rect 10324 15574 10376 15580
rect 10428 14822 10456 15642
rect 10520 15366 10548 18022
rect 10968 17876 11020 17882
rect 10968 17818 11020 17824
rect 10692 17672 10744 17678
rect 10692 17614 10744 17620
rect 10600 17536 10652 17542
rect 10600 17478 10652 17484
rect 10612 17134 10640 17478
rect 10704 17202 10732 17614
rect 10692 17196 10744 17202
rect 10692 17138 10744 17144
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 10612 15910 10640 17070
rect 10704 16726 10732 17138
rect 10980 16998 11008 17818
rect 10968 16992 11020 16998
rect 10968 16934 11020 16940
rect 10692 16720 10744 16726
rect 10692 16662 10744 16668
rect 11072 16522 11100 20198
rect 12728 19922 12756 23582
rect 14002 23582 14136 23610
rect 14002 23520 14058 23582
rect 12956 21788 13252 21808
rect 13012 21786 13036 21788
rect 13092 21786 13116 21788
rect 13172 21786 13196 21788
rect 13034 21734 13036 21786
rect 13098 21734 13110 21786
rect 13172 21734 13174 21786
rect 13012 21732 13036 21734
rect 13092 21732 13116 21734
rect 13172 21732 13196 21734
rect 12956 21712 13252 21732
rect 13728 20800 13780 20806
rect 13728 20742 13780 20748
rect 12956 20700 13252 20720
rect 13012 20698 13036 20700
rect 13092 20698 13116 20700
rect 13172 20698 13196 20700
rect 13034 20646 13036 20698
rect 13098 20646 13110 20698
rect 13172 20646 13174 20698
rect 13012 20644 13036 20646
rect 13092 20644 13116 20646
rect 13172 20644 13196 20646
rect 12956 20624 13252 20644
rect 13544 20052 13596 20058
rect 13544 19994 13596 20000
rect 12716 19916 12768 19922
rect 12716 19858 12768 19864
rect 12072 19372 12124 19378
rect 12072 19314 12124 19320
rect 12084 18290 12112 19314
rect 12728 19310 12756 19858
rect 13360 19712 13412 19718
rect 13360 19654 13412 19660
rect 12956 19612 13252 19632
rect 13012 19610 13036 19612
rect 13092 19610 13116 19612
rect 13172 19610 13196 19612
rect 13034 19558 13036 19610
rect 13098 19558 13110 19610
rect 13172 19558 13174 19610
rect 13012 19556 13036 19558
rect 13092 19556 13116 19558
rect 13172 19556 13196 19558
rect 12956 19536 13252 19556
rect 12716 19304 12768 19310
rect 12716 19246 12768 19252
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 12820 18902 12848 19110
rect 12808 18896 12860 18902
rect 12808 18838 12860 18844
rect 12072 18284 12124 18290
rect 12072 18226 12124 18232
rect 12532 18284 12584 18290
rect 12532 18226 12584 18232
rect 11152 18148 11204 18154
rect 11152 18090 11204 18096
rect 11244 18148 11296 18154
rect 11244 18090 11296 18096
rect 11164 17882 11192 18090
rect 11152 17876 11204 17882
rect 11152 17818 11204 17824
rect 10876 16516 10928 16522
rect 10876 16458 10928 16464
rect 11060 16516 11112 16522
rect 11060 16458 11112 16464
rect 10784 16040 10836 16046
rect 10784 15982 10836 15988
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 10796 15502 10824 15982
rect 10784 15496 10836 15502
rect 10784 15438 10836 15444
rect 10692 15428 10744 15434
rect 10692 15370 10744 15376
rect 10508 15360 10560 15366
rect 10508 15302 10560 15308
rect 10520 14890 10548 15302
rect 10508 14884 10560 14890
rect 10508 14826 10560 14832
rect 10600 14884 10652 14890
rect 10600 14826 10652 14832
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 10428 13734 10456 14758
rect 10612 14414 10640 14826
rect 10704 14482 10732 15370
rect 10796 14550 10824 15438
rect 10784 14544 10836 14550
rect 10784 14486 10836 14492
rect 10692 14476 10744 14482
rect 10692 14418 10744 14424
rect 10600 14408 10652 14414
rect 10600 14350 10652 14356
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 10612 13326 10640 14350
rect 10796 13938 10824 14486
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 10888 13814 10916 16458
rect 10796 13786 10916 13814
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 10692 13456 10744 13462
rect 10692 13398 10744 13404
rect 10600 13320 10652 13326
rect 10600 13262 10652 13268
rect 9864 13184 9916 13190
rect 9784 13144 9864 13172
rect 9864 13126 9916 13132
rect 9876 12986 9904 13126
rect 10612 12986 10640 13262
rect 9864 12980 9916 12986
rect 9864 12922 9916 12928
rect 10600 12980 10652 12986
rect 10600 12922 10652 12928
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 10324 12776 10376 12782
rect 10324 12718 10376 12724
rect 9600 12442 9628 12718
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9864 12640 9916 12646
rect 9864 12582 9916 12588
rect 9588 12436 9640 12442
rect 9588 12378 9640 12384
rect 9416 11614 9536 11642
rect 9600 11626 9628 12378
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9508 11506 9536 11614
rect 9588 11620 9640 11626
rect 9588 11562 9640 11568
rect 8956 11452 9252 11472
rect 9012 11450 9036 11452
rect 9092 11450 9116 11452
rect 9172 11450 9196 11452
rect 9034 11398 9036 11450
rect 9098 11398 9110 11450
rect 9172 11398 9174 11450
rect 9012 11396 9036 11398
rect 9092 11396 9116 11398
rect 9172 11396 9196 11398
rect 8956 11376 9252 11396
rect 8392 10668 8444 10674
rect 8392 10610 8444 10616
rect 8956 10364 9252 10384
rect 9012 10362 9036 10364
rect 9092 10362 9116 10364
rect 9172 10362 9196 10364
rect 9034 10310 9036 10362
rect 9098 10310 9110 10362
rect 9172 10310 9174 10362
rect 9012 10308 9036 10310
rect 9092 10308 9116 10310
rect 9172 10308 9196 10310
rect 8956 10288 9252 10308
rect 8116 9920 8168 9926
rect 8116 9862 8168 9868
rect 8128 9625 8156 9862
rect 8114 9616 8170 9625
rect 8114 9551 8170 9560
rect 8128 9450 8156 9551
rect 8116 9444 8168 9450
rect 8116 9386 8168 9392
rect 8392 9444 8444 9450
rect 8392 9386 8444 9392
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 8404 9178 8432 9386
rect 8956 9276 9252 9296
rect 9012 9274 9036 9276
rect 9092 9274 9116 9276
rect 9172 9274 9196 9276
rect 9034 9222 9036 9274
rect 9098 9222 9110 9274
rect 9172 9222 9174 9274
rect 9012 9220 9036 9222
rect 9092 9220 9116 9222
rect 9172 9220 9196 9222
rect 8956 9200 9252 9220
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 7104 9104 7156 9110
rect 7104 9046 7156 9052
rect 9312 9104 9364 9110
rect 9312 9046 9364 9052
rect 6736 8560 6788 8566
rect 6736 8502 6788 8508
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5920 7478 5948 7822
rect 6184 7744 6236 7750
rect 6184 7686 6236 7692
rect 5908 7472 5960 7478
rect 5908 7414 5960 7420
rect 6092 6792 6144 6798
rect 6092 6734 6144 6740
rect 6104 6118 6132 6734
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 6104 5914 6132 6054
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 6196 5778 6224 7686
rect 6748 7546 6776 8502
rect 7116 8498 7144 9046
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6748 7342 6776 7482
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 7116 6934 7144 8434
rect 7288 8424 7340 8430
rect 7288 8366 7340 8372
rect 7300 8090 7328 8366
rect 7484 8090 7512 8910
rect 9324 8430 9352 9046
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 8220 8294 8248 8366
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8852 8356 8904 8362
rect 8852 8298 8904 8304
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 8220 7750 8248 8230
rect 8496 7954 8524 8298
rect 8864 7954 8892 8298
rect 8956 8188 9252 8208
rect 9012 8186 9036 8188
rect 9092 8186 9116 8188
rect 9172 8186 9196 8188
rect 9034 8134 9036 8186
rect 9098 8134 9110 8186
rect 9172 8134 9174 8186
rect 9012 8132 9036 8134
rect 9092 8132 9116 8134
rect 9172 8132 9196 8134
rect 8956 8112 9252 8132
rect 8484 7948 8536 7954
rect 8484 7890 8536 7896
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7104 6928 7156 6934
rect 7104 6870 7156 6876
rect 7116 6458 7144 6870
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7392 6458 7420 6598
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 6736 6180 6788 6186
rect 6736 6122 6788 6128
rect 6184 5772 6236 5778
rect 6184 5714 6236 5720
rect 5814 5672 5870 5681
rect 5814 5607 5870 5616
rect 6196 5370 6224 5714
rect 6748 5710 6776 6122
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 6184 5364 6236 5370
rect 6184 5306 6236 5312
rect 6196 5166 6224 5306
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 6184 5160 6236 5166
rect 6184 5102 6236 5108
rect 5828 4214 5856 5102
rect 6196 4690 6224 5102
rect 6656 5030 6684 5646
rect 7116 5370 7144 6394
rect 7392 6118 7420 6394
rect 7668 6322 7696 7346
rect 7760 7274 7788 7482
rect 8220 7478 8248 7686
rect 8496 7546 8524 7890
rect 8484 7540 8536 7546
rect 8484 7482 8536 7488
rect 8208 7472 8260 7478
rect 8208 7414 8260 7420
rect 7748 7268 7800 7274
rect 7748 7210 7800 7216
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7668 5914 7696 6258
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7288 5568 7340 5574
rect 7288 5510 7340 5516
rect 7472 5568 7524 5574
rect 7472 5510 7524 5516
rect 7104 5364 7156 5370
rect 7104 5306 7156 5312
rect 7116 5166 7144 5306
rect 7300 5234 7328 5510
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 7484 5098 7512 5510
rect 7564 5296 7616 5302
rect 7562 5264 7564 5273
rect 7616 5264 7618 5273
rect 7562 5199 7618 5208
rect 7472 5092 7524 5098
rect 7472 5034 7524 5040
rect 6644 5024 6696 5030
rect 6644 4966 6696 4972
rect 6092 4684 6144 4690
rect 6092 4626 6144 4632
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 5816 4208 5868 4214
rect 5816 4150 5868 4156
rect 6104 3942 6132 4626
rect 6184 4548 6236 4554
rect 6184 4490 6236 4496
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6196 3670 6224 4490
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 6184 3664 6236 3670
rect 6288 3641 6316 3878
rect 6184 3606 6236 3612
rect 6274 3632 6330 3641
rect 5724 3596 5776 3602
rect 6274 3567 6330 3576
rect 5724 3538 5776 3544
rect 5632 3120 5684 3126
rect 5632 3062 5684 3068
rect 5736 2854 5764 3538
rect 6380 3466 6408 4626
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6564 4282 6592 4558
rect 6552 4276 6604 4282
rect 6552 4218 6604 4224
rect 6460 3732 6512 3738
rect 6460 3674 6512 3680
rect 6368 3460 6420 3466
rect 6368 3402 6420 3408
rect 6380 3194 6408 3402
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 5908 2916 5960 2922
rect 5908 2858 5960 2864
rect 5724 2848 5776 2854
rect 5724 2790 5776 2796
rect 5354 54 5488 82
rect 5920 82 5948 2858
rect 6472 2650 6500 3674
rect 6656 3670 6684 4966
rect 7576 4214 7604 5199
rect 7760 5166 7788 7210
rect 8864 6934 8892 7890
rect 9324 7546 9352 8366
rect 9312 7540 9364 7546
rect 9312 7482 9364 7488
rect 9312 7268 9364 7274
rect 9312 7210 9364 7216
rect 8956 7100 9252 7120
rect 9012 7098 9036 7100
rect 9092 7098 9116 7100
rect 9172 7098 9196 7100
rect 9034 7046 9036 7098
rect 9098 7046 9110 7098
rect 9172 7046 9174 7098
rect 9012 7044 9036 7046
rect 9092 7044 9116 7046
rect 9172 7044 9196 7046
rect 8956 7024 9252 7044
rect 8852 6928 8904 6934
rect 8852 6870 8904 6876
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8220 6458 8248 6802
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8404 6322 8432 6802
rect 9324 6662 9352 7210
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9324 6390 9352 6598
rect 9312 6384 9364 6390
rect 9312 6326 9364 6332
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 8392 6180 8444 6186
rect 8392 6122 8444 6128
rect 8760 6180 8812 6186
rect 8760 6122 8812 6128
rect 8208 5840 8260 5846
rect 8208 5782 8260 5788
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 7656 5092 7708 5098
rect 7656 5034 7708 5040
rect 7668 4826 7696 5034
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7668 4214 7696 4762
rect 8128 4486 8156 5646
rect 8220 5370 8248 5782
rect 8404 5710 8432 6122
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 8220 4826 8248 5306
rect 8300 5092 8352 5098
rect 8300 5034 8352 5040
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8116 4480 8168 4486
rect 8116 4422 8168 4428
rect 7564 4208 7616 4214
rect 7564 4150 7616 4156
rect 7656 4208 7708 4214
rect 7656 4150 7708 4156
rect 7576 4078 7604 4150
rect 7564 4072 7616 4078
rect 7564 4014 7616 4020
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 6644 3664 6696 3670
rect 6644 3606 6696 3612
rect 6656 3058 6684 3606
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6748 3058 6776 3538
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 6182 82 6238 480
rect 5920 54 6238 82
rect 5354 0 5410 54
rect 6182 0 6238 54
rect 7010 82 7066 480
rect 7116 82 7144 3878
rect 8312 3738 8340 5034
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 7760 3058 7788 3674
rect 7932 3596 7984 3602
rect 7932 3538 7984 3544
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 7944 3126 7972 3538
rect 8024 3460 8076 3466
rect 8024 3402 8076 3408
rect 7932 3120 7984 3126
rect 7932 3062 7984 3068
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7208 2961 7236 2994
rect 7194 2952 7250 2961
rect 8036 2938 8064 3402
rect 7760 2922 8064 2938
rect 7194 2887 7250 2896
rect 7748 2916 8064 2922
rect 7800 2910 8064 2916
rect 7748 2858 7800 2864
rect 7656 2848 7708 2854
rect 7654 2816 7656 2825
rect 7932 2848 7984 2854
rect 7708 2816 7710 2825
rect 7932 2790 7984 2796
rect 7654 2751 7710 2760
rect 7668 2514 7696 2751
rect 7944 2650 7972 2790
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 7656 2508 7708 2514
rect 7656 2450 7708 2456
rect 7564 2372 7616 2378
rect 7564 2314 7616 2320
rect 7010 54 7144 82
rect 7576 82 7604 2314
rect 7668 649 7696 2450
rect 8036 2310 8064 2910
rect 8220 2514 8248 3538
rect 8404 3058 8432 5646
rect 8576 5160 8628 5166
rect 8576 5102 8628 5108
rect 8588 4826 8616 5102
rect 8576 4820 8628 4826
rect 8576 4762 8628 4768
rect 8588 4010 8616 4762
rect 8772 4554 8800 6122
rect 8956 6012 9252 6032
rect 9012 6010 9036 6012
rect 9092 6010 9116 6012
rect 9172 6010 9196 6012
rect 9034 5958 9036 6010
rect 9098 5958 9110 6010
rect 9172 5958 9174 6010
rect 9012 5956 9036 5958
rect 9092 5956 9116 5958
rect 9172 5956 9196 5958
rect 8956 5936 9252 5956
rect 8852 5024 8904 5030
rect 8852 4966 8904 4972
rect 8864 4554 8892 4966
rect 8956 4924 9252 4944
rect 9012 4922 9036 4924
rect 9092 4922 9116 4924
rect 9172 4922 9196 4924
rect 9034 4870 9036 4922
rect 9098 4870 9110 4922
rect 9172 4870 9174 4922
rect 9012 4868 9036 4870
rect 9092 4868 9116 4870
rect 9172 4868 9196 4870
rect 8956 4848 9252 4868
rect 8760 4548 8812 4554
rect 8760 4490 8812 4496
rect 8852 4548 8904 4554
rect 8852 4490 8904 4496
rect 9128 4548 9180 4554
rect 9128 4490 9180 4496
rect 8944 4480 8996 4486
rect 8944 4422 8996 4428
rect 8956 4146 8984 4422
rect 9140 4214 9168 4490
rect 9220 4480 9272 4486
rect 9220 4422 9272 4428
rect 9128 4208 9180 4214
rect 9128 4150 9180 4156
rect 9232 4154 9260 4422
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 9232 4126 9352 4154
rect 9232 4010 9260 4126
rect 8576 4004 8628 4010
rect 8576 3946 8628 3952
rect 9220 4004 9272 4010
rect 9220 3946 9272 3952
rect 8956 3836 9252 3856
rect 9012 3834 9036 3836
rect 9092 3834 9116 3836
rect 9172 3834 9196 3836
rect 9034 3782 9036 3834
rect 9098 3782 9110 3834
rect 9172 3782 9174 3834
rect 9012 3780 9036 3782
rect 9092 3780 9116 3782
rect 9172 3780 9196 3782
rect 8956 3760 9252 3780
rect 9324 3097 9352 4126
rect 9416 3738 9444 11494
rect 9508 11478 9628 11506
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9508 10266 9536 10610
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9600 10146 9628 11478
rect 9508 10118 9628 10146
rect 9508 6118 9536 10118
rect 9692 9466 9720 12582
rect 9876 12306 9904 12582
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 9876 11898 9904 12242
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 9956 11212 10008 11218
rect 9956 11154 10008 11160
rect 9772 11076 9824 11082
rect 9772 11018 9824 11024
rect 9784 10674 9812 11018
rect 9968 10810 9996 11154
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 9772 10668 9824 10674
rect 9772 10610 9824 10616
rect 9784 9586 9812 10610
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9692 9438 9812 9466
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9692 9042 9720 9318
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9600 8498 9628 8774
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9600 7342 9628 8026
rect 9692 7954 9720 8978
rect 9784 8498 9812 9438
rect 10336 9178 10364 12718
rect 10704 12646 10732 13398
rect 10796 13376 10824 13786
rect 10796 13348 10916 13376
rect 10784 13252 10836 13258
rect 10784 13194 10836 13200
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10704 12442 10732 12582
rect 10416 12436 10468 12442
rect 10416 12378 10468 12384
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10428 11558 10456 12378
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10796 11286 10824 13194
rect 10784 11280 10836 11286
rect 10784 11222 10836 11228
rect 10692 11144 10744 11150
rect 10692 11086 10744 11092
rect 10416 11076 10468 11082
rect 10416 11018 10468 11024
rect 10428 10470 10456 11018
rect 10704 10470 10732 11086
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 10428 9586 10456 10406
rect 10600 9920 10652 9926
rect 10600 9862 10652 9868
rect 10612 9722 10640 9862
rect 10600 9716 10652 9722
rect 10600 9658 10652 9664
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 10428 9382 10456 9522
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 10324 9172 10376 9178
rect 10324 9114 10376 9120
rect 9864 9036 9916 9042
rect 9864 8978 9916 8984
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9876 8090 9904 8978
rect 10428 8838 10456 9318
rect 10612 9042 10640 9658
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10704 8974 10732 10406
rect 10784 9988 10836 9994
rect 10784 9930 10836 9936
rect 10796 9586 10824 9930
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10784 8900 10836 8906
rect 10784 8842 10836 8848
rect 10416 8832 10468 8838
rect 10416 8774 10468 8780
rect 10428 8294 10456 8774
rect 10796 8566 10824 8842
rect 10784 8560 10836 8566
rect 10784 8502 10836 8508
rect 10416 8288 10468 8294
rect 10416 8230 10468 8236
rect 10692 8288 10744 8294
rect 10692 8230 10744 8236
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 10232 7948 10284 7954
rect 10232 7890 10284 7896
rect 10244 7546 10272 7890
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 9588 7336 9640 7342
rect 9588 7278 9640 7284
rect 9956 7336 10008 7342
rect 9956 7278 10008 7284
rect 9600 7002 9628 7278
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 9968 6458 9996 7278
rect 10152 6866 10180 7482
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9968 5817 9996 6394
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 9954 5808 10010 5817
rect 10060 5778 10088 6258
rect 10152 5914 10180 6802
rect 10428 6730 10456 8230
rect 10704 7800 10732 8230
rect 10796 7954 10824 8502
rect 10784 7948 10836 7954
rect 10784 7890 10836 7896
rect 10784 7812 10836 7818
rect 10704 7772 10784 7800
rect 10784 7754 10836 7760
rect 10796 7206 10824 7754
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 10796 6866 10824 7142
rect 10784 6860 10836 6866
rect 10784 6802 10836 6808
rect 10416 6724 10468 6730
rect 10416 6666 10468 6672
rect 10428 6458 10456 6666
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 10796 6186 10824 6802
rect 10784 6180 10836 6186
rect 10784 6122 10836 6128
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 9954 5743 10010 5752
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 10140 5772 10192 5778
rect 10140 5714 10192 5720
rect 10060 5370 10088 5714
rect 10048 5364 10100 5370
rect 9968 5324 10048 5352
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9680 4276 9732 4282
rect 9680 4218 9732 4224
rect 9692 3777 9720 4218
rect 9784 4214 9812 4626
rect 9968 4321 9996 5324
rect 10048 5306 10100 5312
rect 10152 4690 10180 5714
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10428 5234 10456 5646
rect 10888 5642 10916 13348
rect 10980 11801 11008 13806
rect 11256 13462 11284 18090
rect 12164 18080 12216 18086
rect 12164 18022 12216 18028
rect 11612 17604 11664 17610
rect 11612 17546 11664 17552
rect 11624 16658 11652 17546
rect 12176 17338 12204 18022
rect 12544 17882 12572 18226
rect 12820 17882 12848 18838
rect 13372 18766 13400 19654
rect 13556 19334 13584 19994
rect 13740 19854 13768 20742
rect 14108 20602 14136 23582
rect 15028 23582 15346 23610
rect 15028 21010 15056 23582
rect 15290 23520 15346 23582
rect 16408 23582 16726 23610
rect 15016 21004 15068 21010
rect 15016 20946 15068 20952
rect 15028 20602 15056 20946
rect 16408 20602 16436 23582
rect 16670 23520 16726 23582
rect 17696 23582 18014 23610
rect 16956 21244 17252 21264
rect 17012 21242 17036 21244
rect 17092 21242 17116 21244
rect 17172 21242 17196 21244
rect 17034 21190 17036 21242
rect 17098 21190 17110 21242
rect 17172 21190 17174 21242
rect 17012 21188 17036 21190
rect 17092 21188 17116 21190
rect 17172 21188 17196 21190
rect 16956 21168 17252 21188
rect 14096 20596 14148 20602
rect 14096 20538 14148 20544
rect 15016 20596 15068 20602
rect 15016 20538 15068 20544
rect 16396 20596 16448 20602
rect 16396 20538 16448 20544
rect 14108 20398 14136 20538
rect 14096 20392 14148 20398
rect 14096 20334 14148 20340
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 13728 19848 13780 19854
rect 13728 19790 13780 19796
rect 13832 19334 13860 20198
rect 14108 19446 14136 20334
rect 15384 20256 15436 20262
rect 15384 20198 15436 20204
rect 15396 19854 15424 20198
rect 16956 20156 17252 20176
rect 17012 20154 17036 20156
rect 17092 20154 17116 20156
rect 17172 20154 17196 20156
rect 17034 20102 17036 20154
rect 17098 20102 17110 20154
rect 17172 20102 17174 20154
rect 17012 20100 17036 20102
rect 17092 20100 17116 20102
rect 17172 20100 17196 20102
rect 16956 20080 17252 20100
rect 15476 19984 15528 19990
rect 15476 19926 15528 19932
rect 14280 19848 14332 19854
rect 14280 19790 14332 19796
rect 15384 19848 15436 19854
rect 15384 19790 15436 19796
rect 14096 19440 14148 19446
rect 14096 19382 14148 19388
rect 13556 19306 13676 19334
rect 13740 19310 13860 19334
rect 13648 19174 13676 19306
rect 13728 19306 13860 19310
rect 13728 19304 13780 19306
rect 13728 19246 13780 19252
rect 14096 19236 14148 19242
rect 14096 19178 14148 19184
rect 14188 19236 14240 19242
rect 14188 19178 14240 19184
rect 13452 19168 13504 19174
rect 13452 19110 13504 19116
rect 13636 19168 13688 19174
rect 13636 19110 13688 19116
rect 13464 18902 13492 19110
rect 14108 18970 14136 19178
rect 14096 18964 14148 18970
rect 14096 18906 14148 18912
rect 13452 18896 13504 18902
rect 13452 18838 13504 18844
rect 13728 18896 13780 18902
rect 13728 18838 13780 18844
rect 13360 18760 13412 18766
rect 13360 18702 13412 18708
rect 12956 18524 13252 18544
rect 13012 18522 13036 18524
rect 13092 18522 13116 18524
rect 13172 18522 13196 18524
rect 13034 18470 13036 18522
rect 13098 18470 13110 18522
rect 13172 18470 13174 18522
rect 13012 18468 13036 18470
rect 13092 18468 13116 18470
rect 13172 18468 13196 18470
rect 12956 18448 13252 18468
rect 13464 18086 13492 18838
rect 13452 18080 13504 18086
rect 13452 18022 13504 18028
rect 12532 17876 12584 17882
rect 12532 17818 12584 17824
rect 12808 17876 12860 17882
rect 12808 17818 12860 17824
rect 12716 17740 12768 17746
rect 12716 17682 12768 17688
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 12728 17270 12756 17682
rect 12956 17436 13252 17456
rect 13012 17434 13036 17436
rect 13092 17434 13116 17436
rect 13172 17434 13196 17436
rect 13034 17382 13036 17434
rect 13098 17382 13110 17434
rect 13172 17382 13174 17434
rect 13012 17380 13036 17382
rect 13092 17380 13116 17382
rect 13172 17380 13196 17382
rect 12956 17360 13252 17380
rect 12716 17264 12768 17270
rect 12636 17224 12716 17252
rect 11704 16788 11756 16794
rect 11704 16730 11756 16736
rect 11612 16652 11664 16658
rect 11612 16594 11664 16600
rect 11612 16040 11664 16046
rect 11612 15982 11664 15988
rect 11624 15706 11652 15982
rect 11612 15700 11664 15706
rect 11612 15642 11664 15648
rect 11716 15570 11744 16730
rect 11980 16652 12032 16658
rect 11980 16594 12032 16600
rect 11992 15706 12020 16594
rect 12256 15972 12308 15978
rect 12256 15914 12308 15920
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 11704 15564 11756 15570
rect 11704 15506 11756 15512
rect 11716 15162 11744 15506
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 11992 15026 12020 15642
rect 11428 15020 11480 15026
rect 11428 14962 11480 14968
rect 11980 15020 12032 15026
rect 11980 14962 12032 14968
rect 11244 13456 11296 13462
rect 11244 13398 11296 13404
rect 11256 11898 11284 13398
rect 11440 12986 11468 14962
rect 11796 14476 11848 14482
rect 11796 14418 11848 14424
rect 11808 14074 11836 14418
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11520 13796 11572 13802
rect 11520 13738 11572 13744
rect 11532 13394 11560 13738
rect 12176 13530 12204 14350
rect 12268 14074 12296 15914
rect 12532 15904 12584 15910
rect 12532 15846 12584 15852
rect 12544 15570 12572 15846
rect 12532 15564 12584 15570
rect 12532 15506 12584 15512
rect 12440 15360 12492 15366
rect 12440 15302 12492 15308
rect 12452 14550 12480 15302
rect 12544 14618 12572 15506
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12440 14544 12492 14550
rect 12440 14486 12492 14492
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 12164 13524 12216 13530
rect 12164 13466 12216 13472
rect 11520 13388 11572 13394
rect 11520 13330 11572 13336
rect 11428 12980 11480 12986
rect 11428 12922 11480 12928
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 10966 11792 11022 11801
rect 11022 11750 11100 11778
rect 10966 11727 11022 11736
rect 10968 10124 11020 10130
rect 10968 10066 11020 10072
rect 10980 9382 11008 10066
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 10876 5636 10928 5642
rect 10876 5578 10928 5584
rect 10416 5228 10468 5234
rect 10416 5170 10468 5176
rect 10428 4826 10456 5170
rect 10508 5092 10560 5098
rect 10508 5034 10560 5040
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 10048 4616 10100 4622
rect 10048 4558 10100 4564
rect 9954 4312 10010 4321
rect 9954 4247 10010 4256
rect 9772 4208 9824 4214
rect 9772 4150 9824 4156
rect 9784 4049 9812 4150
rect 9770 4040 9826 4049
rect 9770 3975 9826 3984
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 9678 3768 9734 3777
rect 9404 3732 9456 3738
rect 9678 3703 9734 3712
rect 9404 3674 9456 3680
rect 9310 3088 9366 3097
rect 8392 3052 8444 3058
rect 9310 3023 9366 3032
rect 8392 2994 8444 3000
rect 8208 2508 8260 2514
rect 8208 2450 8260 2456
rect 8404 2446 8432 2994
rect 9416 2990 9444 3674
rect 9404 2984 9456 2990
rect 9404 2926 9456 2932
rect 9404 2848 9456 2854
rect 9404 2790 9456 2796
rect 8956 2748 9252 2768
rect 9012 2746 9036 2748
rect 9092 2746 9116 2748
rect 9172 2746 9196 2748
rect 9034 2694 9036 2746
rect 9098 2694 9110 2746
rect 9172 2694 9174 2746
rect 9012 2692 9036 2694
rect 9092 2692 9116 2694
rect 9172 2692 9196 2694
rect 8956 2672 9252 2692
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 8024 2304 8076 2310
rect 8024 2246 8076 2252
rect 8942 2000 8998 2009
rect 8942 1935 8998 1944
rect 7654 640 7710 649
rect 7654 575 7710 584
rect 7838 82 7894 480
rect 7576 54 7894 82
rect 7010 0 7066 54
rect 7838 0 7894 54
rect 8666 82 8722 480
rect 8956 82 8984 1935
rect 8666 54 8984 82
rect 9416 82 9444 2790
rect 9876 2514 9904 3878
rect 9968 3670 9996 4247
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 10060 3194 10088 4558
rect 10152 4554 10180 4626
rect 10140 4548 10192 4554
rect 10140 4490 10192 4496
rect 10152 4146 10180 4490
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 10140 4004 10192 4010
rect 10140 3946 10192 3952
rect 10152 3738 10180 3946
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 10324 3664 10376 3670
rect 10324 3606 10376 3612
rect 10048 3188 10100 3194
rect 10048 3130 10100 3136
rect 10336 2650 10364 3606
rect 10520 3126 10548 5034
rect 10600 4072 10652 4078
rect 10600 4014 10652 4020
rect 10508 3120 10560 3126
rect 10508 3062 10560 3068
rect 10324 2644 10376 2650
rect 10324 2586 10376 2592
rect 10520 2582 10548 3062
rect 10508 2576 10560 2582
rect 10508 2518 10560 2524
rect 9864 2508 9916 2514
rect 9864 2450 9916 2456
rect 9494 82 9550 480
rect 9416 54 9550 82
rect 8666 0 8722 54
rect 9494 0 9550 54
rect 10322 82 10378 480
rect 10612 82 10640 4014
rect 10980 4010 11008 9318
rect 11072 8022 11100 11750
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11716 11286 11744 11494
rect 11704 11280 11756 11286
rect 11704 11222 11756 11228
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 11256 9042 11284 10746
rect 11624 10470 11652 11086
rect 11716 10810 11744 11222
rect 11808 11014 11836 12718
rect 12268 11898 12296 14010
rect 12452 13530 12480 14486
rect 12636 13870 12664 17224
rect 12716 17206 12768 17212
rect 13268 16652 13320 16658
rect 13268 16594 13320 16600
rect 12956 16348 13252 16368
rect 13012 16346 13036 16348
rect 13092 16346 13116 16348
rect 13172 16346 13196 16348
rect 13034 16294 13036 16346
rect 13098 16294 13110 16346
rect 13172 16294 13174 16346
rect 13012 16292 13036 16294
rect 13092 16292 13116 16294
rect 13172 16292 13196 16294
rect 12956 16272 13252 16292
rect 13280 16114 13308 16594
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 13280 15910 13308 16050
rect 13268 15904 13320 15910
rect 13268 15846 13320 15852
rect 12956 15260 13252 15280
rect 13012 15258 13036 15260
rect 13092 15258 13116 15260
rect 13172 15258 13196 15260
rect 13034 15206 13036 15258
rect 13098 15206 13110 15258
rect 13172 15206 13174 15258
rect 13012 15204 13036 15206
rect 13092 15204 13116 15206
rect 13172 15204 13196 15206
rect 12956 15184 13252 15204
rect 13280 15094 13308 15846
rect 13464 15366 13492 18022
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 13556 17338 13584 17682
rect 13544 17332 13596 17338
rect 13544 17274 13596 17280
rect 13556 17066 13584 17274
rect 13544 17060 13596 17066
rect 13544 17002 13596 17008
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 13636 15156 13688 15162
rect 13636 15098 13688 15104
rect 13268 15088 13320 15094
rect 13268 15030 13320 15036
rect 12716 14816 12768 14822
rect 12716 14758 12768 14764
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12728 14414 12756 14758
rect 12716 14408 12768 14414
rect 12716 14350 12768 14356
rect 12624 13864 12676 13870
rect 12624 13806 12676 13812
rect 12820 13705 12848 14758
rect 12956 14172 13252 14192
rect 13012 14170 13036 14172
rect 13092 14170 13116 14172
rect 13172 14170 13196 14172
rect 13034 14118 13036 14170
rect 13098 14118 13110 14170
rect 13172 14118 13174 14170
rect 13012 14116 13036 14118
rect 13092 14116 13116 14118
rect 13172 14116 13196 14118
rect 12956 14096 13252 14116
rect 12806 13696 12862 13705
rect 12806 13631 12862 13640
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12716 13456 12768 13462
rect 12716 13398 12768 13404
rect 12728 12646 12756 13398
rect 12956 13084 13252 13104
rect 13012 13082 13036 13084
rect 13092 13082 13116 13084
rect 13172 13082 13196 13084
rect 13034 13030 13036 13082
rect 13098 13030 13110 13082
rect 13172 13030 13174 13082
rect 13012 13028 13036 13030
rect 13092 13028 13116 13030
rect 13172 13028 13196 13030
rect 12956 13008 13252 13028
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 12728 12442 12756 12582
rect 12716 12436 12768 12442
rect 12716 12378 12768 12384
rect 12256 11892 12308 11898
rect 12176 11852 12256 11880
rect 11796 11008 11848 11014
rect 11796 10950 11848 10956
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11612 10464 11664 10470
rect 11612 10406 11664 10412
rect 11624 10198 11652 10406
rect 11612 10192 11664 10198
rect 11612 10134 11664 10140
rect 12176 10130 12204 11852
rect 12256 11834 12308 11840
rect 12728 11286 12756 12378
rect 12820 12102 12848 12786
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12820 11762 12848 12038
rect 12956 11996 13252 12016
rect 13012 11994 13036 11996
rect 13092 11994 13116 11996
rect 13172 11994 13196 11996
rect 13034 11942 13036 11994
rect 13098 11942 13110 11994
rect 13172 11942 13174 11994
rect 13012 11940 13036 11942
rect 13092 11940 13116 11942
rect 13172 11940 13196 11942
rect 12956 11920 13252 11940
rect 13280 11778 13308 15030
rect 13452 14952 13504 14958
rect 13452 14894 13504 14900
rect 13464 14278 13492 14894
rect 13648 14890 13676 15098
rect 13636 14884 13688 14890
rect 13636 14826 13688 14832
rect 13544 14408 13596 14414
rect 13544 14350 13596 14356
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13464 13938 13492 14214
rect 13452 13932 13504 13938
rect 13452 13874 13504 13880
rect 13360 12640 13412 12646
rect 13360 12582 13412 12588
rect 13372 12374 13400 12582
rect 13360 12368 13412 12374
rect 13360 12310 13412 12316
rect 13372 11898 13400 12310
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 12808 11756 12860 11762
rect 13280 11750 13492 11778
rect 12808 11698 12860 11704
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 12716 11280 12768 11286
rect 12716 11222 12768 11228
rect 12956 10908 13252 10928
rect 13012 10906 13036 10908
rect 13092 10906 13116 10908
rect 13172 10906 13196 10908
rect 13034 10854 13036 10906
rect 13098 10854 13110 10906
rect 13172 10854 13174 10906
rect 13012 10852 13036 10854
rect 13092 10852 13116 10854
rect 13172 10852 13196 10854
rect 12956 10832 13252 10852
rect 13372 10810 13400 11290
rect 13360 10804 13412 10810
rect 13360 10746 13412 10752
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 11336 10124 11388 10130
rect 11336 10066 11388 10072
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 11348 9722 11376 10066
rect 11336 9716 11388 9722
rect 11336 9658 11388 9664
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 11532 9042 11560 9522
rect 11244 9036 11296 9042
rect 11244 8978 11296 8984
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 11256 8090 11284 8978
rect 11532 8294 11560 8978
rect 11520 8288 11572 8294
rect 11520 8230 11572 8236
rect 11244 8084 11296 8090
rect 11244 8026 11296 8032
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 11152 7948 11204 7954
rect 11152 7890 11204 7896
rect 11796 7948 11848 7954
rect 11796 7890 11848 7896
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11164 7002 11192 7890
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11152 6996 11204 7002
rect 11152 6938 11204 6944
rect 11348 6458 11376 7142
rect 11808 7002 11836 7890
rect 11900 7546 11928 7890
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11796 6996 11848 7002
rect 11796 6938 11848 6944
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 11520 6180 11572 6186
rect 11520 6122 11572 6128
rect 11244 6112 11296 6118
rect 11244 6054 11296 6060
rect 11256 4554 11284 6054
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 11348 4758 11376 4966
rect 11336 4752 11388 4758
rect 11336 4694 11388 4700
rect 11244 4548 11296 4554
rect 11244 4490 11296 4496
rect 10968 4004 11020 4010
rect 10968 3946 11020 3952
rect 11058 3768 11114 3777
rect 11256 3738 11284 4490
rect 11348 4282 11376 4694
rect 11336 4276 11388 4282
rect 11336 4218 11388 4224
rect 11532 4185 11560 6122
rect 11518 4176 11574 4185
rect 11808 4154 11836 6938
rect 11900 6934 11928 7482
rect 11888 6928 11940 6934
rect 11888 6870 11940 6876
rect 11900 5778 11928 6870
rect 12164 6792 12216 6798
rect 12164 6734 12216 6740
rect 12176 6458 12204 6734
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 11900 5370 11928 5714
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 11888 5364 11940 5370
rect 11888 5306 11940 5312
rect 11518 4111 11574 4120
rect 11716 4126 11836 4154
rect 11058 3703 11114 3712
rect 11244 3732 11296 3738
rect 10322 54 10640 82
rect 11072 82 11100 3703
rect 11244 3674 11296 3680
rect 11336 3528 11388 3534
rect 11336 3470 11388 3476
rect 11348 2650 11376 3470
rect 11716 2961 11744 4126
rect 11900 4078 11928 5306
rect 12084 5234 12112 5646
rect 12268 5522 12296 10406
rect 12544 10266 12572 10542
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 12360 9382 12388 10066
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12348 9376 12400 9382
rect 12348 9318 12400 9324
rect 12360 5642 12388 9318
rect 12820 9178 12848 9998
rect 12956 9820 13252 9840
rect 13012 9818 13036 9820
rect 13092 9818 13116 9820
rect 13172 9818 13196 9820
rect 13034 9766 13036 9818
rect 13098 9766 13110 9818
rect 13172 9766 13174 9818
rect 13012 9764 13036 9766
rect 13092 9764 13116 9766
rect 13172 9764 13196 9766
rect 12956 9744 13252 9764
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 13268 9376 13320 9382
rect 13268 9318 13320 9324
rect 13004 9178 13032 9318
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12992 9172 13044 9178
rect 12992 9114 13044 9120
rect 12956 8732 13252 8752
rect 13012 8730 13036 8732
rect 13092 8730 13116 8732
rect 13172 8730 13196 8732
rect 13034 8678 13036 8730
rect 13098 8678 13110 8730
rect 13172 8678 13174 8730
rect 13012 8676 13036 8678
rect 13092 8676 13116 8678
rect 13172 8676 13196 8678
rect 12956 8656 13252 8676
rect 13280 8537 13308 9318
rect 13266 8528 13322 8537
rect 13266 8463 13322 8472
rect 13464 8430 13492 11750
rect 13556 11082 13584 14350
rect 13648 13530 13676 14826
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13636 13388 13688 13394
rect 13636 13330 13688 13336
rect 13648 12986 13676 13330
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13740 12238 13768 18838
rect 14200 18630 14228 19178
rect 14188 18624 14240 18630
rect 14188 18566 14240 18572
rect 13912 17672 13964 17678
rect 13912 17614 13964 17620
rect 13924 17202 13952 17614
rect 13912 17196 13964 17202
rect 13912 17138 13964 17144
rect 13820 17060 13872 17066
rect 13820 17002 13872 17008
rect 13832 16658 13860 17002
rect 13912 16992 13964 16998
rect 13912 16934 13964 16940
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13832 15366 13860 16594
rect 13924 15910 13952 16934
rect 14004 16584 14056 16590
rect 14004 16526 14056 16532
rect 14016 16114 14044 16526
rect 14004 16108 14056 16114
rect 14004 16050 14056 16056
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 14016 15706 14044 16050
rect 14004 15700 14056 15706
rect 14004 15642 14056 15648
rect 13820 15360 13872 15366
rect 13820 15302 13872 15308
rect 13832 15094 13860 15302
rect 13820 15088 13872 15094
rect 13820 15030 13872 15036
rect 14096 14476 14148 14482
rect 14096 14418 14148 14424
rect 14108 13802 14136 14418
rect 14096 13796 14148 13802
rect 14096 13738 14148 13744
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 14016 12986 14044 13126
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 14016 12646 14044 12922
rect 14004 12640 14056 12646
rect 14004 12582 14056 12588
rect 14004 12368 14056 12374
rect 14004 12310 14056 12316
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13740 11898 13768 12174
rect 13728 11892 13780 11898
rect 13728 11834 13780 11840
rect 14016 11286 14044 12310
rect 14004 11280 14056 11286
rect 14004 11222 14056 11228
rect 13544 11076 13596 11082
rect 13544 11018 13596 11024
rect 13556 10742 13584 11018
rect 13544 10736 13596 10742
rect 13544 10678 13596 10684
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13556 9518 13584 9998
rect 13544 9512 13596 9518
rect 13544 9454 13596 9460
rect 13556 8498 13584 9454
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13452 8424 13504 8430
rect 13452 8366 13504 8372
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 12452 7410 12480 7822
rect 12716 7812 12768 7818
rect 12716 7754 12768 7760
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12452 7002 12480 7346
rect 12532 7268 12584 7274
rect 12532 7210 12584 7216
rect 12440 6996 12492 7002
rect 12440 6938 12492 6944
rect 12348 5636 12400 5642
rect 12348 5578 12400 5584
rect 12176 5494 12296 5522
rect 12072 5228 12124 5234
rect 12072 5170 12124 5176
rect 11888 4072 11940 4078
rect 11888 4014 11940 4020
rect 11796 3596 11848 3602
rect 11796 3538 11848 3544
rect 11808 3398 11836 3538
rect 11796 3392 11848 3398
rect 11796 3334 11848 3340
rect 11980 3392 12032 3398
rect 11980 3334 12032 3340
rect 11702 2952 11758 2961
rect 11702 2887 11758 2896
rect 11808 2650 11836 3334
rect 11336 2644 11388 2650
rect 11336 2586 11388 2592
rect 11796 2644 11848 2650
rect 11796 2586 11848 2592
rect 11992 1766 12020 3334
rect 12072 2848 12124 2854
rect 12072 2790 12124 2796
rect 12084 2650 12112 2790
rect 12072 2644 12124 2650
rect 12072 2586 12124 2592
rect 12176 2417 12204 5494
rect 12544 5370 12572 7210
rect 12728 7002 12756 7754
rect 12956 7644 13252 7664
rect 13012 7642 13036 7644
rect 13092 7642 13116 7644
rect 13172 7642 13196 7644
rect 13034 7590 13036 7642
rect 13098 7590 13110 7642
rect 13172 7590 13174 7642
rect 13012 7588 13036 7590
rect 13092 7588 13116 7590
rect 13172 7588 13196 7590
rect 12956 7568 13252 7588
rect 12716 6996 12768 7002
rect 12716 6938 12768 6944
rect 12956 6556 13252 6576
rect 13012 6554 13036 6556
rect 13092 6554 13116 6556
rect 13172 6554 13196 6556
rect 13034 6502 13036 6554
rect 13098 6502 13110 6554
rect 13172 6502 13174 6554
rect 13012 6500 13036 6502
rect 13092 6500 13116 6502
rect 13172 6500 13196 6502
rect 12956 6480 13252 6500
rect 13280 6254 13308 8366
rect 13452 7880 13504 7886
rect 13452 7822 13504 7828
rect 13464 7546 13492 7822
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13360 7200 13412 7206
rect 13360 7142 13412 7148
rect 13372 6934 13400 7142
rect 13728 6996 13780 7002
rect 13728 6938 13780 6944
rect 13360 6928 13412 6934
rect 13360 6870 13412 6876
rect 13372 6458 13400 6870
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13268 6248 13320 6254
rect 13268 6190 13320 6196
rect 13360 5840 13412 5846
rect 13360 5782 13412 5788
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 13268 5704 13320 5710
rect 13268 5646 13320 5652
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 12440 5228 12492 5234
rect 12440 5170 12492 5176
rect 12254 5128 12310 5137
rect 12254 5063 12310 5072
rect 12162 2408 12218 2417
rect 12162 2343 12218 2352
rect 11980 1760 12032 1766
rect 11980 1702 12032 1708
rect 11150 82 11206 480
rect 11072 54 11206 82
rect 10322 0 10378 54
rect 11150 0 11206 54
rect 11978 82 12034 480
rect 12268 82 12296 5063
rect 12452 4826 12480 5170
rect 12820 4826 12848 5646
rect 12956 5468 13252 5488
rect 13012 5466 13036 5468
rect 13092 5466 13116 5468
rect 13172 5466 13196 5468
rect 13034 5414 13036 5466
rect 13098 5414 13110 5466
rect 13172 5414 13174 5466
rect 13012 5412 13036 5414
rect 13092 5412 13116 5414
rect 13172 5412 13196 5414
rect 12956 5392 13252 5412
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 13280 4622 13308 5646
rect 13372 5370 13400 5782
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 13452 4752 13504 4758
rect 13452 4694 13504 4700
rect 13268 4616 13320 4622
rect 13268 4558 13320 4564
rect 12956 4380 13252 4400
rect 13012 4378 13036 4380
rect 13092 4378 13116 4380
rect 13172 4378 13196 4380
rect 13034 4326 13036 4378
rect 13098 4326 13110 4378
rect 13172 4326 13174 4378
rect 13012 4324 13036 4326
rect 13092 4324 13116 4326
rect 13172 4324 13196 4326
rect 12956 4304 13252 4324
rect 12440 4072 12492 4078
rect 12440 4014 12492 4020
rect 12348 3936 12400 3942
rect 12348 3878 12400 3884
rect 12360 2446 12388 3878
rect 12452 3738 12480 4014
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12452 3641 12480 3674
rect 12438 3632 12494 3641
rect 12438 3567 12494 3576
rect 12544 3058 12572 3878
rect 13280 3534 13308 4558
rect 13464 4282 13492 4694
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 13360 3664 13412 3670
rect 13360 3606 13412 3612
rect 13268 3528 13320 3534
rect 13268 3470 13320 3476
rect 12956 3292 13252 3312
rect 13012 3290 13036 3292
rect 13092 3290 13116 3292
rect 13172 3290 13196 3292
rect 13034 3238 13036 3290
rect 13098 3238 13110 3290
rect 13172 3238 13174 3290
rect 13012 3236 13036 3238
rect 13092 3236 13116 3238
rect 13172 3236 13196 3238
rect 12956 3216 13252 3236
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 12348 2440 12400 2446
rect 12348 2382 12400 2388
rect 12438 2408 12494 2417
rect 13280 2378 13308 3470
rect 13372 3194 13400 3606
rect 13648 3466 13676 6734
rect 13740 6254 13768 6938
rect 13832 6798 13860 10678
rect 14016 10674 14044 11222
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 13912 10600 13964 10606
rect 13912 10542 13964 10548
rect 13924 10130 13952 10542
rect 14004 10532 14056 10538
rect 14004 10474 14056 10480
rect 13912 10124 13964 10130
rect 13912 10066 13964 10072
rect 14016 9722 14044 10474
rect 14004 9716 14056 9722
rect 14004 9658 14056 9664
rect 14016 9382 14044 9658
rect 14004 9376 14056 9382
rect 14004 9318 14056 9324
rect 13912 9036 13964 9042
rect 13912 8978 13964 8984
rect 13924 8294 13952 8978
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 13924 7954 13952 8230
rect 14016 8090 14044 9318
rect 14004 8084 14056 8090
rect 14004 8026 14056 8032
rect 13912 7948 13964 7954
rect 13912 7890 13964 7896
rect 14016 7478 14044 8026
rect 14004 7472 14056 7478
rect 14004 7414 14056 7420
rect 13820 6792 13872 6798
rect 13820 6734 13872 6740
rect 13728 6248 13780 6254
rect 13728 6190 13780 6196
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13636 3460 13688 3466
rect 13636 3402 13688 3408
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 13372 2650 13400 3130
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 13728 2576 13780 2582
rect 13728 2518 13780 2524
rect 12438 2343 12494 2352
rect 13268 2372 13320 2378
rect 12452 2310 12480 2343
rect 13268 2314 13320 2320
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 12716 2304 12768 2310
rect 12716 2246 12768 2252
rect 11978 54 12296 82
rect 12728 82 12756 2246
rect 12956 2204 13252 2224
rect 13012 2202 13036 2204
rect 13092 2202 13116 2204
rect 13172 2202 13196 2204
rect 13034 2150 13036 2202
rect 13098 2150 13110 2202
rect 13172 2150 13174 2202
rect 13012 2148 13036 2150
rect 13092 2148 13116 2150
rect 13172 2148 13196 2150
rect 12956 2128 13252 2148
rect 12806 82 12862 480
rect 12728 54 12862 82
rect 11978 0 12034 54
rect 12806 0 12862 54
rect 13634 82 13690 480
rect 13740 82 13768 2518
rect 13832 134 13860 6054
rect 14108 4690 14136 13738
rect 14292 13190 14320 19790
rect 15396 19514 15424 19790
rect 15384 19508 15436 19514
rect 15384 19450 15436 19456
rect 14372 19372 14424 19378
rect 14372 19314 14424 19320
rect 14384 18902 14412 19314
rect 15488 19242 15516 19926
rect 17696 19922 17724 23582
rect 17958 23520 18014 23582
rect 19076 23582 19394 23610
rect 19076 20602 19104 23582
rect 19338 23520 19394 23582
rect 20626 23610 20682 24000
rect 22006 23610 22062 24000
rect 20626 23582 20760 23610
rect 20626 23520 20682 23582
rect 19064 20596 19116 20602
rect 19064 20538 19116 20544
rect 18604 20256 18656 20262
rect 18604 20198 18656 20204
rect 18696 20256 18748 20262
rect 18696 20198 18748 20204
rect 16948 19916 17000 19922
rect 16948 19858 17000 19864
rect 17684 19916 17736 19922
rect 17684 19858 17736 19864
rect 16856 19712 16908 19718
rect 16856 19654 16908 19660
rect 16302 19272 16358 19281
rect 15476 19236 15528 19242
rect 16302 19207 16358 19216
rect 15476 19178 15528 19184
rect 15384 19168 15436 19174
rect 15384 19110 15436 19116
rect 14372 18896 14424 18902
rect 14372 18838 14424 18844
rect 14740 18624 14792 18630
rect 14740 18566 14792 18572
rect 14556 18148 14608 18154
rect 14556 18090 14608 18096
rect 14568 17338 14596 18090
rect 14556 17332 14608 17338
rect 14556 17274 14608 17280
rect 14464 15904 14516 15910
rect 14464 15846 14516 15852
rect 14476 15638 14504 15846
rect 14464 15632 14516 15638
rect 14464 15574 14516 15580
rect 14476 15162 14504 15574
rect 14464 15156 14516 15162
rect 14464 15098 14516 15104
rect 14752 14822 14780 18566
rect 15396 18290 15424 19110
rect 16316 18970 16344 19207
rect 16868 18970 16896 19654
rect 16960 19514 16988 19858
rect 17408 19712 17460 19718
rect 17408 19654 17460 19660
rect 16948 19508 17000 19514
rect 16948 19450 17000 19456
rect 16956 19068 17252 19088
rect 17012 19066 17036 19068
rect 17092 19066 17116 19068
rect 17172 19066 17196 19068
rect 17034 19014 17036 19066
rect 17098 19014 17110 19066
rect 17172 19014 17174 19066
rect 17012 19012 17036 19014
rect 17092 19012 17116 19014
rect 17172 19012 17196 19014
rect 16956 18992 17252 19012
rect 16304 18964 16356 18970
rect 16304 18906 16356 18912
rect 16856 18964 16908 18970
rect 16856 18906 16908 18912
rect 15844 18896 15896 18902
rect 15844 18838 15896 18844
rect 15476 18760 15528 18766
rect 15476 18702 15528 18708
rect 15568 18760 15620 18766
rect 15568 18702 15620 18708
rect 15384 18284 15436 18290
rect 15384 18226 15436 18232
rect 15488 17882 15516 18702
rect 15580 18358 15608 18702
rect 15568 18352 15620 18358
rect 15568 18294 15620 18300
rect 15856 18086 15884 18838
rect 15936 18352 15988 18358
rect 15936 18294 15988 18300
rect 15844 18080 15896 18086
rect 15844 18022 15896 18028
rect 15476 17876 15528 17882
rect 15476 17818 15528 17824
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 15212 16998 15240 17614
rect 15856 16998 15884 18022
rect 15948 17814 15976 18294
rect 16316 18290 16344 18906
rect 16672 18760 16724 18766
rect 16672 18702 16724 18708
rect 16304 18284 16356 18290
rect 16304 18226 16356 18232
rect 15936 17808 15988 17814
rect 15936 17750 15988 17756
rect 15948 17338 15976 17750
rect 15936 17332 15988 17338
rect 15936 17274 15988 17280
rect 16120 17060 16172 17066
rect 16120 17002 16172 17008
rect 15200 16992 15252 16998
rect 15200 16934 15252 16940
rect 15844 16992 15896 16998
rect 15844 16934 15896 16940
rect 15212 16726 15240 16934
rect 15200 16720 15252 16726
rect 15200 16662 15252 16668
rect 15384 16652 15436 16658
rect 15384 16594 15436 16600
rect 15396 16046 15424 16594
rect 15856 16250 15884 16934
rect 16132 16794 16160 17002
rect 16120 16788 16172 16794
rect 16120 16730 16172 16736
rect 16120 16516 16172 16522
rect 16120 16458 16172 16464
rect 16132 16250 16160 16458
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 16120 16244 16172 16250
rect 16172 16204 16252 16232
rect 16120 16186 16172 16192
rect 15384 16040 15436 16046
rect 15384 15982 15436 15988
rect 16120 16040 16172 16046
rect 16120 15982 16172 15988
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 15764 15570 15792 15846
rect 15108 15564 15160 15570
rect 15108 15506 15160 15512
rect 15752 15564 15804 15570
rect 15752 15506 15804 15512
rect 15120 15162 15148 15506
rect 15108 15156 15160 15162
rect 15108 15098 15160 15104
rect 15764 15094 15792 15506
rect 15752 15088 15804 15094
rect 15752 15030 15804 15036
rect 15568 14952 15620 14958
rect 15568 14894 15620 14900
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 14648 14272 14700 14278
rect 14648 14214 14700 14220
rect 14660 13938 14688 14214
rect 14648 13932 14700 13938
rect 14648 13874 14700 13880
rect 14752 13802 14780 14758
rect 15580 14618 15608 14894
rect 15568 14612 15620 14618
rect 15620 14572 15700 14600
rect 15568 14554 15620 14560
rect 15568 14476 15620 14482
rect 15568 14418 15620 14424
rect 14924 14408 14976 14414
rect 14924 14350 14976 14356
rect 14936 13938 14964 14350
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 14740 13796 14792 13802
rect 14740 13738 14792 13744
rect 14752 13530 14780 13738
rect 14740 13524 14792 13530
rect 14740 13466 14792 13472
rect 15200 13388 15252 13394
rect 15200 13330 15252 13336
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 14740 13184 14792 13190
rect 14740 13126 14792 13132
rect 14292 12714 14320 13126
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14280 12708 14332 12714
rect 14280 12650 14332 12656
rect 14292 12170 14320 12650
rect 14464 12640 14516 12646
rect 14464 12582 14516 12588
rect 14280 12164 14332 12170
rect 14280 12106 14332 12112
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 14292 9042 14320 11494
rect 14280 9036 14332 9042
rect 14280 8978 14332 8984
rect 14292 8294 14320 8978
rect 14280 8288 14332 8294
rect 14280 8230 14332 8236
rect 14188 6180 14240 6186
rect 14188 6122 14240 6128
rect 14200 5914 14228 6122
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 14200 5234 14228 5850
rect 14188 5228 14240 5234
rect 14188 5170 14240 5176
rect 14096 4684 14148 4690
rect 14096 4626 14148 4632
rect 14108 4282 14136 4626
rect 14096 4276 14148 4282
rect 14096 4218 14148 4224
rect 14108 3777 14136 4218
rect 14292 3942 14320 8230
rect 14372 7744 14424 7750
rect 14372 7686 14424 7692
rect 14384 7478 14412 7686
rect 14372 7472 14424 7478
rect 14372 7414 14424 7420
rect 14476 6118 14504 12582
rect 14568 12374 14596 12786
rect 14752 12442 14780 13126
rect 15212 12646 15240 13330
rect 15580 13190 15608 14418
rect 15568 13184 15620 13190
rect 15568 13126 15620 13132
rect 15384 12776 15436 12782
rect 15384 12718 15436 12724
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 14740 12436 14792 12442
rect 14740 12378 14792 12384
rect 14556 12368 14608 12374
rect 14556 12310 14608 12316
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 14568 11898 14596 12174
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14752 11626 14780 12378
rect 14740 11620 14792 11626
rect 14740 11562 14792 11568
rect 15396 11558 15424 12718
rect 15476 12368 15528 12374
rect 15476 12310 15528 12316
rect 15488 11626 15516 12310
rect 15672 11898 15700 14572
rect 15764 14550 15792 15030
rect 15752 14544 15804 14550
rect 15752 14486 15804 14492
rect 15936 13728 15988 13734
rect 15936 13670 15988 13676
rect 15752 13252 15804 13258
rect 15752 13194 15804 13200
rect 15764 12782 15792 13194
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15856 12782 15884 13126
rect 15752 12776 15804 12782
rect 15752 12718 15804 12724
rect 15844 12776 15896 12782
rect 15844 12718 15896 12724
rect 15660 11892 15712 11898
rect 15660 11834 15712 11840
rect 15476 11620 15528 11626
rect 15476 11562 15528 11568
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15488 11286 15516 11562
rect 14832 11280 14884 11286
rect 14832 11222 14884 11228
rect 15476 11280 15528 11286
rect 15476 11222 15528 11228
rect 14844 10810 14872 11222
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 14832 10804 14884 10810
rect 14832 10746 14884 10752
rect 14556 9920 14608 9926
rect 14556 9862 14608 9868
rect 14568 7313 14596 9862
rect 14648 9376 14700 9382
rect 14648 9318 14700 9324
rect 14660 8634 14688 9318
rect 14924 9172 14976 9178
rect 14924 9114 14976 9120
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 14660 8362 14688 8570
rect 14830 8528 14886 8537
rect 14936 8498 14964 9114
rect 15016 8968 15068 8974
rect 15016 8910 15068 8916
rect 14830 8463 14886 8472
rect 14924 8492 14976 8498
rect 14648 8356 14700 8362
rect 14648 8298 14700 8304
rect 14740 7472 14792 7478
rect 14740 7414 14792 7420
rect 14554 7304 14610 7313
rect 14752 7274 14780 7414
rect 14554 7239 14610 7248
rect 14740 7268 14792 7274
rect 14740 7210 14792 7216
rect 14556 7200 14608 7206
rect 14556 7142 14608 7148
rect 14568 6662 14596 7142
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14568 6390 14596 6598
rect 14556 6384 14608 6390
rect 14556 6326 14608 6332
rect 14844 6254 14872 8463
rect 14924 8434 14976 8440
rect 15028 8090 15056 8910
rect 15016 8084 15068 8090
rect 15016 8026 15068 8032
rect 14832 6248 14884 6254
rect 14832 6190 14884 6196
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 15108 6112 15160 6118
rect 15108 6054 15160 6060
rect 15120 5710 15148 6054
rect 15108 5704 15160 5710
rect 15108 5646 15160 5652
rect 15120 4826 15148 5646
rect 15108 4820 15160 4826
rect 15108 4762 15160 4768
rect 14556 4480 14608 4486
rect 14556 4422 14608 4428
rect 14568 4010 14596 4422
rect 14556 4004 14608 4010
rect 14556 3946 14608 3952
rect 14648 4004 14700 4010
rect 14648 3946 14700 3952
rect 14280 3936 14332 3942
rect 14280 3878 14332 3884
rect 14094 3768 14150 3777
rect 14094 3703 14150 3712
rect 14568 2582 14596 3946
rect 14660 3738 14688 3946
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 14660 3194 14688 3674
rect 14648 3188 14700 3194
rect 14648 3130 14700 3136
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 14556 2576 14608 2582
rect 14278 2544 14334 2553
rect 14556 2518 14608 2524
rect 14278 2479 14334 2488
rect 14292 2446 14320 2479
rect 15120 2446 15148 3130
rect 14280 2440 14332 2446
rect 14280 2382 14332 2388
rect 15108 2440 15160 2446
rect 15108 2382 15160 2388
rect 13634 54 13768 82
rect 13820 128 13872 134
rect 13820 70 13872 76
rect 14462 128 14518 480
rect 14462 76 14464 128
rect 14516 76 14518 128
rect 13634 0 13690 54
rect 14462 0 14518 76
rect 15212 82 15240 10950
rect 15396 10470 15424 11086
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15672 10266 15700 11834
rect 15752 10464 15804 10470
rect 15752 10406 15804 10412
rect 15660 10260 15712 10266
rect 15660 10202 15712 10208
rect 15764 9994 15792 10406
rect 15844 10124 15896 10130
rect 15844 10066 15896 10072
rect 15752 9988 15804 9994
rect 15752 9930 15804 9936
rect 15856 9926 15884 10066
rect 15844 9920 15896 9926
rect 15844 9862 15896 9868
rect 15856 9654 15884 9862
rect 15844 9648 15896 9654
rect 15844 9590 15896 9596
rect 15568 9512 15620 9518
rect 15568 9454 15620 9460
rect 15580 8362 15608 9454
rect 15660 9172 15712 9178
rect 15660 9114 15712 9120
rect 15672 8498 15700 9114
rect 15660 8492 15712 8498
rect 15660 8434 15712 8440
rect 15568 8356 15620 8362
rect 15568 8298 15620 8304
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 15396 7546 15424 8026
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 15580 7478 15608 8298
rect 15948 7954 15976 13670
rect 16132 10198 16160 15982
rect 16224 15094 16252 16204
rect 16580 16040 16632 16046
rect 16580 15982 16632 15988
rect 16592 15706 16620 15982
rect 16580 15700 16632 15706
rect 16408 15660 16580 15688
rect 16212 15088 16264 15094
rect 16212 15030 16264 15036
rect 16212 11688 16264 11694
rect 16212 11630 16264 11636
rect 16224 10810 16252 11630
rect 16408 11014 16436 15660
rect 16580 15642 16632 15648
rect 16488 14884 16540 14890
rect 16488 14826 16540 14832
rect 16500 14414 16528 14826
rect 16488 14408 16540 14414
rect 16488 14350 16540 14356
rect 16500 13530 16528 14350
rect 16580 14272 16632 14278
rect 16580 14214 16632 14220
rect 16592 13938 16620 14214
rect 16684 13938 16712 18702
rect 16868 18426 16896 18906
rect 17040 18896 17092 18902
rect 17040 18838 17092 18844
rect 16856 18420 16908 18426
rect 16856 18362 16908 18368
rect 17052 18358 17080 18838
rect 17224 18760 17276 18766
rect 17224 18702 17276 18708
rect 17040 18352 17092 18358
rect 17040 18294 17092 18300
rect 17236 18290 17264 18702
rect 17224 18284 17276 18290
rect 17224 18226 17276 18232
rect 17420 18193 17448 19654
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 18156 18970 18184 19110
rect 18144 18964 18196 18970
rect 18144 18906 18196 18912
rect 18156 18290 18184 18906
rect 18236 18352 18288 18358
rect 18236 18294 18288 18300
rect 18144 18284 18196 18290
rect 18144 18226 18196 18232
rect 17406 18184 17462 18193
rect 17406 18119 17462 18128
rect 17592 18080 17644 18086
rect 17592 18022 17644 18028
rect 16956 17980 17252 18000
rect 17012 17978 17036 17980
rect 17092 17978 17116 17980
rect 17172 17978 17196 17980
rect 17034 17926 17036 17978
rect 17098 17926 17110 17978
rect 17172 17926 17174 17978
rect 17012 17924 17036 17926
rect 17092 17924 17116 17926
rect 17172 17924 17196 17926
rect 16956 17904 17252 17924
rect 17604 17814 17632 18022
rect 17592 17808 17644 17814
rect 17592 17750 17644 17756
rect 17316 17672 17368 17678
rect 17316 17614 17368 17620
rect 17328 17338 17356 17614
rect 17316 17332 17368 17338
rect 17316 17274 17368 17280
rect 17604 16998 17632 17750
rect 17868 17604 17920 17610
rect 17868 17546 17920 17552
rect 17880 17066 17908 17546
rect 18248 17202 18276 18294
rect 18328 17536 18380 17542
rect 18328 17478 18380 17484
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 17868 17060 17920 17066
rect 17868 17002 17920 17008
rect 17592 16992 17644 16998
rect 17592 16934 17644 16940
rect 16956 16892 17252 16912
rect 17012 16890 17036 16892
rect 17092 16890 17116 16892
rect 17172 16890 17196 16892
rect 17034 16838 17036 16890
rect 17098 16838 17110 16890
rect 17172 16838 17174 16890
rect 17012 16836 17036 16838
rect 17092 16836 17116 16838
rect 17172 16836 17196 16838
rect 16956 16816 17252 16836
rect 17408 16720 17460 16726
rect 17408 16662 17460 16668
rect 17316 16584 17368 16590
rect 17316 16526 17368 16532
rect 17328 16114 17356 16526
rect 17316 16108 17368 16114
rect 17316 16050 17368 16056
rect 17316 15904 17368 15910
rect 17420 15892 17448 16662
rect 17368 15864 17448 15892
rect 17316 15846 17368 15852
rect 16956 15804 17252 15824
rect 17012 15802 17036 15804
rect 17092 15802 17116 15804
rect 17172 15802 17196 15804
rect 17034 15750 17036 15802
rect 17098 15750 17110 15802
rect 17172 15750 17174 15802
rect 17012 15748 17036 15750
rect 17092 15748 17116 15750
rect 17172 15748 17196 15750
rect 16956 15728 17252 15748
rect 17328 15638 17356 15846
rect 16856 15632 16908 15638
rect 16856 15574 16908 15580
rect 17316 15632 17368 15638
rect 17316 15574 17368 15580
rect 16868 14822 16896 15574
rect 17500 15496 17552 15502
rect 17500 15438 17552 15444
rect 17512 15162 17540 15438
rect 17500 15156 17552 15162
rect 17500 15098 17552 15104
rect 16856 14816 16908 14822
rect 16856 14758 16908 14764
rect 16868 14550 16896 14758
rect 16956 14716 17252 14736
rect 17012 14714 17036 14716
rect 17092 14714 17116 14716
rect 17172 14714 17196 14716
rect 17034 14662 17036 14714
rect 17098 14662 17110 14714
rect 17172 14662 17174 14714
rect 17012 14660 17036 14662
rect 17092 14660 17116 14662
rect 17172 14660 17196 14662
rect 16956 14640 17252 14660
rect 16856 14544 16908 14550
rect 16856 14486 16908 14492
rect 16868 14006 16896 14486
rect 17604 14278 17632 16934
rect 17880 16114 17908 17002
rect 18248 16658 18276 17138
rect 18340 17066 18368 17478
rect 18328 17060 18380 17066
rect 18328 17002 18380 17008
rect 18340 16794 18368 17002
rect 18328 16788 18380 16794
rect 18328 16730 18380 16736
rect 18236 16652 18288 16658
rect 18236 16594 18288 16600
rect 17868 16108 17920 16114
rect 17868 16050 17920 16056
rect 18236 15972 18288 15978
rect 18236 15914 18288 15920
rect 17960 15904 18012 15910
rect 17960 15846 18012 15852
rect 17592 14272 17644 14278
rect 17592 14214 17644 14220
rect 16856 14000 16908 14006
rect 16856 13942 16908 13948
rect 16580 13932 16632 13938
rect 16580 13874 16632 13880
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 16592 13802 16620 13874
rect 16580 13796 16632 13802
rect 16580 13738 16632 13744
rect 16488 13524 16540 13530
rect 16488 13466 16540 13472
rect 16868 13462 16896 13942
rect 17500 13728 17552 13734
rect 17500 13670 17552 13676
rect 16956 13628 17252 13648
rect 17012 13626 17036 13628
rect 17092 13626 17116 13628
rect 17172 13626 17196 13628
rect 17034 13574 17036 13626
rect 17098 13574 17110 13626
rect 17172 13574 17174 13626
rect 17012 13572 17036 13574
rect 17092 13572 17116 13574
rect 17172 13572 17196 13574
rect 16956 13552 17252 13572
rect 16856 13456 16908 13462
rect 16856 13398 16908 13404
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 16684 12850 16712 13262
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16868 12646 16896 13398
rect 17512 12986 17540 13670
rect 17500 12980 17552 12986
rect 17500 12922 17552 12928
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16488 11552 16540 11558
rect 16488 11494 16540 11500
rect 16396 11008 16448 11014
rect 16396 10950 16448 10956
rect 16212 10804 16264 10810
rect 16212 10746 16264 10752
rect 16224 10606 16252 10746
rect 16212 10600 16264 10606
rect 16212 10542 16264 10548
rect 16120 10192 16172 10198
rect 16120 10134 16172 10140
rect 16500 10130 16528 11494
rect 16764 10600 16816 10606
rect 16764 10542 16816 10548
rect 16488 10124 16540 10130
rect 16488 10066 16540 10072
rect 16500 9722 16528 10066
rect 16488 9716 16540 9722
rect 16488 9658 16540 9664
rect 16212 9376 16264 9382
rect 16212 9318 16264 9324
rect 16224 9178 16252 9318
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16776 8430 16804 10542
rect 16868 10538 16896 12582
rect 16956 12540 17252 12560
rect 17012 12538 17036 12540
rect 17092 12538 17116 12540
rect 17172 12538 17196 12540
rect 17034 12486 17036 12538
rect 17098 12486 17110 12538
rect 17172 12486 17174 12538
rect 17012 12484 17036 12486
rect 17092 12484 17116 12486
rect 17172 12484 17196 12486
rect 16956 12464 17252 12484
rect 16956 11452 17252 11472
rect 17012 11450 17036 11452
rect 17092 11450 17116 11452
rect 17172 11450 17196 11452
rect 17034 11398 17036 11450
rect 17098 11398 17110 11450
rect 17172 11398 17174 11450
rect 17012 11396 17036 11398
rect 17092 11396 17116 11398
rect 17172 11396 17196 11398
rect 16956 11376 17252 11396
rect 17316 11008 17368 11014
rect 17316 10950 17368 10956
rect 17328 10606 17356 10950
rect 17972 10742 18000 15846
rect 18248 15706 18276 15914
rect 18236 15700 18288 15706
rect 18236 15642 18288 15648
rect 18328 13864 18380 13870
rect 18328 13806 18380 13812
rect 18340 13308 18368 13806
rect 18512 13320 18564 13326
rect 18340 13280 18512 13308
rect 18512 13262 18564 13268
rect 18524 12918 18552 13262
rect 18512 12912 18564 12918
rect 18512 12854 18564 12860
rect 18616 10742 18644 20198
rect 18708 18737 18736 20198
rect 20732 19514 20760 23582
rect 21744 23582 22062 23610
rect 20956 21788 21252 21808
rect 21012 21786 21036 21788
rect 21092 21786 21116 21788
rect 21172 21786 21196 21788
rect 21034 21734 21036 21786
rect 21098 21734 21110 21786
rect 21172 21734 21174 21786
rect 21012 21732 21036 21734
rect 21092 21732 21116 21734
rect 21172 21732 21196 21734
rect 20956 21712 21252 21732
rect 21454 21448 21510 21457
rect 21454 21383 21510 21392
rect 20956 20700 21252 20720
rect 21012 20698 21036 20700
rect 21092 20698 21116 20700
rect 21172 20698 21196 20700
rect 21034 20646 21036 20698
rect 21098 20646 21110 20698
rect 21172 20646 21174 20698
rect 21012 20644 21036 20646
rect 21092 20644 21116 20646
rect 21172 20644 21196 20646
rect 20956 20624 21252 20644
rect 21468 20602 21496 21383
rect 21456 20596 21508 20602
rect 21456 20538 21508 20544
rect 21468 20398 21496 20538
rect 21456 20392 21508 20398
rect 21456 20334 21508 20340
rect 21178 20224 21234 20233
rect 21178 20159 21234 20168
rect 21192 19922 21220 20159
rect 21180 19916 21232 19922
rect 21232 19876 21312 19904
rect 21180 19858 21232 19864
rect 20956 19612 21252 19632
rect 21012 19610 21036 19612
rect 21092 19610 21116 19612
rect 21172 19610 21196 19612
rect 21034 19558 21036 19610
rect 21098 19558 21110 19610
rect 21172 19558 21174 19610
rect 21012 19556 21036 19558
rect 21092 19556 21116 19558
rect 21172 19556 21196 19558
rect 20956 19536 21252 19556
rect 21284 19514 21312 19876
rect 21744 19514 21772 23582
rect 22006 23520 22062 23582
rect 22100 23588 22152 23594
rect 22100 23530 22152 23536
rect 23294 23588 23350 24000
rect 23294 23536 23296 23588
rect 23348 23536 23350 23588
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 21272 19508 21324 19514
rect 21272 19450 21324 19456
rect 21732 19508 21784 19514
rect 21732 19450 21784 19456
rect 18972 19168 19024 19174
rect 18972 19110 19024 19116
rect 20812 19168 20864 19174
rect 20812 19110 20864 19116
rect 18984 18873 19012 19110
rect 18970 18864 19026 18873
rect 18970 18799 19026 18808
rect 20626 18864 20682 18873
rect 20626 18799 20682 18808
rect 18694 18728 18750 18737
rect 18694 18663 18750 18672
rect 18696 17196 18748 17202
rect 18696 17138 18748 17144
rect 18708 16182 18736 17138
rect 18696 16176 18748 16182
rect 18696 16118 18748 16124
rect 18708 13326 18736 16118
rect 19340 14884 19392 14890
rect 19340 14826 19392 14832
rect 18880 13456 18932 13462
rect 18880 13398 18932 13404
rect 18696 13320 18748 13326
rect 18696 13262 18748 13268
rect 18708 12782 18736 13262
rect 18892 12986 18920 13398
rect 18880 12980 18932 12986
rect 18880 12922 18932 12928
rect 18696 12776 18748 12782
rect 18696 12718 18748 12724
rect 18696 11280 18748 11286
rect 18696 11222 18748 11228
rect 17960 10736 18012 10742
rect 17960 10678 18012 10684
rect 18604 10736 18656 10742
rect 18604 10678 18656 10684
rect 17316 10600 17368 10606
rect 17316 10542 17368 10548
rect 16856 10532 16908 10538
rect 16856 10474 16908 10480
rect 16868 10266 16896 10474
rect 16956 10364 17252 10384
rect 17012 10362 17036 10364
rect 17092 10362 17116 10364
rect 17172 10362 17196 10364
rect 17034 10310 17036 10362
rect 17098 10310 17110 10362
rect 17172 10310 17174 10362
rect 17012 10308 17036 10310
rect 17092 10308 17116 10310
rect 17172 10308 17196 10310
rect 16956 10288 17252 10308
rect 16856 10260 16908 10266
rect 16856 10202 16908 10208
rect 16868 9382 16896 10202
rect 17328 9586 17356 10542
rect 18616 10538 18644 10678
rect 18708 10674 18736 11222
rect 18788 11144 18840 11150
rect 18788 11086 18840 11092
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 17776 10532 17828 10538
rect 17776 10474 17828 10480
rect 18604 10532 18656 10538
rect 18604 10474 18656 10480
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17420 9926 17448 10406
rect 17788 10062 17816 10474
rect 18708 10266 18736 10610
rect 18800 10538 18828 11086
rect 19156 11076 19208 11082
rect 19156 11018 19208 11024
rect 18880 10736 18932 10742
rect 18880 10678 18932 10684
rect 18788 10532 18840 10538
rect 18788 10474 18840 10480
rect 18892 10470 18920 10678
rect 18880 10464 18932 10470
rect 18880 10406 18932 10412
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 18328 10192 18380 10198
rect 18328 10134 18380 10140
rect 17776 10056 17828 10062
rect 17776 9998 17828 10004
rect 17408 9920 17460 9926
rect 17408 9862 17460 9868
rect 17316 9580 17368 9586
rect 17316 9522 17368 9528
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16956 9276 17252 9296
rect 17012 9274 17036 9276
rect 17092 9274 17116 9276
rect 17172 9274 17196 9276
rect 17034 9222 17036 9274
rect 17098 9222 17110 9274
rect 17172 9222 17174 9274
rect 17012 9220 17036 9222
rect 17092 9220 17116 9222
rect 17172 9220 17196 9222
rect 16956 9200 17252 9220
rect 16764 8424 16816 8430
rect 16764 8366 16816 8372
rect 16212 8288 16264 8294
rect 16212 8230 16264 8236
rect 16224 8022 16252 8230
rect 16776 8090 16804 8366
rect 16956 8188 17252 8208
rect 17012 8186 17036 8188
rect 17092 8186 17116 8188
rect 17172 8186 17196 8188
rect 17034 8134 17036 8186
rect 17098 8134 17110 8186
rect 17172 8134 17174 8186
rect 17012 8132 17036 8134
rect 17092 8132 17116 8134
rect 17172 8132 17196 8134
rect 16956 8112 17252 8132
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 16212 8016 16264 8022
rect 16212 7958 16264 7964
rect 15936 7948 15988 7954
rect 15936 7890 15988 7896
rect 16856 7948 16908 7954
rect 16856 7890 16908 7896
rect 15660 7880 15712 7886
rect 15660 7822 15712 7828
rect 15672 7546 15700 7822
rect 15660 7540 15712 7546
rect 15660 7482 15712 7488
rect 15568 7472 15620 7478
rect 15568 7414 15620 7420
rect 15948 7410 15976 7890
rect 16488 7744 16540 7750
rect 16488 7686 16540 7692
rect 16500 7410 16528 7686
rect 15936 7404 15988 7410
rect 15764 7364 15936 7392
rect 15292 6316 15344 6322
rect 15292 6258 15344 6264
rect 15304 2514 15332 6258
rect 15476 5840 15528 5846
rect 15476 5782 15528 5788
rect 15488 5030 15516 5782
rect 15658 5400 15714 5409
rect 15658 5335 15714 5344
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 15384 4820 15436 4826
rect 15384 4762 15436 4768
rect 15396 3602 15424 4762
rect 15672 4758 15700 5335
rect 15660 4752 15712 4758
rect 15660 4694 15712 4700
rect 15476 4684 15528 4690
rect 15476 4626 15528 4632
rect 15568 4684 15620 4690
rect 15568 4626 15620 4632
rect 15488 3942 15516 4626
rect 15580 4282 15608 4626
rect 15568 4276 15620 4282
rect 15568 4218 15620 4224
rect 15476 3936 15528 3942
rect 15476 3878 15528 3884
rect 15384 3596 15436 3602
rect 15384 3538 15436 3544
rect 15396 2650 15424 3538
rect 15476 3392 15528 3398
rect 15476 3334 15528 3340
rect 15384 2644 15436 2650
rect 15384 2586 15436 2592
rect 15292 2508 15344 2514
rect 15292 2450 15344 2456
rect 15488 2009 15516 3334
rect 15580 3194 15608 4218
rect 15764 4214 15792 7364
rect 15936 7346 15988 7352
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 16304 7268 16356 7274
rect 16304 7210 16356 7216
rect 16028 7200 16080 7206
rect 15948 7160 16028 7188
rect 15948 6866 15976 7160
rect 16028 7142 16080 7148
rect 16316 6934 16344 7210
rect 16500 7002 16528 7346
rect 16868 7206 16896 7890
rect 16856 7200 16908 7206
rect 16856 7142 16908 7148
rect 16956 7100 17252 7120
rect 17012 7098 17036 7100
rect 17092 7098 17116 7100
rect 17172 7098 17196 7100
rect 17034 7046 17036 7098
rect 17098 7046 17110 7098
rect 17172 7046 17174 7098
rect 17012 7044 17036 7046
rect 17092 7044 17116 7046
rect 17172 7044 17196 7046
rect 16956 7024 17252 7044
rect 16488 6996 16540 7002
rect 16488 6938 16540 6944
rect 16304 6928 16356 6934
rect 16304 6870 16356 6876
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 17132 6860 17184 6866
rect 17132 6802 17184 6808
rect 15948 6118 15976 6802
rect 16028 6656 16080 6662
rect 16028 6598 16080 6604
rect 16488 6656 16540 6662
rect 16488 6598 16540 6604
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15752 4208 15804 4214
rect 15752 4150 15804 4156
rect 15752 3664 15804 3670
rect 15752 3606 15804 3612
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 15764 2922 15792 3606
rect 15752 2916 15804 2922
rect 15752 2858 15804 2864
rect 15764 2582 15792 2858
rect 15752 2576 15804 2582
rect 15752 2518 15804 2524
rect 15474 2000 15530 2009
rect 15474 1935 15530 1944
rect 15290 82 15346 480
rect 15212 54 15346 82
rect 15948 82 15976 6054
rect 16040 5914 16068 6598
rect 16500 6254 16528 6598
rect 16120 6248 16172 6254
rect 16120 6190 16172 6196
rect 16488 6248 16540 6254
rect 16488 6190 16540 6196
rect 16028 5908 16080 5914
rect 16028 5850 16080 5856
rect 16040 5234 16068 5850
rect 16132 5642 16160 6190
rect 16120 5636 16172 5642
rect 16120 5578 16172 5584
rect 16396 5568 16448 5574
rect 16396 5510 16448 5516
rect 16028 5228 16080 5234
rect 16028 5170 16080 5176
rect 16408 5098 16436 5510
rect 16396 5092 16448 5098
rect 16396 5034 16448 5040
rect 16500 4758 16528 6190
rect 16580 5704 16632 5710
rect 16580 5646 16632 5652
rect 16592 5234 16620 5646
rect 16580 5228 16632 5234
rect 16580 5170 16632 5176
rect 16488 4752 16540 4758
rect 16488 4694 16540 4700
rect 16304 4480 16356 4486
rect 16304 4422 16356 4428
rect 16212 4208 16264 4214
rect 16212 4150 16264 4156
rect 16120 4004 16172 4010
rect 16120 3946 16172 3952
rect 16132 3670 16160 3946
rect 16120 3664 16172 3670
rect 16120 3606 16172 3612
rect 16224 2990 16252 4150
rect 16316 4010 16344 4422
rect 16304 4004 16356 4010
rect 16304 3946 16356 3952
rect 16316 3738 16344 3946
rect 16304 3732 16356 3738
rect 16304 3674 16356 3680
rect 16592 3670 16620 5170
rect 16580 3664 16632 3670
rect 16580 3606 16632 3612
rect 16684 3602 16712 6598
rect 17144 6458 17172 6802
rect 16764 6452 16816 6458
rect 16764 6394 16816 6400
rect 17132 6452 17184 6458
rect 17132 6394 17184 6400
rect 16776 4146 16804 6394
rect 16856 6180 16908 6186
rect 16856 6122 16908 6128
rect 16868 5778 16896 6122
rect 16956 6012 17252 6032
rect 17012 6010 17036 6012
rect 17092 6010 17116 6012
rect 17172 6010 17196 6012
rect 17034 5958 17036 6010
rect 17098 5958 17110 6010
rect 17172 5958 17174 6010
rect 17012 5956 17036 5958
rect 17092 5956 17116 5958
rect 17172 5956 17196 5958
rect 16956 5936 17252 5956
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 16868 4826 16896 5714
rect 16956 4924 17252 4944
rect 17012 4922 17036 4924
rect 17092 4922 17116 4924
rect 17172 4922 17196 4924
rect 17034 4870 17036 4922
rect 17098 4870 17110 4922
rect 17172 4870 17174 4922
rect 17012 4868 17036 4870
rect 17092 4868 17116 4870
rect 17172 4868 17196 4870
rect 16956 4848 17252 4868
rect 16856 4820 16908 4826
rect 17328 4808 17356 9522
rect 17420 6934 17448 9862
rect 17788 9722 17816 9998
rect 17776 9716 17828 9722
rect 17776 9658 17828 9664
rect 18052 9444 18104 9450
rect 18052 9386 18104 9392
rect 18064 9110 18092 9386
rect 18340 9382 18368 10134
rect 19064 9648 19116 9654
rect 19168 9636 19196 11018
rect 19248 11008 19300 11014
rect 19248 10950 19300 10956
rect 19116 9608 19196 9636
rect 19064 9590 19116 9596
rect 18328 9376 18380 9382
rect 18328 9318 18380 9324
rect 18052 9104 18104 9110
rect 18052 9046 18104 9052
rect 17960 8968 18012 8974
rect 17960 8910 18012 8916
rect 17972 8566 18000 8910
rect 18064 8634 18092 9046
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 17960 8560 18012 8566
rect 17960 8502 18012 8508
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17512 8294 17540 8434
rect 18052 8424 18104 8430
rect 18052 8366 18104 8372
rect 17500 8288 17552 8294
rect 17500 8230 17552 8236
rect 17408 6928 17460 6934
rect 17408 6870 17460 6876
rect 17408 5840 17460 5846
rect 17512 5828 17540 8230
rect 18064 8090 18092 8366
rect 18340 8362 18368 9318
rect 18604 8968 18656 8974
rect 18418 8936 18474 8945
rect 18604 8910 18656 8916
rect 18418 8871 18474 8880
rect 18328 8356 18380 8362
rect 18328 8298 18380 8304
rect 18052 8084 18104 8090
rect 18052 8026 18104 8032
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17880 7546 17908 7958
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 18236 7336 18288 7342
rect 18236 7278 18288 7284
rect 17460 5800 17540 5828
rect 17408 5782 17460 5788
rect 17420 5030 17448 5782
rect 17408 5024 17460 5030
rect 17408 4966 17460 4972
rect 16856 4762 16908 4768
rect 17052 4780 17356 4808
rect 17052 4690 17080 4780
rect 17040 4684 17092 4690
rect 17040 4626 17092 4632
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 17052 4214 17080 4626
rect 17328 4282 17356 4626
rect 17316 4276 17368 4282
rect 17316 4218 17368 4224
rect 17040 4208 17092 4214
rect 17040 4150 17092 4156
rect 17420 4154 17448 4966
rect 17592 4616 17644 4622
rect 17592 4558 17644 4564
rect 17500 4548 17552 4554
rect 17500 4490 17552 4496
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 17328 4126 17448 4154
rect 17328 3942 17356 4126
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 16956 3836 17252 3856
rect 17012 3834 17036 3836
rect 17092 3834 17116 3836
rect 17172 3834 17196 3836
rect 17034 3782 17036 3834
rect 17098 3782 17110 3834
rect 17172 3782 17174 3834
rect 17012 3780 17036 3782
rect 17092 3780 17116 3782
rect 17172 3780 17196 3782
rect 16956 3760 17252 3780
rect 16672 3596 16724 3602
rect 16672 3538 16724 3544
rect 16212 2984 16264 2990
rect 16212 2926 16264 2932
rect 16956 2748 17252 2768
rect 17012 2746 17036 2748
rect 17092 2746 17116 2748
rect 17172 2746 17196 2748
rect 17034 2694 17036 2746
rect 17098 2694 17110 2746
rect 17172 2694 17174 2746
rect 17012 2692 17036 2694
rect 17092 2692 17116 2694
rect 17172 2692 17196 2694
rect 16956 2672 17252 2692
rect 17328 2582 17356 3878
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 17420 3097 17448 3334
rect 17406 3088 17462 3097
rect 17406 3023 17462 3032
rect 17316 2576 17368 2582
rect 17316 2518 17368 2524
rect 17040 1760 17092 1766
rect 17040 1702 17092 1708
rect 16118 82 16174 480
rect 15948 54 16174 82
rect 15290 0 15346 54
rect 16118 0 16174 54
rect 16946 82 17002 480
rect 17052 82 17080 1702
rect 16946 54 17080 82
rect 17512 82 17540 4490
rect 17604 4146 17632 4558
rect 17592 4140 17644 4146
rect 17592 4082 17644 4088
rect 18052 4140 18104 4146
rect 18052 4082 18104 4088
rect 18064 3738 18092 4082
rect 18052 3732 18104 3738
rect 18052 3674 18104 3680
rect 17868 2848 17920 2854
rect 17868 2790 17920 2796
rect 17880 2650 17908 2790
rect 17868 2644 17920 2650
rect 17868 2586 17920 2592
rect 18248 2378 18276 7278
rect 18328 6248 18380 6254
rect 18432 6236 18460 8871
rect 18616 8498 18644 8910
rect 18604 8492 18656 8498
rect 18604 8434 18656 8440
rect 18616 7970 18644 8434
rect 18972 8288 19024 8294
rect 18972 8230 19024 8236
rect 18984 8022 19012 8230
rect 19168 8022 19196 9608
rect 19260 9586 19288 10950
rect 19248 9580 19300 9586
rect 19248 9522 19300 9528
rect 19260 9178 19288 9522
rect 19248 9172 19300 9178
rect 19248 9114 19300 9120
rect 18972 8016 19024 8022
rect 18524 7942 18736 7970
rect 18972 7958 19024 7964
rect 19156 8016 19208 8022
rect 19156 7958 19208 7964
rect 18524 7886 18552 7942
rect 18512 7880 18564 7886
rect 18512 7822 18564 7828
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 18512 6928 18564 6934
rect 18512 6870 18564 6876
rect 18380 6208 18460 6236
rect 18328 6190 18380 6196
rect 18340 5273 18368 6190
rect 18420 6112 18472 6118
rect 18420 6054 18472 6060
rect 18326 5264 18382 5273
rect 18432 5234 18460 6054
rect 18524 5914 18552 6870
rect 18616 6798 18644 7822
rect 18708 6798 18736 7942
rect 19248 7404 19300 7410
rect 19352 7392 19380 14826
rect 19892 12640 19944 12646
rect 19892 12582 19944 12588
rect 19904 12306 19932 12582
rect 19892 12300 19944 12306
rect 19892 12242 19944 12248
rect 19892 10464 19944 10470
rect 19892 10406 19944 10412
rect 19904 9450 19932 10406
rect 20168 9988 20220 9994
rect 20168 9930 20220 9936
rect 19892 9444 19944 9450
rect 19892 9386 19944 9392
rect 19524 8288 19576 8294
rect 19524 8230 19576 8236
rect 19800 8288 19852 8294
rect 19800 8230 19852 8236
rect 19536 8090 19564 8230
rect 19524 8084 19576 8090
rect 19524 8026 19576 8032
rect 19432 7744 19484 7750
rect 19432 7686 19484 7692
rect 19300 7364 19380 7392
rect 19248 7346 19300 7352
rect 19444 7274 19472 7686
rect 19536 7478 19564 8026
rect 19812 7750 19840 8230
rect 19800 7744 19852 7750
rect 19800 7686 19852 7692
rect 19812 7546 19840 7686
rect 19800 7540 19852 7546
rect 19800 7482 19852 7488
rect 19524 7472 19576 7478
rect 19524 7414 19576 7420
rect 19536 7274 19564 7414
rect 19904 7410 19932 9386
rect 19984 8356 20036 8362
rect 19984 8298 20036 8304
rect 19996 8090 20024 8298
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 19892 7404 19944 7410
rect 19892 7346 19944 7352
rect 19432 7268 19484 7274
rect 19432 7210 19484 7216
rect 19524 7268 19576 7274
rect 19524 7210 19576 7216
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 18696 6792 18748 6798
rect 18696 6734 18748 6740
rect 18616 6458 18644 6734
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 19248 6316 19300 6322
rect 19248 6258 19300 6264
rect 18512 5908 18564 5914
rect 18512 5850 18564 5856
rect 18512 5704 18564 5710
rect 18512 5646 18564 5652
rect 18524 5370 18552 5646
rect 18512 5364 18564 5370
rect 18512 5306 18564 5312
rect 19260 5302 19288 6258
rect 19352 6186 19380 6598
rect 19340 6180 19392 6186
rect 19340 6122 19392 6128
rect 19352 5914 19380 6122
rect 19444 5914 19472 7210
rect 19616 7200 19668 7206
rect 19616 7142 19668 7148
rect 19340 5908 19392 5914
rect 19340 5850 19392 5856
rect 19432 5908 19484 5914
rect 19432 5850 19484 5856
rect 19352 5760 19380 5850
rect 19352 5732 19472 5760
rect 19340 5636 19392 5642
rect 19340 5578 19392 5584
rect 19248 5296 19300 5302
rect 19248 5238 19300 5244
rect 18326 5199 18382 5208
rect 18420 5228 18472 5234
rect 18420 5170 18472 5176
rect 18788 5092 18840 5098
rect 18788 5034 18840 5040
rect 18800 4758 18828 5034
rect 19260 4842 19288 5238
rect 19076 4814 19288 4842
rect 18788 4752 18840 4758
rect 18788 4694 18840 4700
rect 18800 4282 18828 4694
rect 18696 4276 18748 4282
rect 18696 4218 18748 4224
rect 18788 4276 18840 4282
rect 18788 4218 18840 4224
rect 18604 4072 18656 4078
rect 18604 4014 18656 4020
rect 18420 3664 18472 3670
rect 18420 3606 18472 3612
rect 18432 3194 18460 3606
rect 18420 3188 18472 3194
rect 18420 3130 18472 3136
rect 18616 2922 18644 4014
rect 18708 3194 18736 4218
rect 19076 4146 19104 4814
rect 19352 4758 19380 5578
rect 19444 5370 19472 5732
rect 19628 5710 19656 7142
rect 19616 5704 19668 5710
rect 19616 5646 19668 5652
rect 19432 5364 19484 5370
rect 19432 5306 19484 5312
rect 19892 5092 19944 5098
rect 19892 5034 19944 5040
rect 19340 4752 19392 4758
rect 19392 4712 19472 4740
rect 19340 4694 19392 4700
rect 19444 4154 19472 4712
rect 18788 4140 18840 4146
rect 18788 4082 18840 4088
rect 19064 4140 19116 4146
rect 19064 4082 19116 4088
rect 19352 4126 19472 4154
rect 19708 4208 19760 4214
rect 19708 4150 19760 4156
rect 18800 3534 18828 4082
rect 19352 4078 19380 4126
rect 19340 4072 19392 4078
rect 19340 4014 19392 4020
rect 18880 4004 18932 4010
rect 18880 3946 18932 3952
rect 18892 3534 18920 3946
rect 18972 3936 19024 3942
rect 18972 3878 19024 3884
rect 19156 3936 19208 3942
rect 19156 3878 19208 3884
rect 18984 3670 19012 3878
rect 18972 3664 19024 3670
rect 18972 3606 19024 3612
rect 18788 3528 18840 3534
rect 18788 3470 18840 3476
rect 18880 3528 18932 3534
rect 18880 3470 18932 3476
rect 18696 3188 18748 3194
rect 18696 3130 18748 3136
rect 18800 3126 18828 3470
rect 18788 3120 18840 3126
rect 18788 3062 18840 3068
rect 18892 3058 18920 3470
rect 18880 3052 18932 3058
rect 18880 2994 18932 3000
rect 18604 2916 18656 2922
rect 18604 2858 18656 2864
rect 19064 2916 19116 2922
rect 19064 2858 19116 2864
rect 18616 2378 18644 2858
rect 19076 2582 19104 2858
rect 19168 2582 19196 3878
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 19352 2961 19380 2994
rect 19338 2952 19394 2961
rect 19338 2887 19394 2896
rect 19064 2576 19116 2582
rect 19064 2518 19116 2524
rect 19156 2576 19208 2582
rect 19156 2518 19208 2524
rect 19064 2440 19116 2446
rect 19168 2428 19196 2518
rect 19116 2400 19196 2428
rect 19064 2382 19116 2388
rect 18236 2372 18288 2378
rect 18236 2314 18288 2320
rect 18604 2372 18656 2378
rect 18604 2314 18656 2320
rect 18880 2304 18932 2310
rect 18880 2246 18932 2252
rect 17774 82 17830 480
rect 17512 54 17830 82
rect 16946 0 17002 54
rect 17774 0 17830 54
rect 18602 82 18658 480
rect 18892 82 18920 2246
rect 18602 54 18920 82
rect 19430 82 19486 480
rect 19720 82 19748 4150
rect 19904 4010 19932 5034
rect 20180 4282 20208 9930
rect 20444 6860 20496 6866
rect 20444 6802 20496 6808
rect 20456 6186 20484 6802
rect 20640 6458 20668 18799
rect 20824 18329 20852 19110
rect 20956 18524 21252 18544
rect 21012 18522 21036 18524
rect 21092 18522 21116 18524
rect 21172 18522 21196 18524
rect 21034 18470 21036 18522
rect 21098 18470 21110 18522
rect 21172 18470 21174 18522
rect 21012 18468 21036 18470
rect 21092 18468 21116 18470
rect 21172 18468 21196 18470
rect 20956 18448 21252 18468
rect 20810 18320 20866 18329
rect 20810 18255 20866 18264
rect 21270 17640 21326 17649
rect 21270 17575 21326 17584
rect 20956 17436 21252 17456
rect 21012 17434 21036 17436
rect 21092 17434 21116 17436
rect 21172 17434 21196 17436
rect 21034 17382 21036 17434
rect 21098 17382 21110 17434
rect 21172 17382 21174 17434
rect 21012 17380 21036 17382
rect 21092 17380 21116 17382
rect 21172 17380 21196 17382
rect 20956 17360 21252 17380
rect 21284 17338 21312 17575
rect 21272 17332 21324 17338
rect 21272 17274 21324 17280
rect 20812 17128 20864 17134
rect 20812 17070 20864 17076
rect 20824 16250 20852 17070
rect 21454 16416 21510 16425
rect 20956 16348 21252 16368
rect 21454 16351 21510 16360
rect 21012 16346 21036 16348
rect 21092 16346 21116 16348
rect 21172 16346 21196 16348
rect 21034 16294 21036 16346
rect 21098 16294 21110 16346
rect 21172 16294 21174 16346
rect 21012 16292 21036 16294
rect 21092 16292 21116 16294
rect 21172 16292 21196 16294
rect 20956 16272 21252 16292
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 21468 15706 21496 16351
rect 21456 15700 21508 15706
rect 21456 15642 21508 15648
rect 20812 15564 20864 15570
rect 20812 15506 20864 15512
rect 20824 14890 20852 15506
rect 21270 15464 21326 15473
rect 21270 15399 21326 15408
rect 20956 15260 21252 15280
rect 21012 15258 21036 15260
rect 21092 15258 21116 15260
rect 21172 15258 21196 15260
rect 21034 15206 21036 15258
rect 21098 15206 21110 15258
rect 21172 15206 21174 15258
rect 21012 15204 21036 15206
rect 21092 15204 21116 15206
rect 21172 15204 21196 15206
rect 20956 15184 21252 15204
rect 21284 15162 21312 15399
rect 21272 15156 21324 15162
rect 21272 15098 21324 15104
rect 20812 14884 20864 14890
rect 20812 14826 20864 14832
rect 20956 14172 21252 14192
rect 21012 14170 21036 14172
rect 21092 14170 21116 14172
rect 21172 14170 21196 14172
rect 21034 14118 21036 14170
rect 21098 14118 21110 14170
rect 21172 14118 21174 14170
rect 21012 14116 21036 14118
rect 21092 14116 21116 14118
rect 21172 14116 21196 14118
rect 20956 14096 21252 14116
rect 21086 13968 21142 13977
rect 21086 13903 21142 13912
rect 21100 13530 21128 13903
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 20812 13388 20864 13394
rect 20812 13330 20864 13336
rect 20824 12918 20852 13330
rect 20956 13084 21252 13104
rect 21012 13082 21036 13084
rect 21092 13082 21116 13084
rect 21172 13082 21196 13084
rect 21034 13030 21036 13082
rect 21098 13030 21110 13082
rect 21172 13030 21174 13082
rect 21012 13028 21036 13030
rect 21092 13028 21116 13030
rect 21172 13028 21196 13030
rect 20956 13008 21252 13028
rect 20812 12912 20864 12918
rect 20812 12854 20864 12860
rect 20720 12776 20772 12782
rect 20720 12718 20772 12724
rect 20732 11665 20760 12718
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 20824 11898 20852 12242
rect 20956 11996 21252 12016
rect 21012 11994 21036 11996
rect 21092 11994 21116 11996
rect 21172 11994 21196 11996
rect 21034 11942 21036 11994
rect 21098 11942 21110 11994
rect 21172 11942 21174 11994
rect 21012 11940 21036 11942
rect 21092 11940 21116 11942
rect 21172 11940 21196 11942
rect 20956 11920 21252 11940
rect 20812 11892 20864 11898
rect 20812 11834 20864 11840
rect 20718 11656 20774 11665
rect 20718 11591 20774 11600
rect 22112 11218 22140 23530
rect 23294 23520 23350 23536
rect 23308 23499 23336 23520
rect 22466 22672 22522 22681
rect 22466 22607 22522 22616
rect 22480 19514 22508 22607
rect 22468 19508 22520 19514
rect 22468 19450 22520 19456
rect 23572 12096 23624 12102
rect 23572 12038 23624 12044
rect 23584 11937 23612 12038
rect 23570 11928 23626 11937
rect 23570 11863 23626 11872
rect 20812 11212 20864 11218
rect 20812 11154 20864 11160
rect 22100 11212 22152 11218
rect 22100 11154 22152 11160
rect 20824 10810 20852 11154
rect 20956 10908 21252 10928
rect 21012 10906 21036 10908
rect 21092 10906 21116 10908
rect 21172 10906 21196 10908
rect 21034 10854 21036 10906
rect 21098 10854 21110 10906
rect 21172 10854 21174 10906
rect 21012 10852 21036 10854
rect 21092 10852 21116 10854
rect 21172 10852 21196 10854
rect 20956 10832 21252 10852
rect 20812 10804 20864 10810
rect 20812 10746 20864 10752
rect 21086 10296 21142 10305
rect 21086 10231 21142 10240
rect 20720 10124 20772 10130
rect 20720 10066 20772 10072
rect 20732 9382 20760 10066
rect 21100 9994 21128 10231
rect 21088 9988 21140 9994
rect 21088 9930 21140 9936
rect 20956 9820 21252 9840
rect 21012 9818 21036 9820
rect 21092 9818 21116 9820
rect 21172 9818 21196 9820
rect 21034 9766 21036 9818
rect 21098 9766 21110 9818
rect 21172 9766 21174 9818
rect 21012 9764 21036 9766
rect 21092 9764 21116 9766
rect 21172 9764 21196 9766
rect 20956 9744 21252 9764
rect 20810 9616 20866 9625
rect 20810 9551 20866 9560
rect 20720 9376 20772 9382
rect 20720 9318 20772 9324
rect 20628 6452 20680 6458
rect 20628 6394 20680 6400
rect 20444 6180 20496 6186
rect 20444 6122 20496 6128
rect 20456 5234 20484 6122
rect 20732 5409 20760 9318
rect 20824 9110 20852 9551
rect 20812 9104 20864 9110
rect 20812 9046 20864 9052
rect 21272 9036 21324 9042
rect 21272 8978 21324 8984
rect 20956 8732 21252 8752
rect 21012 8730 21036 8732
rect 21092 8730 21116 8732
rect 21172 8730 21196 8732
rect 21034 8678 21036 8730
rect 21098 8678 21110 8730
rect 21172 8678 21174 8730
rect 21012 8676 21036 8678
rect 21092 8676 21116 8678
rect 21172 8676 21196 8678
rect 20956 8656 21252 8676
rect 21284 8294 21312 8978
rect 21272 8288 21324 8294
rect 21272 8230 21324 8236
rect 23204 8288 23256 8294
rect 23204 8230 23256 8236
rect 20956 7644 21252 7664
rect 21012 7642 21036 7644
rect 21092 7642 21116 7644
rect 21172 7642 21196 7644
rect 21034 7590 21036 7642
rect 21098 7590 21110 7642
rect 21172 7590 21174 7642
rect 21012 7588 21036 7590
rect 21092 7588 21116 7590
rect 21172 7588 21196 7590
rect 20956 7568 21252 7588
rect 21362 7576 21418 7585
rect 21362 7511 21418 7520
rect 21376 7002 21404 7511
rect 21364 6996 21416 7002
rect 21364 6938 21416 6944
rect 20956 6556 21252 6576
rect 21012 6554 21036 6556
rect 21092 6554 21116 6556
rect 21172 6554 21196 6556
rect 21034 6502 21036 6554
rect 21098 6502 21110 6554
rect 21172 6502 21174 6554
rect 21012 6500 21036 6502
rect 21092 6500 21116 6502
rect 21172 6500 21196 6502
rect 20956 6480 21252 6500
rect 21454 5808 21510 5817
rect 21454 5743 21510 5752
rect 21548 5772 21600 5778
rect 20956 5468 21252 5488
rect 21012 5466 21036 5468
rect 21092 5466 21116 5468
rect 21172 5466 21196 5468
rect 21034 5414 21036 5466
rect 21098 5414 21110 5466
rect 21172 5414 21174 5466
rect 21012 5412 21036 5414
rect 21092 5412 21116 5414
rect 21172 5412 21196 5414
rect 20718 5400 20774 5409
rect 20956 5392 21252 5412
rect 20718 5335 20774 5344
rect 20444 5228 20496 5234
rect 20444 5170 20496 5176
rect 20628 5228 20680 5234
rect 20628 5170 20680 5176
rect 20168 4276 20220 4282
rect 20168 4218 20220 4224
rect 19892 4004 19944 4010
rect 19892 3946 19944 3952
rect 19904 3738 19932 3946
rect 19892 3732 19944 3738
rect 19892 3674 19944 3680
rect 20076 2984 20128 2990
rect 20076 2926 20128 2932
rect 20088 2582 20116 2926
rect 20168 2848 20220 2854
rect 20168 2790 20220 2796
rect 20180 2650 20208 2790
rect 20168 2644 20220 2650
rect 20168 2586 20220 2592
rect 20076 2576 20128 2582
rect 20076 2518 20128 2524
rect 20456 2514 20484 5170
rect 20536 5160 20588 5166
rect 20640 5137 20668 5170
rect 20536 5102 20588 5108
rect 20626 5128 20682 5137
rect 20444 2508 20496 2514
rect 20444 2450 20496 2456
rect 19430 54 19748 82
rect 20258 82 20314 480
rect 20548 82 20576 5102
rect 20626 5063 20682 5072
rect 20720 5092 20772 5098
rect 20720 5034 20772 5040
rect 20626 4312 20682 4321
rect 20626 4247 20682 4256
rect 20640 3641 20668 4247
rect 20626 3632 20682 3641
rect 20626 3567 20682 3576
rect 20732 2922 20760 5034
rect 21468 4865 21496 5743
rect 21548 5714 21600 5720
rect 21560 5030 21588 5714
rect 21548 5024 21600 5030
rect 21548 4966 21600 4972
rect 21454 4856 21510 4865
rect 21454 4791 21510 4800
rect 20812 4684 20864 4690
rect 20812 4626 20864 4632
rect 20824 4214 20852 4626
rect 20956 4380 21252 4400
rect 21012 4378 21036 4380
rect 21092 4378 21116 4380
rect 21172 4378 21196 4380
rect 21034 4326 21036 4378
rect 21098 4326 21110 4378
rect 21172 4326 21174 4378
rect 21012 4324 21036 4326
rect 21092 4324 21116 4326
rect 21172 4324 21196 4326
rect 20956 4304 21252 4324
rect 20812 4208 20864 4214
rect 20812 4150 20864 4156
rect 21364 3936 21416 3942
rect 21364 3878 21416 3884
rect 21272 3596 21324 3602
rect 21272 3538 21324 3544
rect 20956 3292 21252 3312
rect 21012 3290 21036 3292
rect 21092 3290 21116 3292
rect 21172 3290 21196 3292
rect 21034 3238 21036 3290
rect 21098 3238 21110 3290
rect 21172 3238 21174 3290
rect 21012 3236 21036 3238
rect 21092 3236 21116 3238
rect 21172 3236 21196 3238
rect 20956 3216 21252 3236
rect 20720 2916 20772 2922
rect 20720 2858 20772 2864
rect 21284 2854 21312 3538
rect 21272 2848 21324 2854
rect 21272 2790 21324 2796
rect 20956 2204 21252 2224
rect 21012 2202 21036 2204
rect 21092 2202 21116 2204
rect 21172 2202 21196 2204
rect 21034 2150 21036 2202
rect 21098 2150 21110 2202
rect 21172 2150 21174 2202
rect 21012 2148 21036 2150
rect 21092 2148 21116 2150
rect 21172 2148 21196 2150
rect 20956 2128 21252 2148
rect 20258 54 20576 82
rect 21086 82 21142 480
rect 21376 82 21404 3878
rect 21086 54 21404 82
rect 21560 82 21588 4966
rect 22468 2848 22520 2854
rect 22468 2790 22520 2796
rect 21914 82 21970 480
rect 21560 54 21970 82
rect 22480 82 22508 2790
rect 22742 82 22798 480
rect 22480 54 22798 82
rect 23216 82 23244 8230
rect 23570 6896 23626 6905
rect 23570 6831 23626 6840
rect 23386 5672 23442 5681
rect 23584 5658 23612 6831
rect 23442 5630 23612 5658
rect 23386 5607 23442 5616
rect 23570 82 23626 480
rect 23216 54 23626 82
rect 18602 0 18658 54
rect 19430 0 19486 54
rect 20258 0 20314 54
rect 21086 0 21142 54
rect 21914 0 21970 54
rect 22742 0 22798 54
rect 23570 0 23626 54
<< via2 >>
rect 1582 22616 1638 22672
rect 110 20304 166 20360
rect 1858 21256 1914 21312
rect 110 18944 166 19000
rect 110 17584 166 17640
rect 110 16088 166 16144
rect 2502 19216 2558 19272
rect 110 13368 166 13424
rect 1582 11328 1638 11384
rect 1582 10240 1638 10296
rect 1582 8608 1638 8664
rect 1490 7248 1546 7304
rect 1858 7112 1914 7168
rect 110 2080 166 2136
rect 1582 4392 1638 4448
rect 4956 21786 5012 21788
rect 5036 21786 5092 21788
rect 5116 21786 5172 21788
rect 5196 21786 5252 21788
rect 4956 21734 4982 21786
rect 4982 21734 5012 21786
rect 5036 21734 5046 21786
rect 5046 21734 5092 21786
rect 5116 21734 5162 21786
rect 5162 21734 5172 21786
rect 5196 21734 5226 21786
rect 5226 21734 5252 21786
rect 4956 21732 5012 21734
rect 5036 21732 5092 21734
rect 5116 21732 5172 21734
rect 5196 21732 5252 21734
rect 4956 20698 5012 20700
rect 5036 20698 5092 20700
rect 5116 20698 5172 20700
rect 5196 20698 5252 20700
rect 4956 20646 4982 20698
rect 4982 20646 5012 20698
rect 5036 20646 5046 20698
rect 5046 20646 5092 20698
rect 5116 20646 5162 20698
rect 5162 20646 5172 20698
rect 5196 20646 5226 20698
rect 5226 20646 5252 20698
rect 4956 20644 5012 20646
rect 5036 20644 5092 20646
rect 5116 20644 5172 20646
rect 5196 20644 5252 20646
rect 3422 14184 3478 14240
rect 4956 19610 5012 19612
rect 5036 19610 5092 19612
rect 5116 19610 5172 19612
rect 5196 19610 5252 19612
rect 4956 19558 4982 19610
rect 4982 19558 5012 19610
rect 5036 19558 5046 19610
rect 5046 19558 5092 19610
rect 5116 19558 5162 19610
rect 5162 19558 5172 19610
rect 5196 19558 5226 19610
rect 5226 19558 5252 19610
rect 4956 19556 5012 19558
rect 5036 19556 5092 19558
rect 5116 19556 5172 19558
rect 5196 19556 5252 19558
rect 4956 18522 5012 18524
rect 5036 18522 5092 18524
rect 5116 18522 5172 18524
rect 5196 18522 5252 18524
rect 4956 18470 4982 18522
rect 4982 18470 5012 18522
rect 5036 18470 5046 18522
rect 5046 18470 5092 18522
rect 5116 18470 5162 18522
rect 5162 18470 5172 18522
rect 5196 18470 5226 18522
rect 5226 18470 5252 18522
rect 4956 18468 5012 18470
rect 5036 18468 5092 18470
rect 5116 18468 5172 18470
rect 5196 18468 5252 18470
rect 3698 11736 3754 11792
rect 4956 17434 5012 17436
rect 5036 17434 5092 17436
rect 5116 17434 5172 17436
rect 5196 17434 5252 17436
rect 4956 17382 4982 17434
rect 4982 17382 5012 17434
rect 5036 17382 5046 17434
rect 5046 17382 5092 17434
rect 5116 17382 5162 17434
rect 5162 17382 5172 17434
rect 5196 17382 5226 17434
rect 5226 17382 5252 17434
rect 4956 17380 5012 17382
rect 5036 17380 5092 17382
rect 5116 17380 5172 17382
rect 5196 17380 5252 17382
rect 4956 16346 5012 16348
rect 5036 16346 5092 16348
rect 5116 16346 5172 16348
rect 5196 16346 5252 16348
rect 4956 16294 4982 16346
rect 4982 16294 5012 16346
rect 5036 16294 5046 16346
rect 5046 16294 5092 16346
rect 5116 16294 5162 16346
rect 5162 16294 5172 16346
rect 5196 16294 5226 16346
rect 5226 16294 5252 16346
rect 4956 16292 5012 16294
rect 5036 16292 5092 16294
rect 5116 16292 5172 16294
rect 5196 16292 5252 16294
rect 4956 15258 5012 15260
rect 5036 15258 5092 15260
rect 5116 15258 5172 15260
rect 5196 15258 5252 15260
rect 4956 15206 4982 15258
rect 4982 15206 5012 15258
rect 5036 15206 5046 15258
rect 5046 15206 5092 15258
rect 5116 15206 5162 15258
rect 5162 15206 5172 15258
rect 5196 15206 5226 15258
rect 5226 15206 5252 15258
rect 4956 15204 5012 15206
rect 5036 15204 5092 15206
rect 5116 15204 5172 15206
rect 5196 15204 5252 15206
rect 4956 14170 5012 14172
rect 5036 14170 5092 14172
rect 5116 14170 5172 14172
rect 5196 14170 5252 14172
rect 4956 14118 4982 14170
rect 4982 14118 5012 14170
rect 5036 14118 5046 14170
rect 5046 14118 5092 14170
rect 5116 14118 5162 14170
rect 5162 14118 5172 14170
rect 5196 14118 5226 14170
rect 5226 14118 5252 14170
rect 4956 14116 5012 14118
rect 5036 14116 5092 14118
rect 5116 14116 5172 14118
rect 5196 14116 5252 14118
rect 4956 13082 5012 13084
rect 5036 13082 5092 13084
rect 5116 13082 5172 13084
rect 5196 13082 5252 13084
rect 4956 13030 4982 13082
rect 4982 13030 5012 13082
rect 5036 13030 5046 13082
rect 5046 13030 5092 13082
rect 5116 13030 5162 13082
rect 5162 13030 5172 13082
rect 5196 13030 5226 13082
rect 5226 13030 5252 13082
rect 4956 13028 5012 13030
rect 5036 13028 5092 13030
rect 5116 13028 5172 13030
rect 5196 13028 5252 13030
rect 6826 18808 6882 18864
rect 8956 21242 9012 21244
rect 9036 21242 9092 21244
rect 9116 21242 9172 21244
rect 9196 21242 9252 21244
rect 8956 21190 8982 21242
rect 8982 21190 9012 21242
rect 9036 21190 9046 21242
rect 9046 21190 9092 21242
rect 9116 21190 9162 21242
rect 9162 21190 9172 21242
rect 9196 21190 9226 21242
rect 9226 21190 9252 21242
rect 8956 21188 9012 21190
rect 9036 21188 9092 21190
rect 9116 21188 9172 21190
rect 9196 21188 9252 21190
rect 7378 18264 7434 18320
rect 4956 11994 5012 11996
rect 5036 11994 5092 11996
rect 5116 11994 5172 11996
rect 5196 11994 5252 11996
rect 4956 11942 4982 11994
rect 4982 11942 5012 11994
rect 5036 11942 5046 11994
rect 5046 11942 5092 11994
rect 5116 11942 5162 11994
rect 5162 11942 5172 11994
rect 5196 11942 5226 11994
rect 5226 11942 5252 11994
rect 4956 11940 5012 11942
rect 5036 11940 5092 11942
rect 5116 11940 5172 11942
rect 5196 11940 5252 11942
rect 5446 11600 5502 11656
rect 4956 10906 5012 10908
rect 5036 10906 5092 10908
rect 5116 10906 5172 10908
rect 5196 10906 5252 10908
rect 4956 10854 4982 10906
rect 4982 10854 5012 10906
rect 5036 10854 5046 10906
rect 5046 10854 5092 10906
rect 5116 10854 5162 10906
rect 5162 10854 5172 10906
rect 5196 10854 5226 10906
rect 5226 10854 5252 10906
rect 4956 10852 5012 10854
rect 5036 10852 5092 10854
rect 5116 10852 5172 10854
rect 5196 10852 5252 10854
rect 4066 9560 4122 9616
rect 3422 8472 3478 8528
rect 2226 6840 2282 6896
rect 1582 3168 1638 3224
rect 2042 2488 2098 2544
rect 1950 1264 2006 1320
rect 3974 3984 4030 4040
rect 4956 9818 5012 9820
rect 5036 9818 5092 9820
rect 5116 9818 5172 9820
rect 5196 9818 5252 9820
rect 4956 9766 4982 9818
rect 4982 9766 5012 9818
rect 5036 9766 5046 9818
rect 5046 9766 5092 9818
rect 5116 9766 5162 9818
rect 5162 9766 5172 9818
rect 5196 9766 5226 9818
rect 5226 9766 5252 9818
rect 4956 9764 5012 9766
rect 5036 9764 5092 9766
rect 5116 9764 5172 9766
rect 5196 9764 5252 9766
rect 5814 9560 5870 9616
rect 4956 8730 5012 8732
rect 5036 8730 5092 8732
rect 5116 8730 5172 8732
rect 5196 8730 5252 8732
rect 4956 8678 4982 8730
rect 4982 8678 5012 8730
rect 5036 8678 5046 8730
rect 5046 8678 5092 8730
rect 5116 8678 5162 8730
rect 5162 8678 5172 8730
rect 5196 8678 5226 8730
rect 5226 8678 5252 8730
rect 4956 8676 5012 8678
rect 5036 8676 5092 8678
rect 5116 8676 5172 8678
rect 5196 8676 5252 8678
rect 4956 7642 5012 7644
rect 5036 7642 5092 7644
rect 5116 7642 5172 7644
rect 5196 7642 5252 7644
rect 4956 7590 4982 7642
rect 4982 7590 5012 7642
rect 5036 7590 5046 7642
rect 5046 7590 5092 7642
rect 5116 7590 5162 7642
rect 5162 7590 5172 7642
rect 5196 7590 5226 7642
rect 5226 7590 5252 7642
rect 4956 7588 5012 7590
rect 5036 7588 5092 7590
rect 5116 7588 5172 7590
rect 5196 7588 5252 7590
rect 4956 6554 5012 6556
rect 5036 6554 5092 6556
rect 5116 6554 5172 6556
rect 5196 6554 5252 6556
rect 4956 6502 4982 6554
rect 4982 6502 5012 6554
rect 5036 6502 5046 6554
rect 5046 6502 5092 6554
rect 5116 6502 5162 6554
rect 5162 6502 5172 6554
rect 5196 6502 5226 6554
rect 5226 6502 5252 6554
rect 4956 6500 5012 6502
rect 5036 6500 5092 6502
rect 5116 6500 5172 6502
rect 5196 6500 5252 6502
rect 4956 5466 5012 5468
rect 5036 5466 5092 5468
rect 5116 5466 5172 5468
rect 5196 5466 5252 5468
rect 4956 5414 4982 5466
rect 4982 5414 5012 5466
rect 5036 5414 5046 5466
rect 5046 5414 5092 5466
rect 5116 5414 5162 5466
rect 5162 5414 5172 5466
rect 5196 5414 5226 5466
rect 5226 5414 5252 5466
rect 4956 5412 5012 5414
rect 5036 5412 5092 5414
rect 5116 5412 5172 5414
rect 5196 5412 5252 5414
rect 4956 4378 5012 4380
rect 5036 4378 5092 4380
rect 5116 4378 5172 4380
rect 5196 4378 5252 4380
rect 4956 4326 4982 4378
rect 4982 4326 5012 4378
rect 5036 4326 5046 4378
rect 5046 4326 5092 4378
rect 5116 4326 5162 4378
rect 5162 4326 5172 4378
rect 5196 4326 5226 4378
rect 5226 4326 5252 4378
rect 4956 4324 5012 4326
rect 5036 4324 5092 4326
rect 5116 4324 5172 4326
rect 5196 4324 5252 4326
rect 4434 2488 4490 2544
rect 4956 3290 5012 3292
rect 5036 3290 5092 3292
rect 5116 3290 5172 3292
rect 5196 3290 5252 3292
rect 4956 3238 4982 3290
rect 4982 3238 5012 3290
rect 5036 3238 5046 3290
rect 5046 3238 5092 3290
rect 5116 3238 5162 3290
rect 5162 3238 5172 3290
rect 5196 3238 5226 3290
rect 5226 3238 5252 3290
rect 4956 3236 5012 3238
rect 5036 3236 5092 3238
rect 5116 3236 5172 3238
rect 5196 3236 5252 3238
rect 4894 2796 4896 2816
rect 4896 2796 4948 2816
rect 4948 2796 4950 2816
rect 4894 2760 4950 2796
rect 4956 2202 5012 2204
rect 5036 2202 5092 2204
rect 5116 2202 5172 2204
rect 5196 2202 5252 2204
rect 4956 2150 4982 2202
rect 4982 2150 5012 2202
rect 5036 2150 5046 2202
rect 5046 2150 5092 2202
rect 5116 2150 5162 2202
rect 5162 2150 5172 2202
rect 5196 2150 5226 2202
rect 5226 2150 5252 2202
rect 4956 2148 5012 2150
rect 5036 2148 5092 2150
rect 5116 2148 5172 2150
rect 5196 2148 5252 2150
rect 5538 4256 5594 4312
rect 8956 20154 9012 20156
rect 9036 20154 9092 20156
rect 9116 20154 9172 20156
rect 9196 20154 9252 20156
rect 8956 20102 8982 20154
rect 8982 20102 9012 20154
rect 9036 20102 9046 20154
rect 9046 20102 9092 20154
rect 9116 20102 9162 20154
rect 9162 20102 9172 20154
rect 9196 20102 9226 20154
rect 9226 20102 9252 20154
rect 8956 20100 9012 20102
rect 9036 20100 9092 20102
rect 9116 20100 9172 20102
rect 9196 20100 9252 20102
rect 8956 19066 9012 19068
rect 9036 19066 9092 19068
rect 9116 19066 9172 19068
rect 9196 19066 9252 19068
rect 8956 19014 8982 19066
rect 8982 19014 9012 19066
rect 9036 19014 9046 19066
rect 9046 19014 9092 19066
rect 9116 19014 9162 19066
rect 9162 19014 9172 19066
rect 9196 19014 9226 19066
rect 9226 19014 9252 19066
rect 8956 19012 9012 19014
rect 9036 19012 9092 19014
rect 9116 19012 9172 19014
rect 9196 19012 9252 19014
rect 8956 17978 9012 17980
rect 9036 17978 9092 17980
rect 9116 17978 9172 17980
rect 9196 17978 9252 17980
rect 8956 17926 8982 17978
rect 8982 17926 9012 17978
rect 9036 17926 9046 17978
rect 9046 17926 9092 17978
rect 9116 17926 9162 17978
rect 9162 17926 9172 17978
rect 9196 17926 9226 17978
rect 9226 17926 9252 17978
rect 8956 17924 9012 17926
rect 9036 17924 9092 17926
rect 9116 17924 9172 17926
rect 9196 17924 9252 17926
rect 9954 18672 10010 18728
rect 8956 16890 9012 16892
rect 9036 16890 9092 16892
rect 9116 16890 9172 16892
rect 9196 16890 9252 16892
rect 8956 16838 8982 16890
rect 8982 16838 9012 16890
rect 9036 16838 9046 16890
rect 9046 16838 9092 16890
rect 9116 16838 9162 16890
rect 9162 16838 9172 16890
rect 9196 16838 9226 16890
rect 9226 16838 9252 16890
rect 8956 16836 9012 16838
rect 9036 16836 9092 16838
rect 9116 16836 9172 16838
rect 9196 16836 9252 16838
rect 8956 15802 9012 15804
rect 9036 15802 9092 15804
rect 9116 15802 9172 15804
rect 9196 15802 9252 15804
rect 8956 15750 8982 15802
rect 8982 15750 9012 15802
rect 9036 15750 9046 15802
rect 9046 15750 9092 15802
rect 9116 15750 9162 15802
rect 9162 15750 9172 15802
rect 9196 15750 9226 15802
rect 9226 15750 9252 15802
rect 8956 15748 9012 15750
rect 9036 15748 9092 15750
rect 9116 15748 9172 15750
rect 9196 15748 9252 15750
rect 8956 14714 9012 14716
rect 9036 14714 9092 14716
rect 9116 14714 9172 14716
rect 9196 14714 9252 14716
rect 8956 14662 8982 14714
rect 8982 14662 9012 14714
rect 9036 14662 9046 14714
rect 9046 14662 9092 14714
rect 9116 14662 9162 14714
rect 9162 14662 9172 14714
rect 9196 14662 9226 14714
rect 9226 14662 9252 14714
rect 8956 14660 9012 14662
rect 9036 14660 9092 14662
rect 9116 14660 9172 14662
rect 9196 14660 9252 14662
rect 10874 18128 10930 18184
rect 8956 13626 9012 13628
rect 9036 13626 9092 13628
rect 9116 13626 9172 13628
rect 9196 13626 9252 13628
rect 8956 13574 8982 13626
rect 8982 13574 9012 13626
rect 9036 13574 9046 13626
rect 9046 13574 9092 13626
rect 9116 13574 9162 13626
rect 9162 13574 9172 13626
rect 9196 13574 9226 13626
rect 9226 13574 9252 13626
rect 8956 13572 9012 13574
rect 9036 13572 9092 13574
rect 9116 13572 9172 13574
rect 9196 13572 9252 13574
rect 9126 12824 9182 12880
rect 9402 13640 9458 13696
rect 8956 12538 9012 12540
rect 9036 12538 9092 12540
rect 9116 12538 9172 12540
rect 9196 12538 9252 12540
rect 8956 12486 8982 12538
rect 8982 12486 9012 12538
rect 9036 12486 9046 12538
rect 9046 12486 9092 12538
rect 9116 12486 9162 12538
rect 9162 12486 9172 12538
rect 9196 12486 9226 12538
rect 9226 12486 9252 12538
rect 8956 12484 9012 12486
rect 9036 12484 9092 12486
rect 9116 12484 9172 12486
rect 9196 12484 9252 12486
rect 12956 21786 13012 21788
rect 13036 21786 13092 21788
rect 13116 21786 13172 21788
rect 13196 21786 13252 21788
rect 12956 21734 12982 21786
rect 12982 21734 13012 21786
rect 13036 21734 13046 21786
rect 13046 21734 13092 21786
rect 13116 21734 13162 21786
rect 13162 21734 13172 21786
rect 13196 21734 13226 21786
rect 13226 21734 13252 21786
rect 12956 21732 13012 21734
rect 13036 21732 13092 21734
rect 13116 21732 13172 21734
rect 13196 21732 13252 21734
rect 12956 20698 13012 20700
rect 13036 20698 13092 20700
rect 13116 20698 13172 20700
rect 13196 20698 13252 20700
rect 12956 20646 12982 20698
rect 12982 20646 13012 20698
rect 13036 20646 13046 20698
rect 13046 20646 13092 20698
rect 13116 20646 13162 20698
rect 13162 20646 13172 20698
rect 13196 20646 13226 20698
rect 13226 20646 13252 20698
rect 12956 20644 13012 20646
rect 13036 20644 13092 20646
rect 13116 20644 13172 20646
rect 13196 20644 13252 20646
rect 12956 19610 13012 19612
rect 13036 19610 13092 19612
rect 13116 19610 13172 19612
rect 13196 19610 13252 19612
rect 12956 19558 12982 19610
rect 12982 19558 13012 19610
rect 13036 19558 13046 19610
rect 13046 19558 13092 19610
rect 13116 19558 13162 19610
rect 13162 19558 13172 19610
rect 13196 19558 13226 19610
rect 13226 19558 13252 19610
rect 12956 19556 13012 19558
rect 13036 19556 13092 19558
rect 13116 19556 13172 19558
rect 13196 19556 13252 19558
rect 8956 11450 9012 11452
rect 9036 11450 9092 11452
rect 9116 11450 9172 11452
rect 9196 11450 9252 11452
rect 8956 11398 8982 11450
rect 8982 11398 9012 11450
rect 9036 11398 9046 11450
rect 9046 11398 9092 11450
rect 9116 11398 9162 11450
rect 9162 11398 9172 11450
rect 9196 11398 9226 11450
rect 9226 11398 9252 11450
rect 8956 11396 9012 11398
rect 9036 11396 9092 11398
rect 9116 11396 9172 11398
rect 9196 11396 9252 11398
rect 8956 10362 9012 10364
rect 9036 10362 9092 10364
rect 9116 10362 9172 10364
rect 9196 10362 9252 10364
rect 8956 10310 8982 10362
rect 8982 10310 9012 10362
rect 9036 10310 9046 10362
rect 9046 10310 9092 10362
rect 9116 10310 9162 10362
rect 9162 10310 9172 10362
rect 9196 10310 9226 10362
rect 9226 10310 9252 10362
rect 8956 10308 9012 10310
rect 9036 10308 9092 10310
rect 9116 10308 9172 10310
rect 9196 10308 9252 10310
rect 8114 9560 8170 9616
rect 8956 9274 9012 9276
rect 9036 9274 9092 9276
rect 9116 9274 9172 9276
rect 9196 9274 9252 9276
rect 8956 9222 8982 9274
rect 8982 9222 9012 9274
rect 9036 9222 9046 9274
rect 9046 9222 9092 9274
rect 9116 9222 9162 9274
rect 9162 9222 9172 9274
rect 9196 9222 9226 9274
rect 9226 9222 9252 9274
rect 8956 9220 9012 9222
rect 9036 9220 9092 9222
rect 9116 9220 9172 9222
rect 9196 9220 9252 9222
rect 8956 8186 9012 8188
rect 9036 8186 9092 8188
rect 9116 8186 9172 8188
rect 9196 8186 9252 8188
rect 8956 8134 8982 8186
rect 8982 8134 9012 8186
rect 9036 8134 9046 8186
rect 9046 8134 9092 8186
rect 9116 8134 9162 8186
rect 9162 8134 9172 8186
rect 9196 8134 9226 8186
rect 9226 8134 9252 8186
rect 8956 8132 9012 8134
rect 9036 8132 9092 8134
rect 9116 8132 9172 8134
rect 9196 8132 9252 8134
rect 5814 5616 5870 5672
rect 7562 5244 7564 5264
rect 7564 5244 7616 5264
rect 7616 5244 7618 5264
rect 7562 5208 7618 5244
rect 6274 3576 6330 3632
rect 8956 7098 9012 7100
rect 9036 7098 9092 7100
rect 9116 7098 9172 7100
rect 9196 7098 9252 7100
rect 8956 7046 8982 7098
rect 8982 7046 9012 7098
rect 9036 7046 9046 7098
rect 9046 7046 9092 7098
rect 9116 7046 9162 7098
rect 9162 7046 9172 7098
rect 9196 7046 9226 7098
rect 9226 7046 9252 7098
rect 8956 7044 9012 7046
rect 9036 7044 9092 7046
rect 9116 7044 9172 7046
rect 9196 7044 9252 7046
rect 7194 2896 7250 2952
rect 7654 2796 7656 2816
rect 7656 2796 7708 2816
rect 7708 2796 7710 2816
rect 7654 2760 7710 2796
rect 8956 6010 9012 6012
rect 9036 6010 9092 6012
rect 9116 6010 9172 6012
rect 9196 6010 9252 6012
rect 8956 5958 8982 6010
rect 8982 5958 9012 6010
rect 9036 5958 9046 6010
rect 9046 5958 9092 6010
rect 9116 5958 9162 6010
rect 9162 5958 9172 6010
rect 9196 5958 9226 6010
rect 9226 5958 9252 6010
rect 8956 5956 9012 5958
rect 9036 5956 9092 5958
rect 9116 5956 9172 5958
rect 9196 5956 9252 5958
rect 8956 4922 9012 4924
rect 9036 4922 9092 4924
rect 9116 4922 9172 4924
rect 9196 4922 9252 4924
rect 8956 4870 8982 4922
rect 8982 4870 9012 4922
rect 9036 4870 9046 4922
rect 9046 4870 9092 4922
rect 9116 4870 9162 4922
rect 9162 4870 9172 4922
rect 9196 4870 9226 4922
rect 9226 4870 9252 4922
rect 8956 4868 9012 4870
rect 9036 4868 9092 4870
rect 9116 4868 9172 4870
rect 9196 4868 9252 4870
rect 8956 3834 9012 3836
rect 9036 3834 9092 3836
rect 9116 3834 9172 3836
rect 9196 3834 9252 3836
rect 8956 3782 8982 3834
rect 8982 3782 9012 3834
rect 9036 3782 9046 3834
rect 9046 3782 9092 3834
rect 9116 3782 9162 3834
rect 9162 3782 9172 3834
rect 9196 3782 9226 3834
rect 9226 3782 9252 3834
rect 8956 3780 9012 3782
rect 9036 3780 9092 3782
rect 9116 3780 9172 3782
rect 9196 3780 9252 3782
rect 9954 5752 10010 5808
rect 16956 21242 17012 21244
rect 17036 21242 17092 21244
rect 17116 21242 17172 21244
rect 17196 21242 17252 21244
rect 16956 21190 16982 21242
rect 16982 21190 17012 21242
rect 17036 21190 17046 21242
rect 17046 21190 17092 21242
rect 17116 21190 17162 21242
rect 17162 21190 17172 21242
rect 17196 21190 17226 21242
rect 17226 21190 17252 21242
rect 16956 21188 17012 21190
rect 17036 21188 17092 21190
rect 17116 21188 17172 21190
rect 17196 21188 17252 21190
rect 16956 20154 17012 20156
rect 17036 20154 17092 20156
rect 17116 20154 17172 20156
rect 17196 20154 17252 20156
rect 16956 20102 16982 20154
rect 16982 20102 17012 20154
rect 17036 20102 17046 20154
rect 17046 20102 17092 20154
rect 17116 20102 17162 20154
rect 17162 20102 17172 20154
rect 17196 20102 17226 20154
rect 17226 20102 17252 20154
rect 16956 20100 17012 20102
rect 17036 20100 17092 20102
rect 17116 20100 17172 20102
rect 17196 20100 17252 20102
rect 12956 18522 13012 18524
rect 13036 18522 13092 18524
rect 13116 18522 13172 18524
rect 13196 18522 13252 18524
rect 12956 18470 12982 18522
rect 12982 18470 13012 18522
rect 13036 18470 13046 18522
rect 13046 18470 13092 18522
rect 13116 18470 13162 18522
rect 13162 18470 13172 18522
rect 13196 18470 13226 18522
rect 13226 18470 13252 18522
rect 12956 18468 13012 18470
rect 13036 18468 13092 18470
rect 13116 18468 13172 18470
rect 13196 18468 13252 18470
rect 12956 17434 13012 17436
rect 13036 17434 13092 17436
rect 13116 17434 13172 17436
rect 13196 17434 13252 17436
rect 12956 17382 12982 17434
rect 12982 17382 13012 17434
rect 13036 17382 13046 17434
rect 13046 17382 13092 17434
rect 13116 17382 13162 17434
rect 13162 17382 13172 17434
rect 13196 17382 13226 17434
rect 13226 17382 13252 17434
rect 12956 17380 13012 17382
rect 13036 17380 13092 17382
rect 13116 17380 13172 17382
rect 13196 17380 13252 17382
rect 10966 11736 11022 11792
rect 9954 4256 10010 4312
rect 9770 3984 9826 4040
rect 9678 3712 9734 3768
rect 9310 3032 9366 3088
rect 8956 2746 9012 2748
rect 9036 2746 9092 2748
rect 9116 2746 9172 2748
rect 9196 2746 9252 2748
rect 8956 2694 8982 2746
rect 8982 2694 9012 2746
rect 9036 2694 9046 2746
rect 9046 2694 9092 2746
rect 9116 2694 9162 2746
rect 9162 2694 9172 2746
rect 9196 2694 9226 2746
rect 9226 2694 9252 2746
rect 8956 2692 9012 2694
rect 9036 2692 9092 2694
rect 9116 2692 9172 2694
rect 9196 2692 9252 2694
rect 8942 1944 8998 2000
rect 7654 584 7710 640
rect 12956 16346 13012 16348
rect 13036 16346 13092 16348
rect 13116 16346 13172 16348
rect 13196 16346 13252 16348
rect 12956 16294 12982 16346
rect 12982 16294 13012 16346
rect 13036 16294 13046 16346
rect 13046 16294 13092 16346
rect 13116 16294 13162 16346
rect 13162 16294 13172 16346
rect 13196 16294 13226 16346
rect 13226 16294 13252 16346
rect 12956 16292 13012 16294
rect 13036 16292 13092 16294
rect 13116 16292 13172 16294
rect 13196 16292 13252 16294
rect 12956 15258 13012 15260
rect 13036 15258 13092 15260
rect 13116 15258 13172 15260
rect 13196 15258 13252 15260
rect 12956 15206 12982 15258
rect 12982 15206 13012 15258
rect 13036 15206 13046 15258
rect 13046 15206 13092 15258
rect 13116 15206 13162 15258
rect 13162 15206 13172 15258
rect 13196 15206 13226 15258
rect 13226 15206 13252 15258
rect 12956 15204 13012 15206
rect 13036 15204 13092 15206
rect 13116 15204 13172 15206
rect 13196 15204 13252 15206
rect 12956 14170 13012 14172
rect 13036 14170 13092 14172
rect 13116 14170 13172 14172
rect 13196 14170 13252 14172
rect 12956 14118 12982 14170
rect 12982 14118 13012 14170
rect 13036 14118 13046 14170
rect 13046 14118 13092 14170
rect 13116 14118 13162 14170
rect 13162 14118 13172 14170
rect 13196 14118 13226 14170
rect 13226 14118 13252 14170
rect 12956 14116 13012 14118
rect 13036 14116 13092 14118
rect 13116 14116 13172 14118
rect 13196 14116 13252 14118
rect 12806 13640 12862 13696
rect 12956 13082 13012 13084
rect 13036 13082 13092 13084
rect 13116 13082 13172 13084
rect 13196 13082 13252 13084
rect 12956 13030 12982 13082
rect 12982 13030 13012 13082
rect 13036 13030 13046 13082
rect 13046 13030 13092 13082
rect 13116 13030 13162 13082
rect 13162 13030 13172 13082
rect 13196 13030 13226 13082
rect 13226 13030 13252 13082
rect 12956 13028 13012 13030
rect 13036 13028 13092 13030
rect 13116 13028 13172 13030
rect 13196 13028 13252 13030
rect 12956 11994 13012 11996
rect 13036 11994 13092 11996
rect 13116 11994 13172 11996
rect 13196 11994 13252 11996
rect 12956 11942 12982 11994
rect 12982 11942 13012 11994
rect 13036 11942 13046 11994
rect 13046 11942 13092 11994
rect 13116 11942 13162 11994
rect 13162 11942 13172 11994
rect 13196 11942 13226 11994
rect 13226 11942 13252 11994
rect 12956 11940 13012 11942
rect 13036 11940 13092 11942
rect 13116 11940 13172 11942
rect 13196 11940 13252 11942
rect 12956 10906 13012 10908
rect 13036 10906 13092 10908
rect 13116 10906 13172 10908
rect 13196 10906 13252 10908
rect 12956 10854 12982 10906
rect 12982 10854 13012 10906
rect 13036 10854 13046 10906
rect 13046 10854 13092 10906
rect 13116 10854 13162 10906
rect 13162 10854 13172 10906
rect 13196 10854 13226 10906
rect 13226 10854 13252 10906
rect 12956 10852 13012 10854
rect 13036 10852 13092 10854
rect 13116 10852 13172 10854
rect 13196 10852 13252 10854
rect 11058 3712 11114 3768
rect 11518 4120 11574 4176
rect 12956 9818 13012 9820
rect 13036 9818 13092 9820
rect 13116 9818 13172 9820
rect 13196 9818 13252 9820
rect 12956 9766 12982 9818
rect 12982 9766 13012 9818
rect 13036 9766 13046 9818
rect 13046 9766 13092 9818
rect 13116 9766 13162 9818
rect 13162 9766 13172 9818
rect 13196 9766 13226 9818
rect 13226 9766 13252 9818
rect 12956 9764 13012 9766
rect 13036 9764 13092 9766
rect 13116 9764 13172 9766
rect 13196 9764 13252 9766
rect 12956 8730 13012 8732
rect 13036 8730 13092 8732
rect 13116 8730 13172 8732
rect 13196 8730 13252 8732
rect 12956 8678 12982 8730
rect 12982 8678 13012 8730
rect 13036 8678 13046 8730
rect 13046 8678 13092 8730
rect 13116 8678 13162 8730
rect 13162 8678 13172 8730
rect 13196 8678 13226 8730
rect 13226 8678 13252 8730
rect 12956 8676 13012 8678
rect 13036 8676 13092 8678
rect 13116 8676 13172 8678
rect 13196 8676 13252 8678
rect 13266 8472 13322 8528
rect 11702 2896 11758 2952
rect 12956 7642 13012 7644
rect 13036 7642 13092 7644
rect 13116 7642 13172 7644
rect 13196 7642 13252 7644
rect 12956 7590 12982 7642
rect 12982 7590 13012 7642
rect 13036 7590 13046 7642
rect 13046 7590 13092 7642
rect 13116 7590 13162 7642
rect 13162 7590 13172 7642
rect 13196 7590 13226 7642
rect 13226 7590 13252 7642
rect 12956 7588 13012 7590
rect 13036 7588 13092 7590
rect 13116 7588 13172 7590
rect 13196 7588 13252 7590
rect 12956 6554 13012 6556
rect 13036 6554 13092 6556
rect 13116 6554 13172 6556
rect 13196 6554 13252 6556
rect 12956 6502 12982 6554
rect 12982 6502 13012 6554
rect 13036 6502 13046 6554
rect 13046 6502 13092 6554
rect 13116 6502 13162 6554
rect 13162 6502 13172 6554
rect 13196 6502 13226 6554
rect 13226 6502 13252 6554
rect 12956 6500 13012 6502
rect 13036 6500 13092 6502
rect 13116 6500 13172 6502
rect 13196 6500 13252 6502
rect 12254 5072 12310 5128
rect 12162 2352 12218 2408
rect 12956 5466 13012 5468
rect 13036 5466 13092 5468
rect 13116 5466 13172 5468
rect 13196 5466 13252 5468
rect 12956 5414 12982 5466
rect 12982 5414 13012 5466
rect 13036 5414 13046 5466
rect 13046 5414 13092 5466
rect 13116 5414 13162 5466
rect 13162 5414 13172 5466
rect 13196 5414 13226 5466
rect 13226 5414 13252 5466
rect 12956 5412 13012 5414
rect 13036 5412 13092 5414
rect 13116 5412 13172 5414
rect 13196 5412 13252 5414
rect 12956 4378 13012 4380
rect 13036 4378 13092 4380
rect 13116 4378 13172 4380
rect 13196 4378 13252 4380
rect 12956 4326 12982 4378
rect 12982 4326 13012 4378
rect 13036 4326 13046 4378
rect 13046 4326 13092 4378
rect 13116 4326 13162 4378
rect 13162 4326 13172 4378
rect 13196 4326 13226 4378
rect 13226 4326 13252 4378
rect 12956 4324 13012 4326
rect 13036 4324 13092 4326
rect 13116 4324 13172 4326
rect 13196 4324 13252 4326
rect 12438 3576 12494 3632
rect 12956 3290 13012 3292
rect 13036 3290 13092 3292
rect 13116 3290 13172 3292
rect 13196 3290 13252 3292
rect 12956 3238 12982 3290
rect 12982 3238 13012 3290
rect 13036 3238 13046 3290
rect 13046 3238 13092 3290
rect 13116 3238 13162 3290
rect 13162 3238 13172 3290
rect 13196 3238 13226 3290
rect 13226 3238 13252 3290
rect 12956 3236 13012 3238
rect 13036 3236 13092 3238
rect 13116 3236 13172 3238
rect 13196 3236 13252 3238
rect 12438 2352 12494 2408
rect 12956 2202 13012 2204
rect 13036 2202 13092 2204
rect 13116 2202 13172 2204
rect 13196 2202 13252 2204
rect 12956 2150 12982 2202
rect 12982 2150 13012 2202
rect 13036 2150 13046 2202
rect 13046 2150 13092 2202
rect 13116 2150 13162 2202
rect 13162 2150 13172 2202
rect 13196 2150 13226 2202
rect 13226 2150 13252 2202
rect 12956 2148 13012 2150
rect 13036 2148 13092 2150
rect 13116 2148 13172 2150
rect 13196 2148 13252 2150
rect 16302 19216 16358 19272
rect 16956 19066 17012 19068
rect 17036 19066 17092 19068
rect 17116 19066 17172 19068
rect 17196 19066 17252 19068
rect 16956 19014 16982 19066
rect 16982 19014 17012 19066
rect 17036 19014 17046 19066
rect 17046 19014 17092 19066
rect 17116 19014 17162 19066
rect 17162 19014 17172 19066
rect 17196 19014 17226 19066
rect 17226 19014 17252 19066
rect 16956 19012 17012 19014
rect 17036 19012 17092 19014
rect 17116 19012 17172 19014
rect 17196 19012 17252 19014
rect 14830 8472 14886 8528
rect 14554 7248 14610 7304
rect 14094 3712 14150 3768
rect 14278 2488 14334 2544
rect 17406 18128 17462 18184
rect 16956 17978 17012 17980
rect 17036 17978 17092 17980
rect 17116 17978 17172 17980
rect 17196 17978 17252 17980
rect 16956 17926 16982 17978
rect 16982 17926 17012 17978
rect 17036 17926 17046 17978
rect 17046 17926 17092 17978
rect 17116 17926 17162 17978
rect 17162 17926 17172 17978
rect 17196 17926 17226 17978
rect 17226 17926 17252 17978
rect 16956 17924 17012 17926
rect 17036 17924 17092 17926
rect 17116 17924 17172 17926
rect 17196 17924 17252 17926
rect 16956 16890 17012 16892
rect 17036 16890 17092 16892
rect 17116 16890 17172 16892
rect 17196 16890 17252 16892
rect 16956 16838 16982 16890
rect 16982 16838 17012 16890
rect 17036 16838 17046 16890
rect 17046 16838 17092 16890
rect 17116 16838 17162 16890
rect 17162 16838 17172 16890
rect 17196 16838 17226 16890
rect 17226 16838 17252 16890
rect 16956 16836 17012 16838
rect 17036 16836 17092 16838
rect 17116 16836 17172 16838
rect 17196 16836 17252 16838
rect 16956 15802 17012 15804
rect 17036 15802 17092 15804
rect 17116 15802 17172 15804
rect 17196 15802 17252 15804
rect 16956 15750 16982 15802
rect 16982 15750 17012 15802
rect 17036 15750 17046 15802
rect 17046 15750 17092 15802
rect 17116 15750 17162 15802
rect 17162 15750 17172 15802
rect 17196 15750 17226 15802
rect 17226 15750 17252 15802
rect 16956 15748 17012 15750
rect 17036 15748 17092 15750
rect 17116 15748 17172 15750
rect 17196 15748 17252 15750
rect 16956 14714 17012 14716
rect 17036 14714 17092 14716
rect 17116 14714 17172 14716
rect 17196 14714 17252 14716
rect 16956 14662 16982 14714
rect 16982 14662 17012 14714
rect 17036 14662 17046 14714
rect 17046 14662 17092 14714
rect 17116 14662 17162 14714
rect 17162 14662 17172 14714
rect 17196 14662 17226 14714
rect 17226 14662 17252 14714
rect 16956 14660 17012 14662
rect 17036 14660 17092 14662
rect 17116 14660 17172 14662
rect 17196 14660 17252 14662
rect 16956 13626 17012 13628
rect 17036 13626 17092 13628
rect 17116 13626 17172 13628
rect 17196 13626 17252 13628
rect 16956 13574 16982 13626
rect 16982 13574 17012 13626
rect 17036 13574 17046 13626
rect 17046 13574 17092 13626
rect 17116 13574 17162 13626
rect 17162 13574 17172 13626
rect 17196 13574 17226 13626
rect 17226 13574 17252 13626
rect 16956 13572 17012 13574
rect 17036 13572 17092 13574
rect 17116 13572 17172 13574
rect 17196 13572 17252 13574
rect 16956 12538 17012 12540
rect 17036 12538 17092 12540
rect 17116 12538 17172 12540
rect 17196 12538 17252 12540
rect 16956 12486 16982 12538
rect 16982 12486 17012 12538
rect 17036 12486 17046 12538
rect 17046 12486 17092 12538
rect 17116 12486 17162 12538
rect 17162 12486 17172 12538
rect 17196 12486 17226 12538
rect 17226 12486 17252 12538
rect 16956 12484 17012 12486
rect 17036 12484 17092 12486
rect 17116 12484 17172 12486
rect 17196 12484 17252 12486
rect 16956 11450 17012 11452
rect 17036 11450 17092 11452
rect 17116 11450 17172 11452
rect 17196 11450 17252 11452
rect 16956 11398 16982 11450
rect 16982 11398 17012 11450
rect 17036 11398 17046 11450
rect 17046 11398 17092 11450
rect 17116 11398 17162 11450
rect 17162 11398 17172 11450
rect 17196 11398 17226 11450
rect 17226 11398 17252 11450
rect 16956 11396 17012 11398
rect 17036 11396 17092 11398
rect 17116 11396 17172 11398
rect 17196 11396 17252 11398
rect 20956 21786 21012 21788
rect 21036 21786 21092 21788
rect 21116 21786 21172 21788
rect 21196 21786 21252 21788
rect 20956 21734 20982 21786
rect 20982 21734 21012 21786
rect 21036 21734 21046 21786
rect 21046 21734 21092 21786
rect 21116 21734 21162 21786
rect 21162 21734 21172 21786
rect 21196 21734 21226 21786
rect 21226 21734 21252 21786
rect 20956 21732 21012 21734
rect 21036 21732 21092 21734
rect 21116 21732 21172 21734
rect 21196 21732 21252 21734
rect 21454 21392 21510 21448
rect 20956 20698 21012 20700
rect 21036 20698 21092 20700
rect 21116 20698 21172 20700
rect 21196 20698 21252 20700
rect 20956 20646 20982 20698
rect 20982 20646 21012 20698
rect 21036 20646 21046 20698
rect 21046 20646 21092 20698
rect 21116 20646 21162 20698
rect 21162 20646 21172 20698
rect 21196 20646 21226 20698
rect 21226 20646 21252 20698
rect 20956 20644 21012 20646
rect 21036 20644 21092 20646
rect 21116 20644 21172 20646
rect 21196 20644 21252 20646
rect 21178 20168 21234 20224
rect 20956 19610 21012 19612
rect 21036 19610 21092 19612
rect 21116 19610 21172 19612
rect 21196 19610 21252 19612
rect 20956 19558 20982 19610
rect 20982 19558 21012 19610
rect 21036 19558 21046 19610
rect 21046 19558 21092 19610
rect 21116 19558 21162 19610
rect 21162 19558 21172 19610
rect 21196 19558 21226 19610
rect 21226 19558 21252 19610
rect 20956 19556 21012 19558
rect 21036 19556 21092 19558
rect 21116 19556 21172 19558
rect 21196 19556 21252 19558
rect 18970 18808 19026 18864
rect 20626 18808 20682 18864
rect 18694 18672 18750 18728
rect 16956 10362 17012 10364
rect 17036 10362 17092 10364
rect 17116 10362 17172 10364
rect 17196 10362 17252 10364
rect 16956 10310 16982 10362
rect 16982 10310 17012 10362
rect 17036 10310 17046 10362
rect 17046 10310 17092 10362
rect 17116 10310 17162 10362
rect 17162 10310 17172 10362
rect 17196 10310 17226 10362
rect 17226 10310 17252 10362
rect 16956 10308 17012 10310
rect 17036 10308 17092 10310
rect 17116 10308 17172 10310
rect 17196 10308 17252 10310
rect 16956 9274 17012 9276
rect 17036 9274 17092 9276
rect 17116 9274 17172 9276
rect 17196 9274 17252 9276
rect 16956 9222 16982 9274
rect 16982 9222 17012 9274
rect 17036 9222 17046 9274
rect 17046 9222 17092 9274
rect 17116 9222 17162 9274
rect 17162 9222 17172 9274
rect 17196 9222 17226 9274
rect 17226 9222 17252 9274
rect 16956 9220 17012 9222
rect 17036 9220 17092 9222
rect 17116 9220 17172 9222
rect 17196 9220 17252 9222
rect 16956 8186 17012 8188
rect 17036 8186 17092 8188
rect 17116 8186 17172 8188
rect 17196 8186 17252 8188
rect 16956 8134 16982 8186
rect 16982 8134 17012 8186
rect 17036 8134 17046 8186
rect 17046 8134 17092 8186
rect 17116 8134 17162 8186
rect 17162 8134 17172 8186
rect 17196 8134 17226 8186
rect 17226 8134 17252 8186
rect 16956 8132 17012 8134
rect 17036 8132 17092 8134
rect 17116 8132 17172 8134
rect 17196 8132 17252 8134
rect 15658 5344 15714 5400
rect 16956 7098 17012 7100
rect 17036 7098 17092 7100
rect 17116 7098 17172 7100
rect 17196 7098 17252 7100
rect 16956 7046 16982 7098
rect 16982 7046 17012 7098
rect 17036 7046 17046 7098
rect 17046 7046 17092 7098
rect 17116 7046 17162 7098
rect 17162 7046 17172 7098
rect 17196 7046 17226 7098
rect 17226 7046 17252 7098
rect 16956 7044 17012 7046
rect 17036 7044 17092 7046
rect 17116 7044 17172 7046
rect 17196 7044 17252 7046
rect 15474 1944 15530 2000
rect 16956 6010 17012 6012
rect 17036 6010 17092 6012
rect 17116 6010 17172 6012
rect 17196 6010 17252 6012
rect 16956 5958 16982 6010
rect 16982 5958 17012 6010
rect 17036 5958 17046 6010
rect 17046 5958 17092 6010
rect 17116 5958 17162 6010
rect 17162 5958 17172 6010
rect 17196 5958 17226 6010
rect 17226 5958 17252 6010
rect 16956 5956 17012 5958
rect 17036 5956 17092 5958
rect 17116 5956 17172 5958
rect 17196 5956 17252 5958
rect 16956 4922 17012 4924
rect 17036 4922 17092 4924
rect 17116 4922 17172 4924
rect 17196 4922 17252 4924
rect 16956 4870 16982 4922
rect 16982 4870 17012 4922
rect 17036 4870 17046 4922
rect 17046 4870 17092 4922
rect 17116 4870 17162 4922
rect 17162 4870 17172 4922
rect 17196 4870 17226 4922
rect 17226 4870 17252 4922
rect 16956 4868 17012 4870
rect 17036 4868 17092 4870
rect 17116 4868 17172 4870
rect 17196 4868 17252 4870
rect 18418 8880 18474 8936
rect 16956 3834 17012 3836
rect 17036 3834 17092 3836
rect 17116 3834 17172 3836
rect 17196 3834 17252 3836
rect 16956 3782 16982 3834
rect 16982 3782 17012 3834
rect 17036 3782 17046 3834
rect 17046 3782 17092 3834
rect 17116 3782 17162 3834
rect 17162 3782 17172 3834
rect 17196 3782 17226 3834
rect 17226 3782 17252 3834
rect 16956 3780 17012 3782
rect 17036 3780 17092 3782
rect 17116 3780 17172 3782
rect 17196 3780 17252 3782
rect 16956 2746 17012 2748
rect 17036 2746 17092 2748
rect 17116 2746 17172 2748
rect 17196 2746 17252 2748
rect 16956 2694 16982 2746
rect 16982 2694 17012 2746
rect 17036 2694 17046 2746
rect 17046 2694 17092 2746
rect 17116 2694 17162 2746
rect 17162 2694 17172 2746
rect 17196 2694 17226 2746
rect 17226 2694 17252 2746
rect 16956 2692 17012 2694
rect 17036 2692 17092 2694
rect 17116 2692 17172 2694
rect 17196 2692 17252 2694
rect 17406 3032 17462 3088
rect 18326 5208 18382 5264
rect 19338 2896 19394 2952
rect 20956 18522 21012 18524
rect 21036 18522 21092 18524
rect 21116 18522 21172 18524
rect 21196 18522 21252 18524
rect 20956 18470 20982 18522
rect 20982 18470 21012 18522
rect 21036 18470 21046 18522
rect 21046 18470 21092 18522
rect 21116 18470 21162 18522
rect 21162 18470 21172 18522
rect 21196 18470 21226 18522
rect 21226 18470 21252 18522
rect 20956 18468 21012 18470
rect 21036 18468 21092 18470
rect 21116 18468 21172 18470
rect 21196 18468 21252 18470
rect 20810 18264 20866 18320
rect 21270 17584 21326 17640
rect 20956 17434 21012 17436
rect 21036 17434 21092 17436
rect 21116 17434 21172 17436
rect 21196 17434 21252 17436
rect 20956 17382 20982 17434
rect 20982 17382 21012 17434
rect 21036 17382 21046 17434
rect 21046 17382 21092 17434
rect 21116 17382 21162 17434
rect 21162 17382 21172 17434
rect 21196 17382 21226 17434
rect 21226 17382 21252 17434
rect 20956 17380 21012 17382
rect 21036 17380 21092 17382
rect 21116 17380 21172 17382
rect 21196 17380 21252 17382
rect 21454 16360 21510 16416
rect 20956 16346 21012 16348
rect 21036 16346 21092 16348
rect 21116 16346 21172 16348
rect 21196 16346 21252 16348
rect 20956 16294 20982 16346
rect 20982 16294 21012 16346
rect 21036 16294 21046 16346
rect 21046 16294 21092 16346
rect 21116 16294 21162 16346
rect 21162 16294 21172 16346
rect 21196 16294 21226 16346
rect 21226 16294 21252 16346
rect 20956 16292 21012 16294
rect 21036 16292 21092 16294
rect 21116 16292 21172 16294
rect 21196 16292 21252 16294
rect 21270 15408 21326 15464
rect 20956 15258 21012 15260
rect 21036 15258 21092 15260
rect 21116 15258 21172 15260
rect 21196 15258 21252 15260
rect 20956 15206 20982 15258
rect 20982 15206 21012 15258
rect 21036 15206 21046 15258
rect 21046 15206 21092 15258
rect 21116 15206 21162 15258
rect 21162 15206 21172 15258
rect 21196 15206 21226 15258
rect 21226 15206 21252 15258
rect 20956 15204 21012 15206
rect 21036 15204 21092 15206
rect 21116 15204 21172 15206
rect 21196 15204 21252 15206
rect 20956 14170 21012 14172
rect 21036 14170 21092 14172
rect 21116 14170 21172 14172
rect 21196 14170 21252 14172
rect 20956 14118 20982 14170
rect 20982 14118 21012 14170
rect 21036 14118 21046 14170
rect 21046 14118 21092 14170
rect 21116 14118 21162 14170
rect 21162 14118 21172 14170
rect 21196 14118 21226 14170
rect 21226 14118 21252 14170
rect 20956 14116 21012 14118
rect 21036 14116 21092 14118
rect 21116 14116 21172 14118
rect 21196 14116 21252 14118
rect 21086 13912 21142 13968
rect 20956 13082 21012 13084
rect 21036 13082 21092 13084
rect 21116 13082 21172 13084
rect 21196 13082 21252 13084
rect 20956 13030 20982 13082
rect 20982 13030 21012 13082
rect 21036 13030 21046 13082
rect 21046 13030 21092 13082
rect 21116 13030 21162 13082
rect 21162 13030 21172 13082
rect 21196 13030 21226 13082
rect 21226 13030 21252 13082
rect 20956 13028 21012 13030
rect 21036 13028 21092 13030
rect 21116 13028 21172 13030
rect 21196 13028 21252 13030
rect 20956 11994 21012 11996
rect 21036 11994 21092 11996
rect 21116 11994 21172 11996
rect 21196 11994 21252 11996
rect 20956 11942 20982 11994
rect 20982 11942 21012 11994
rect 21036 11942 21046 11994
rect 21046 11942 21092 11994
rect 21116 11942 21162 11994
rect 21162 11942 21172 11994
rect 21196 11942 21226 11994
rect 21226 11942 21252 11994
rect 20956 11940 21012 11942
rect 21036 11940 21092 11942
rect 21116 11940 21172 11942
rect 21196 11940 21252 11942
rect 20718 11600 20774 11656
rect 22466 22616 22522 22672
rect 23570 11872 23626 11928
rect 20956 10906 21012 10908
rect 21036 10906 21092 10908
rect 21116 10906 21172 10908
rect 21196 10906 21252 10908
rect 20956 10854 20982 10906
rect 20982 10854 21012 10906
rect 21036 10854 21046 10906
rect 21046 10854 21092 10906
rect 21116 10854 21162 10906
rect 21162 10854 21172 10906
rect 21196 10854 21226 10906
rect 21226 10854 21252 10906
rect 20956 10852 21012 10854
rect 21036 10852 21092 10854
rect 21116 10852 21172 10854
rect 21196 10852 21252 10854
rect 21086 10240 21142 10296
rect 20956 9818 21012 9820
rect 21036 9818 21092 9820
rect 21116 9818 21172 9820
rect 21196 9818 21252 9820
rect 20956 9766 20982 9818
rect 20982 9766 21012 9818
rect 21036 9766 21046 9818
rect 21046 9766 21092 9818
rect 21116 9766 21162 9818
rect 21162 9766 21172 9818
rect 21196 9766 21226 9818
rect 21226 9766 21252 9818
rect 20956 9764 21012 9766
rect 21036 9764 21092 9766
rect 21116 9764 21172 9766
rect 21196 9764 21252 9766
rect 20810 9560 20866 9616
rect 20956 8730 21012 8732
rect 21036 8730 21092 8732
rect 21116 8730 21172 8732
rect 21196 8730 21252 8732
rect 20956 8678 20982 8730
rect 20982 8678 21012 8730
rect 21036 8678 21046 8730
rect 21046 8678 21092 8730
rect 21116 8678 21162 8730
rect 21162 8678 21172 8730
rect 21196 8678 21226 8730
rect 21226 8678 21252 8730
rect 20956 8676 21012 8678
rect 21036 8676 21092 8678
rect 21116 8676 21172 8678
rect 21196 8676 21252 8678
rect 20956 7642 21012 7644
rect 21036 7642 21092 7644
rect 21116 7642 21172 7644
rect 21196 7642 21252 7644
rect 20956 7590 20982 7642
rect 20982 7590 21012 7642
rect 21036 7590 21046 7642
rect 21046 7590 21092 7642
rect 21116 7590 21162 7642
rect 21162 7590 21172 7642
rect 21196 7590 21226 7642
rect 21226 7590 21252 7642
rect 20956 7588 21012 7590
rect 21036 7588 21092 7590
rect 21116 7588 21172 7590
rect 21196 7588 21252 7590
rect 21362 7520 21418 7576
rect 20956 6554 21012 6556
rect 21036 6554 21092 6556
rect 21116 6554 21172 6556
rect 21196 6554 21252 6556
rect 20956 6502 20982 6554
rect 20982 6502 21012 6554
rect 21036 6502 21046 6554
rect 21046 6502 21092 6554
rect 21116 6502 21162 6554
rect 21162 6502 21172 6554
rect 21196 6502 21226 6554
rect 21226 6502 21252 6554
rect 20956 6500 21012 6502
rect 21036 6500 21092 6502
rect 21116 6500 21172 6502
rect 21196 6500 21252 6502
rect 21454 5752 21510 5808
rect 20956 5466 21012 5468
rect 21036 5466 21092 5468
rect 21116 5466 21172 5468
rect 21196 5466 21252 5468
rect 20956 5414 20982 5466
rect 20982 5414 21012 5466
rect 21036 5414 21046 5466
rect 21046 5414 21092 5466
rect 21116 5414 21162 5466
rect 21162 5414 21172 5466
rect 21196 5414 21226 5466
rect 21226 5414 21252 5466
rect 20956 5412 21012 5414
rect 21036 5412 21092 5414
rect 21116 5412 21172 5414
rect 21196 5412 21252 5414
rect 20718 5344 20774 5400
rect 20626 5072 20682 5128
rect 20626 4256 20682 4312
rect 20626 3576 20682 3632
rect 21454 4800 21510 4856
rect 20956 4378 21012 4380
rect 21036 4378 21092 4380
rect 21116 4378 21172 4380
rect 21196 4378 21252 4380
rect 20956 4326 20982 4378
rect 20982 4326 21012 4378
rect 21036 4326 21046 4378
rect 21046 4326 21092 4378
rect 21116 4326 21162 4378
rect 21162 4326 21172 4378
rect 21196 4326 21226 4378
rect 21226 4326 21252 4378
rect 20956 4324 21012 4326
rect 21036 4324 21092 4326
rect 21116 4324 21172 4326
rect 21196 4324 21252 4326
rect 20956 3290 21012 3292
rect 21036 3290 21092 3292
rect 21116 3290 21172 3292
rect 21196 3290 21252 3292
rect 20956 3238 20982 3290
rect 20982 3238 21012 3290
rect 21036 3238 21046 3290
rect 21046 3238 21092 3290
rect 21116 3238 21162 3290
rect 21162 3238 21172 3290
rect 21196 3238 21226 3290
rect 21226 3238 21252 3290
rect 20956 3236 21012 3238
rect 21036 3236 21092 3238
rect 21116 3236 21172 3238
rect 21196 3236 21252 3238
rect 20956 2202 21012 2204
rect 21036 2202 21092 2204
rect 21116 2202 21172 2204
rect 21196 2202 21252 2204
rect 20956 2150 20982 2202
rect 20982 2150 21012 2202
rect 21036 2150 21046 2202
rect 21046 2150 21092 2202
rect 21116 2150 21162 2202
rect 21162 2150 21172 2202
rect 21196 2150 21226 2202
rect 21226 2150 21252 2202
rect 20956 2148 21012 2150
rect 21036 2148 21092 2150
rect 21116 2148 21172 2150
rect 21196 2148 21252 2150
rect 23570 6840 23626 6896
rect 23386 5616 23442 5672
<< metal3 >>
rect 0 23128 480 23248
rect 23520 23128 24000 23248
rect 62 22674 122 23128
rect 1577 22674 1643 22677
rect 62 22672 1643 22674
rect 62 22616 1582 22672
rect 1638 22616 1643 22672
rect 62 22614 1643 22616
rect 1577 22611 1643 22614
rect 22461 22674 22527 22677
rect 23614 22674 23674 23128
rect 22461 22672 23674 22674
rect 22461 22616 22466 22672
rect 22522 22616 23674 22672
rect 22461 22614 23674 22616
rect 22461 22611 22527 22614
rect 23520 21904 24000 22024
rect 0 21768 480 21888
rect 4944 21792 5264 21793
rect 62 21314 122 21768
rect 4944 21728 4952 21792
rect 5016 21728 5032 21792
rect 5096 21728 5112 21792
rect 5176 21728 5192 21792
rect 5256 21728 5264 21792
rect 4944 21727 5264 21728
rect 12944 21792 13264 21793
rect 12944 21728 12952 21792
rect 13016 21728 13032 21792
rect 13096 21728 13112 21792
rect 13176 21728 13192 21792
rect 13256 21728 13264 21792
rect 12944 21727 13264 21728
rect 20944 21792 21264 21793
rect 20944 21728 20952 21792
rect 21016 21728 21032 21792
rect 21096 21728 21112 21792
rect 21176 21728 21192 21792
rect 21256 21728 21264 21792
rect 20944 21727 21264 21728
rect 21449 21450 21515 21453
rect 23614 21450 23674 21904
rect 21449 21448 23674 21450
rect 21449 21392 21454 21448
rect 21510 21392 23674 21448
rect 21449 21390 23674 21392
rect 21449 21387 21515 21390
rect 1853 21314 1919 21317
rect 62 21312 1919 21314
rect 62 21256 1858 21312
rect 1914 21256 1919 21312
rect 62 21254 1919 21256
rect 1853 21251 1919 21254
rect 8944 21248 9264 21249
rect 8944 21184 8952 21248
rect 9016 21184 9032 21248
rect 9096 21184 9112 21248
rect 9176 21184 9192 21248
rect 9256 21184 9264 21248
rect 8944 21183 9264 21184
rect 16944 21248 17264 21249
rect 16944 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17264 21248
rect 16944 21183 17264 21184
rect 4944 20704 5264 20705
rect 4944 20640 4952 20704
rect 5016 20640 5032 20704
rect 5096 20640 5112 20704
rect 5176 20640 5192 20704
rect 5256 20640 5264 20704
rect 4944 20639 5264 20640
rect 12944 20704 13264 20705
rect 12944 20640 12952 20704
rect 13016 20640 13032 20704
rect 13096 20640 13112 20704
rect 13176 20640 13192 20704
rect 13256 20640 13264 20704
rect 12944 20639 13264 20640
rect 20944 20704 21264 20705
rect 20944 20640 20952 20704
rect 21016 20640 21032 20704
rect 21096 20640 21112 20704
rect 21176 20640 21192 20704
rect 21256 20640 21264 20704
rect 23520 20680 24000 20800
rect 20944 20639 21264 20640
rect 0 20360 480 20392
rect 0 20304 110 20360
rect 166 20304 480 20360
rect 0 20272 480 20304
rect 21173 20226 21239 20229
rect 23614 20226 23674 20680
rect 21173 20224 23674 20226
rect 21173 20168 21178 20224
rect 21234 20168 23674 20224
rect 21173 20166 23674 20168
rect 21173 20163 21239 20166
rect 8944 20160 9264 20161
rect 8944 20096 8952 20160
rect 9016 20096 9032 20160
rect 9096 20096 9112 20160
rect 9176 20096 9192 20160
rect 9256 20096 9264 20160
rect 8944 20095 9264 20096
rect 16944 20160 17264 20161
rect 16944 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17264 20160
rect 16944 20095 17264 20096
rect 4944 19616 5264 19617
rect 4944 19552 4952 19616
rect 5016 19552 5032 19616
rect 5096 19552 5112 19616
rect 5176 19552 5192 19616
rect 5256 19552 5264 19616
rect 4944 19551 5264 19552
rect 12944 19616 13264 19617
rect 12944 19552 12952 19616
rect 13016 19552 13032 19616
rect 13096 19552 13112 19616
rect 13176 19552 13192 19616
rect 13256 19552 13264 19616
rect 12944 19551 13264 19552
rect 20944 19616 21264 19617
rect 20944 19552 20952 19616
rect 21016 19552 21032 19616
rect 21096 19552 21112 19616
rect 21176 19552 21192 19616
rect 21256 19552 21264 19616
rect 20944 19551 21264 19552
rect 23520 19320 24000 19440
rect 2497 19274 2563 19277
rect 16297 19274 16363 19277
rect 2497 19272 16363 19274
rect 2497 19216 2502 19272
rect 2558 19216 16302 19272
rect 16358 19216 16363 19272
rect 2497 19214 16363 19216
rect 2497 19211 2563 19214
rect 16297 19211 16363 19214
rect 8944 19072 9264 19073
rect 0 19000 480 19032
rect 8944 19008 8952 19072
rect 9016 19008 9032 19072
rect 9096 19008 9112 19072
rect 9176 19008 9192 19072
rect 9256 19008 9264 19072
rect 8944 19007 9264 19008
rect 16944 19072 17264 19073
rect 16944 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17264 19072
rect 16944 19007 17264 19008
rect 0 18944 110 19000
rect 166 18944 480 19000
rect 0 18912 480 18944
rect 6821 18866 6887 18869
rect 18965 18866 19031 18869
rect 6821 18864 19031 18866
rect 6821 18808 6826 18864
rect 6882 18808 18970 18864
rect 19026 18808 19031 18864
rect 6821 18806 19031 18808
rect 6821 18803 6887 18806
rect 18965 18803 19031 18806
rect 20621 18866 20687 18869
rect 23614 18866 23674 19320
rect 20621 18864 23674 18866
rect 20621 18808 20626 18864
rect 20682 18808 23674 18864
rect 20621 18806 23674 18808
rect 20621 18803 20687 18806
rect 9949 18730 10015 18733
rect 18689 18730 18755 18733
rect 9949 18728 18755 18730
rect 9949 18672 9954 18728
rect 10010 18672 18694 18728
rect 18750 18672 18755 18728
rect 9949 18670 18755 18672
rect 9949 18667 10015 18670
rect 18689 18667 18755 18670
rect 4944 18528 5264 18529
rect 4944 18464 4952 18528
rect 5016 18464 5032 18528
rect 5096 18464 5112 18528
rect 5176 18464 5192 18528
rect 5256 18464 5264 18528
rect 4944 18463 5264 18464
rect 12944 18528 13264 18529
rect 12944 18464 12952 18528
rect 13016 18464 13032 18528
rect 13096 18464 13112 18528
rect 13176 18464 13192 18528
rect 13256 18464 13264 18528
rect 12944 18463 13264 18464
rect 20944 18528 21264 18529
rect 20944 18464 20952 18528
rect 21016 18464 21032 18528
rect 21096 18464 21112 18528
rect 21176 18464 21192 18528
rect 21256 18464 21264 18528
rect 20944 18463 21264 18464
rect 7373 18322 7439 18325
rect 20805 18322 20871 18325
rect 7373 18320 20871 18322
rect 7373 18264 7378 18320
rect 7434 18264 20810 18320
rect 20866 18264 20871 18320
rect 7373 18262 20871 18264
rect 7373 18259 7439 18262
rect 20805 18259 20871 18262
rect 10869 18186 10935 18189
rect 17401 18186 17467 18189
rect 10869 18184 17467 18186
rect 10869 18128 10874 18184
rect 10930 18128 17406 18184
rect 17462 18128 17467 18184
rect 10869 18126 17467 18128
rect 10869 18123 10935 18126
rect 17401 18123 17467 18126
rect 23520 18096 24000 18216
rect 8944 17984 9264 17985
rect 8944 17920 8952 17984
rect 9016 17920 9032 17984
rect 9096 17920 9112 17984
rect 9176 17920 9192 17984
rect 9256 17920 9264 17984
rect 8944 17919 9264 17920
rect 16944 17984 17264 17985
rect 16944 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17264 17984
rect 16944 17919 17264 17920
rect 0 17640 480 17672
rect 0 17584 110 17640
rect 166 17584 480 17640
rect 0 17552 480 17584
rect 21265 17642 21331 17645
rect 23614 17642 23674 18096
rect 21265 17640 23674 17642
rect 21265 17584 21270 17640
rect 21326 17584 23674 17640
rect 21265 17582 23674 17584
rect 21265 17579 21331 17582
rect 4944 17440 5264 17441
rect 4944 17376 4952 17440
rect 5016 17376 5032 17440
rect 5096 17376 5112 17440
rect 5176 17376 5192 17440
rect 5256 17376 5264 17440
rect 4944 17375 5264 17376
rect 12944 17440 13264 17441
rect 12944 17376 12952 17440
rect 13016 17376 13032 17440
rect 13096 17376 13112 17440
rect 13176 17376 13192 17440
rect 13256 17376 13264 17440
rect 12944 17375 13264 17376
rect 20944 17440 21264 17441
rect 20944 17376 20952 17440
rect 21016 17376 21032 17440
rect 21096 17376 21112 17440
rect 21176 17376 21192 17440
rect 21256 17376 21264 17440
rect 20944 17375 21264 17376
rect 8944 16896 9264 16897
rect 8944 16832 8952 16896
rect 9016 16832 9032 16896
rect 9096 16832 9112 16896
rect 9176 16832 9192 16896
rect 9256 16832 9264 16896
rect 8944 16831 9264 16832
rect 16944 16896 17264 16897
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 23520 16872 24000 16992
rect 16944 16831 17264 16832
rect 21449 16418 21515 16421
rect 23614 16418 23674 16872
rect 21449 16416 23674 16418
rect 21449 16360 21454 16416
rect 21510 16360 23674 16416
rect 21449 16358 23674 16360
rect 21449 16355 21515 16358
rect 4944 16352 5264 16353
rect 4944 16288 4952 16352
rect 5016 16288 5032 16352
rect 5096 16288 5112 16352
rect 5176 16288 5192 16352
rect 5256 16288 5264 16352
rect 4944 16287 5264 16288
rect 12944 16352 13264 16353
rect 12944 16288 12952 16352
rect 13016 16288 13032 16352
rect 13096 16288 13112 16352
rect 13176 16288 13192 16352
rect 13256 16288 13264 16352
rect 12944 16287 13264 16288
rect 20944 16352 21264 16353
rect 20944 16288 20952 16352
rect 21016 16288 21032 16352
rect 21096 16288 21112 16352
rect 21176 16288 21192 16352
rect 21256 16288 21264 16352
rect 20944 16287 21264 16288
rect 0 16144 480 16176
rect 0 16088 110 16144
rect 166 16088 480 16144
rect 0 16056 480 16088
rect 8944 15808 9264 15809
rect 8944 15744 8952 15808
rect 9016 15744 9032 15808
rect 9096 15744 9112 15808
rect 9176 15744 9192 15808
rect 9256 15744 9264 15808
rect 8944 15743 9264 15744
rect 16944 15808 17264 15809
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 16944 15743 17264 15744
rect 23520 15648 24000 15768
rect 21265 15466 21331 15469
rect 23614 15466 23674 15648
rect 21265 15464 23674 15466
rect 21265 15408 21270 15464
rect 21326 15408 23674 15464
rect 21265 15406 23674 15408
rect 21265 15403 21331 15406
rect 4944 15264 5264 15265
rect 4944 15200 4952 15264
rect 5016 15200 5032 15264
rect 5096 15200 5112 15264
rect 5176 15200 5192 15264
rect 5256 15200 5264 15264
rect 4944 15199 5264 15200
rect 12944 15264 13264 15265
rect 12944 15200 12952 15264
rect 13016 15200 13032 15264
rect 13096 15200 13112 15264
rect 13176 15200 13192 15264
rect 13256 15200 13264 15264
rect 12944 15199 13264 15200
rect 20944 15264 21264 15265
rect 20944 15200 20952 15264
rect 21016 15200 21032 15264
rect 21096 15200 21112 15264
rect 21176 15200 21192 15264
rect 21256 15200 21264 15264
rect 20944 15199 21264 15200
rect 0 14696 480 14816
rect 8944 14720 9264 14721
rect 62 14242 122 14696
rect 8944 14656 8952 14720
rect 9016 14656 9032 14720
rect 9096 14656 9112 14720
rect 9176 14656 9192 14720
rect 9256 14656 9264 14720
rect 8944 14655 9264 14656
rect 16944 14720 17264 14721
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 16944 14655 17264 14656
rect 23520 14288 24000 14408
rect 3417 14242 3483 14245
rect 62 14240 3483 14242
rect 62 14184 3422 14240
rect 3478 14184 3483 14240
rect 62 14182 3483 14184
rect 3417 14179 3483 14182
rect 4944 14176 5264 14177
rect 4944 14112 4952 14176
rect 5016 14112 5032 14176
rect 5096 14112 5112 14176
rect 5176 14112 5192 14176
rect 5256 14112 5264 14176
rect 4944 14111 5264 14112
rect 12944 14176 13264 14177
rect 12944 14112 12952 14176
rect 13016 14112 13032 14176
rect 13096 14112 13112 14176
rect 13176 14112 13192 14176
rect 13256 14112 13264 14176
rect 12944 14111 13264 14112
rect 20944 14176 21264 14177
rect 20944 14112 20952 14176
rect 21016 14112 21032 14176
rect 21096 14112 21112 14176
rect 21176 14112 21192 14176
rect 21256 14112 21264 14176
rect 20944 14111 21264 14112
rect 21081 13970 21147 13973
rect 23614 13970 23674 14288
rect 21081 13968 23674 13970
rect 21081 13912 21086 13968
rect 21142 13912 23674 13968
rect 21081 13910 23674 13912
rect 21081 13907 21147 13910
rect 9397 13698 9463 13701
rect 12801 13698 12867 13701
rect 9397 13696 12867 13698
rect 9397 13640 9402 13696
rect 9458 13640 12806 13696
rect 12862 13640 12867 13696
rect 9397 13638 12867 13640
rect 9397 13635 9463 13638
rect 12801 13635 12867 13638
rect 8944 13632 9264 13633
rect 8944 13568 8952 13632
rect 9016 13568 9032 13632
rect 9096 13568 9112 13632
rect 9176 13568 9192 13632
rect 9256 13568 9264 13632
rect 8944 13567 9264 13568
rect 16944 13632 17264 13633
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 16944 13567 17264 13568
rect 0 13424 480 13456
rect 0 13368 110 13424
rect 166 13368 480 13424
rect 0 13336 480 13368
rect 4944 13088 5264 13089
rect 4944 13024 4952 13088
rect 5016 13024 5032 13088
rect 5096 13024 5112 13088
rect 5176 13024 5192 13088
rect 5256 13024 5264 13088
rect 4944 13023 5264 13024
rect 12944 13088 13264 13089
rect 12944 13024 12952 13088
rect 13016 13024 13032 13088
rect 13096 13024 13112 13088
rect 13176 13024 13192 13088
rect 13256 13024 13264 13088
rect 12944 13023 13264 13024
rect 20944 13088 21264 13089
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 23520 13064 24000 13184
rect 20944 13023 21264 13024
rect 9121 12882 9187 12885
rect 23614 12882 23674 13064
rect 9121 12880 23674 12882
rect 9121 12824 9126 12880
rect 9182 12824 23674 12880
rect 9121 12822 23674 12824
rect 9121 12819 9187 12822
rect 8944 12544 9264 12545
rect 8944 12480 8952 12544
rect 9016 12480 9032 12544
rect 9096 12480 9112 12544
rect 9176 12480 9192 12544
rect 9256 12480 9264 12544
rect 8944 12479 9264 12480
rect 16944 12544 17264 12545
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 16944 12479 17264 12480
rect 4944 12000 5264 12001
rect 0 11840 480 11960
rect 4944 11936 4952 12000
rect 5016 11936 5032 12000
rect 5096 11936 5112 12000
rect 5176 11936 5192 12000
rect 5256 11936 5264 12000
rect 4944 11935 5264 11936
rect 12944 12000 13264 12001
rect 12944 11936 12952 12000
rect 13016 11936 13032 12000
rect 13096 11936 13112 12000
rect 13176 11936 13192 12000
rect 13256 11936 13264 12000
rect 12944 11935 13264 11936
rect 20944 12000 21264 12001
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 11935 21264 11936
rect 23520 11930 24000 11960
rect 23484 11928 24000 11930
rect 23484 11872 23570 11928
rect 23626 11872 24000 11928
rect 23484 11870 24000 11872
rect 23520 11840 24000 11870
rect 62 11386 122 11840
rect 3693 11794 3759 11797
rect 10961 11794 11027 11797
rect 3693 11792 11027 11794
rect 3693 11736 3698 11792
rect 3754 11736 10966 11792
rect 11022 11736 11027 11792
rect 3693 11734 11027 11736
rect 3693 11731 3759 11734
rect 10961 11731 11027 11734
rect 5441 11658 5507 11661
rect 20713 11658 20779 11661
rect 5441 11656 20779 11658
rect 5441 11600 5446 11656
rect 5502 11600 20718 11656
rect 20774 11600 20779 11656
rect 5441 11598 20779 11600
rect 5441 11595 5507 11598
rect 20713 11595 20779 11598
rect 8944 11456 9264 11457
rect 8944 11392 8952 11456
rect 9016 11392 9032 11456
rect 9096 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9264 11456
rect 8944 11391 9264 11392
rect 16944 11456 17264 11457
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 11391 17264 11392
rect 1577 11386 1643 11389
rect 62 11384 1643 11386
rect 62 11328 1582 11384
rect 1638 11328 1643 11384
rect 62 11326 1643 11328
rect 1577 11323 1643 11326
rect 4944 10912 5264 10913
rect 4944 10848 4952 10912
rect 5016 10848 5032 10912
rect 5096 10848 5112 10912
rect 5176 10848 5192 10912
rect 5256 10848 5264 10912
rect 4944 10847 5264 10848
rect 12944 10912 13264 10913
rect 12944 10848 12952 10912
rect 13016 10848 13032 10912
rect 13096 10848 13112 10912
rect 13176 10848 13192 10912
rect 13256 10848 13264 10912
rect 12944 10847 13264 10848
rect 20944 10912 21264 10913
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 10847 21264 10848
rect 23520 10616 24000 10736
rect 0 10480 480 10600
rect 62 10298 122 10480
rect 8944 10368 9264 10369
rect 8944 10304 8952 10368
rect 9016 10304 9032 10368
rect 9096 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9264 10368
rect 8944 10303 9264 10304
rect 16944 10368 17264 10369
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 16944 10303 17264 10304
rect 1577 10298 1643 10301
rect 62 10296 1643 10298
rect 62 10240 1582 10296
rect 1638 10240 1643 10296
rect 62 10238 1643 10240
rect 1577 10235 1643 10238
rect 21081 10298 21147 10301
rect 23614 10298 23674 10616
rect 21081 10296 23674 10298
rect 21081 10240 21086 10296
rect 21142 10240 23674 10296
rect 21081 10238 23674 10240
rect 21081 10235 21147 10238
rect 4944 9824 5264 9825
rect 4944 9760 4952 9824
rect 5016 9760 5032 9824
rect 5096 9760 5112 9824
rect 5176 9760 5192 9824
rect 5256 9760 5264 9824
rect 4944 9759 5264 9760
rect 12944 9824 13264 9825
rect 12944 9760 12952 9824
rect 13016 9760 13032 9824
rect 13096 9760 13112 9824
rect 13176 9760 13192 9824
rect 13256 9760 13264 9824
rect 12944 9759 13264 9760
rect 20944 9824 21264 9825
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 9759 21264 9760
rect 4061 9618 4127 9621
rect 5809 9618 5875 9621
rect 4061 9616 5875 9618
rect 4061 9560 4066 9616
rect 4122 9560 5814 9616
rect 5870 9560 5875 9616
rect 4061 9558 5875 9560
rect 4061 9555 4127 9558
rect 5809 9555 5875 9558
rect 8109 9618 8175 9621
rect 20805 9618 20871 9621
rect 8109 9616 20871 9618
rect 8109 9560 8114 9616
rect 8170 9560 20810 9616
rect 20866 9560 20871 9616
rect 8109 9558 20871 9560
rect 8109 9555 8175 9558
rect 20805 9555 20871 9558
rect 8944 9280 9264 9281
rect 0 9120 480 9240
rect 8944 9216 8952 9280
rect 9016 9216 9032 9280
rect 9096 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9264 9280
rect 8944 9215 9264 9216
rect 16944 9280 17264 9281
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 23520 9256 24000 9376
rect 16944 9215 17264 9216
rect 62 8666 122 9120
rect 18413 8938 18479 8941
rect 23614 8938 23674 9256
rect 18413 8936 23674 8938
rect 18413 8880 18418 8936
rect 18474 8880 23674 8936
rect 18413 8878 23674 8880
rect 18413 8875 18479 8878
rect 4944 8736 5264 8737
rect 4944 8672 4952 8736
rect 5016 8672 5032 8736
rect 5096 8672 5112 8736
rect 5176 8672 5192 8736
rect 5256 8672 5264 8736
rect 4944 8671 5264 8672
rect 12944 8736 13264 8737
rect 12944 8672 12952 8736
rect 13016 8672 13032 8736
rect 13096 8672 13112 8736
rect 13176 8672 13192 8736
rect 13256 8672 13264 8736
rect 12944 8671 13264 8672
rect 20944 8736 21264 8737
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 8671 21264 8672
rect 1577 8666 1643 8669
rect 62 8664 1643 8666
rect 62 8608 1582 8664
rect 1638 8608 1643 8664
rect 62 8606 1643 8608
rect 1577 8603 1643 8606
rect 3417 8530 3483 8533
rect 13261 8530 13327 8533
rect 14825 8530 14891 8533
rect 3417 8528 14891 8530
rect 3417 8472 3422 8528
rect 3478 8472 13266 8528
rect 13322 8472 14830 8528
rect 14886 8472 14891 8528
rect 3417 8470 14891 8472
rect 3417 8467 3483 8470
rect 13261 8467 13327 8470
rect 14825 8467 14891 8470
rect 8944 8192 9264 8193
rect 8944 8128 8952 8192
rect 9016 8128 9032 8192
rect 9096 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9264 8192
rect 8944 8127 9264 8128
rect 16944 8192 17264 8193
rect 16944 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17264 8192
rect 16944 8127 17264 8128
rect 23520 8032 24000 8152
rect 0 7624 480 7744
rect 4944 7648 5264 7649
rect 62 7170 122 7624
rect 4944 7584 4952 7648
rect 5016 7584 5032 7648
rect 5096 7584 5112 7648
rect 5176 7584 5192 7648
rect 5256 7584 5264 7648
rect 4944 7583 5264 7584
rect 12944 7648 13264 7649
rect 12944 7584 12952 7648
rect 13016 7584 13032 7648
rect 13096 7584 13112 7648
rect 13176 7584 13192 7648
rect 13256 7584 13264 7648
rect 12944 7583 13264 7584
rect 20944 7648 21264 7649
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 7583 21264 7584
rect 21357 7578 21423 7581
rect 23614 7578 23674 8032
rect 21357 7576 23674 7578
rect 21357 7520 21362 7576
rect 21418 7520 23674 7576
rect 21357 7518 23674 7520
rect 21357 7515 21423 7518
rect 1485 7306 1551 7309
rect 14549 7306 14615 7309
rect 1485 7304 14615 7306
rect 1485 7248 1490 7304
rect 1546 7248 14554 7304
rect 14610 7248 14615 7304
rect 1485 7246 14615 7248
rect 1485 7243 1551 7246
rect 14549 7243 14615 7246
rect 1853 7170 1919 7173
rect 62 7168 1919 7170
rect 62 7112 1858 7168
rect 1914 7112 1919 7168
rect 62 7110 1919 7112
rect 1853 7107 1919 7110
rect 8944 7104 9264 7105
rect 8944 7040 8952 7104
rect 9016 7040 9032 7104
rect 9096 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9264 7104
rect 8944 7039 9264 7040
rect 16944 7104 17264 7105
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16944 7039 17264 7040
rect 2221 6898 2287 6901
rect 23520 6898 24000 6928
rect 62 6896 2287 6898
rect 62 6840 2226 6896
rect 2282 6840 2287 6896
rect 62 6838 2287 6840
rect 23484 6896 24000 6898
rect 23484 6840 23570 6896
rect 23626 6840 24000 6896
rect 23484 6838 24000 6840
rect 62 6384 122 6838
rect 2221 6835 2287 6838
rect 23520 6808 24000 6838
rect 4944 6560 5264 6561
rect 4944 6496 4952 6560
rect 5016 6496 5032 6560
rect 5096 6496 5112 6560
rect 5176 6496 5192 6560
rect 5256 6496 5264 6560
rect 4944 6495 5264 6496
rect 12944 6560 13264 6561
rect 12944 6496 12952 6560
rect 13016 6496 13032 6560
rect 13096 6496 13112 6560
rect 13176 6496 13192 6560
rect 13256 6496 13264 6560
rect 12944 6495 13264 6496
rect 20944 6560 21264 6561
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 6495 21264 6496
rect 0 6264 480 6384
rect 8944 6016 9264 6017
rect 8944 5952 8952 6016
rect 9016 5952 9032 6016
rect 9096 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9264 6016
rect 8944 5951 9264 5952
rect 16944 6016 17264 6017
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 16944 5951 17264 5952
rect 9949 5810 10015 5813
rect 21449 5810 21515 5813
rect 9949 5808 21515 5810
rect 9949 5752 9954 5808
rect 10010 5752 21454 5808
rect 21510 5752 21515 5808
rect 9949 5750 21515 5752
rect 9949 5747 10015 5750
rect 21449 5747 21515 5750
rect 5809 5674 5875 5677
rect 23381 5674 23447 5677
rect 5809 5672 23447 5674
rect 5809 5616 5814 5672
rect 5870 5616 23386 5672
rect 23442 5616 23447 5672
rect 5809 5614 23447 5616
rect 5809 5611 5875 5614
rect 23381 5611 23447 5614
rect 23520 5584 24000 5704
rect 4944 5472 5264 5473
rect 4944 5408 4952 5472
rect 5016 5408 5032 5472
rect 5096 5408 5112 5472
rect 5176 5408 5192 5472
rect 5256 5408 5264 5472
rect 4944 5407 5264 5408
rect 12944 5472 13264 5473
rect 12944 5408 12952 5472
rect 13016 5408 13032 5472
rect 13096 5408 13112 5472
rect 13176 5408 13192 5472
rect 13256 5408 13264 5472
rect 12944 5407 13264 5408
rect 20944 5472 21264 5473
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 5407 21264 5408
rect 15653 5402 15719 5405
rect 20713 5402 20779 5405
rect 15653 5400 20779 5402
rect 15653 5344 15658 5400
rect 15714 5344 20718 5400
rect 20774 5344 20779 5400
rect 15653 5342 20779 5344
rect 15653 5339 15719 5342
rect 20670 5339 20779 5342
rect 7557 5266 7623 5269
rect 18321 5266 18387 5269
rect 7557 5264 18387 5266
rect 7557 5208 7562 5264
rect 7618 5208 18326 5264
rect 18382 5208 18387 5264
rect 7557 5206 18387 5208
rect 20670 5266 20730 5339
rect 23614 5266 23674 5584
rect 20670 5206 23674 5266
rect 7557 5203 7623 5206
rect 18321 5203 18387 5206
rect 12249 5130 12315 5133
rect 20621 5130 20687 5133
rect 12249 5128 20687 5130
rect 12249 5072 12254 5128
rect 12310 5072 20626 5128
rect 20682 5072 20687 5128
rect 12249 5070 20687 5072
rect 12249 5067 12315 5070
rect 20621 5067 20687 5070
rect 0 4904 480 5024
rect 8944 4928 9264 4929
rect 62 4450 122 4904
rect 8944 4864 8952 4928
rect 9016 4864 9032 4928
rect 9096 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9264 4928
rect 8944 4863 9264 4864
rect 16944 4928 17264 4929
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 16944 4863 17264 4864
rect 21449 4858 21515 4861
rect 21449 4856 23674 4858
rect 21449 4800 21454 4856
rect 21510 4800 23674 4856
rect 21449 4798 23674 4800
rect 21449 4795 21515 4798
rect 1577 4450 1643 4453
rect 62 4448 1643 4450
rect 62 4392 1582 4448
rect 1638 4392 1643 4448
rect 62 4390 1643 4392
rect 1577 4387 1643 4390
rect 4944 4384 5264 4385
rect 4944 4320 4952 4384
rect 5016 4320 5032 4384
rect 5096 4320 5112 4384
rect 5176 4320 5192 4384
rect 5256 4320 5264 4384
rect 4944 4319 5264 4320
rect 12944 4384 13264 4385
rect 12944 4320 12952 4384
rect 13016 4320 13032 4384
rect 13096 4320 13112 4384
rect 13176 4320 13192 4384
rect 13256 4320 13264 4384
rect 12944 4319 13264 4320
rect 20944 4384 21264 4385
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 23614 4344 23674 4798
rect 20944 4319 21264 4320
rect 5533 4314 5599 4317
rect 9949 4314 10015 4317
rect 20621 4314 20687 4317
rect 5533 4312 10015 4314
rect 5533 4256 5538 4312
rect 5594 4256 9954 4312
rect 10010 4256 10015 4312
rect 5533 4254 10015 4256
rect 5533 4251 5599 4254
rect 9949 4251 10015 4254
rect 13770 4312 20687 4314
rect 13770 4256 20626 4312
rect 20682 4256 20687 4312
rect 13770 4254 20687 4256
rect 11513 4178 11579 4181
rect 13770 4178 13830 4254
rect 20621 4251 20687 4254
rect 23520 4224 24000 4344
rect 11513 4176 13830 4178
rect 11513 4120 11518 4176
rect 11574 4120 13830 4176
rect 11513 4118 13830 4120
rect 11513 4115 11579 4118
rect 3969 4042 4035 4045
rect 9765 4042 9831 4045
rect 3969 4040 9831 4042
rect 3969 3984 3974 4040
rect 4030 3984 9770 4040
rect 9826 3984 9831 4040
rect 3969 3982 9831 3984
rect 3969 3979 4035 3982
rect 9765 3979 9831 3982
rect 8944 3840 9264 3841
rect 8944 3776 8952 3840
rect 9016 3776 9032 3840
rect 9096 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9264 3840
rect 8944 3775 9264 3776
rect 16944 3840 17264 3841
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16944 3775 17264 3776
rect 9673 3770 9739 3773
rect 11053 3770 11119 3773
rect 14089 3770 14155 3773
rect 9673 3768 14155 3770
rect 9673 3712 9678 3768
rect 9734 3712 11058 3768
rect 11114 3712 14094 3768
rect 14150 3712 14155 3768
rect 9673 3710 14155 3712
rect 9673 3707 9739 3710
rect 11053 3707 11119 3710
rect 14089 3707 14155 3710
rect 6269 3634 6335 3637
rect 12433 3634 12499 3637
rect 6269 3632 12499 3634
rect 6269 3576 6274 3632
rect 6330 3576 12438 3632
rect 12494 3576 12499 3632
rect 6269 3574 12499 3576
rect 6269 3571 6335 3574
rect 12433 3571 12499 3574
rect 20621 3634 20687 3637
rect 20621 3632 23674 3634
rect 20621 3576 20626 3632
rect 20682 3576 23674 3632
rect 20621 3574 23674 3576
rect 20621 3571 20687 3574
rect 0 3500 480 3528
rect 0 3436 60 3500
rect 124 3436 480 3500
rect 0 3408 480 3436
rect 4944 3296 5264 3297
rect 4944 3232 4952 3296
rect 5016 3232 5032 3296
rect 5096 3232 5112 3296
rect 5176 3232 5192 3296
rect 5256 3232 5264 3296
rect 4944 3231 5264 3232
rect 12944 3296 13264 3297
rect 12944 3232 12952 3296
rect 13016 3232 13032 3296
rect 13096 3232 13112 3296
rect 13176 3232 13192 3296
rect 13256 3232 13264 3296
rect 12944 3231 13264 3232
rect 20944 3296 21264 3297
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 3231 21264 3232
rect 54 3164 60 3228
rect 124 3226 130 3228
rect 1577 3226 1643 3229
rect 124 3224 1643 3226
rect 124 3168 1582 3224
rect 1638 3168 1643 3224
rect 124 3166 1643 3168
rect 124 3164 130 3166
rect 1577 3163 1643 3166
rect 23614 3120 23674 3574
rect 9305 3090 9371 3093
rect 17401 3090 17467 3093
rect 9305 3088 17467 3090
rect 9305 3032 9310 3088
rect 9366 3032 17406 3088
rect 17462 3032 17467 3088
rect 9305 3030 17467 3032
rect 9305 3027 9371 3030
rect 17401 3027 17467 3030
rect 23520 3000 24000 3120
rect 7189 2954 7255 2957
rect 11697 2954 11763 2957
rect 19333 2954 19399 2957
rect 7189 2952 19399 2954
rect 7189 2896 7194 2952
rect 7250 2896 11702 2952
rect 11758 2896 19338 2952
rect 19394 2896 19399 2952
rect 7189 2894 19399 2896
rect 7189 2891 7255 2894
rect 11697 2891 11763 2894
rect 19333 2891 19399 2894
rect 4889 2818 4955 2821
rect 7649 2818 7715 2821
rect 4889 2816 7715 2818
rect 4889 2760 4894 2816
rect 4950 2760 7654 2816
rect 7710 2760 7715 2816
rect 4889 2758 7715 2760
rect 4889 2755 4955 2758
rect 7649 2755 7715 2758
rect 8944 2752 9264 2753
rect 8944 2688 8952 2752
rect 9016 2688 9032 2752
rect 9096 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9264 2752
rect 8944 2687 9264 2688
rect 16944 2752 17264 2753
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 16944 2687 17264 2688
rect 2037 2546 2103 2549
rect 4429 2546 4495 2549
rect 14273 2546 14339 2549
rect 2037 2544 4170 2546
rect 2037 2488 2042 2544
rect 2098 2488 4170 2544
rect 2037 2486 4170 2488
rect 2037 2483 2103 2486
rect 4110 2410 4170 2486
rect 4429 2544 14339 2546
rect 4429 2488 4434 2544
rect 4490 2488 14278 2544
rect 14334 2488 14339 2544
rect 4429 2486 14339 2488
rect 4429 2483 4495 2486
rect 14273 2483 14339 2486
rect 12157 2410 12223 2413
rect 4110 2408 12223 2410
rect 4110 2352 12162 2408
rect 12218 2352 12223 2408
rect 4110 2350 12223 2352
rect 12157 2347 12223 2350
rect 12433 2410 12499 2413
rect 12433 2408 23674 2410
rect 12433 2352 12438 2408
rect 12494 2352 23674 2408
rect 12433 2350 23674 2352
rect 12433 2347 12499 2350
rect 4944 2208 5264 2209
rect 0 2136 480 2168
rect 4944 2144 4952 2208
rect 5016 2144 5032 2208
rect 5096 2144 5112 2208
rect 5176 2144 5192 2208
rect 5256 2144 5264 2208
rect 4944 2143 5264 2144
rect 12944 2208 13264 2209
rect 12944 2144 12952 2208
rect 13016 2144 13032 2208
rect 13096 2144 13112 2208
rect 13176 2144 13192 2208
rect 13256 2144 13264 2208
rect 12944 2143 13264 2144
rect 20944 2208 21264 2209
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2143 21264 2144
rect 0 2080 110 2136
rect 166 2080 480 2136
rect 0 2048 480 2080
rect 8937 2002 9003 2005
rect 15469 2002 15535 2005
rect 8937 2000 15535 2002
rect 8937 1944 8942 2000
rect 8998 1944 15474 2000
rect 15530 1944 15535 2000
rect 8937 1942 15535 1944
rect 8937 1939 9003 1942
rect 15469 1939 15535 1942
rect 23614 1896 23674 2350
rect 23520 1776 24000 1896
rect 1945 1322 2011 1325
rect 62 1320 2011 1322
rect 62 1264 1950 1320
rect 2006 1264 2011 1320
rect 62 1262 2011 1264
rect 62 808 122 1262
rect 1945 1259 2011 1262
rect 0 688 480 808
rect 7649 642 7715 645
rect 23520 642 24000 672
rect 7649 640 24000 642
rect 7649 584 7654 640
rect 7710 584 24000 640
rect 7649 582 24000 584
rect 7649 579 7715 582
rect 23520 552 24000 582
<< via3 >>
rect 4952 21788 5016 21792
rect 4952 21732 4956 21788
rect 4956 21732 5012 21788
rect 5012 21732 5016 21788
rect 4952 21728 5016 21732
rect 5032 21788 5096 21792
rect 5032 21732 5036 21788
rect 5036 21732 5092 21788
rect 5092 21732 5096 21788
rect 5032 21728 5096 21732
rect 5112 21788 5176 21792
rect 5112 21732 5116 21788
rect 5116 21732 5172 21788
rect 5172 21732 5176 21788
rect 5112 21728 5176 21732
rect 5192 21788 5256 21792
rect 5192 21732 5196 21788
rect 5196 21732 5252 21788
rect 5252 21732 5256 21788
rect 5192 21728 5256 21732
rect 12952 21788 13016 21792
rect 12952 21732 12956 21788
rect 12956 21732 13012 21788
rect 13012 21732 13016 21788
rect 12952 21728 13016 21732
rect 13032 21788 13096 21792
rect 13032 21732 13036 21788
rect 13036 21732 13092 21788
rect 13092 21732 13096 21788
rect 13032 21728 13096 21732
rect 13112 21788 13176 21792
rect 13112 21732 13116 21788
rect 13116 21732 13172 21788
rect 13172 21732 13176 21788
rect 13112 21728 13176 21732
rect 13192 21788 13256 21792
rect 13192 21732 13196 21788
rect 13196 21732 13252 21788
rect 13252 21732 13256 21788
rect 13192 21728 13256 21732
rect 20952 21788 21016 21792
rect 20952 21732 20956 21788
rect 20956 21732 21012 21788
rect 21012 21732 21016 21788
rect 20952 21728 21016 21732
rect 21032 21788 21096 21792
rect 21032 21732 21036 21788
rect 21036 21732 21092 21788
rect 21092 21732 21096 21788
rect 21032 21728 21096 21732
rect 21112 21788 21176 21792
rect 21112 21732 21116 21788
rect 21116 21732 21172 21788
rect 21172 21732 21176 21788
rect 21112 21728 21176 21732
rect 21192 21788 21256 21792
rect 21192 21732 21196 21788
rect 21196 21732 21252 21788
rect 21252 21732 21256 21788
rect 21192 21728 21256 21732
rect 8952 21244 9016 21248
rect 8952 21188 8956 21244
rect 8956 21188 9012 21244
rect 9012 21188 9016 21244
rect 8952 21184 9016 21188
rect 9032 21244 9096 21248
rect 9032 21188 9036 21244
rect 9036 21188 9092 21244
rect 9092 21188 9096 21244
rect 9032 21184 9096 21188
rect 9112 21244 9176 21248
rect 9112 21188 9116 21244
rect 9116 21188 9172 21244
rect 9172 21188 9176 21244
rect 9112 21184 9176 21188
rect 9192 21244 9256 21248
rect 9192 21188 9196 21244
rect 9196 21188 9252 21244
rect 9252 21188 9256 21244
rect 9192 21184 9256 21188
rect 16952 21244 17016 21248
rect 16952 21188 16956 21244
rect 16956 21188 17012 21244
rect 17012 21188 17016 21244
rect 16952 21184 17016 21188
rect 17032 21244 17096 21248
rect 17032 21188 17036 21244
rect 17036 21188 17092 21244
rect 17092 21188 17096 21244
rect 17032 21184 17096 21188
rect 17112 21244 17176 21248
rect 17112 21188 17116 21244
rect 17116 21188 17172 21244
rect 17172 21188 17176 21244
rect 17112 21184 17176 21188
rect 17192 21244 17256 21248
rect 17192 21188 17196 21244
rect 17196 21188 17252 21244
rect 17252 21188 17256 21244
rect 17192 21184 17256 21188
rect 4952 20700 5016 20704
rect 4952 20644 4956 20700
rect 4956 20644 5012 20700
rect 5012 20644 5016 20700
rect 4952 20640 5016 20644
rect 5032 20700 5096 20704
rect 5032 20644 5036 20700
rect 5036 20644 5092 20700
rect 5092 20644 5096 20700
rect 5032 20640 5096 20644
rect 5112 20700 5176 20704
rect 5112 20644 5116 20700
rect 5116 20644 5172 20700
rect 5172 20644 5176 20700
rect 5112 20640 5176 20644
rect 5192 20700 5256 20704
rect 5192 20644 5196 20700
rect 5196 20644 5252 20700
rect 5252 20644 5256 20700
rect 5192 20640 5256 20644
rect 12952 20700 13016 20704
rect 12952 20644 12956 20700
rect 12956 20644 13012 20700
rect 13012 20644 13016 20700
rect 12952 20640 13016 20644
rect 13032 20700 13096 20704
rect 13032 20644 13036 20700
rect 13036 20644 13092 20700
rect 13092 20644 13096 20700
rect 13032 20640 13096 20644
rect 13112 20700 13176 20704
rect 13112 20644 13116 20700
rect 13116 20644 13172 20700
rect 13172 20644 13176 20700
rect 13112 20640 13176 20644
rect 13192 20700 13256 20704
rect 13192 20644 13196 20700
rect 13196 20644 13252 20700
rect 13252 20644 13256 20700
rect 13192 20640 13256 20644
rect 20952 20700 21016 20704
rect 20952 20644 20956 20700
rect 20956 20644 21012 20700
rect 21012 20644 21016 20700
rect 20952 20640 21016 20644
rect 21032 20700 21096 20704
rect 21032 20644 21036 20700
rect 21036 20644 21092 20700
rect 21092 20644 21096 20700
rect 21032 20640 21096 20644
rect 21112 20700 21176 20704
rect 21112 20644 21116 20700
rect 21116 20644 21172 20700
rect 21172 20644 21176 20700
rect 21112 20640 21176 20644
rect 21192 20700 21256 20704
rect 21192 20644 21196 20700
rect 21196 20644 21252 20700
rect 21252 20644 21256 20700
rect 21192 20640 21256 20644
rect 8952 20156 9016 20160
rect 8952 20100 8956 20156
rect 8956 20100 9012 20156
rect 9012 20100 9016 20156
rect 8952 20096 9016 20100
rect 9032 20156 9096 20160
rect 9032 20100 9036 20156
rect 9036 20100 9092 20156
rect 9092 20100 9096 20156
rect 9032 20096 9096 20100
rect 9112 20156 9176 20160
rect 9112 20100 9116 20156
rect 9116 20100 9172 20156
rect 9172 20100 9176 20156
rect 9112 20096 9176 20100
rect 9192 20156 9256 20160
rect 9192 20100 9196 20156
rect 9196 20100 9252 20156
rect 9252 20100 9256 20156
rect 9192 20096 9256 20100
rect 16952 20156 17016 20160
rect 16952 20100 16956 20156
rect 16956 20100 17012 20156
rect 17012 20100 17016 20156
rect 16952 20096 17016 20100
rect 17032 20156 17096 20160
rect 17032 20100 17036 20156
rect 17036 20100 17092 20156
rect 17092 20100 17096 20156
rect 17032 20096 17096 20100
rect 17112 20156 17176 20160
rect 17112 20100 17116 20156
rect 17116 20100 17172 20156
rect 17172 20100 17176 20156
rect 17112 20096 17176 20100
rect 17192 20156 17256 20160
rect 17192 20100 17196 20156
rect 17196 20100 17252 20156
rect 17252 20100 17256 20156
rect 17192 20096 17256 20100
rect 4952 19612 5016 19616
rect 4952 19556 4956 19612
rect 4956 19556 5012 19612
rect 5012 19556 5016 19612
rect 4952 19552 5016 19556
rect 5032 19612 5096 19616
rect 5032 19556 5036 19612
rect 5036 19556 5092 19612
rect 5092 19556 5096 19612
rect 5032 19552 5096 19556
rect 5112 19612 5176 19616
rect 5112 19556 5116 19612
rect 5116 19556 5172 19612
rect 5172 19556 5176 19612
rect 5112 19552 5176 19556
rect 5192 19612 5256 19616
rect 5192 19556 5196 19612
rect 5196 19556 5252 19612
rect 5252 19556 5256 19612
rect 5192 19552 5256 19556
rect 12952 19612 13016 19616
rect 12952 19556 12956 19612
rect 12956 19556 13012 19612
rect 13012 19556 13016 19612
rect 12952 19552 13016 19556
rect 13032 19612 13096 19616
rect 13032 19556 13036 19612
rect 13036 19556 13092 19612
rect 13092 19556 13096 19612
rect 13032 19552 13096 19556
rect 13112 19612 13176 19616
rect 13112 19556 13116 19612
rect 13116 19556 13172 19612
rect 13172 19556 13176 19612
rect 13112 19552 13176 19556
rect 13192 19612 13256 19616
rect 13192 19556 13196 19612
rect 13196 19556 13252 19612
rect 13252 19556 13256 19612
rect 13192 19552 13256 19556
rect 20952 19612 21016 19616
rect 20952 19556 20956 19612
rect 20956 19556 21012 19612
rect 21012 19556 21016 19612
rect 20952 19552 21016 19556
rect 21032 19612 21096 19616
rect 21032 19556 21036 19612
rect 21036 19556 21092 19612
rect 21092 19556 21096 19612
rect 21032 19552 21096 19556
rect 21112 19612 21176 19616
rect 21112 19556 21116 19612
rect 21116 19556 21172 19612
rect 21172 19556 21176 19612
rect 21112 19552 21176 19556
rect 21192 19612 21256 19616
rect 21192 19556 21196 19612
rect 21196 19556 21252 19612
rect 21252 19556 21256 19612
rect 21192 19552 21256 19556
rect 8952 19068 9016 19072
rect 8952 19012 8956 19068
rect 8956 19012 9012 19068
rect 9012 19012 9016 19068
rect 8952 19008 9016 19012
rect 9032 19068 9096 19072
rect 9032 19012 9036 19068
rect 9036 19012 9092 19068
rect 9092 19012 9096 19068
rect 9032 19008 9096 19012
rect 9112 19068 9176 19072
rect 9112 19012 9116 19068
rect 9116 19012 9172 19068
rect 9172 19012 9176 19068
rect 9112 19008 9176 19012
rect 9192 19068 9256 19072
rect 9192 19012 9196 19068
rect 9196 19012 9252 19068
rect 9252 19012 9256 19068
rect 9192 19008 9256 19012
rect 16952 19068 17016 19072
rect 16952 19012 16956 19068
rect 16956 19012 17012 19068
rect 17012 19012 17016 19068
rect 16952 19008 17016 19012
rect 17032 19068 17096 19072
rect 17032 19012 17036 19068
rect 17036 19012 17092 19068
rect 17092 19012 17096 19068
rect 17032 19008 17096 19012
rect 17112 19068 17176 19072
rect 17112 19012 17116 19068
rect 17116 19012 17172 19068
rect 17172 19012 17176 19068
rect 17112 19008 17176 19012
rect 17192 19068 17256 19072
rect 17192 19012 17196 19068
rect 17196 19012 17252 19068
rect 17252 19012 17256 19068
rect 17192 19008 17256 19012
rect 4952 18524 5016 18528
rect 4952 18468 4956 18524
rect 4956 18468 5012 18524
rect 5012 18468 5016 18524
rect 4952 18464 5016 18468
rect 5032 18524 5096 18528
rect 5032 18468 5036 18524
rect 5036 18468 5092 18524
rect 5092 18468 5096 18524
rect 5032 18464 5096 18468
rect 5112 18524 5176 18528
rect 5112 18468 5116 18524
rect 5116 18468 5172 18524
rect 5172 18468 5176 18524
rect 5112 18464 5176 18468
rect 5192 18524 5256 18528
rect 5192 18468 5196 18524
rect 5196 18468 5252 18524
rect 5252 18468 5256 18524
rect 5192 18464 5256 18468
rect 12952 18524 13016 18528
rect 12952 18468 12956 18524
rect 12956 18468 13012 18524
rect 13012 18468 13016 18524
rect 12952 18464 13016 18468
rect 13032 18524 13096 18528
rect 13032 18468 13036 18524
rect 13036 18468 13092 18524
rect 13092 18468 13096 18524
rect 13032 18464 13096 18468
rect 13112 18524 13176 18528
rect 13112 18468 13116 18524
rect 13116 18468 13172 18524
rect 13172 18468 13176 18524
rect 13112 18464 13176 18468
rect 13192 18524 13256 18528
rect 13192 18468 13196 18524
rect 13196 18468 13252 18524
rect 13252 18468 13256 18524
rect 13192 18464 13256 18468
rect 20952 18524 21016 18528
rect 20952 18468 20956 18524
rect 20956 18468 21012 18524
rect 21012 18468 21016 18524
rect 20952 18464 21016 18468
rect 21032 18524 21096 18528
rect 21032 18468 21036 18524
rect 21036 18468 21092 18524
rect 21092 18468 21096 18524
rect 21032 18464 21096 18468
rect 21112 18524 21176 18528
rect 21112 18468 21116 18524
rect 21116 18468 21172 18524
rect 21172 18468 21176 18524
rect 21112 18464 21176 18468
rect 21192 18524 21256 18528
rect 21192 18468 21196 18524
rect 21196 18468 21252 18524
rect 21252 18468 21256 18524
rect 21192 18464 21256 18468
rect 8952 17980 9016 17984
rect 8952 17924 8956 17980
rect 8956 17924 9012 17980
rect 9012 17924 9016 17980
rect 8952 17920 9016 17924
rect 9032 17980 9096 17984
rect 9032 17924 9036 17980
rect 9036 17924 9092 17980
rect 9092 17924 9096 17980
rect 9032 17920 9096 17924
rect 9112 17980 9176 17984
rect 9112 17924 9116 17980
rect 9116 17924 9172 17980
rect 9172 17924 9176 17980
rect 9112 17920 9176 17924
rect 9192 17980 9256 17984
rect 9192 17924 9196 17980
rect 9196 17924 9252 17980
rect 9252 17924 9256 17980
rect 9192 17920 9256 17924
rect 16952 17980 17016 17984
rect 16952 17924 16956 17980
rect 16956 17924 17012 17980
rect 17012 17924 17016 17980
rect 16952 17920 17016 17924
rect 17032 17980 17096 17984
rect 17032 17924 17036 17980
rect 17036 17924 17092 17980
rect 17092 17924 17096 17980
rect 17032 17920 17096 17924
rect 17112 17980 17176 17984
rect 17112 17924 17116 17980
rect 17116 17924 17172 17980
rect 17172 17924 17176 17980
rect 17112 17920 17176 17924
rect 17192 17980 17256 17984
rect 17192 17924 17196 17980
rect 17196 17924 17252 17980
rect 17252 17924 17256 17980
rect 17192 17920 17256 17924
rect 4952 17436 5016 17440
rect 4952 17380 4956 17436
rect 4956 17380 5012 17436
rect 5012 17380 5016 17436
rect 4952 17376 5016 17380
rect 5032 17436 5096 17440
rect 5032 17380 5036 17436
rect 5036 17380 5092 17436
rect 5092 17380 5096 17436
rect 5032 17376 5096 17380
rect 5112 17436 5176 17440
rect 5112 17380 5116 17436
rect 5116 17380 5172 17436
rect 5172 17380 5176 17436
rect 5112 17376 5176 17380
rect 5192 17436 5256 17440
rect 5192 17380 5196 17436
rect 5196 17380 5252 17436
rect 5252 17380 5256 17436
rect 5192 17376 5256 17380
rect 12952 17436 13016 17440
rect 12952 17380 12956 17436
rect 12956 17380 13012 17436
rect 13012 17380 13016 17436
rect 12952 17376 13016 17380
rect 13032 17436 13096 17440
rect 13032 17380 13036 17436
rect 13036 17380 13092 17436
rect 13092 17380 13096 17436
rect 13032 17376 13096 17380
rect 13112 17436 13176 17440
rect 13112 17380 13116 17436
rect 13116 17380 13172 17436
rect 13172 17380 13176 17436
rect 13112 17376 13176 17380
rect 13192 17436 13256 17440
rect 13192 17380 13196 17436
rect 13196 17380 13252 17436
rect 13252 17380 13256 17436
rect 13192 17376 13256 17380
rect 20952 17436 21016 17440
rect 20952 17380 20956 17436
rect 20956 17380 21012 17436
rect 21012 17380 21016 17436
rect 20952 17376 21016 17380
rect 21032 17436 21096 17440
rect 21032 17380 21036 17436
rect 21036 17380 21092 17436
rect 21092 17380 21096 17436
rect 21032 17376 21096 17380
rect 21112 17436 21176 17440
rect 21112 17380 21116 17436
rect 21116 17380 21172 17436
rect 21172 17380 21176 17436
rect 21112 17376 21176 17380
rect 21192 17436 21256 17440
rect 21192 17380 21196 17436
rect 21196 17380 21252 17436
rect 21252 17380 21256 17436
rect 21192 17376 21256 17380
rect 8952 16892 9016 16896
rect 8952 16836 8956 16892
rect 8956 16836 9012 16892
rect 9012 16836 9016 16892
rect 8952 16832 9016 16836
rect 9032 16892 9096 16896
rect 9032 16836 9036 16892
rect 9036 16836 9092 16892
rect 9092 16836 9096 16892
rect 9032 16832 9096 16836
rect 9112 16892 9176 16896
rect 9112 16836 9116 16892
rect 9116 16836 9172 16892
rect 9172 16836 9176 16892
rect 9112 16832 9176 16836
rect 9192 16892 9256 16896
rect 9192 16836 9196 16892
rect 9196 16836 9252 16892
rect 9252 16836 9256 16892
rect 9192 16832 9256 16836
rect 16952 16892 17016 16896
rect 16952 16836 16956 16892
rect 16956 16836 17012 16892
rect 17012 16836 17016 16892
rect 16952 16832 17016 16836
rect 17032 16892 17096 16896
rect 17032 16836 17036 16892
rect 17036 16836 17092 16892
rect 17092 16836 17096 16892
rect 17032 16832 17096 16836
rect 17112 16892 17176 16896
rect 17112 16836 17116 16892
rect 17116 16836 17172 16892
rect 17172 16836 17176 16892
rect 17112 16832 17176 16836
rect 17192 16892 17256 16896
rect 17192 16836 17196 16892
rect 17196 16836 17252 16892
rect 17252 16836 17256 16892
rect 17192 16832 17256 16836
rect 4952 16348 5016 16352
rect 4952 16292 4956 16348
rect 4956 16292 5012 16348
rect 5012 16292 5016 16348
rect 4952 16288 5016 16292
rect 5032 16348 5096 16352
rect 5032 16292 5036 16348
rect 5036 16292 5092 16348
rect 5092 16292 5096 16348
rect 5032 16288 5096 16292
rect 5112 16348 5176 16352
rect 5112 16292 5116 16348
rect 5116 16292 5172 16348
rect 5172 16292 5176 16348
rect 5112 16288 5176 16292
rect 5192 16348 5256 16352
rect 5192 16292 5196 16348
rect 5196 16292 5252 16348
rect 5252 16292 5256 16348
rect 5192 16288 5256 16292
rect 12952 16348 13016 16352
rect 12952 16292 12956 16348
rect 12956 16292 13012 16348
rect 13012 16292 13016 16348
rect 12952 16288 13016 16292
rect 13032 16348 13096 16352
rect 13032 16292 13036 16348
rect 13036 16292 13092 16348
rect 13092 16292 13096 16348
rect 13032 16288 13096 16292
rect 13112 16348 13176 16352
rect 13112 16292 13116 16348
rect 13116 16292 13172 16348
rect 13172 16292 13176 16348
rect 13112 16288 13176 16292
rect 13192 16348 13256 16352
rect 13192 16292 13196 16348
rect 13196 16292 13252 16348
rect 13252 16292 13256 16348
rect 13192 16288 13256 16292
rect 20952 16348 21016 16352
rect 20952 16292 20956 16348
rect 20956 16292 21012 16348
rect 21012 16292 21016 16348
rect 20952 16288 21016 16292
rect 21032 16348 21096 16352
rect 21032 16292 21036 16348
rect 21036 16292 21092 16348
rect 21092 16292 21096 16348
rect 21032 16288 21096 16292
rect 21112 16348 21176 16352
rect 21112 16292 21116 16348
rect 21116 16292 21172 16348
rect 21172 16292 21176 16348
rect 21112 16288 21176 16292
rect 21192 16348 21256 16352
rect 21192 16292 21196 16348
rect 21196 16292 21252 16348
rect 21252 16292 21256 16348
rect 21192 16288 21256 16292
rect 8952 15804 9016 15808
rect 8952 15748 8956 15804
rect 8956 15748 9012 15804
rect 9012 15748 9016 15804
rect 8952 15744 9016 15748
rect 9032 15804 9096 15808
rect 9032 15748 9036 15804
rect 9036 15748 9092 15804
rect 9092 15748 9096 15804
rect 9032 15744 9096 15748
rect 9112 15804 9176 15808
rect 9112 15748 9116 15804
rect 9116 15748 9172 15804
rect 9172 15748 9176 15804
rect 9112 15744 9176 15748
rect 9192 15804 9256 15808
rect 9192 15748 9196 15804
rect 9196 15748 9252 15804
rect 9252 15748 9256 15804
rect 9192 15744 9256 15748
rect 16952 15804 17016 15808
rect 16952 15748 16956 15804
rect 16956 15748 17012 15804
rect 17012 15748 17016 15804
rect 16952 15744 17016 15748
rect 17032 15804 17096 15808
rect 17032 15748 17036 15804
rect 17036 15748 17092 15804
rect 17092 15748 17096 15804
rect 17032 15744 17096 15748
rect 17112 15804 17176 15808
rect 17112 15748 17116 15804
rect 17116 15748 17172 15804
rect 17172 15748 17176 15804
rect 17112 15744 17176 15748
rect 17192 15804 17256 15808
rect 17192 15748 17196 15804
rect 17196 15748 17252 15804
rect 17252 15748 17256 15804
rect 17192 15744 17256 15748
rect 4952 15260 5016 15264
rect 4952 15204 4956 15260
rect 4956 15204 5012 15260
rect 5012 15204 5016 15260
rect 4952 15200 5016 15204
rect 5032 15260 5096 15264
rect 5032 15204 5036 15260
rect 5036 15204 5092 15260
rect 5092 15204 5096 15260
rect 5032 15200 5096 15204
rect 5112 15260 5176 15264
rect 5112 15204 5116 15260
rect 5116 15204 5172 15260
rect 5172 15204 5176 15260
rect 5112 15200 5176 15204
rect 5192 15260 5256 15264
rect 5192 15204 5196 15260
rect 5196 15204 5252 15260
rect 5252 15204 5256 15260
rect 5192 15200 5256 15204
rect 12952 15260 13016 15264
rect 12952 15204 12956 15260
rect 12956 15204 13012 15260
rect 13012 15204 13016 15260
rect 12952 15200 13016 15204
rect 13032 15260 13096 15264
rect 13032 15204 13036 15260
rect 13036 15204 13092 15260
rect 13092 15204 13096 15260
rect 13032 15200 13096 15204
rect 13112 15260 13176 15264
rect 13112 15204 13116 15260
rect 13116 15204 13172 15260
rect 13172 15204 13176 15260
rect 13112 15200 13176 15204
rect 13192 15260 13256 15264
rect 13192 15204 13196 15260
rect 13196 15204 13252 15260
rect 13252 15204 13256 15260
rect 13192 15200 13256 15204
rect 20952 15260 21016 15264
rect 20952 15204 20956 15260
rect 20956 15204 21012 15260
rect 21012 15204 21016 15260
rect 20952 15200 21016 15204
rect 21032 15260 21096 15264
rect 21032 15204 21036 15260
rect 21036 15204 21092 15260
rect 21092 15204 21096 15260
rect 21032 15200 21096 15204
rect 21112 15260 21176 15264
rect 21112 15204 21116 15260
rect 21116 15204 21172 15260
rect 21172 15204 21176 15260
rect 21112 15200 21176 15204
rect 21192 15260 21256 15264
rect 21192 15204 21196 15260
rect 21196 15204 21252 15260
rect 21252 15204 21256 15260
rect 21192 15200 21256 15204
rect 8952 14716 9016 14720
rect 8952 14660 8956 14716
rect 8956 14660 9012 14716
rect 9012 14660 9016 14716
rect 8952 14656 9016 14660
rect 9032 14716 9096 14720
rect 9032 14660 9036 14716
rect 9036 14660 9092 14716
rect 9092 14660 9096 14716
rect 9032 14656 9096 14660
rect 9112 14716 9176 14720
rect 9112 14660 9116 14716
rect 9116 14660 9172 14716
rect 9172 14660 9176 14716
rect 9112 14656 9176 14660
rect 9192 14716 9256 14720
rect 9192 14660 9196 14716
rect 9196 14660 9252 14716
rect 9252 14660 9256 14716
rect 9192 14656 9256 14660
rect 16952 14716 17016 14720
rect 16952 14660 16956 14716
rect 16956 14660 17012 14716
rect 17012 14660 17016 14716
rect 16952 14656 17016 14660
rect 17032 14716 17096 14720
rect 17032 14660 17036 14716
rect 17036 14660 17092 14716
rect 17092 14660 17096 14716
rect 17032 14656 17096 14660
rect 17112 14716 17176 14720
rect 17112 14660 17116 14716
rect 17116 14660 17172 14716
rect 17172 14660 17176 14716
rect 17112 14656 17176 14660
rect 17192 14716 17256 14720
rect 17192 14660 17196 14716
rect 17196 14660 17252 14716
rect 17252 14660 17256 14716
rect 17192 14656 17256 14660
rect 4952 14172 5016 14176
rect 4952 14116 4956 14172
rect 4956 14116 5012 14172
rect 5012 14116 5016 14172
rect 4952 14112 5016 14116
rect 5032 14172 5096 14176
rect 5032 14116 5036 14172
rect 5036 14116 5092 14172
rect 5092 14116 5096 14172
rect 5032 14112 5096 14116
rect 5112 14172 5176 14176
rect 5112 14116 5116 14172
rect 5116 14116 5172 14172
rect 5172 14116 5176 14172
rect 5112 14112 5176 14116
rect 5192 14172 5256 14176
rect 5192 14116 5196 14172
rect 5196 14116 5252 14172
rect 5252 14116 5256 14172
rect 5192 14112 5256 14116
rect 12952 14172 13016 14176
rect 12952 14116 12956 14172
rect 12956 14116 13012 14172
rect 13012 14116 13016 14172
rect 12952 14112 13016 14116
rect 13032 14172 13096 14176
rect 13032 14116 13036 14172
rect 13036 14116 13092 14172
rect 13092 14116 13096 14172
rect 13032 14112 13096 14116
rect 13112 14172 13176 14176
rect 13112 14116 13116 14172
rect 13116 14116 13172 14172
rect 13172 14116 13176 14172
rect 13112 14112 13176 14116
rect 13192 14172 13256 14176
rect 13192 14116 13196 14172
rect 13196 14116 13252 14172
rect 13252 14116 13256 14172
rect 13192 14112 13256 14116
rect 20952 14172 21016 14176
rect 20952 14116 20956 14172
rect 20956 14116 21012 14172
rect 21012 14116 21016 14172
rect 20952 14112 21016 14116
rect 21032 14172 21096 14176
rect 21032 14116 21036 14172
rect 21036 14116 21092 14172
rect 21092 14116 21096 14172
rect 21032 14112 21096 14116
rect 21112 14172 21176 14176
rect 21112 14116 21116 14172
rect 21116 14116 21172 14172
rect 21172 14116 21176 14172
rect 21112 14112 21176 14116
rect 21192 14172 21256 14176
rect 21192 14116 21196 14172
rect 21196 14116 21252 14172
rect 21252 14116 21256 14172
rect 21192 14112 21256 14116
rect 8952 13628 9016 13632
rect 8952 13572 8956 13628
rect 8956 13572 9012 13628
rect 9012 13572 9016 13628
rect 8952 13568 9016 13572
rect 9032 13628 9096 13632
rect 9032 13572 9036 13628
rect 9036 13572 9092 13628
rect 9092 13572 9096 13628
rect 9032 13568 9096 13572
rect 9112 13628 9176 13632
rect 9112 13572 9116 13628
rect 9116 13572 9172 13628
rect 9172 13572 9176 13628
rect 9112 13568 9176 13572
rect 9192 13628 9256 13632
rect 9192 13572 9196 13628
rect 9196 13572 9252 13628
rect 9252 13572 9256 13628
rect 9192 13568 9256 13572
rect 16952 13628 17016 13632
rect 16952 13572 16956 13628
rect 16956 13572 17012 13628
rect 17012 13572 17016 13628
rect 16952 13568 17016 13572
rect 17032 13628 17096 13632
rect 17032 13572 17036 13628
rect 17036 13572 17092 13628
rect 17092 13572 17096 13628
rect 17032 13568 17096 13572
rect 17112 13628 17176 13632
rect 17112 13572 17116 13628
rect 17116 13572 17172 13628
rect 17172 13572 17176 13628
rect 17112 13568 17176 13572
rect 17192 13628 17256 13632
rect 17192 13572 17196 13628
rect 17196 13572 17252 13628
rect 17252 13572 17256 13628
rect 17192 13568 17256 13572
rect 4952 13084 5016 13088
rect 4952 13028 4956 13084
rect 4956 13028 5012 13084
rect 5012 13028 5016 13084
rect 4952 13024 5016 13028
rect 5032 13084 5096 13088
rect 5032 13028 5036 13084
rect 5036 13028 5092 13084
rect 5092 13028 5096 13084
rect 5032 13024 5096 13028
rect 5112 13084 5176 13088
rect 5112 13028 5116 13084
rect 5116 13028 5172 13084
rect 5172 13028 5176 13084
rect 5112 13024 5176 13028
rect 5192 13084 5256 13088
rect 5192 13028 5196 13084
rect 5196 13028 5252 13084
rect 5252 13028 5256 13084
rect 5192 13024 5256 13028
rect 12952 13084 13016 13088
rect 12952 13028 12956 13084
rect 12956 13028 13012 13084
rect 13012 13028 13016 13084
rect 12952 13024 13016 13028
rect 13032 13084 13096 13088
rect 13032 13028 13036 13084
rect 13036 13028 13092 13084
rect 13092 13028 13096 13084
rect 13032 13024 13096 13028
rect 13112 13084 13176 13088
rect 13112 13028 13116 13084
rect 13116 13028 13172 13084
rect 13172 13028 13176 13084
rect 13112 13024 13176 13028
rect 13192 13084 13256 13088
rect 13192 13028 13196 13084
rect 13196 13028 13252 13084
rect 13252 13028 13256 13084
rect 13192 13024 13256 13028
rect 20952 13084 21016 13088
rect 20952 13028 20956 13084
rect 20956 13028 21012 13084
rect 21012 13028 21016 13084
rect 20952 13024 21016 13028
rect 21032 13084 21096 13088
rect 21032 13028 21036 13084
rect 21036 13028 21092 13084
rect 21092 13028 21096 13084
rect 21032 13024 21096 13028
rect 21112 13084 21176 13088
rect 21112 13028 21116 13084
rect 21116 13028 21172 13084
rect 21172 13028 21176 13084
rect 21112 13024 21176 13028
rect 21192 13084 21256 13088
rect 21192 13028 21196 13084
rect 21196 13028 21252 13084
rect 21252 13028 21256 13084
rect 21192 13024 21256 13028
rect 8952 12540 9016 12544
rect 8952 12484 8956 12540
rect 8956 12484 9012 12540
rect 9012 12484 9016 12540
rect 8952 12480 9016 12484
rect 9032 12540 9096 12544
rect 9032 12484 9036 12540
rect 9036 12484 9092 12540
rect 9092 12484 9096 12540
rect 9032 12480 9096 12484
rect 9112 12540 9176 12544
rect 9112 12484 9116 12540
rect 9116 12484 9172 12540
rect 9172 12484 9176 12540
rect 9112 12480 9176 12484
rect 9192 12540 9256 12544
rect 9192 12484 9196 12540
rect 9196 12484 9252 12540
rect 9252 12484 9256 12540
rect 9192 12480 9256 12484
rect 16952 12540 17016 12544
rect 16952 12484 16956 12540
rect 16956 12484 17012 12540
rect 17012 12484 17016 12540
rect 16952 12480 17016 12484
rect 17032 12540 17096 12544
rect 17032 12484 17036 12540
rect 17036 12484 17092 12540
rect 17092 12484 17096 12540
rect 17032 12480 17096 12484
rect 17112 12540 17176 12544
rect 17112 12484 17116 12540
rect 17116 12484 17172 12540
rect 17172 12484 17176 12540
rect 17112 12480 17176 12484
rect 17192 12540 17256 12544
rect 17192 12484 17196 12540
rect 17196 12484 17252 12540
rect 17252 12484 17256 12540
rect 17192 12480 17256 12484
rect 4952 11996 5016 12000
rect 4952 11940 4956 11996
rect 4956 11940 5012 11996
rect 5012 11940 5016 11996
rect 4952 11936 5016 11940
rect 5032 11996 5096 12000
rect 5032 11940 5036 11996
rect 5036 11940 5092 11996
rect 5092 11940 5096 11996
rect 5032 11936 5096 11940
rect 5112 11996 5176 12000
rect 5112 11940 5116 11996
rect 5116 11940 5172 11996
rect 5172 11940 5176 11996
rect 5112 11936 5176 11940
rect 5192 11996 5256 12000
rect 5192 11940 5196 11996
rect 5196 11940 5252 11996
rect 5252 11940 5256 11996
rect 5192 11936 5256 11940
rect 12952 11996 13016 12000
rect 12952 11940 12956 11996
rect 12956 11940 13012 11996
rect 13012 11940 13016 11996
rect 12952 11936 13016 11940
rect 13032 11996 13096 12000
rect 13032 11940 13036 11996
rect 13036 11940 13092 11996
rect 13092 11940 13096 11996
rect 13032 11936 13096 11940
rect 13112 11996 13176 12000
rect 13112 11940 13116 11996
rect 13116 11940 13172 11996
rect 13172 11940 13176 11996
rect 13112 11936 13176 11940
rect 13192 11996 13256 12000
rect 13192 11940 13196 11996
rect 13196 11940 13252 11996
rect 13252 11940 13256 11996
rect 13192 11936 13256 11940
rect 20952 11996 21016 12000
rect 20952 11940 20956 11996
rect 20956 11940 21012 11996
rect 21012 11940 21016 11996
rect 20952 11936 21016 11940
rect 21032 11996 21096 12000
rect 21032 11940 21036 11996
rect 21036 11940 21092 11996
rect 21092 11940 21096 11996
rect 21032 11936 21096 11940
rect 21112 11996 21176 12000
rect 21112 11940 21116 11996
rect 21116 11940 21172 11996
rect 21172 11940 21176 11996
rect 21112 11936 21176 11940
rect 21192 11996 21256 12000
rect 21192 11940 21196 11996
rect 21196 11940 21252 11996
rect 21252 11940 21256 11996
rect 21192 11936 21256 11940
rect 8952 11452 9016 11456
rect 8952 11396 8956 11452
rect 8956 11396 9012 11452
rect 9012 11396 9016 11452
rect 8952 11392 9016 11396
rect 9032 11452 9096 11456
rect 9032 11396 9036 11452
rect 9036 11396 9092 11452
rect 9092 11396 9096 11452
rect 9032 11392 9096 11396
rect 9112 11452 9176 11456
rect 9112 11396 9116 11452
rect 9116 11396 9172 11452
rect 9172 11396 9176 11452
rect 9112 11392 9176 11396
rect 9192 11452 9256 11456
rect 9192 11396 9196 11452
rect 9196 11396 9252 11452
rect 9252 11396 9256 11452
rect 9192 11392 9256 11396
rect 16952 11452 17016 11456
rect 16952 11396 16956 11452
rect 16956 11396 17012 11452
rect 17012 11396 17016 11452
rect 16952 11392 17016 11396
rect 17032 11452 17096 11456
rect 17032 11396 17036 11452
rect 17036 11396 17092 11452
rect 17092 11396 17096 11452
rect 17032 11392 17096 11396
rect 17112 11452 17176 11456
rect 17112 11396 17116 11452
rect 17116 11396 17172 11452
rect 17172 11396 17176 11452
rect 17112 11392 17176 11396
rect 17192 11452 17256 11456
rect 17192 11396 17196 11452
rect 17196 11396 17252 11452
rect 17252 11396 17256 11452
rect 17192 11392 17256 11396
rect 4952 10908 5016 10912
rect 4952 10852 4956 10908
rect 4956 10852 5012 10908
rect 5012 10852 5016 10908
rect 4952 10848 5016 10852
rect 5032 10908 5096 10912
rect 5032 10852 5036 10908
rect 5036 10852 5092 10908
rect 5092 10852 5096 10908
rect 5032 10848 5096 10852
rect 5112 10908 5176 10912
rect 5112 10852 5116 10908
rect 5116 10852 5172 10908
rect 5172 10852 5176 10908
rect 5112 10848 5176 10852
rect 5192 10908 5256 10912
rect 5192 10852 5196 10908
rect 5196 10852 5252 10908
rect 5252 10852 5256 10908
rect 5192 10848 5256 10852
rect 12952 10908 13016 10912
rect 12952 10852 12956 10908
rect 12956 10852 13012 10908
rect 13012 10852 13016 10908
rect 12952 10848 13016 10852
rect 13032 10908 13096 10912
rect 13032 10852 13036 10908
rect 13036 10852 13092 10908
rect 13092 10852 13096 10908
rect 13032 10848 13096 10852
rect 13112 10908 13176 10912
rect 13112 10852 13116 10908
rect 13116 10852 13172 10908
rect 13172 10852 13176 10908
rect 13112 10848 13176 10852
rect 13192 10908 13256 10912
rect 13192 10852 13196 10908
rect 13196 10852 13252 10908
rect 13252 10852 13256 10908
rect 13192 10848 13256 10852
rect 20952 10908 21016 10912
rect 20952 10852 20956 10908
rect 20956 10852 21012 10908
rect 21012 10852 21016 10908
rect 20952 10848 21016 10852
rect 21032 10908 21096 10912
rect 21032 10852 21036 10908
rect 21036 10852 21092 10908
rect 21092 10852 21096 10908
rect 21032 10848 21096 10852
rect 21112 10908 21176 10912
rect 21112 10852 21116 10908
rect 21116 10852 21172 10908
rect 21172 10852 21176 10908
rect 21112 10848 21176 10852
rect 21192 10908 21256 10912
rect 21192 10852 21196 10908
rect 21196 10852 21252 10908
rect 21252 10852 21256 10908
rect 21192 10848 21256 10852
rect 8952 10364 9016 10368
rect 8952 10308 8956 10364
rect 8956 10308 9012 10364
rect 9012 10308 9016 10364
rect 8952 10304 9016 10308
rect 9032 10364 9096 10368
rect 9032 10308 9036 10364
rect 9036 10308 9092 10364
rect 9092 10308 9096 10364
rect 9032 10304 9096 10308
rect 9112 10364 9176 10368
rect 9112 10308 9116 10364
rect 9116 10308 9172 10364
rect 9172 10308 9176 10364
rect 9112 10304 9176 10308
rect 9192 10364 9256 10368
rect 9192 10308 9196 10364
rect 9196 10308 9252 10364
rect 9252 10308 9256 10364
rect 9192 10304 9256 10308
rect 16952 10364 17016 10368
rect 16952 10308 16956 10364
rect 16956 10308 17012 10364
rect 17012 10308 17016 10364
rect 16952 10304 17016 10308
rect 17032 10364 17096 10368
rect 17032 10308 17036 10364
rect 17036 10308 17092 10364
rect 17092 10308 17096 10364
rect 17032 10304 17096 10308
rect 17112 10364 17176 10368
rect 17112 10308 17116 10364
rect 17116 10308 17172 10364
rect 17172 10308 17176 10364
rect 17112 10304 17176 10308
rect 17192 10364 17256 10368
rect 17192 10308 17196 10364
rect 17196 10308 17252 10364
rect 17252 10308 17256 10364
rect 17192 10304 17256 10308
rect 4952 9820 5016 9824
rect 4952 9764 4956 9820
rect 4956 9764 5012 9820
rect 5012 9764 5016 9820
rect 4952 9760 5016 9764
rect 5032 9820 5096 9824
rect 5032 9764 5036 9820
rect 5036 9764 5092 9820
rect 5092 9764 5096 9820
rect 5032 9760 5096 9764
rect 5112 9820 5176 9824
rect 5112 9764 5116 9820
rect 5116 9764 5172 9820
rect 5172 9764 5176 9820
rect 5112 9760 5176 9764
rect 5192 9820 5256 9824
rect 5192 9764 5196 9820
rect 5196 9764 5252 9820
rect 5252 9764 5256 9820
rect 5192 9760 5256 9764
rect 12952 9820 13016 9824
rect 12952 9764 12956 9820
rect 12956 9764 13012 9820
rect 13012 9764 13016 9820
rect 12952 9760 13016 9764
rect 13032 9820 13096 9824
rect 13032 9764 13036 9820
rect 13036 9764 13092 9820
rect 13092 9764 13096 9820
rect 13032 9760 13096 9764
rect 13112 9820 13176 9824
rect 13112 9764 13116 9820
rect 13116 9764 13172 9820
rect 13172 9764 13176 9820
rect 13112 9760 13176 9764
rect 13192 9820 13256 9824
rect 13192 9764 13196 9820
rect 13196 9764 13252 9820
rect 13252 9764 13256 9820
rect 13192 9760 13256 9764
rect 20952 9820 21016 9824
rect 20952 9764 20956 9820
rect 20956 9764 21012 9820
rect 21012 9764 21016 9820
rect 20952 9760 21016 9764
rect 21032 9820 21096 9824
rect 21032 9764 21036 9820
rect 21036 9764 21092 9820
rect 21092 9764 21096 9820
rect 21032 9760 21096 9764
rect 21112 9820 21176 9824
rect 21112 9764 21116 9820
rect 21116 9764 21172 9820
rect 21172 9764 21176 9820
rect 21112 9760 21176 9764
rect 21192 9820 21256 9824
rect 21192 9764 21196 9820
rect 21196 9764 21252 9820
rect 21252 9764 21256 9820
rect 21192 9760 21256 9764
rect 8952 9276 9016 9280
rect 8952 9220 8956 9276
rect 8956 9220 9012 9276
rect 9012 9220 9016 9276
rect 8952 9216 9016 9220
rect 9032 9276 9096 9280
rect 9032 9220 9036 9276
rect 9036 9220 9092 9276
rect 9092 9220 9096 9276
rect 9032 9216 9096 9220
rect 9112 9276 9176 9280
rect 9112 9220 9116 9276
rect 9116 9220 9172 9276
rect 9172 9220 9176 9276
rect 9112 9216 9176 9220
rect 9192 9276 9256 9280
rect 9192 9220 9196 9276
rect 9196 9220 9252 9276
rect 9252 9220 9256 9276
rect 9192 9216 9256 9220
rect 16952 9276 17016 9280
rect 16952 9220 16956 9276
rect 16956 9220 17012 9276
rect 17012 9220 17016 9276
rect 16952 9216 17016 9220
rect 17032 9276 17096 9280
rect 17032 9220 17036 9276
rect 17036 9220 17092 9276
rect 17092 9220 17096 9276
rect 17032 9216 17096 9220
rect 17112 9276 17176 9280
rect 17112 9220 17116 9276
rect 17116 9220 17172 9276
rect 17172 9220 17176 9276
rect 17112 9216 17176 9220
rect 17192 9276 17256 9280
rect 17192 9220 17196 9276
rect 17196 9220 17252 9276
rect 17252 9220 17256 9276
rect 17192 9216 17256 9220
rect 4952 8732 5016 8736
rect 4952 8676 4956 8732
rect 4956 8676 5012 8732
rect 5012 8676 5016 8732
rect 4952 8672 5016 8676
rect 5032 8732 5096 8736
rect 5032 8676 5036 8732
rect 5036 8676 5092 8732
rect 5092 8676 5096 8732
rect 5032 8672 5096 8676
rect 5112 8732 5176 8736
rect 5112 8676 5116 8732
rect 5116 8676 5172 8732
rect 5172 8676 5176 8732
rect 5112 8672 5176 8676
rect 5192 8732 5256 8736
rect 5192 8676 5196 8732
rect 5196 8676 5252 8732
rect 5252 8676 5256 8732
rect 5192 8672 5256 8676
rect 12952 8732 13016 8736
rect 12952 8676 12956 8732
rect 12956 8676 13012 8732
rect 13012 8676 13016 8732
rect 12952 8672 13016 8676
rect 13032 8732 13096 8736
rect 13032 8676 13036 8732
rect 13036 8676 13092 8732
rect 13092 8676 13096 8732
rect 13032 8672 13096 8676
rect 13112 8732 13176 8736
rect 13112 8676 13116 8732
rect 13116 8676 13172 8732
rect 13172 8676 13176 8732
rect 13112 8672 13176 8676
rect 13192 8732 13256 8736
rect 13192 8676 13196 8732
rect 13196 8676 13252 8732
rect 13252 8676 13256 8732
rect 13192 8672 13256 8676
rect 20952 8732 21016 8736
rect 20952 8676 20956 8732
rect 20956 8676 21012 8732
rect 21012 8676 21016 8732
rect 20952 8672 21016 8676
rect 21032 8732 21096 8736
rect 21032 8676 21036 8732
rect 21036 8676 21092 8732
rect 21092 8676 21096 8732
rect 21032 8672 21096 8676
rect 21112 8732 21176 8736
rect 21112 8676 21116 8732
rect 21116 8676 21172 8732
rect 21172 8676 21176 8732
rect 21112 8672 21176 8676
rect 21192 8732 21256 8736
rect 21192 8676 21196 8732
rect 21196 8676 21252 8732
rect 21252 8676 21256 8732
rect 21192 8672 21256 8676
rect 8952 8188 9016 8192
rect 8952 8132 8956 8188
rect 8956 8132 9012 8188
rect 9012 8132 9016 8188
rect 8952 8128 9016 8132
rect 9032 8188 9096 8192
rect 9032 8132 9036 8188
rect 9036 8132 9092 8188
rect 9092 8132 9096 8188
rect 9032 8128 9096 8132
rect 9112 8188 9176 8192
rect 9112 8132 9116 8188
rect 9116 8132 9172 8188
rect 9172 8132 9176 8188
rect 9112 8128 9176 8132
rect 9192 8188 9256 8192
rect 9192 8132 9196 8188
rect 9196 8132 9252 8188
rect 9252 8132 9256 8188
rect 9192 8128 9256 8132
rect 16952 8188 17016 8192
rect 16952 8132 16956 8188
rect 16956 8132 17012 8188
rect 17012 8132 17016 8188
rect 16952 8128 17016 8132
rect 17032 8188 17096 8192
rect 17032 8132 17036 8188
rect 17036 8132 17092 8188
rect 17092 8132 17096 8188
rect 17032 8128 17096 8132
rect 17112 8188 17176 8192
rect 17112 8132 17116 8188
rect 17116 8132 17172 8188
rect 17172 8132 17176 8188
rect 17112 8128 17176 8132
rect 17192 8188 17256 8192
rect 17192 8132 17196 8188
rect 17196 8132 17252 8188
rect 17252 8132 17256 8188
rect 17192 8128 17256 8132
rect 4952 7644 5016 7648
rect 4952 7588 4956 7644
rect 4956 7588 5012 7644
rect 5012 7588 5016 7644
rect 4952 7584 5016 7588
rect 5032 7644 5096 7648
rect 5032 7588 5036 7644
rect 5036 7588 5092 7644
rect 5092 7588 5096 7644
rect 5032 7584 5096 7588
rect 5112 7644 5176 7648
rect 5112 7588 5116 7644
rect 5116 7588 5172 7644
rect 5172 7588 5176 7644
rect 5112 7584 5176 7588
rect 5192 7644 5256 7648
rect 5192 7588 5196 7644
rect 5196 7588 5252 7644
rect 5252 7588 5256 7644
rect 5192 7584 5256 7588
rect 12952 7644 13016 7648
rect 12952 7588 12956 7644
rect 12956 7588 13012 7644
rect 13012 7588 13016 7644
rect 12952 7584 13016 7588
rect 13032 7644 13096 7648
rect 13032 7588 13036 7644
rect 13036 7588 13092 7644
rect 13092 7588 13096 7644
rect 13032 7584 13096 7588
rect 13112 7644 13176 7648
rect 13112 7588 13116 7644
rect 13116 7588 13172 7644
rect 13172 7588 13176 7644
rect 13112 7584 13176 7588
rect 13192 7644 13256 7648
rect 13192 7588 13196 7644
rect 13196 7588 13252 7644
rect 13252 7588 13256 7644
rect 13192 7584 13256 7588
rect 20952 7644 21016 7648
rect 20952 7588 20956 7644
rect 20956 7588 21012 7644
rect 21012 7588 21016 7644
rect 20952 7584 21016 7588
rect 21032 7644 21096 7648
rect 21032 7588 21036 7644
rect 21036 7588 21092 7644
rect 21092 7588 21096 7644
rect 21032 7584 21096 7588
rect 21112 7644 21176 7648
rect 21112 7588 21116 7644
rect 21116 7588 21172 7644
rect 21172 7588 21176 7644
rect 21112 7584 21176 7588
rect 21192 7644 21256 7648
rect 21192 7588 21196 7644
rect 21196 7588 21252 7644
rect 21252 7588 21256 7644
rect 21192 7584 21256 7588
rect 8952 7100 9016 7104
rect 8952 7044 8956 7100
rect 8956 7044 9012 7100
rect 9012 7044 9016 7100
rect 8952 7040 9016 7044
rect 9032 7100 9096 7104
rect 9032 7044 9036 7100
rect 9036 7044 9092 7100
rect 9092 7044 9096 7100
rect 9032 7040 9096 7044
rect 9112 7100 9176 7104
rect 9112 7044 9116 7100
rect 9116 7044 9172 7100
rect 9172 7044 9176 7100
rect 9112 7040 9176 7044
rect 9192 7100 9256 7104
rect 9192 7044 9196 7100
rect 9196 7044 9252 7100
rect 9252 7044 9256 7100
rect 9192 7040 9256 7044
rect 16952 7100 17016 7104
rect 16952 7044 16956 7100
rect 16956 7044 17012 7100
rect 17012 7044 17016 7100
rect 16952 7040 17016 7044
rect 17032 7100 17096 7104
rect 17032 7044 17036 7100
rect 17036 7044 17092 7100
rect 17092 7044 17096 7100
rect 17032 7040 17096 7044
rect 17112 7100 17176 7104
rect 17112 7044 17116 7100
rect 17116 7044 17172 7100
rect 17172 7044 17176 7100
rect 17112 7040 17176 7044
rect 17192 7100 17256 7104
rect 17192 7044 17196 7100
rect 17196 7044 17252 7100
rect 17252 7044 17256 7100
rect 17192 7040 17256 7044
rect 4952 6556 5016 6560
rect 4952 6500 4956 6556
rect 4956 6500 5012 6556
rect 5012 6500 5016 6556
rect 4952 6496 5016 6500
rect 5032 6556 5096 6560
rect 5032 6500 5036 6556
rect 5036 6500 5092 6556
rect 5092 6500 5096 6556
rect 5032 6496 5096 6500
rect 5112 6556 5176 6560
rect 5112 6500 5116 6556
rect 5116 6500 5172 6556
rect 5172 6500 5176 6556
rect 5112 6496 5176 6500
rect 5192 6556 5256 6560
rect 5192 6500 5196 6556
rect 5196 6500 5252 6556
rect 5252 6500 5256 6556
rect 5192 6496 5256 6500
rect 12952 6556 13016 6560
rect 12952 6500 12956 6556
rect 12956 6500 13012 6556
rect 13012 6500 13016 6556
rect 12952 6496 13016 6500
rect 13032 6556 13096 6560
rect 13032 6500 13036 6556
rect 13036 6500 13092 6556
rect 13092 6500 13096 6556
rect 13032 6496 13096 6500
rect 13112 6556 13176 6560
rect 13112 6500 13116 6556
rect 13116 6500 13172 6556
rect 13172 6500 13176 6556
rect 13112 6496 13176 6500
rect 13192 6556 13256 6560
rect 13192 6500 13196 6556
rect 13196 6500 13252 6556
rect 13252 6500 13256 6556
rect 13192 6496 13256 6500
rect 20952 6556 21016 6560
rect 20952 6500 20956 6556
rect 20956 6500 21012 6556
rect 21012 6500 21016 6556
rect 20952 6496 21016 6500
rect 21032 6556 21096 6560
rect 21032 6500 21036 6556
rect 21036 6500 21092 6556
rect 21092 6500 21096 6556
rect 21032 6496 21096 6500
rect 21112 6556 21176 6560
rect 21112 6500 21116 6556
rect 21116 6500 21172 6556
rect 21172 6500 21176 6556
rect 21112 6496 21176 6500
rect 21192 6556 21256 6560
rect 21192 6500 21196 6556
rect 21196 6500 21252 6556
rect 21252 6500 21256 6556
rect 21192 6496 21256 6500
rect 8952 6012 9016 6016
rect 8952 5956 8956 6012
rect 8956 5956 9012 6012
rect 9012 5956 9016 6012
rect 8952 5952 9016 5956
rect 9032 6012 9096 6016
rect 9032 5956 9036 6012
rect 9036 5956 9092 6012
rect 9092 5956 9096 6012
rect 9032 5952 9096 5956
rect 9112 6012 9176 6016
rect 9112 5956 9116 6012
rect 9116 5956 9172 6012
rect 9172 5956 9176 6012
rect 9112 5952 9176 5956
rect 9192 6012 9256 6016
rect 9192 5956 9196 6012
rect 9196 5956 9252 6012
rect 9252 5956 9256 6012
rect 9192 5952 9256 5956
rect 16952 6012 17016 6016
rect 16952 5956 16956 6012
rect 16956 5956 17012 6012
rect 17012 5956 17016 6012
rect 16952 5952 17016 5956
rect 17032 6012 17096 6016
rect 17032 5956 17036 6012
rect 17036 5956 17092 6012
rect 17092 5956 17096 6012
rect 17032 5952 17096 5956
rect 17112 6012 17176 6016
rect 17112 5956 17116 6012
rect 17116 5956 17172 6012
rect 17172 5956 17176 6012
rect 17112 5952 17176 5956
rect 17192 6012 17256 6016
rect 17192 5956 17196 6012
rect 17196 5956 17252 6012
rect 17252 5956 17256 6012
rect 17192 5952 17256 5956
rect 4952 5468 5016 5472
rect 4952 5412 4956 5468
rect 4956 5412 5012 5468
rect 5012 5412 5016 5468
rect 4952 5408 5016 5412
rect 5032 5468 5096 5472
rect 5032 5412 5036 5468
rect 5036 5412 5092 5468
rect 5092 5412 5096 5468
rect 5032 5408 5096 5412
rect 5112 5468 5176 5472
rect 5112 5412 5116 5468
rect 5116 5412 5172 5468
rect 5172 5412 5176 5468
rect 5112 5408 5176 5412
rect 5192 5468 5256 5472
rect 5192 5412 5196 5468
rect 5196 5412 5252 5468
rect 5252 5412 5256 5468
rect 5192 5408 5256 5412
rect 12952 5468 13016 5472
rect 12952 5412 12956 5468
rect 12956 5412 13012 5468
rect 13012 5412 13016 5468
rect 12952 5408 13016 5412
rect 13032 5468 13096 5472
rect 13032 5412 13036 5468
rect 13036 5412 13092 5468
rect 13092 5412 13096 5468
rect 13032 5408 13096 5412
rect 13112 5468 13176 5472
rect 13112 5412 13116 5468
rect 13116 5412 13172 5468
rect 13172 5412 13176 5468
rect 13112 5408 13176 5412
rect 13192 5468 13256 5472
rect 13192 5412 13196 5468
rect 13196 5412 13252 5468
rect 13252 5412 13256 5468
rect 13192 5408 13256 5412
rect 20952 5468 21016 5472
rect 20952 5412 20956 5468
rect 20956 5412 21012 5468
rect 21012 5412 21016 5468
rect 20952 5408 21016 5412
rect 21032 5468 21096 5472
rect 21032 5412 21036 5468
rect 21036 5412 21092 5468
rect 21092 5412 21096 5468
rect 21032 5408 21096 5412
rect 21112 5468 21176 5472
rect 21112 5412 21116 5468
rect 21116 5412 21172 5468
rect 21172 5412 21176 5468
rect 21112 5408 21176 5412
rect 21192 5468 21256 5472
rect 21192 5412 21196 5468
rect 21196 5412 21252 5468
rect 21252 5412 21256 5468
rect 21192 5408 21256 5412
rect 8952 4924 9016 4928
rect 8952 4868 8956 4924
rect 8956 4868 9012 4924
rect 9012 4868 9016 4924
rect 8952 4864 9016 4868
rect 9032 4924 9096 4928
rect 9032 4868 9036 4924
rect 9036 4868 9092 4924
rect 9092 4868 9096 4924
rect 9032 4864 9096 4868
rect 9112 4924 9176 4928
rect 9112 4868 9116 4924
rect 9116 4868 9172 4924
rect 9172 4868 9176 4924
rect 9112 4864 9176 4868
rect 9192 4924 9256 4928
rect 9192 4868 9196 4924
rect 9196 4868 9252 4924
rect 9252 4868 9256 4924
rect 9192 4864 9256 4868
rect 16952 4924 17016 4928
rect 16952 4868 16956 4924
rect 16956 4868 17012 4924
rect 17012 4868 17016 4924
rect 16952 4864 17016 4868
rect 17032 4924 17096 4928
rect 17032 4868 17036 4924
rect 17036 4868 17092 4924
rect 17092 4868 17096 4924
rect 17032 4864 17096 4868
rect 17112 4924 17176 4928
rect 17112 4868 17116 4924
rect 17116 4868 17172 4924
rect 17172 4868 17176 4924
rect 17112 4864 17176 4868
rect 17192 4924 17256 4928
rect 17192 4868 17196 4924
rect 17196 4868 17252 4924
rect 17252 4868 17256 4924
rect 17192 4864 17256 4868
rect 4952 4380 5016 4384
rect 4952 4324 4956 4380
rect 4956 4324 5012 4380
rect 5012 4324 5016 4380
rect 4952 4320 5016 4324
rect 5032 4380 5096 4384
rect 5032 4324 5036 4380
rect 5036 4324 5092 4380
rect 5092 4324 5096 4380
rect 5032 4320 5096 4324
rect 5112 4380 5176 4384
rect 5112 4324 5116 4380
rect 5116 4324 5172 4380
rect 5172 4324 5176 4380
rect 5112 4320 5176 4324
rect 5192 4380 5256 4384
rect 5192 4324 5196 4380
rect 5196 4324 5252 4380
rect 5252 4324 5256 4380
rect 5192 4320 5256 4324
rect 12952 4380 13016 4384
rect 12952 4324 12956 4380
rect 12956 4324 13012 4380
rect 13012 4324 13016 4380
rect 12952 4320 13016 4324
rect 13032 4380 13096 4384
rect 13032 4324 13036 4380
rect 13036 4324 13092 4380
rect 13092 4324 13096 4380
rect 13032 4320 13096 4324
rect 13112 4380 13176 4384
rect 13112 4324 13116 4380
rect 13116 4324 13172 4380
rect 13172 4324 13176 4380
rect 13112 4320 13176 4324
rect 13192 4380 13256 4384
rect 13192 4324 13196 4380
rect 13196 4324 13252 4380
rect 13252 4324 13256 4380
rect 13192 4320 13256 4324
rect 20952 4380 21016 4384
rect 20952 4324 20956 4380
rect 20956 4324 21012 4380
rect 21012 4324 21016 4380
rect 20952 4320 21016 4324
rect 21032 4380 21096 4384
rect 21032 4324 21036 4380
rect 21036 4324 21092 4380
rect 21092 4324 21096 4380
rect 21032 4320 21096 4324
rect 21112 4380 21176 4384
rect 21112 4324 21116 4380
rect 21116 4324 21172 4380
rect 21172 4324 21176 4380
rect 21112 4320 21176 4324
rect 21192 4380 21256 4384
rect 21192 4324 21196 4380
rect 21196 4324 21252 4380
rect 21252 4324 21256 4380
rect 21192 4320 21256 4324
rect 8952 3836 9016 3840
rect 8952 3780 8956 3836
rect 8956 3780 9012 3836
rect 9012 3780 9016 3836
rect 8952 3776 9016 3780
rect 9032 3836 9096 3840
rect 9032 3780 9036 3836
rect 9036 3780 9092 3836
rect 9092 3780 9096 3836
rect 9032 3776 9096 3780
rect 9112 3836 9176 3840
rect 9112 3780 9116 3836
rect 9116 3780 9172 3836
rect 9172 3780 9176 3836
rect 9112 3776 9176 3780
rect 9192 3836 9256 3840
rect 9192 3780 9196 3836
rect 9196 3780 9252 3836
rect 9252 3780 9256 3836
rect 9192 3776 9256 3780
rect 16952 3836 17016 3840
rect 16952 3780 16956 3836
rect 16956 3780 17012 3836
rect 17012 3780 17016 3836
rect 16952 3776 17016 3780
rect 17032 3836 17096 3840
rect 17032 3780 17036 3836
rect 17036 3780 17092 3836
rect 17092 3780 17096 3836
rect 17032 3776 17096 3780
rect 17112 3836 17176 3840
rect 17112 3780 17116 3836
rect 17116 3780 17172 3836
rect 17172 3780 17176 3836
rect 17112 3776 17176 3780
rect 17192 3836 17256 3840
rect 17192 3780 17196 3836
rect 17196 3780 17252 3836
rect 17252 3780 17256 3836
rect 17192 3776 17256 3780
rect 60 3436 124 3500
rect 4952 3292 5016 3296
rect 4952 3236 4956 3292
rect 4956 3236 5012 3292
rect 5012 3236 5016 3292
rect 4952 3232 5016 3236
rect 5032 3292 5096 3296
rect 5032 3236 5036 3292
rect 5036 3236 5092 3292
rect 5092 3236 5096 3292
rect 5032 3232 5096 3236
rect 5112 3292 5176 3296
rect 5112 3236 5116 3292
rect 5116 3236 5172 3292
rect 5172 3236 5176 3292
rect 5112 3232 5176 3236
rect 5192 3292 5256 3296
rect 5192 3236 5196 3292
rect 5196 3236 5252 3292
rect 5252 3236 5256 3292
rect 5192 3232 5256 3236
rect 12952 3292 13016 3296
rect 12952 3236 12956 3292
rect 12956 3236 13012 3292
rect 13012 3236 13016 3292
rect 12952 3232 13016 3236
rect 13032 3292 13096 3296
rect 13032 3236 13036 3292
rect 13036 3236 13092 3292
rect 13092 3236 13096 3292
rect 13032 3232 13096 3236
rect 13112 3292 13176 3296
rect 13112 3236 13116 3292
rect 13116 3236 13172 3292
rect 13172 3236 13176 3292
rect 13112 3232 13176 3236
rect 13192 3292 13256 3296
rect 13192 3236 13196 3292
rect 13196 3236 13252 3292
rect 13252 3236 13256 3292
rect 13192 3232 13256 3236
rect 20952 3292 21016 3296
rect 20952 3236 20956 3292
rect 20956 3236 21012 3292
rect 21012 3236 21016 3292
rect 20952 3232 21016 3236
rect 21032 3292 21096 3296
rect 21032 3236 21036 3292
rect 21036 3236 21092 3292
rect 21092 3236 21096 3292
rect 21032 3232 21096 3236
rect 21112 3292 21176 3296
rect 21112 3236 21116 3292
rect 21116 3236 21172 3292
rect 21172 3236 21176 3292
rect 21112 3232 21176 3236
rect 21192 3292 21256 3296
rect 21192 3236 21196 3292
rect 21196 3236 21252 3292
rect 21252 3236 21256 3292
rect 21192 3232 21256 3236
rect 60 3164 124 3228
rect 8952 2748 9016 2752
rect 8952 2692 8956 2748
rect 8956 2692 9012 2748
rect 9012 2692 9016 2748
rect 8952 2688 9016 2692
rect 9032 2748 9096 2752
rect 9032 2692 9036 2748
rect 9036 2692 9092 2748
rect 9092 2692 9096 2748
rect 9032 2688 9096 2692
rect 9112 2748 9176 2752
rect 9112 2692 9116 2748
rect 9116 2692 9172 2748
rect 9172 2692 9176 2748
rect 9112 2688 9176 2692
rect 9192 2748 9256 2752
rect 9192 2692 9196 2748
rect 9196 2692 9252 2748
rect 9252 2692 9256 2748
rect 9192 2688 9256 2692
rect 16952 2748 17016 2752
rect 16952 2692 16956 2748
rect 16956 2692 17012 2748
rect 17012 2692 17016 2748
rect 16952 2688 17016 2692
rect 17032 2748 17096 2752
rect 17032 2692 17036 2748
rect 17036 2692 17092 2748
rect 17092 2692 17096 2748
rect 17032 2688 17096 2692
rect 17112 2748 17176 2752
rect 17112 2692 17116 2748
rect 17116 2692 17172 2748
rect 17172 2692 17176 2748
rect 17112 2688 17176 2692
rect 17192 2748 17256 2752
rect 17192 2692 17196 2748
rect 17196 2692 17252 2748
rect 17252 2692 17256 2748
rect 17192 2688 17256 2692
rect 4952 2204 5016 2208
rect 4952 2148 4956 2204
rect 4956 2148 5012 2204
rect 5012 2148 5016 2204
rect 4952 2144 5016 2148
rect 5032 2204 5096 2208
rect 5032 2148 5036 2204
rect 5036 2148 5092 2204
rect 5092 2148 5096 2204
rect 5032 2144 5096 2148
rect 5112 2204 5176 2208
rect 5112 2148 5116 2204
rect 5116 2148 5172 2204
rect 5172 2148 5176 2204
rect 5112 2144 5176 2148
rect 5192 2204 5256 2208
rect 5192 2148 5196 2204
rect 5196 2148 5252 2204
rect 5252 2148 5256 2204
rect 5192 2144 5256 2148
rect 12952 2204 13016 2208
rect 12952 2148 12956 2204
rect 12956 2148 13012 2204
rect 13012 2148 13016 2204
rect 12952 2144 13016 2148
rect 13032 2204 13096 2208
rect 13032 2148 13036 2204
rect 13036 2148 13092 2204
rect 13092 2148 13096 2204
rect 13032 2144 13096 2148
rect 13112 2204 13176 2208
rect 13112 2148 13116 2204
rect 13116 2148 13172 2204
rect 13172 2148 13176 2204
rect 13112 2144 13176 2148
rect 13192 2204 13256 2208
rect 13192 2148 13196 2204
rect 13196 2148 13252 2204
rect 13252 2148 13256 2204
rect 13192 2144 13256 2148
rect 20952 2204 21016 2208
rect 20952 2148 20956 2204
rect 20956 2148 21012 2204
rect 21012 2148 21016 2204
rect 20952 2144 21016 2148
rect 21032 2204 21096 2208
rect 21032 2148 21036 2204
rect 21036 2148 21092 2204
rect 21092 2148 21096 2204
rect 21032 2144 21096 2148
rect 21112 2204 21176 2208
rect 21112 2148 21116 2204
rect 21116 2148 21172 2204
rect 21172 2148 21176 2204
rect 21112 2144 21176 2148
rect 21192 2204 21256 2208
rect 21192 2148 21196 2204
rect 21196 2148 21252 2204
rect 21252 2148 21256 2204
rect 21192 2144 21256 2148
<< metal4 >>
rect 4944 21792 5264 21808
rect 4944 21728 4952 21792
rect 5016 21728 5032 21792
rect 5096 21728 5112 21792
rect 5176 21728 5192 21792
rect 5256 21728 5264 21792
rect 4944 20704 5264 21728
rect 4944 20640 4952 20704
rect 5016 20640 5032 20704
rect 5096 20640 5112 20704
rect 5176 20640 5192 20704
rect 5256 20640 5264 20704
rect 4944 19616 5264 20640
rect 4944 19552 4952 19616
rect 5016 19552 5032 19616
rect 5096 19552 5112 19616
rect 5176 19552 5192 19616
rect 5256 19552 5264 19616
rect 4944 18528 5264 19552
rect 4944 18464 4952 18528
rect 5016 18464 5032 18528
rect 5096 18464 5112 18528
rect 5176 18464 5192 18528
rect 5256 18464 5264 18528
rect 4944 17440 5264 18464
rect 4944 17376 4952 17440
rect 5016 17376 5032 17440
rect 5096 17376 5112 17440
rect 5176 17376 5192 17440
rect 5256 17376 5264 17440
rect 4944 16352 5264 17376
rect 4944 16288 4952 16352
rect 5016 16288 5032 16352
rect 5096 16288 5112 16352
rect 5176 16288 5192 16352
rect 5256 16288 5264 16352
rect 4944 15264 5264 16288
rect 4944 15200 4952 15264
rect 5016 15200 5032 15264
rect 5096 15200 5112 15264
rect 5176 15200 5192 15264
rect 5256 15200 5264 15264
rect 4944 14176 5264 15200
rect 4944 14112 4952 14176
rect 5016 14112 5032 14176
rect 5096 14112 5112 14176
rect 5176 14112 5192 14176
rect 5256 14112 5264 14176
rect 4944 13088 5264 14112
rect 4944 13024 4952 13088
rect 5016 13024 5032 13088
rect 5096 13024 5112 13088
rect 5176 13024 5192 13088
rect 5256 13024 5264 13088
rect 4944 12000 5264 13024
rect 4944 11936 4952 12000
rect 5016 11936 5032 12000
rect 5096 11936 5112 12000
rect 5176 11936 5192 12000
rect 5256 11936 5264 12000
rect 4944 10912 5264 11936
rect 4944 10848 4952 10912
rect 5016 10848 5032 10912
rect 5096 10848 5112 10912
rect 5176 10848 5192 10912
rect 5256 10848 5264 10912
rect 4944 9824 5264 10848
rect 4944 9760 4952 9824
rect 5016 9760 5032 9824
rect 5096 9760 5112 9824
rect 5176 9760 5192 9824
rect 5256 9760 5264 9824
rect 4944 8736 5264 9760
rect 4944 8672 4952 8736
rect 5016 8672 5032 8736
rect 5096 8672 5112 8736
rect 5176 8672 5192 8736
rect 5256 8672 5264 8736
rect 4944 7648 5264 8672
rect 4944 7584 4952 7648
rect 5016 7584 5032 7648
rect 5096 7584 5112 7648
rect 5176 7584 5192 7648
rect 5256 7584 5264 7648
rect 4944 6560 5264 7584
rect 4944 6496 4952 6560
rect 5016 6496 5032 6560
rect 5096 6496 5112 6560
rect 5176 6496 5192 6560
rect 5256 6496 5264 6560
rect 4944 5472 5264 6496
rect 4944 5408 4952 5472
rect 5016 5408 5032 5472
rect 5096 5408 5112 5472
rect 5176 5408 5192 5472
rect 5256 5408 5264 5472
rect 4944 4384 5264 5408
rect 4944 4320 4952 4384
rect 5016 4320 5032 4384
rect 5096 4320 5112 4384
rect 5176 4320 5192 4384
rect 5256 4320 5264 4384
rect 59 3500 125 3501
rect 59 3436 60 3500
rect 124 3436 125 3500
rect 59 3435 125 3436
rect 62 3229 122 3435
rect 4944 3296 5264 4320
rect 4944 3232 4952 3296
rect 5016 3232 5032 3296
rect 5096 3232 5112 3296
rect 5176 3232 5192 3296
rect 5256 3232 5264 3296
rect 59 3228 125 3229
rect 59 3164 60 3228
rect 124 3164 125 3228
rect 59 3163 125 3164
rect 4944 2208 5264 3232
rect 4944 2144 4952 2208
rect 5016 2144 5032 2208
rect 5096 2144 5112 2208
rect 5176 2144 5192 2208
rect 5256 2144 5264 2208
rect 4944 2128 5264 2144
rect 8944 21248 9264 21808
rect 8944 21184 8952 21248
rect 9016 21184 9032 21248
rect 9096 21184 9112 21248
rect 9176 21184 9192 21248
rect 9256 21184 9264 21248
rect 8944 20160 9264 21184
rect 8944 20096 8952 20160
rect 9016 20096 9032 20160
rect 9096 20096 9112 20160
rect 9176 20096 9192 20160
rect 9256 20096 9264 20160
rect 8944 19072 9264 20096
rect 8944 19008 8952 19072
rect 9016 19008 9032 19072
rect 9096 19008 9112 19072
rect 9176 19008 9192 19072
rect 9256 19008 9264 19072
rect 8944 17984 9264 19008
rect 8944 17920 8952 17984
rect 9016 17920 9032 17984
rect 9096 17920 9112 17984
rect 9176 17920 9192 17984
rect 9256 17920 9264 17984
rect 8944 16896 9264 17920
rect 8944 16832 8952 16896
rect 9016 16832 9032 16896
rect 9096 16832 9112 16896
rect 9176 16832 9192 16896
rect 9256 16832 9264 16896
rect 8944 15808 9264 16832
rect 8944 15744 8952 15808
rect 9016 15744 9032 15808
rect 9096 15744 9112 15808
rect 9176 15744 9192 15808
rect 9256 15744 9264 15808
rect 8944 14720 9264 15744
rect 8944 14656 8952 14720
rect 9016 14656 9032 14720
rect 9096 14656 9112 14720
rect 9176 14656 9192 14720
rect 9256 14656 9264 14720
rect 8944 13632 9264 14656
rect 8944 13568 8952 13632
rect 9016 13568 9032 13632
rect 9096 13568 9112 13632
rect 9176 13568 9192 13632
rect 9256 13568 9264 13632
rect 8944 12544 9264 13568
rect 8944 12480 8952 12544
rect 9016 12480 9032 12544
rect 9096 12480 9112 12544
rect 9176 12480 9192 12544
rect 9256 12480 9264 12544
rect 8944 11456 9264 12480
rect 8944 11392 8952 11456
rect 9016 11392 9032 11456
rect 9096 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9264 11456
rect 8944 10368 9264 11392
rect 8944 10304 8952 10368
rect 9016 10304 9032 10368
rect 9096 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9264 10368
rect 8944 9280 9264 10304
rect 8944 9216 8952 9280
rect 9016 9216 9032 9280
rect 9096 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9264 9280
rect 8944 8192 9264 9216
rect 8944 8128 8952 8192
rect 9016 8128 9032 8192
rect 9096 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9264 8192
rect 8944 7104 9264 8128
rect 8944 7040 8952 7104
rect 9016 7040 9032 7104
rect 9096 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9264 7104
rect 8944 6016 9264 7040
rect 8944 5952 8952 6016
rect 9016 5952 9032 6016
rect 9096 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9264 6016
rect 8944 4928 9264 5952
rect 8944 4864 8952 4928
rect 9016 4864 9032 4928
rect 9096 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9264 4928
rect 8944 3840 9264 4864
rect 8944 3776 8952 3840
rect 9016 3776 9032 3840
rect 9096 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9264 3840
rect 8944 2752 9264 3776
rect 8944 2688 8952 2752
rect 9016 2688 9032 2752
rect 9096 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9264 2752
rect 8944 2128 9264 2688
rect 12944 21792 13264 21808
rect 12944 21728 12952 21792
rect 13016 21728 13032 21792
rect 13096 21728 13112 21792
rect 13176 21728 13192 21792
rect 13256 21728 13264 21792
rect 12944 20704 13264 21728
rect 12944 20640 12952 20704
rect 13016 20640 13032 20704
rect 13096 20640 13112 20704
rect 13176 20640 13192 20704
rect 13256 20640 13264 20704
rect 12944 19616 13264 20640
rect 12944 19552 12952 19616
rect 13016 19552 13032 19616
rect 13096 19552 13112 19616
rect 13176 19552 13192 19616
rect 13256 19552 13264 19616
rect 12944 18528 13264 19552
rect 12944 18464 12952 18528
rect 13016 18464 13032 18528
rect 13096 18464 13112 18528
rect 13176 18464 13192 18528
rect 13256 18464 13264 18528
rect 12944 17440 13264 18464
rect 12944 17376 12952 17440
rect 13016 17376 13032 17440
rect 13096 17376 13112 17440
rect 13176 17376 13192 17440
rect 13256 17376 13264 17440
rect 12944 16352 13264 17376
rect 12944 16288 12952 16352
rect 13016 16288 13032 16352
rect 13096 16288 13112 16352
rect 13176 16288 13192 16352
rect 13256 16288 13264 16352
rect 12944 15264 13264 16288
rect 12944 15200 12952 15264
rect 13016 15200 13032 15264
rect 13096 15200 13112 15264
rect 13176 15200 13192 15264
rect 13256 15200 13264 15264
rect 12944 14176 13264 15200
rect 12944 14112 12952 14176
rect 13016 14112 13032 14176
rect 13096 14112 13112 14176
rect 13176 14112 13192 14176
rect 13256 14112 13264 14176
rect 12944 13088 13264 14112
rect 12944 13024 12952 13088
rect 13016 13024 13032 13088
rect 13096 13024 13112 13088
rect 13176 13024 13192 13088
rect 13256 13024 13264 13088
rect 12944 12000 13264 13024
rect 12944 11936 12952 12000
rect 13016 11936 13032 12000
rect 13096 11936 13112 12000
rect 13176 11936 13192 12000
rect 13256 11936 13264 12000
rect 12944 10912 13264 11936
rect 12944 10848 12952 10912
rect 13016 10848 13032 10912
rect 13096 10848 13112 10912
rect 13176 10848 13192 10912
rect 13256 10848 13264 10912
rect 12944 9824 13264 10848
rect 12944 9760 12952 9824
rect 13016 9760 13032 9824
rect 13096 9760 13112 9824
rect 13176 9760 13192 9824
rect 13256 9760 13264 9824
rect 12944 8736 13264 9760
rect 12944 8672 12952 8736
rect 13016 8672 13032 8736
rect 13096 8672 13112 8736
rect 13176 8672 13192 8736
rect 13256 8672 13264 8736
rect 12944 7648 13264 8672
rect 12944 7584 12952 7648
rect 13016 7584 13032 7648
rect 13096 7584 13112 7648
rect 13176 7584 13192 7648
rect 13256 7584 13264 7648
rect 12944 6560 13264 7584
rect 12944 6496 12952 6560
rect 13016 6496 13032 6560
rect 13096 6496 13112 6560
rect 13176 6496 13192 6560
rect 13256 6496 13264 6560
rect 12944 5472 13264 6496
rect 12944 5408 12952 5472
rect 13016 5408 13032 5472
rect 13096 5408 13112 5472
rect 13176 5408 13192 5472
rect 13256 5408 13264 5472
rect 12944 4384 13264 5408
rect 12944 4320 12952 4384
rect 13016 4320 13032 4384
rect 13096 4320 13112 4384
rect 13176 4320 13192 4384
rect 13256 4320 13264 4384
rect 12944 3296 13264 4320
rect 12944 3232 12952 3296
rect 13016 3232 13032 3296
rect 13096 3232 13112 3296
rect 13176 3232 13192 3296
rect 13256 3232 13264 3296
rect 12944 2208 13264 3232
rect 12944 2144 12952 2208
rect 13016 2144 13032 2208
rect 13096 2144 13112 2208
rect 13176 2144 13192 2208
rect 13256 2144 13264 2208
rect 12944 2128 13264 2144
rect 16944 21248 17264 21808
rect 16944 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17264 21248
rect 16944 20160 17264 21184
rect 16944 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17264 20160
rect 16944 19072 17264 20096
rect 16944 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17264 19072
rect 16944 17984 17264 19008
rect 16944 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17264 17984
rect 16944 16896 17264 17920
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 16944 15808 17264 16832
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 16944 14720 17264 15744
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 16944 13632 17264 14656
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 16944 12544 17264 13568
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 16944 11456 17264 12480
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 10368 17264 11392
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 16944 9280 17264 10304
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 16944 8192 17264 9216
rect 16944 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17264 8192
rect 16944 7104 17264 8128
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16944 6016 17264 7040
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 16944 4928 17264 5952
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 16944 3840 17264 4864
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16944 2752 17264 3776
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 16944 2128 17264 2688
rect 20944 21792 21264 21808
rect 20944 21728 20952 21792
rect 21016 21728 21032 21792
rect 21096 21728 21112 21792
rect 21176 21728 21192 21792
rect 21256 21728 21264 21792
rect 20944 20704 21264 21728
rect 20944 20640 20952 20704
rect 21016 20640 21032 20704
rect 21096 20640 21112 20704
rect 21176 20640 21192 20704
rect 21256 20640 21264 20704
rect 20944 19616 21264 20640
rect 20944 19552 20952 19616
rect 21016 19552 21032 19616
rect 21096 19552 21112 19616
rect 21176 19552 21192 19616
rect 21256 19552 21264 19616
rect 20944 18528 21264 19552
rect 20944 18464 20952 18528
rect 21016 18464 21032 18528
rect 21096 18464 21112 18528
rect 21176 18464 21192 18528
rect 21256 18464 21264 18528
rect 20944 17440 21264 18464
rect 20944 17376 20952 17440
rect 21016 17376 21032 17440
rect 21096 17376 21112 17440
rect 21176 17376 21192 17440
rect 21256 17376 21264 17440
rect 20944 16352 21264 17376
rect 20944 16288 20952 16352
rect 21016 16288 21032 16352
rect 21096 16288 21112 16352
rect 21176 16288 21192 16352
rect 21256 16288 21264 16352
rect 20944 15264 21264 16288
rect 20944 15200 20952 15264
rect 21016 15200 21032 15264
rect 21096 15200 21112 15264
rect 21176 15200 21192 15264
rect 21256 15200 21264 15264
rect 20944 14176 21264 15200
rect 20944 14112 20952 14176
rect 21016 14112 21032 14176
rect 21096 14112 21112 14176
rect 21176 14112 21192 14176
rect 21256 14112 21264 14176
rect 20944 13088 21264 14112
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 12000 21264 13024
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 10912 21264 11936
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 9824 21264 10848
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 8736 21264 9760
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 7648 21264 8672
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 6560 21264 7584
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 5472 21264 6496
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 4384 21264 5408
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 3296 21264 4320
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 2208 21264 3232
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2128 21264 2144
use scs8hd_decap_6  FILLER_1_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_7
timestamp 1586364061
transform 1 0 1748 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1564 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_buf_2  _144_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_16
timestamp 1586364061
transform 1 0 2576 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_13 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2300 0 1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_11 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2116 0 -1 2720
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2392 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__049__A
timestamp 1586364061
transform 1 0 2760 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _141_
timestamp 1586364061
transform 1 0 2852 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_34
timestamp 1586364061
transform 1 0 4232 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_29
timestamp 1586364061
transform 1 0 3772 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__B
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__A
timestamp 1586364061
transform 1 0 4232 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__A
timestamp 1586364061
transform 1 0 4048 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_72 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_8  _049_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2944 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__058__C
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_1_51
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_47
timestamp 1586364061
transform 1 0 5428 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_53
timestamp 1586364061
transform 1 0 5980 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_49
timestamp 1586364061
transform 1 0 5612 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_45
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__C
timestamp 1586364061
transform 1 0 5796 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__B
timestamp 1586364061
transform 1 0 5428 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__048__A
timestamp 1586364061
transform 1 0 5612 0 1 2720
box -38 -48 222 592
use scs8hd_or3_4  _058_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 866 592
use scs8hd_or3_4  _054_
timestamp 1586364061
transform 1 0 4416 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_59
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_66
timestamp 1586364061
transform 1 0 7176 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 6992 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 7452 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_5_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6992 0 -1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_80
timestamp 1586364061
transform 1 0 8464 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_79
timestamp 1586364061
transform 1 0 8372 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__B
timestamp 1586364061
transform 1 0 8188 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_84
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__C
timestamp 1586364061
transform 1 0 8648 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _136_
timestamp 1586364061
transform 1 0 9200 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_96
timestamp 1586364061
transform 1 0 9936 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_92 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9568 0 1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_99
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_105
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_109
timestamp 1586364061
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11316 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11500 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_138
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_134
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_138
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _148_
timestamp 1586364061
transform 1 0 14168 0 -1 2720
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_0_146
timestamp 1586364061
transform 1 0 14536 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_150
timestamp 1586364061
transform 1 0 14904 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 14720 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_153
timestamp 1586364061
transform 1 0 15180 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_157
timestamp 1586364061
transform 1 0 15548 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 15364 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_159
timestamp 1586364061
transform 1 0 15732 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_163
timestamp 1586364061
transform 1 0 16100 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15916 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_174
timestamp 1586364061
transform 1 0 17112 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_170
timestamp 1586364061
transform 1 0 16744 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_178
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 16928 0 1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 16468 0 -1 2720
box -38 -48 1050 592
use scs8hd_nor2_4  _095_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15916 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18308 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_191
timestamp 1586364061
transform 1 0 18676 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18768 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18952 0 -1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _091_
timestamp 1586364061
transform 1 0 20056 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 19872 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 20056 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19504 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_203
timestamp 1586364061
transform 1 0 19780 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_0_208
timestamp 1586364061
transform 1 0 20240 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_198
timestamp 1586364061
transform 1 0 19320 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_202
timestamp 1586364061
transform 1 0 19688 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_215
timestamp 1586364061
transform 1 0 20884 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_222
timestamp 1586364061
transform 1 0 21528 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_216
timestamp 1586364061
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21068 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _159_
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_231
timestamp 1586364061
transform 1 0 22356 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_226
timestamp 1586364061
transform 1 0 21896 0 -1 2720
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 21712 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_219 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 21252 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 22816 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 22816 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_232
timestamp 1586364061
transform 1 0 22448 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _143_
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 2392 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_7
timestamp 1586364061
transform 1 0 1748 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_13
timestamp 1586364061
transform 1 0 2300 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_16
timestamp 1586364061
transform 1 0 2576 0 -1 3808
box -38 -48 406 592
use scs8hd_inv_8  _048_
timestamp 1586364061
transform 1 0 4232 0 -1 3808
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__064__B
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__060__A
timestamp 1586364061
transform 1 0 5244 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_43
timestamp 1586364061
transform 1 0 5060 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_47
timestamp 1586364061
transform 1 0 5428 0 -1 3808
box -38 -48 774 592
use scs8hd_nor2_4  _106_
timestamp 1586364061
transform 1 0 6348 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_55
timestamp 1586364061
transform 1 0 6164 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_66
timestamp 1586364061
transform 1 0 7176 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_70
timestamp 1586364061
transform 1 0 7544 0 -1 3808
box -38 -48 130 592
use scs8hd_or3_4  _066_
timestamp 1586364061
transform 1 0 7912 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_73
timestamp 1586364061
transform 1 0 7820 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_83
timestamp 1586364061
transform 1 0 8740 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_87
timestamp 1586364061
transform 1 0 9108 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 9844 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_90
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_97
timestamp 1586364061
transform 1 0 10028 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_107
timestamp 1586364061
transform 1 0 10948 0 -1 3808
box -38 -48 314 592
use scs8hd_buf_2  _162_
timestamp 1586364061
transform 1 0 11776 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 11592 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_112
timestamp 1586364061
transform 1 0 11408 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_120
timestamp 1586364061
transform 1 0 12144 0 -1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12880 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13892 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_125
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_137
timestamp 1586364061
transform 1 0 13708 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_147
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 590 592
use scs8hd_buf_2  _140_
timestamp 1586364061
transform 1 0 17020 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_165
timestamp 1586364061
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_169
timestamp 1586364061
transform 1 0 16652 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_177
timestamp 1586364061
transform 1 0 17388 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 17572 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_181
timestamp 1586364061
transform 1 0 17756 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_186
timestamp 1586364061
transform 1 0 18216 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_198
timestamp 1586364061
transform 1 0 19320 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_205
timestamp 1586364061
transform 1 0 19964 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_213
timestamp 1586364061
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_218
timestamp 1586364061
transform 1 0 21160 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_2_230
timestamp 1586364061
transform 1 0 22264 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 22816 0 -1 3808
box -38 -48 314 592
use scs8hd_buf_2  _139_
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__062__C
timestamp 1586364061
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__B
timestamp 1586364061
transform 1 0 2024 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_12
timestamp 1586364061
transform 1 0 2208 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_16
timestamp 1586364061
transform 1 0 2576 0 1 3808
box -38 -48 406 592
use scs8hd_or3_4  _064_
timestamp 1586364061
transform 1 0 3220 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__047__A
timestamp 1586364061
transform 1 0 4232 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_20
timestamp 1586364061
transform 1 0 2944 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_32
timestamp 1586364061
transform 1 0 4048 0 1 3808
box -38 -48 222 592
use scs8hd_or3_4  _060_
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__060__B
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_36
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_49
timestamp 1586364061
transform 1 0 5612 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _142_
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 7360 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_66
timestamp 1586364061
transform 1 0 7176 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_70
timestamp 1586364061
transform 1 0 7544 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7728 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 9200 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 9752 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 9568 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_90
timestamp 1586364061
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_103
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_107
timestamp 1586364061
transform 1 0 10948 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 14076 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_136
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_140
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14444 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_143
timestamp 1586364061
transform 1 0 14260 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_154
timestamp 1586364061
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_158
timestamp 1586364061
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__092__B
timestamp 1586364061
transform 1 0 17020 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_175
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_195
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_199
timestamp 1586364061
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_212
timestamp 1586364061
transform 1 0 20608 0 1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21804 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_217
timestamp 1586364061
transform 1 0 21068 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_223
timestamp 1586364061
transform 1 0 21620 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_227
timestamp 1586364061
transform 1 0 21988 0 1 3808
box -38 -48 590 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 22816 0 1 3808
box -38 -48 314 592
use scs8hd_or3_4  _062_
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_7
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_13
timestamp 1586364061
transform 1 0 2300 0 -1 4896
box -38 -48 130 592
use scs8hd_inv_8  _047_
timestamp 1586364061
transform 1 0 4232 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__064__C
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _108_
timestamp 1586364061
transform 1 0 5796 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__060__C
timestamp 1586364061
transform 1 0 5244 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_43
timestamp 1586364061
transform 1 0 5060 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_47
timestamp 1586364061
transform 1 0 5428 0 -1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_60
timestamp 1586364061
transform 1 0 6624 0 -1 4896
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_79
timestamp 1586364061
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_83
timestamp 1586364061
transform 1 0 8740 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_87
timestamp 1586364061
transform 1 0 9108 0 -1 4896
box -38 -48 406 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_91
timestamp 1586364061
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_106
timestamp 1586364061
transform 1 0 10856 0 -1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_119
timestamp 1586364061
transform 1 0 12052 0 -1 4896
box -38 -48 406 592
use scs8hd_buf_2  _160_
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13064 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12880 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_125
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_133
timestamp 1586364061
transform 1 0 13340 0 -1 4896
box -38 -48 774 592
use scs8hd_nor2_4  _093_
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _092_
timestamp 1586364061
transform 1 0 16836 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16652 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16284 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_163
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_167
timestamp 1586364061
transform 1 0 16468 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18400 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_180
timestamp 1586364061
transform 1 0 17664 0 -1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_199
timestamp 1586364061
transform 1 0 19412 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_4_211
timestamp 1586364061
transform 1 0 20516 0 -1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_218
timestamp 1586364061
transform 1 0 21160 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_4_230
timestamp 1586364061
transform 1 0 22264 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 22816 0 -1 4896
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 2576 0 1 4896
box -38 -48 1050 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 2392 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2024 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_9
timestamp 1586364061
transform 1 0 1932 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_12
timestamp 1586364061
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3772 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 4140 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_31
timestamp 1586364061
transform 1 0 3956 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_35
timestamp 1586364061
transform 1 0 4324 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 4508 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7268 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7084 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use scs8hd_conb_1  _131_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 8832 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8464 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_78
timestamp 1586364061
transform 1 0 8280 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_82
timestamp 1586364061
transform 1 0 8648 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_89
timestamp 1586364061
transform 1 0 9292 0 1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10396 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 9752 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_93
timestamp 1586364061
transform 1 0 9660 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_5_96
timestamp 1586364061
transform 1 0 9936 0 1 4896
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_112
timestamp 1586364061
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_116
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 14168 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13984 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_134
timestamp 1586364061
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_138
timestamp 1586364061
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15364 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_153
timestamp 1586364061
transform 1 0 15180 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_157
timestamp 1586364061
transform 1 0 15548 0 1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16192 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_161
timestamp 1586364061
transform 1 0 15916 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_173
timestamp 1586364061
transform 1 0 17020 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_177
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18400 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20148 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20608 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19964 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_199
timestamp 1586364061
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_203
timestamp 1586364061
transform 1 0 19780 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_210
timestamp 1586364061
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_214
timestamp 1586364061
transform 1 0 20792 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_221
timestamp 1586364061
transform 1 0 21436 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_225
timestamp 1586364061
transform 1 0 21804 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 22816 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_6
timestamp 1586364061
transform 1 0 1656 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_16
timestamp 1586364061
transform 1 0 2576 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_10
timestamp 1586364061
transform 1 0 2024 0 1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_6_16
timestamp 1586364061
transform 1 0 2576 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_6_11
timestamp 1586364061
transform 1 0 2116 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 2392 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_34
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_28
timestamp 1586364061
transform 1 0 3680 0 1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2852 0 1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _109_
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use scs8hd_decap_3  FILLER_6_41
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4508 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_52
timestamp 1586364061
transform 1 0 5888 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_48
timestamp 1586364061
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_50
timestamp 1586364061
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_46
timestamp 1586364061
transform 1 0 5336 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5520 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5704 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 5796 0 -1 5984
box -38 -48 866 592
use scs8hd_decap_4  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_60
timestamp 1586364061
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_56
timestamp 1586364061
transform 1 0 6256 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_60
timestamp 1586364061
transform 1 0 6624 0 -1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6440 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_66
timestamp 1586364061
transform 1 0 7176 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_69
timestamp 1586364061
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_66
timestamp 1586364061
transform 1 0 7176 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7268 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7268 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 8464 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__050__A
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 8832 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_73
timestamp 1586364061
transform 1 0 7820 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_78
timestamp 1586364061
transform 1 0 8280 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_82
timestamp 1586364061
transform 1 0 8648 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_103
timestamp 1586364061
transform 1 0 10580 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_99
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_107
timestamp 1586364061
transform 1 0 10948 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_103
timestamp 1586364061
transform 1 0 10580 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__C
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 10764 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10948 0 1 5984
box -38 -48 314 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 9752 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_8  _050_
timestamp 1586364061
transform 1 0 9384 0 1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 11316 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 11132 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_120
timestamp 1586364061
transform 1 0 12144 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 590 592
use scs8hd_nor2_4  _096_
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12880 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14168 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_137
timestamp 1586364061
transform 1 0 13708 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_126
timestamp 1586364061
transform 1 0 12696 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_130
timestamp 1586364061
transform 1 0 13064 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_143
timestamp 1586364061
transform 1 0 14260 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_144
timestamp 1586364061
transform 1 0 14352 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14996 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_158
timestamp 1586364061
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_154
timestamp 1586364061
transform 1 0 15272 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_152
timestamp 1586364061
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_1  FILLER_7_162
timestamp 1586364061
transform 1 0 16008 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_167
timestamp 1586364061
transform 1 0 16468 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 16284 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_176
timestamp 1586364061
transform 1 0 17296 0 1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_172
timestamp 1586364061
transform 1 0 16928 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17112 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_2_.latch
timestamp 1586364061
transform 1 0 16836 0 -1 5984
box -38 -48 1050 592
use scs8hd_nor2_4  _094_
timestamp 1586364061
transform 1 0 16100 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_187
timestamp 1586364061
transform 1 0 18308 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_182
timestamp 1586364061
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_6_182
timestamp 1586364061
transform 1 0 17848 0 -1 5984
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_191
timestamp 1586364061
transform 1 0 18676 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18400 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20608 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20056 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_200
timestamp 1586364061
transform 1 0 19504 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_6_212
timestamp 1586364061
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_204
timestamp 1586364061
transform 1 0 19872 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 21068 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21436 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_218
timestamp 1586364061
transform 1 0 21160 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_6_230
timestamp 1586364061
transform 1 0 22264 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_215
timestamp 1586364061
transform 1 0 20884 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_219
timestamp 1586364061
transform 1 0 21252 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_223
timestamp 1586364061
transform 1 0 21620 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_231
timestamp 1586364061
transform 1 0 22356 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 22816 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 22816 0 1 5984
box -38 -48 314 592
use scs8hd_nor2_4  _110_
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 1564 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_7
timestamp 1586364061
transform 1 0 1748 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_13
timestamp 1586364061
transform 1 0 2300 0 -1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__105__D
timestamp 1586364061
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_43
timestamp 1586364061
transform 1 0 5060 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_47
timestamp 1586364061
transform 1 0 5428 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_50
timestamp 1586364061
transform 1 0 5704 0 -1 7072
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6440 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_8_69
timestamp 1586364061
transform 1 0 7452 0 -1 7072
box -38 -48 774 592
use scs8hd_or2_4  _082_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8188 0 -1 7072
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__055__A
timestamp 1586364061
transform 1 0 9292 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 130 592
use scs8hd_or3_4  _118_
timestamp 1586364061
transform 1 0 10120 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__090__C
timestamp 1586364061
transform 1 0 9936 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_91
timestamp 1586364061
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_107
timestamp 1586364061
transform 1 0 10948 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 11132 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 11776 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_111
timestamp 1586364061
transform 1 0 11316 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_115
timestamp 1586364061
transform 1 0 11684 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_118
timestamp 1586364061
transform 1 0 11960 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_122
timestamp 1586364061
transform 1 0 12328 0 -1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__096__B
timestamp 1586364061
transform 1 0 13800 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_125
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_136
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_140
timestamp 1586364061
transform 1 0 13984 0 -1 7072
box -38 -48 590 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15640 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15456 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_148
timestamp 1586364061
transform 1 0 14720 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_152
timestamp 1586364061
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16652 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__094__B
timestamp 1586364061
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16468 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_161
timestamp 1586364061
transform 1 0 15916 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_165
timestamp 1586364061
transform 1 0 16284 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_172
timestamp 1586364061
transform 1 0 16928 0 -1 7072
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18400 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_184
timestamp 1586364061
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19412 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_197
timestamp 1586364061
transform 1 0 19228 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_201
timestamp 1586364061
transform 1 0 19596 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_8_213
timestamp 1586364061
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_2  _138_
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_219
timestamp 1586364061
transform 1 0 21252 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_8_231
timestamp 1586364061
transform 1 0 22356 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 22816 0 -1 7072
box -38 -48 314 592
use scs8hd_buf_2  _153_
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__053__A
timestamp 1586364061
transform 1 0 2024 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__C
timestamp 1586364061
transform 1 0 2392 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_7
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_12
timestamp 1586364061
transform 1 0 2208 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_16
timestamp 1586364061
transform 1 0 2576 0 1 7072
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4140 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_24
timestamp 1586364061
transform 1 0 3312 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_29
timestamp 1586364061
transform 1 0 3772 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 5520 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__C
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_42
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_46
timestamp 1586364061
transform 1 0 5336 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7544 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6992 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_66
timestamp 1586364061
transform 1 0 7176 0 1 7072
box -38 -48 222 592
use scs8hd_nand3_4  _055_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9292 0 1 7072
box -38 -48 1326 592
use scs8hd_diode_2  ANTENNA__055__B
timestamp 1586364061
transform 1 0 9108 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__051__A
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_79
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_83
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_103
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_107
timestamp 1586364061
transform 1 0 10948 0 1 7072
box -38 -48 222 592
use scs8hd_conb_1  _133_
timestamp 1586364061
transform 1 0 11316 0 1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__D
timestamp 1586364061
transform 1 0 11132 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_134
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_138
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_142
timestamp 1586364061
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14536 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 15548 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14352 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_155
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_159
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17112 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__065__B
timestamp 1586364061
transform 1 0 15916 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_172
timestamp 1586364061
transform 1 0 16928 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_176
timestamp 1586364061
transform 1 0 17296 0 1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18308 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18768 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_180
timestamp 1586364061
transform 1 0 17664 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_190
timestamp 1586364061
transform 1 0 18584 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_194
timestamp 1586364061
transform 1 0 18952 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19320 0 1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_9_207
timestamp 1586364061
transform 1 0 20148 0 1 7072
box -38 -48 774 592
use scs8hd_conb_1  _127_
timestamp 1586364061
transform 1 0 20884 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_218
timestamp 1586364061
transform 1 0 21160 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_9_230
timestamp 1586364061
transform 1 0 22264 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 22816 0 1 7072
box -38 -48 314 592
use scs8hd_inv_8  _053_
timestamp 1586364061
transform 1 0 2024 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_7
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__116__D
timestamp 1586364061
transform 1 0 3036 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_19
timestamp 1586364061
transform 1 0 2852 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_or4_4  _105_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5520 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 5244 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_47
timestamp 1586364061
transform 1 0 5428 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_57
timestamp 1586364061
transform 1 0 6348 0 -1 8160
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_10_71
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_8  _051_
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__055__C
timestamp 1586364061
transform 1 0 9292 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_82
timestamp 1586364061
transform 1 0 8648 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 130 592
use scs8hd_or4_4  _090_
timestamp 1586364061
transform 1 0 10212 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__097__C
timestamp 1586364061
transform 1 0 9844 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_91
timestamp 1586364061
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_97
timestamp 1586364061
transform 1 0 10028 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 11776 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__056__B
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__056__C
timestamp 1586364061
transform 1 0 11592 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_108
timestamp 1586364061
transform 1 0 11040 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_112
timestamp 1586364061
transform 1 0 11408 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_125
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_133
timestamp 1586364061
transform 1 0 13340 0 -1 8160
box -38 -48 130 592
use scs8hd_nor2_4  _065_
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__057__B
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_163
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_10_168
timestamp 1586364061
transform 1 0 16560 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_174
timestamp 1586364061
transform 1 0 17112 0 -1 8160
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18400 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18032 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_182
timestamp 1586364061
transform 1 0 17848 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_186
timestamp 1586364061
transform 1 0 18216 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_197
timestamp 1586364061
transform 1 0 19228 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_201
timestamp 1586364061
transform 1 0 19596 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_205
timestamp 1586364061
transform 1 0 19964 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_213
timestamp 1586364061
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use scs8hd_conb_1  _128_
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_218
timestamp 1586364061
transform 1 0 21160 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_10_230
timestamp 1586364061
transform 1 0 22264 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 22816 0 -1 8160
box -38 -48 314 592
use scs8hd_nor4_4  _115_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 1 8160
box -38 -48 1602 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__115__D
timestamp 1586364061
transform 1 0 1656 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__C
timestamp 1586364061
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 3956 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_25
timestamp 1586364061
transform 1 0 3404 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_29
timestamp 1586364061
transform 1 0 3772 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_33
timestamp 1586364061
transform 1 0 4140 0 1 8160
box -38 -48 222 592
use scs8hd_or2_4  _104_
timestamp 1586364061
transform 1 0 5244 0 1 8160
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__113__D
timestamp 1586364061
transform 1 0 5060 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_37
timestamp 1586364061
transform 1 0 4508 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_41
timestamp 1586364061
transform 1 0 4876 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_52
timestamp 1586364061
transform 1 0 5888 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_60
timestamp 1586364061
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_56
timestamp 1586364061
transform 1 0 6256 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 6440 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 6072 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_66
timestamp 1586364061
transform 1 0 7176 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6992 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__052__A
timestamp 1586364061
transform 1 0 7360 0 1 8160
box -38 -48 222 592
use scs8hd_inv_8  _052_
timestamp 1586364061
transform 1 0 7544 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__097__D
timestamp 1586364061
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 8832 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_79
timestamp 1586364061
transform 1 0 8372 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_83
timestamp 1586364061
transform 1 0 8740 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 222 592
use scs8hd_or3_4  _075_
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10948 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__B
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_99
timestamp 1586364061
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_103
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__056__A
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_110
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _067_
timestamp 1586364061
transform 1 0 12788 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__067__B
timestamp 1586364061
transform 1 0 12604 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__061__A
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__061__B
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_136
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_140
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14812 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 15824 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_144
timestamp 1586364061
transform 1 0 14352 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_158
timestamp 1586364061
transform 1 0 15640 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _057_
timestamp 1586364061
transform 1 0 16376 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__057__A
timestamp 1586364061
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_162
timestamp 1586364061
transform 1 0 16008 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_175
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_195
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_199
timestamp 1586364061
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_212
timestamp 1586364061
transform 1 0 20608 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_217
timestamp 1586364061
transform 1 0 21068 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_11_229
timestamp 1586364061
transform 1 0 22172 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 22816 0 1 8160
box -38 -48 314 592
use scs8hd_nor4_4  _116_
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 1602 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__114__D
timestamp 1586364061
transform 1 0 4232 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use scs8hd_nor4_4  _113_
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 4692 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_36
timestamp 1586364061
transform 1 0 4416 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_12_41
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7452 0 -1 9248
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_12_61
timestamp 1586364061
transform 1 0 6716 0 -1 9248
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__075__C
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_2  FILLER_12_88
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use scs8hd_or4_4  _097_
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 774 592
use scs8hd_or3_4  _056_
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_12_119
timestamp 1586364061
transform 1 0 12052 0 -1 9248
box -38 -48 774 592
use scs8hd_nor2_4  _061_
timestamp 1586364061
transform 1 0 13616 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__087__B
timestamp 1586364061
transform 1 0 12880 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_127
timestamp 1586364061
transform 1 0 12788 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_12_130
timestamp 1586364061
transform 1 0 13064 0 -1 9248
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_151
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_165
timestamp 1586364061
transform 1 0 16284 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_12_177
timestamp 1586364061
transform 1 0 17388 0 -1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17848 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_181
timestamp 1586364061
transform 1 0 17756 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_191
timestamp 1586364061
transform 1 0 18676 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_197
timestamp 1586364061
transform 1 0 19228 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_12_209
timestamp 1586364061
transform 1 0 20332 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_213
timestamp 1586364061
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_218
timestamp 1586364061
transform 1 0 21160 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_12_230
timestamp 1586364061
transform 1 0 22264 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 22816 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_7
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__117__D
timestamp 1586364061
transform 1 0 1656 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_buf_2  _150_
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_11
timestamp 1586364061
transform 1 0 2116 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__C
timestamp 1586364061
transform 1 0 2300 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 1932 0 -1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 314 592
use scs8hd_nor4_4  _117_
timestamp 1586364061
transform 1 0 1840 0 1 9248
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_14_26
timestamp 1586364061
transform 1 0 3496 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_22
timestamp 1586364061
transform 1 0 3128 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_18
timestamp 1586364061
transform 1 0 2760 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_25
timestamp 1586364061
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 3312 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 2944 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_30
timestamp 1586364061
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_29
timestamp 1586364061
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3680 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 4232 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__C
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_nor4_4  _114_
timestamp 1586364061
transform 1 0 4140 0 1 9248
box -38 -48 1602 592
use scs8hd_nor4_4  _112_
timestamp 1586364061
transform 1 0 4692 0 -1 10336
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__112__C
timestamp 1586364061
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_50
timestamp 1586364061
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_36
timestamp 1586364061
transform 1 0 4416 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_58
timestamp 1586364061
transform 1 0 6440 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_54
timestamp 1586364061
transform 1 0 6072 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__D
timestamp 1586364061
transform 1 0 6256 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_70
timestamp 1586364061
transform 1 0 7544 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_66
timestamp 1586364061
transform 1 0 7176 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7360 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6992 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6992 0 -1 10336
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_84
timestamp 1586364061
transform 1 0 8832 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_75
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_79
timestamp 1586364061
transform 1 0 8372 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_14_87
timestamp 1586364061
transform 1 0 9108 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_6  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_95
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_92
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__D
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_101
timestamp 1586364061
transform 1 0 10396 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__C
timestamp 1586364061
transform 1 0 10580 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 10212 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _085_
timestamp 1586364061
transform 1 0 10856 0 -1 10336
box -38 -48 866 592
use scs8hd_or4_4  _083_
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_14_115
timestamp 1586364061
transform 1 0 11684 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_112
timestamp 1586364061
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_108
timestamp 1586364061
transform 1 0 11040 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_116
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_128
timestamp 1586364061
transform 1 0 12880 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13064 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_137
timestamp 1586364061
transform 1 0 13708 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13892 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 1050 592
use scs8hd_nor2_4  _087_
timestamp 1586364061
transform 1 0 12880 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_8  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_13_151
timestamp 1586364061
transform 1 0 14996 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_147
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14260 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_157
timestamp 1586364061
transform 1 0 15548 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_154
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15732 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15088 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 1 9248
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 16468 0 -1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 16652 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17020 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_167
timestamp 1586364061
transform 1 0 16468 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_171
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 590 592
use scs8hd_decap_6  FILLER_14_161
timestamp 1586364061
transform 1 0 15916 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_8  FILLER_14_178
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 18216 0 -1 10336
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 18216 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_188
timestamp 1586364061
transform 1 0 18400 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_192
timestamp 1586364061
transform 1 0 18768 0 1 9248
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_204
timestamp 1586364061
transform 1 0 19872 0 1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_13_212
timestamp 1586364061
transform 1 0 20608 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_197
timestamp 1586364061
transform 1 0 19228 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_209
timestamp 1586364061
transform 1 0 20332 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_213
timestamp 1586364061
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_2  _151_
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_217
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_13_229
timestamp 1586364061
transform 1 0 22172 0 1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_219
timestamp 1586364061
transform 1 0 21252 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_231
timestamp 1586364061
transform 1 0 22356 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 22816 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 22816 0 -1 10336
box -38 -48 314 592
use scs8hd_buf_2  _146_
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2300 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_11
timestamp 1586364061
transform 1 0 2116 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_26
timestamp 1586364061
transform 1 0 3496 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_22
timestamp 1586364061
transform 1 0 3128 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_18
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3312 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_34
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_30
timestamp 1586364061
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__043__A
timestamp 1586364061
transform 1 0 3680 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use scs8hd_inv_8  _043_
timestamp 1586364061
transform 1 0 4324 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5336 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_44
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_48
timestamp 1586364061
transform 1 0 5520 0 1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_54
timestamp 1586364061
transform 1 0 6072 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_65
timestamp 1586364061
transform 1 0 7084 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_69
timestamp 1586364061
transform 1 0 7452 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9200 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_82
timestamp 1586364061
transform 1 0 8648 0 1 10336
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9384 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__068__B
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_99
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_103
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_107
timestamp 1586364061
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__C
timestamp 1586364061
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11868 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_111
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_115
timestamp 1586364061
transform 1 0 11684 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_119
timestamp 1586364061
transform 1 0 12052 0 1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 13892 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 13708 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12880 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_126
timestamp 1586364061
transform 1 0 12696 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_130
timestamp 1586364061
transform 1 0 13064 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_134
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_150
timestamp 1586364061
transform 1 0 14904 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_156
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_160
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 406 592
use scs8hd_nor2_4  _059_
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__059__A
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18308 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19504 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19872 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_198
timestamp 1586364061
transform 1 0 19320 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_202
timestamp 1586364061
transform 1 0 19688 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_206
timestamp 1586364061
transform 1 0 20056 0 1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_15_214
timestamp 1586364061
transform 1 0 20792 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_217
timestamp 1586364061
transform 1 0 21068 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_15_229
timestamp 1586364061
transform 1 0 22172 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 22816 0 1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 1050 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_18
timestamp 1586364061
transform 1 0 2760 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_22
timestamp 1586364061
transform 1 0 3128 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_30
timestamp 1586364061
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use scs8hd_conb_1  _135_
timestamp 1586364061
transform 1 0 5796 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_43
timestamp 1586364061
transform 1 0 5060 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_54
timestamp 1586364061
transform 1 0 6072 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_62
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 130 592
use scs8hd_conb_1  _134_
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7912 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_72
timestamp 1586364061
transform 1 0 7728 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_76
timestamp 1586364061
transform 1 0 8096 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_16_83
timestamp 1586364061
transform 1 0 8740 0 -1 11424
box -38 -48 774 592
use scs8hd_or3_4  _068_
timestamp 1586364061
transform 1 0 9936 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_91
timestamp 1586364061
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 11500 0 -1 11424
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_16_124
timestamp 1586364061
transform 1 0 12512 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13248 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_6  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_149
timestamp 1586364061
transform 1 0 14812 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__B
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_163
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_168
timestamp 1586364061
transform 1 0 16560 0 -1 11424
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_180
timestamp 1586364061
transform 1 0 17664 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_188
timestamp 1586364061
transform 1 0 18400 0 -1 11424
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_198
timestamp 1586364061
transform 1 0 19320 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_16_210
timestamp 1586364061
transform 1 0 20424 0 -1 11424
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_218
timestamp 1586364061
transform 1 0 21160 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_16_230
timestamp 1586364061
transform 1 0 22264 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 22816 0 -1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2208 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_6
timestamp 1586364061
transform 1 0 1656 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_10
timestamp 1586364061
transform 1 0 2024 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4232 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3404 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_23
timestamp 1586364061
transform 1 0 3220 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_31
timestamp 1586364061
transform 1 0 3956 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5244 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_43
timestamp 1586364061
transform 1 0 5060 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_47
timestamp 1586364061
transform 1 0 5428 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__042__A
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_73
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_77
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9936 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10948 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_90
timestamp 1586364061
transform 1 0 9384 0 1 11424
box -38 -48 590 592
use scs8hd_fill_2  FILLER_17_101
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_105
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _086_
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_109
timestamp 1586364061
transform 1 0 11132 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_115
timestamp 1586364061
transform 1 0 11684 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_132
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_136
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_140
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__063__B
timestamp 1586364061
transform 1 0 15640 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_144
timestamp 1586364061
transform 1 0 14352 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_156
timestamp 1586364061
transform 1 0 15456 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_160
timestamp 1586364061
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _063_
timestamp 1586364061
transform 1 0 16192 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 16008 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_173
timestamp 1586364061
transform 1 0 17020 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_181
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_214
timestamp 1586364061
transform 1 0 20792 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_217
timestamp 1586364061
transform 1 0 21068 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_17_229
timestamp 1586364061
transform 1 0 22172 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 22816 0 1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2300 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 1564 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2116 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_7
timestamp 1586364061
transform 1 0 1748 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4232 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_22
timestamp 1586364061
transform 1 0 3128 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_30
timestamp 1586364061
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4784 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_4  FILLER_18_36
timestamp 1586364061
transform 1 0 4416 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_18_49
timestamp 1586364061
transform 1 0 5612 0 -1 12512
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6348 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__041__A
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7176 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_59
timestamp 1586364061
transform 1 0 6532 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_64
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 406 592
use scs8hd_inv_8  _042_
timestamp 1586364061
transform 1 0 7728 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_81
timestamp 1586364061
transform 1 0 8556 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_85
timestamp 1586364061
transform 1 0 8924 0 -1 12512
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 10028 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_91
timestamp 1586364061
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_108
timestamp 1586364061
transform 1 0 11040 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_18_120
timestamp 1586364061
transform 1 0 12144 0 -1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13248 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12788 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_125
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_129
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_6  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_149
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 406 592
use scs8hd_conb_1  _125_
timestamp 1586364061
transform 1 0 16836 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_163
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_18_174
timestamp 1586364061
transform 1 0 17112 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_186
timestamp 1586364061
transform 1 0 18216 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_198
timestamp 1586364061
transform 1 0 19320 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_18_210
timestamp 1586364061
transform 1 0 20424 0 -1 12512
box -38 -48 406 592
use scs8hd_buf_2  _149_
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_219
timestamp 1586364061
transform 1 0 21252 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_18_231
timestamp 1586364061
transform 1 0 22356 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 22816 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__044__A
timestamp 1586364061
transform 1 0 1840 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_buf_2  _145_
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_11
timestamp 1586364061
transform 1 0 2116 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2300 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 1932 0 -1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 314 592
use scs8hd_inv_8  _044_
timestamp 1586364061
transform 1 0 2024 0 1 12512
box -38 -48 866 592
use scs8hd_decap_4  FILLER_19_23
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_19
timestamp 1586364061
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_30
timestamp 1586364061
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_29
timestamp 1586364061
transform 1 0 3772 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 3956 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_18
timestamp 1586364061
transform 1 0 2760 0 -1 13600
box -38 -48 1142 592
use scs8hd_nor2_4  _076_
timestamp 1586364061
transform 1 0 4140 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_42
timestamp 1586364061
transform 1 0 4968 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_40
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_36
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_50
timestamp 1586364061
transform 1 0 5704 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_46
timestamp 1586364061
transform 1 0 5336 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5520 0 -1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _078_
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use scs8hd_inv_8  _041_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 6348 0 -1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7544 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_71
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_68
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_72
timestamp 1586364061
transform 1 0 7728 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_3  FILLER_19_78
timestamp 1586364061
transform 1 0 8280 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_19_75
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8096 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8096 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_6  FILLER_20_79
timestamp 1586364061
transform 1 0 8372 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_84
timestamp 1586364061
transform 1 0 8832 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 -1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_87
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_88
timestamp 1586364061
transform 1 0 9200 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_97
timestamp 1586364061
transform 1 0 10028 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_91
timestamp 1586364061
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 9384 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_101
timestamp 1586364061
transform 1 0 10396 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_105
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_101
timestamp 1586364061
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10948 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 866 592
use scs8hd_nor2_4  _100_
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_20_111
timestamp 1586364061
transform 1 0 11316 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_112
timestamp 1586364061
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11132 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_121
timestamp 1586364061
transform 1 0 12236 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_116
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_134
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_138
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_136
timestamp 1586364061
transform 1 0 13616 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_4  FILLER_20_148
timestamp 1586364061
transform 1 0 14720 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_144
timestamp 1586364061
transform 1 0 14352 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_151
timestamp 1586364061
transform 1 0 14996 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14536 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_157
timestamp 1586364061
transform 1 0 15548 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_152
timestamp 1586364061
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_19_156
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__071__B
timestamp 1586364061
transform 1 0 15732 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use scs8hd_nor2_4  _071_
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_165
timestamp 1586364061
transform 1 0 16284 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_161
timestamp 1586364061
transform 1 0 15916 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_168
timestamp 1586364061
transform 1 0 16560 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16468 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_176
timestamp 1586364061
transform 1 0 17296 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_172
timestamp 1586364061
transform 1 0 16928 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17112 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 16744 0 1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 16652 0 -1 13600
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_20_180
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_187
timestamp 1586364061
transform 1 0 18308 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_182
timestamp 1586364061
transform 1 0 17848 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_195
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_191
timestamp 1586364061
transform 1 0 18676 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18400 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_203
timestamp 1586364061
transform 1 0 19780 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_199
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19964 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19504 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_213
timestamp 1586364061
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_209
timestamp 1586364061
transform 1 0 20332 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_214
timestamp 1586364061
transform 1 0 20792 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_207
timestamp 1586364061
transform 1 0 20148 0 1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20516 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_197
timestamp 1586364061
transform 1 0 19228 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_2  _158_
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20976 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_218
timestamp 1586364061
transform 1 0 21160 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_222
timestamp 1586364061
transform 1 0 21528 0 1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_19_230
timestamp 1586364061
transform 1 0 22264 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_219
timestamp 1586364061
transform 1 0 21252 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_20_231
timestamp 1586364061
transform 1 0 22356 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 22816 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 22816 0 -1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 1564 0 1 13600
box -38 -48 1050 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_16
timestamp 1586364061
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 4232 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3128 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_20
timestamp 1586364061
transform 1 0 2944 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_24
timestamp 1586364061
transform 1 0 3312 0 1 13600
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5428 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_45
timestamp 1586364061
transform 1 0 5244 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_49
timestamp 1586364061
transform 1 0 5612 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6440 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6072 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_56
timestamp 1586364061
transform 1 0 6256 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_60
timestamp 1586364061
transform 1 0 6624 0 1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8924 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8740 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_72
timestamp 1586364061
transform 1 0 7728 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_77
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_81
timestamp 1586364061
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _084_
timestamp 1586364061
transform 1 0 10764 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__084__B
timestamp 1586364061
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_96
timestamp 1586364061
transform 1 0 9936 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_100
timestamp 1586364061
transform 1 0 10304 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 12696 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14168 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 13708 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_135
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_139
timestamp 1586364061
transform 1 0 13892 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14536 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_144
timestamp 1586364061
transform 1 0 14352 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_155
timestamp 1586364061
transform 1 0 15364 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_159
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 16192 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_162
timestamp 1586364061
transform 1 0 16008 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_175
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_196
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 22816 0 1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_21_232
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 1656 0 -1 14688
box -38 -48 1050 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_17
timestamp 1586364061
transform 1 0 2668 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_29
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4876 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4600 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_36
timestamp 1586364061
transform 1 0 4416 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_40
timestamp 1586364061
transform 1 0 4784 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_6  FILLER_22_50
timestamp 1586364061
transform 1 0 5704 0 -1 14688
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6440 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7452 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_67
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_71
timestamp 1586364061
transform 1 0 7636 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_102
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_107
timestamp 1586364061
transform 1 0 10948 0 -1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_113
timestamp 1586364061
transform 1 0 11500 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_121
timestamp 1586364061
transform 1 0 12236 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13616 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_134
timestamp 1586364061
transform 1 0 13432 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_138
timestamp 1586364061
transform 1 0 13800 0 -1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__069__B
timestamp 1586364061
transform 1 0 15548 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_149
timestamp 1586364061
transform 1 0 14812 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_3  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_159
timestamp 1586364061
transform 1 0 15732 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 16192 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 15916 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_163
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_175
timestamp 1586364061
transform 1 0 17204 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_187
timestamp 1586364061
transform 1 0 18308 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_199
timestamp 1586364061
transform 1 0 19412 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_22_211
timestamp 1586364061
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 590 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 22816 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_16
timestamp 1586364061
transform 1 0 2576 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3312 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3772 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4140 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__046__A
timestamp 1586364061
transform 1 0 2760 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3128 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_20
timestamp 1586364061
transform 1 0 2944 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_31
timestamp 1586364061
transform 1 0 3956 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_35
timestamp 1586364061
transform 1 0 4324 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_49
timestamp 1586364061
transform 1 0 5612 0 1 14688
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use scs8hd_nor2_4  _103_
timestamp 1586364061
transform 1 0 8648 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_74
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_79
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_91
timestamp 1586364061
transform 1 0 9476 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_95
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_99
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11316 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_109
timestamp 1586364061
transform 1 0 11132 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_113
timestamp 1586364061
transform 1 0 11500 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_117
timestamp 1586364061
transform 1 0 11868 0 1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13340 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_126
timestamp 1586364061
transform 1 0 12696 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_130
timestamp 1586364061
transform 1 0 13064 0 1 14688
box -38 -48 314 592
use scs8hd_nor2_4  _072_
timestamp 1586364061
transform 1 0 15548 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__072__B
timestamp 1586364061
transform 1 0 15364 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 14996 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_146
timestamp 1586364061
transform 1 0 14536 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_150
timestamp 1586364061
transform 1 0 14904 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_153
timestamp 1586364061
transform 1 0 15180 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 17112 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17480 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_166
timestamp 1586364061
transform 1 0 16376 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_176
timestamp 1586364061
transform 1 0 17296 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_23_180
timestamp 1586364061
transform 1 0 17664 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_196
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 20700 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_212
timestamp 1586364061
transform 1 0 20608 0 1 14688
box -38 -48 130 592
use scs8hd_buf_2  _157_
timestamp 1586364061
transform 1 0 20884 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 21436 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_219
timestamp 1586364061
transform 1 0 21252 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_223
timestamp 1586364061
transform 1 0 21620 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_231
timestamp 1586364061
transform 1 0 22356 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 22816 0 1 14688
box -38 -48 314 592
use scs8hd_inv_8  _046_
timestamp 1586364061
transform 1 0 1656 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2668 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4140 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_19
timestamp 1586364061
transform 1 0 2852 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_42
timestamp 1586364061
transform 1 0 4968 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_46
timestamp 1586364061
transform 1 0 5336 0 -1 15776
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6624 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_58
timestamp 1586364061
transform 1 0 6440 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_69
timestamp 1586364061
transform 1 0 7452 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8188 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 8648 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_73
timestamp 1586364061
transform 1 0 7820 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10028 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 9844 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12420 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 11592 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 11224 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 11960 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_108
timestamp 1586364061
transform 1 0 11040 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_112
timestamp 1586364061
transform 1 0 11408 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_116
timestamp 1586364061
transform 1 0 11776 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_120
timestamp 1586364061
transform 1 0 12144 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__074__B
timestamp 1586364061
transform 1 0 13616 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14076 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_134
timestamp 1586364061
transform 1 0 13432 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_138
timestamp 1586364061
transform 1 0 13800 0 -1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _069_
timestamp 1586364061
transform 1 0 15548 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_143
timestamp 1586364061
transform 1 0 14260 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_151
timestamp 1586364061
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 17112 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 16560 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_166
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_170
timestamp 1586364061
transform 1 0 16744 0 -1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18308 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_185
timestamp 1586364061
transform 1 0 18124 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_189
timestamp 1586364061
transform 1 0 18492 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_201
timestamp 1586364061
transform 1 0 19596 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_24_213
timestamp 1586364061
transform 1 0 20700 0 -1 15776
box -38 -48 130 592
use scs8hd_buf_2  _156_
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_219
timestamp 1586364061
transform 1 0 21252 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_24_231
timestamp 1586364061
transform 1 0 22356 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 22816 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 4232 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 3864 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 3496 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_18
timestamp 1586364061
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_22
timestamp 1586364061
transform 1 0 3128 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_28
timestamp 1586364061
transform 1 0 3680 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_32
timestamp 1586364061
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4416 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5612 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_47
timestamp 1586364061
transform 1 0 5428 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _081_
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_55
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_71
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8924 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8740 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_75
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 774 592
use scs8hd_nor2_4  _098_
timestamp 1586364061
transform 1 0 10488 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 10028 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_94
timestamp 1586364061
transform 1 0 9752 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_25_99
timestamp 1586364061
transform 1 0 10212 0 1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _089_
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_111
timestamp 1586364061
transform 1 0 11316 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_115
timestamp 1586364061
transform 1 0 11684 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 14076 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13892 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_132
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_136
timestamp 1586364061
transform 1 0 13616 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__B
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_152
timestamp 1586364061
transform 1 0 15088 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_156
timestamp 1586364061
transform 1 0 15456 0 1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _070_
timestamp 1586364061
transform 1 0 16284 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16100 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 17296 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_161
timestamp 1586364061
transform 1 0 15916 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_174
timestamp 1586364061
transform 1 0 17112 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_178
timestamp 1586364061
transform 1 0 17480 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17664 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_182
timestamp 1586364061
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_193
timestamp 1586364061
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19964 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20424 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_197
timestamp 1586364061
transform 1 0 19228 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_208
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_212
timestamp 1586364061
transform 1 0 20608 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_224
timestamp 1586364061
transform 1 0 21712 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 22816 0 1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_25_232
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_7
timestamp 1586364061
transform 1 0 1748 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_14
timestamp 1586364061
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_25
timestamp 1586364061
transform 1 0 3404 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_18
timestamp 1586364061
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_22
timestamp 1586364061
transform 1 0 3128 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_26_18
timestamp 1586364061
transform 1 0 2760 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__045__A
timestamp 1586364061
transform 1 0 2944 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3128 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_29
timestamp 1586364061
transform 1 0 3772 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_28
timestamp 1586364061
transform 1 0 3680 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__079__B
timestamp 1586364061
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4232 0 1 16864
box -38 -48 1050 592
use scs8hd_nor2_4  _080_
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5980 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 5612 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_41
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_45
timestamp 1586364061
transform 1 0 5244 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_4  FILLER_27_45
timestamp 1586364061
transform 1 0 5244 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _077_
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__081__B
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__B
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 590 592
use scs8hd_decap_4  FILLER_27_55
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_27_71
timestamp 1586364061
transform 1 0 7636 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_77
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_79
timestamp 1586364061
transform 1 0 8372 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_75
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 8188 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_87
timestamp 1586364061
transform 1 0 9108 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_83
timestamp 1586364061
transform 1 0 8740 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8556 0 -1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_27_97
timestamp 1586364061
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_92
timestamp 1586364061
transform 1 0 9568 0 1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_91
timestamp 1586364061
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 9844 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_106
timestamp 1586364061
transform 1 0 10856 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 1050 592
use scs8hd_nor2_4  _099_
timestamp 1586364061
transform 1 0 10028 0 -1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 11592 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 11040 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_110
timestamp 1586364061
transform 1 0 11224 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_8  FILLER_26_123
timestamp 1586364061
transform 1 0 12420 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_112
timestamp 1586364061
transform 1 0 11408 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_116
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 590 592
use scs8hd_decap_3  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_128
timestamp 1586364061
transform 1 0 12880 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_131
timestamp 1586364061
transform 1 0 13156 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 12696 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__B
timestamp 1586364061
transform 1 0 13064 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_136
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13708 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_141
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13892 0 1 16864
box -38 -48 1050 592
use scs8hd_nor2_4  _074_
timestamp 1586364061
transform 1 0 13248 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15088 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_157
timestamp 1586364061
transform 1 0 15548 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_150
timestamp 1586364061
transform 1 0 14904 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_154
timestamp 1586364061
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_158
timestamp 1586364061
transform 1 0 15640 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_168
timestamp 1586364061
transform 1 0 16560 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_26_164
timestamp 1586364061
transform 1 0 16192 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_161
timestamp 1586364061
transform 1 0 15916 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16008 0 -1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16284 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_177
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_171
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 17296 0 -1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18124 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18492 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_187
timestamp 1586364061
transform 1 0 18308 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_191
timestamp 1586364061
transform 1 0 18676 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_181
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_194
timestamp 1586364061
transform 1 0 18952 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_203
timestamp 1586364061
transform 1 0 19780 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_26_211
timestamp 1586364061
transform 1 0 20516 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_27_206
timestamp 1586364061
transform 1 0 20056 0 1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_27_214
timestamp 1586364061
transform 1 0 20792 0 1 16864
box -38 -48 130 592
use scs8hd_buf_2  _154_
timestamp 1586364061
transform 1 0 20884 0 1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 21436 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_219
timestamp 1586364061
transform 1 0 21252 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_27_223
timestamp 1586364061
transform 1 0 21620 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_231
timestamp 1586364061
transform 1 0 22356 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 22816 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 22816 0 1 16864
box -38 -48 314 592
use scs8hd_inv_8  _045_
timestamp 1586364061
transform 1 0 1656 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_nor2_4  _079_
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 5612 0 -1 17952
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_28_41
timestamp 1586364061
transform 1 0 4876 0 -1 17952
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 6808 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7176 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7544 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_60
timestamp 1586364061
transform 1 0 6624 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_64
timestamp 1586364061
transform 1 0 6992 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _102_
timestamp 1586364061
transform 1 0 8004 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_72
timestamp 1586364061
transform 1 0 7728 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_84
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_88
timestamp 1586364061
transform 1 0 9200 0 -1 17952
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 10672 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10396 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_28_103
timestamp 1586364061
transform 1 0 10580 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_115
timestamp 1586364061
transform 1 0 11684 0 -1 17952
box -38 -48 774 592
use scs8hd_nor2_4  _073_
timestamp 1586364061
transform 1 0 13064 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12880 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_125
timestamp 1586364061
transform 1 0 12604 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_139
timestamp 1586364061
transform 1 0 13892 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15456 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_143
timestamp 1586364061
transform 1 0 14260 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_151
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17204 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_8  FILLER_28_167
timestamp 1586364061
transform 1 0 16468 0 -1 17952
box -38 -48 774 592
use scs8hd_conb_1  _130_
timestamp 1586364061
transform 1 0 18768 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18216 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_184
timestamp 1586364061
transform 1 0 18032 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_188
timestamp 1586364061
transform 1 0 18400 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_195
timestamp 1586364061
transform 1 0 19044 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_28_207
timestamp 1586364061
transform 1 0 20148 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_213
timestamp 1586364061
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 590 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 22816 0 -1 17952
box -38 -48 314 592
use scs8hd_buf_2  _161_
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 2300 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_7
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_11
timestamp 1586364061
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_18
timestamp 1586364061
transform 1 0 2760 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_22
timestamp 1586364061
transform 1 0 3128 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_29_34
timestamp 1586364061
transform 1 0 4232 0 1 17952
box -38 -48 314 592
use scs8hd_conb_1  _129_
timestamp 1586364061
transform 1 0 4508 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5520 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_40
timestamp 1586364061
transform 1 0 4784 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_46
timestamp 1586364061
transform 1 0 5336 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_50
timestamp 1586364061
transform 1 0 5704 0 1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_54
timestamp 1586364061
transform 1 0 6072 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_71
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8648 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_76
timestamp 1586364061
transform 1 0 8096 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_80
timestamp 1586364061
transform 1 0 8464 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_91
timestamp 1586364061
transform 1 0 9476 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_97
timestamp 1586364061
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_101
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14168 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_132
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_136
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_140
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14352 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15364 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_153
timestamp 1586364061
transform 1 0 15180 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_157
timestamp 1586364061
transform 1 0 15548 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16928 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17296 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_170
timestamp 1586364061
transform 1 0 16744 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_174
timestamp 1586364061
transform 1 0 17112 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_178
timestamp 1586364061
transform 1 0 17480 0 1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_193
timestamp 1586364061
transform 1 0 18860 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_205
timestamp 1586364061
transform 1 0 19964 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_217
timestamp 1586364061
transform 1 0 21068 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_29_229
timestamp 1586364061
transform 1 0 22172 0 1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 22816 0 1 17952
box -38 -48 314 592
use scs8hd_conb_1  _132_
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 314 592
use scs8hd_buf_2  _155_
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_7
timestamp 1586364061
transform 1 0 1748 0 -1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_18
timestamp 1586364061
transform 1 0 2760 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_30_30
timestamp 1586364061
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_8  FILLER_30_53
timestamp 1586364061
transform 1 0 5980 0 -1 19040
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6716 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_8  FILLER_30_70
timestamp 1586364061
transform 1 0 7544 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8280 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8740 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_81
timestamp 1586364061
transform 1 0 8556 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_85
timestamp 1586364061
transform 1 0 8924 0 -1 19040
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_91
timestamp 1586364061
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_97
timestamp 1586364061
transform 1 0 10028 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_114
timestamp 1586364061
transform 1 0 11592 0 -1 19040
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12880 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_126
timestamp 1586364061
transform 1 0 12696 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_137
timestamp 1586364061
transform 1 0 13708 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_142
timestamp 1586364061
transform 1 0 14168 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14352 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_146
timestamp 1586364061
transform 1 0 14536 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_152
timestamp 1586364061
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_163
timestamp 1586364061
transform 1 0 16100 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_167
timestamp 1586364061
transform 1 0 16468 0 -1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_180
timestamp 1586364061
transform 1 0 17664 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_186
timestamp 1586364061
transform 1 0 18216 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_198
timestamp 1586364061
transform 1 0 19320 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_30_210
timestamp 1586364061
transform 1 0 20424 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 590 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 22816 0 -1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2024 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_6
timestamp 1586364061
transform 1 0 1656 0 1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_31_12
timestamp 1586364061
transform 1 0 2208 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_24
timestamp 1586364061
transform 1 0 3312 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_36
timestamp 1586364061
transform 1 0 4416 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_48
timestamp 1586364061
transform 1 0 5520 0 1 19040
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_56
timestamp 1586364061
transform 1 0 6256 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_71
timestamp 1586364061
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8740 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8464 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_75
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_79
timestamp 1586364061
transform 1 0 8372 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_82
timestamp 1586364061
transform 1 0 8648 0 1 19040
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_92
timestamp 1586364061
transform 1 0 9568 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_96
timestamp 1586364061
transform 1 0 9936 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12512 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_109
timestamp 1586364061
transform 1 0 11132 0 1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_31_121
timestamp 1586364061
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13984 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12972 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13340 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13708 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_127
timestamp 1586364061
transform 1 0 12788 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_131
timestamp 1586364061
transform 1 0 13156 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_139
timestamp 1586364061
transform 1 0 13892 0 1 19040
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15548 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_149
timestamp 1586364061
transform 1 0 14812 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_153
timestamp 1586364061
transform 1 0 15180 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_156
timestamp 1586364061
transform 1 0 15456 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_160
timestamp 1586364061
transform 1 0 15824 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16008 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_164
timestamp 1586364061
transform 1 0 16192 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_168
timestamp 1586364061
transform 1 0 16560 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_173
timestamp 1586364061
transform 1 0 17020 0 1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18676 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_181
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_31_190
timestamp 1586364061
transform 1 0 18584 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_194
timestamp 1586364061
transform 1 0 18952 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20516 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_198
timestamp 1586364061
transform 1 0 19320 0 1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_31_210
timestamp 1586364061
transform 1 0 20424 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_214
timestamp 1586364061
transform 1 0 20792 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21528 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20976 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21988 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_218
timestamp 1586364061
transform 1 0 21160 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_225
timestamp 1586364061
transform 1 0 21804 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_229
timestamp 1586364061
transform 1 0 22172 0 1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 22816 0 1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2024 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_7
timestamp 1586364061
transform 1 0 1748 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_13
timestamp 1586364061
transform 1 0 2300 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_6  FILLER_32_25
timestamp 1586364061
transform 1 0 3404 0 -1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7452 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6808 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 590 592
use scs8hd_decap_4  FILLER_32_64
timestamp 1586364061
transform 1 0 6992 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_72
timestamp 1586364061
transform 1 0 7728 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_32_83
timestamp 1586364061
transform 1 0 8740 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_87
timestamp 1586364061
transform 1 0 9108 0 -1 20128
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9844 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_91
timestamp 1586364061
transform 1 0 9476 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_104
timestamp 1586364061
transform 1 0 10672 0 -1 20128
box -38 -48 774 592
use scs8hd_conb_1  _126_
timestamp 1586364061
transform 1 0 11408 0 -1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12512 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_115
timestamp 1586364061
transform 1 0 11684 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_123
timestamp 1586364061
transform 1 0 12420 0 -1 20128
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13340 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_127
timestamp 1586364061
transform 1 0 12788 0 -1 20128
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_144
timestamp 1586364061
transform 1 0 14352 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_152
timestamp 1586364061
transform 1 0 15088 0 -1 20128
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_163
timestamp 1586364061
transform 1 0 16100 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_32_174
timestamp 1586364061
transform 1 0 17112 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_186
timestamp 1586364061
transform 1 0 18216 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_198
timestamp 1586364061
transform 1 0 19320 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_32_210
timestamp 1586364061
transform 1 0 20424 0 -1 20128
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_218
timestamp 1586364061
transform 1 0 21160 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_32_230
timestamp 1586364061
transform 1 0 22264 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 22816 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_6
timestamp 1586364061
transform 1 0 1656 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_33_14
timestamp 1586364061
transform 1 0 2392 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_10
timestamp 1586364061
transform 1 0 2024 0 1 20128
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_33_26
timestamp 1586364061
transform 1 0 3496 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_22
timestamp 1586364061
transform 1 0 3128 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_18
timestamp 1586364061
transform 1 0 2760 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_31
timestamp 1586364061
transform 1 0 3956 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 4140 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_buf_2  _137_
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_35
timestamp 1586364061
transform 1 0 4324 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_47
timestamp 1586364061
transform 1 0 5428 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7544 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8004 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8556 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_73
timestamp 1586364061
transform 1 0 7820 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_77
timestamp 1586364061
transform 1 0 8188 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_34_83
timestamp 1586364061
transform 1 0 8740 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_6  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_34_91
timestamp 1586364061
transform 1 0 9476 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_90
timestamp 1586364061
transform 1 0 9384 0 1 20128
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_buf_2  _152_
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_99
timestamp 1586364061
transform 1 0 10212 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_106
timestamp 1586364061
transform 1 0 10856 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_102
timestamp 1586364061
transform 1 0 10488 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 10672 0 1 20128
box -38 -48 222 592
use scs8hd_buf_2  _147_
timestamp 1586364061
transform 1 0 10304 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_104
timestamp 1586364061
transform 1 0 10672 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 11040 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_116
timestamp 1586364061
transform 1 0 11776 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13708 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13984 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_138
timestamp 1586364061
transform 1 0 13800 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_142
timestamp 1586364061
transform 1 0 14168 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_128
timestamp 1586364061
transform 1 0 12880 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_136
timestamp 1586364061
transform 1 0 13616 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_140
timestamp 1586364061
transform 1 0 13984 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15088 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15548 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14352 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_146
timestamp 1586364061
transform 1 0 14536 0 1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_33_155
timestamp 1586364061
transform 1 0 15364 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_159
timestamp 1586364061
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_152
timestamp 1586364061
transform 1 0 15088 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_171
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18308 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18768 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_190
timestamp 1586364061
transform 1 0 18584 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_194
timestamp 1586364061
transform 1 0 18952 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_206
timestamp 1586364061
transform 1 0 20056 0 1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_33_214
timestamp 1586364061
transform 1 0 20792 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_218
timestamp 1586364061
transform 1 0 21160 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_222
timestamp 1586364061
transform 1 0 21528 0 1 20128
box -38 -48 774 592
use scs8hd_decap_3  FILLER_33_230
timestamp 1586364061
transform 1 0 22264 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 590 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 22816 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 22816 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 3956 0 1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_35_32
timestamp 1586364061
transform 1 0 4048 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_44
timestamp 1586364061
transform 1 0 5152 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_56
timestamp 1586364061
transform 1 0 6256 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_63
timestamp 1586364061
transform 1 0 6900 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_75
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_87
timestamp 1586364061
transform 1 0 9108 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 9660 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_94
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_106
timestamp 1586364061
transform 1 0 10856 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_125
timestamp 1586364061
transform 1 0 12604 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_137
timestamp 1586364061
transform 1 0 13708 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_149
timestamp 1586364061
transform 1 0 14812 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_156
timestamp 1586364061
transform 1 0 15456 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_168
timestamp 1586364061
transform 1 0 16560 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 18216 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_180
timestamp 1586364061
transform 1 0 17664 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_187
timestamp 1586364061
transform 1 0 18308 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_199
timestamp 1586364061
transform 1 0 19412 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_211
timestamp 1586364061
transform 1 0 20516 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_218
timestamp 1586364061
transform 1 0 21160 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_35_230
timestamp 1586364061
transform 1 0 22264 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 22816 0 1 21216
box -38 -48 314 592
<< labels >>
rlabel metal2 s 2042 0 2098 480 6 address[0]
port 0 nsew default input
rlabel metal3 s 23520 552 24000 672 6 address[1]
port 1 nsew default input
rlabel metal3 s 23520 1776 24000 1896 6 address[2]
port 2 nsew default input
rlabel metal2 s 2870 0 2926 480 6 address[3]
port 3 nsew default input
rlabel metal3 s 23520 3000 24000 3120 6 address[4]
port 4 nsew default input
rlabel metal3 s 23520 4224 24000 4344 6 address[5]
port 5 nsew default input
rlabel metal2 s 3698 0 3754 480 6 address[6]
port 6 nsew default input
rlabel metal2 s 662 23520 718 24000 6 chanx_left_in[0]
port 7 nsew default input
rlabel metal3 s 23520 5584 24000 5704 6 chanx_left_in[1]
port 8 nsew default input
rlabel metal3 s 23520 6808 24000 6928 6 chanx_left_in[2]
port 9 nsew default input
rlabel metal2 s 1950 23520 2006 24000 6 chanx_left_in[3]
port 10 nsew default input
rlabel metal2 s 4526 0 4582 480 6 chanx_left_in[4]
port 11 nsew default input
rlabel metal2 s 5354 0 5410 480 6 chanx_left_in[5]
port 12 nsew default input
rlabel metal3 s 0 688 480 808 6 chanx_left_in[6]
port 13 nsew default input
rlabel metal2 s 6182 0 6238 480 6 chanx_left_in[7]
port 14 nsew default input
rlabel metal2 s 3330 23520 3386 24000 6 chanx_left_in[8]
port 15 nsew default input
rlabel metal3 s 0 2048 480 2168 6 chanx_left_out[0]
port 16 nsew default tristate
rlabel metal3 s 0 3408 480 3528 6 chanx_left_out[1]
port 17 nsew default tristate
rlabel metal2 s 7010 0 7066 480 6 chanx_left_out[2]
port 18 nsew default tristate
rlabel metal2 s 7838 0 7894 480 6 chanx_left_out[3]
port 19 nsew default tristate
rlabel metal2 s 8666 0 8722 480 6 chanx_left_out[4]
port 20 nsew default tristate
rlabel metal3 s 0 4904 480 5024 6 chanx_left_out[5]
port 21 nsew default tristate
rlabel metal3 s 23520 8032 24000 8152 6 chanx_left_out[6]
port 22 nsew default tristate
rlabel metal2 s 4618 23520 4674 24000 6 chanx_left_out[7]
port 23 nsew default tristate
rlabel metal2 s 9494 0 9550 480 6 chanx_left_out[8]
port 24 nsew default tristate
rlabel metal2 s 5998 23520 6054 24000 6 chanx_right_in[0]
port 25 nsew default input
rlabel metal3 s 23520 9256 24000 9376 6 chanx_right_in[1]
port 26 nsew default input
rlabel metal2 s 7286 23520 7342 24000 6 chanx_right_in[2]
port 27 nsew default input
rlabel metal2 s 10322 0 10378 480 6 chanx_right_in[3]
port 28 nsew default input
rlabel metal2 s 11150 0 11206 480 6 chanx_right_in[4]
port 29 nsew default input
rlabel metal2 s 11978 0 12034 480 6 chanx_right_in[5]
port 30 nsew default input
rlabel metal3 s 0 6264 480 6384 6 chanx_right_in[6]
port 31 nsew default input
rlabel metal3 s 0 7624 480 7744 6 chanx_right_in[7]
port 32 nsew default input
rlabel metal2 s 8666 23520 8722 24000 6 chanx_right_in[8]
port 33 nsew default input
rlabel metal3 s 0 9120 480 9240 6 chanx_right_out[0]
port 34 nsew default tristate
rlabel metal2 s 9954 23520 10010 24000 6 chanx_right_out[1]
port 35 nsew default tristate
rlabel metal3 s 23520 10616 24000 10736 6 chanx_right_out[2]
port 36 nsew default tristate
rlabel metal3 s 0 10480 480 10600 6 chanx_right_out[3]
port 37 nsew default tristate
rlabel metal3 s 23520 11840 24000 11960 6 chanx_right_out[4]
port 38 nsew default tristate
rlabel metal2 s 12806 0 12862 480 6 chanx_right_out[5]
port 39 nsew default tristate
rlabel metal2 s 11334 23520 11390 24000 6 chanx_right_out[6]
port 40 nsew default tristate
rlabel metal3 s 0 11840 480 11960 6 chanx_right_out[7]
port 41 nsew default tristate
rlabel metal3 s 0 13336 480 13456 6 chanx_right_out[8]
port 42 nsew default tristate
rlabel metal2 s 12622 23520 12678 24000 6 chany_top_in[0]
port 43 nsew default input
rlabel metal3 s 23520 13064 24000 13184 6 chany_top_in[1]
port 44 nsew default input
rlabel metal3 s 0 14696 480 14816 6 chany_top_in[2]
port 45 nsew default input
rlabel metal2 s 14002 23520 14058 24000 6 chany_top_in[3]
port 46 nsew default input
rlabel metal3 s 0 16056 480 16176 6 chany_top_in[4]
port 47 nsew default input
rlabel metal2 s 13634 0 13690 480 6 chany_top_in[5]
port 48 nsew default input
rlabel metal2 s 14462 0 14518 480 6 chany_top_in[6]
port 49 nsew default input
rlabel metal2 s 15290 0 15346 480 6 chany_top_in[7]
port 50 nsew default input
rlabel metal2 s 16118 0 16174 480 6 chany_top_in[8]
port 51 nsew default input
rlabel metal2 s 16946 0 17002 480 6 chany_top_out[0]
port 52 nsew default tristate
rlabel metal3 s 0 17552 480 17672 6 chany_top_out[1]
port 53 nsew default tristate
rlabel metal2 s 17774 0 17830 480 6 chany_top_out[2]
port 54 nsew default tristate
rlabel metal2 s 18602 0 18658 480 6 chany_top_out[3]
port 55 nsew default tristate
rlabel metal3 s 23520 14288 24000 14408 6 chany_top_out[4]
port 56 nsew default tristate
rlabel metal3 s 23520 15648 24000 15768 6 chany_top_out[5]
port 57 nsew default tristate
rlabel metal3 s 23520 16872 24000 16992 6 chany_top_out[6]
port 58 nsew default tristate
rlabel metal3 s 0 18912 480 19032 6 chany_top_out[7]
port 59 nsew default tristate
rlabel metal3 s 23520 18096 24000 18216 6 chany_top_out[8]
port 60 nsew default tristate
rlabel metal2 s 1214 0 1270 480 6 data_in
port 61 nsew default input
rlabel metal2 s 386 0 442 480 6 enable
port 62 nsew default input
rlabel metal2 s 16670 23520 16726 24000 6 left_bottom_grid_pin_11_
port 63 nsew default input
rlabel metal2 s 20258 0 20314 480 6 left_bottom_grid_pin_13_
port 64 nsew default input
rlabel metal3 s 23520 21904 24000 22024 6 left_bottom_grid_pin_15_
port 65 nsew default input
rlabel metal3 s 23520 19320 24000 19440 6 left_bottom_grid_pin_1_
port 66 nsew default input
rlabel metal3 s 23520 20680 24000 20800 6 left_bottom_grid_pin_3_
port 67 nsew default input
rlabel metal2 s 15290 23520 15346 24000 6 left_bottom_grid_pin_5_
port 68 nsew default input
rlabel metal2 s 19430 0 19486 480 6 left_bottom_grid_pin_7_
port 69 nsew default input
rlabel metal3 s 0 20272 480 20392 6 left_bottom_grid_pin_9_
port 70 nsew default input
rlabel metal2 s 21086 0 21142 480 6 left_top_grid_pin_10_
port 71 nsew default input
rlabel metal2 s 19338 23520 19394 24000 6 right_bottom_grid_pin_11_
port 72 nsew default input
rlabel metal2 s 20626 23520 20682 24000 6 right_bottom_grid_pin_13_
port 73 nsew default input
rlabel metal2 s 22006 23520 22062 24000 6 right_bottom_grid_pin_15_
port 74 nsew default input
rlabel metal3 s 0 21768 480 21888 6 right_bottom_grid_pin_1_
port 75 nsew default input
rlabel metal3 s 0 23128 480 23248 6 right_bottom_grid_pin_3_
port 76 nsew default input
rlabel metal2 s 21914 0 21970 480 6 right_bottom_grid_pin_5_
port 77 nsew default input
rlabel metal2 s 17958 23520 18014 24000 6 right_bottom_grid_pin_7_
port 78 nsew default input
rlabel metal3 s 23520 23128 24000 23248 6 right_bottom_grid_pin_9_
port 79 nsew default input
rlabel metal2 s 23294 23520 23350 24000 6 right_top_grid_pin_10_
port 80 nsew default input
rlabel metal2 s 22742 0 22798 480 6 top_left_grid_pin_13_
port 81 nsew default input
rlabel metal2 s 23570 0 23626 480 6 top_right_grid_pin_11_
port 82 nsew default input
rlabel metal4 s 4944 2128 5264 21808 6 vpwr
port 83 nsew default input
rlabel metal4 s 8944 2128 9264 21808 6 vgnd
port 84 nsew default input
<< end >>
