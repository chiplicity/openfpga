magic
tech EFS8A
magscale 1 2
timestamp 1602523286
<< locali >>
rect 18705 12631 18739 12733
rect 9631 12257 9758 12291
rect 10735 12257 10770 12291
rect 15703 12257 15830 12291
rect 23523 12257 23558 12291
rect 8677 11679 8711 11849
rect 11069 11543 11103 11645
rect 14105 11611 14139 11713
rect 4663 11169 4698 11203
rect 11805 11169 11966 11203
rect 17601 11169 17762 11203
rect 26467 11169 26594 11203
rect 30975 11169 31102 11203
rect 33275 11169 33402 11203
rect 11805 10999 11839 11169
rect 17601 10999 17635 11169
rect 35299 10081 35334 10115
rect 13277 9911 13311 10081
rect 28089 9367 28123 9469
rect 2599 9129 2605 9163
rect 7291 9129 7297 9163
rect 13823 9129 13829 9163
rect 23483 9129 23489 9163
rect 32499 9129 32505 9163
rect 2599 9061 2633 9129
rect 7291 9061 7325 9129
rect 13823 9061 13857 9129
rect 23483 9061 23517 9129
rect 32499 9061 32533 9129
rect 18613 8415 18647 8585
rect 2599 8279 2633 8347
rect 14743 8279 14777 8347
rect 29923 8279 29957 8347
rect 2599 8245 2605 8279
rect 14743 8245 14749 8279
rect 29923 8245 29929 8279
rect 5819 8041 5825 8075
rect 32499 8041 32505 8075
rect 5819 7973 5853 8041
rect 32499 7973 32533 8041
rect 30659 6953 30665 6987
rect 30659 6885 30693 6953
rect 21315 6817 21350 6851
rect 29923 5865 29929 5899
rect 29923 5797 29957 5865
rect 13179 5015 13213 5083
rect 21643 5015 21677 5083
rect 13179 4981 13185 5015
rect 21643 4981 21649 5015
rect 22011 4777 22017 4811
rect 2547 4709 2592 4743
rect 22011 4709 22045 4777
rect 16589 4641 16703 4675
rect 24995 4641 25030 4675
rect 16589 4607 16623 4641
rect 12081 3927 12115 4029
rect 16037 3927 16071 4029
rect 25455 3553 25490 3587
rect 8309 2839 8343 3145
rect 9321 3145 9413 3179
rect 9229 2839 9263 3009
rect 9321 2975 9355 3145
rect 14013 2839 14047 3145
rect 20085 2907 20119 3077
rect 26893 2839 26927 3009
rect 7021 2363 7055 2601
rect 21131 2465 21211 2499
rect 10701 2295 10735 2465
rect 26709 2295 26743 2465
<< viali >>
rect 18521 12937 18555 12971
rect 28273 12937 28307 12971
rect 31953 12937 31987 12971
rect 35633 12937 35667 12971
rect 1409 12733 1443 12767
rect 7297 12733 7331 12767
rect 8344 12733 8378 12767
rect 8769 12733 8803 12767
rect 18337 12733 18371 12767
rect 18705 12733 18739 12767
rect 28089 12733 28123 12767
rect 31769 12733 31803 12767
rect 32321 12733 32355 12767
rect 35449 12733 35483 12767
rect 36001 12733 36035 12767
rect 7849 12665 7883 12699
rect 1593 12597 1627 12631
rect 1961 12597 1995 12631
rect 7481 12597 7515 12631
rect 8447 12597 8481 12631
rect 18705 12597 18739 12631
rect 18981 12597 19015 12631
rect 28733 12597 28767 12631
rect 1409 12257 1443 12291
rect 6688 12257 6722 12291
rect 7732 12257 7766 12291
rect 9597 12257 9631 12291
rect 10701 12257 10735 12291
rect 15669 12257 15703 12291
rect 16840 12257 16874 12291
rect 18864 12257 18898 12291
rect 19809 12257 19843 12291
rect 23489 12257 23523 12291
rect 24501 12257 24535 12291
rect 27353 12257 27387 12291
rect 2697 12189 2731 12223
rect 17785 12189 17819 12223
rect 1593 12121 1627 12155
rect 15899 12121 15933 12155
rect 6791 12053 6825 12087
rect 7803 12053 7837 12087
rect 9827 12053 9861 12087
rect 10839 12053 10873 12087
rect 16911 12053 16945 12087
rect 18935 12053 18969 12087
rect 19993 12053 20027 12087
rect 23627 12053 23661 12087
rect 24685 12053 24719 12087
rect 27537 12053 27571 12087
rect 1593 11849 1627 11883
rect 2697 11849 2731 11883
rect 8677 11849 8711 11883
rect 8861 11849 8895 11883
rect 17049 11849 17083 11883
rect 23029 11849 23063 11883
rect 35633 11849 35667 11883
rect 6561 11781 6595 11815
rect 2053 11713 2087 11747
rect 20545 11781 20579 11815
rect 25559 11781 25593 11815
rect 9873 11713 9907 11747
rect 14105 11713 14139 11747
rect 15853 11713 15887 11747
rect 25329 11713 25363 11747
rect 1409 11645 1443 11679
rect 2513 11645 2547 11679
rect 7021 11645 7055 11679
rect 7389 11645 7423 11679
rect 8468 11645 8502 11679
rect 8677 11645 8711 11679
rect 9448 11645 9482 11679
rect 10241 11645 10275 11679
rect 10492 11645 10526 11679
rect 11069 11645 11103 11679
rect 13896 11645 13930 11679
rect 6285 11577 6319 11611
rect 18245 11645 18279 11679
rect 18705 11645 18739 11679
rect 19752 11645 19786 11679
rect 20177 11645 20211 11679
rect 22636 11645 22670 11679
rect 24409 11645 24443 11679
rect 25488 11645 25522 11679
rect 35449 11645 35483 11679
rect 36001 11645 36035 11679
rect 14105 11577 14139 11611
rect 14381 11577 14415 11611
rect 17877 11577 17911 11611
rect 19855 11577 19889 11611
rect 25973 11577 26007 11611
rect 3065 11509 3099 11543
rect 7113 11509 7147 11543
rect 7941 11509 7975 11543
rect 8539 11509 8573 11543
rect 9551 11509 9585 11543
rect 10563 11509 10597 11543
rect 10885 11509 10919 11543
rect 11069 11509 11103 11543
rect 11345 11509 11379 11543
rect 13967 11509 14001 11543
rect 14841 11509 14875 11543
rect 16589 11509 16623 11543
rect 18245 11509 18279 11543
rect 19257 11509 19291 11543
rect 22707 11509 22741 11543
rect 23857 11509 23891 11543
rect 24593 11509 24627 11543
rect 24961 11509 24995 11543
rect 27353 11509 27387 11543
rect 27905 11509 27939 11543
rect 1685 11305 1719 11339
rect 4767 11305 4801 11339
rect 5733 11305 5767 11339
rect 8861 11305 8895 11339
rect 15761 11305 15795 11339
rect 16727 11305 16761 11339
rect 19257 11305 19291 11339
rect 23765 11305 23799 11339
rect 24501 11305 24535 11339
rect 33471 11305 33505 11339
rect 8033 11237 8067 11271
rect 17831 11237 17865 11271
rect 2421 11169 2455 11203
rect 2697 11169 2731 11203
rect 4629 11169 4663 11203
rect 5917 11169 5951 11203
rect 6193 11169 6227 11203
rect 9724 11169 9758 11203
rect 10736 11169 10770 11203
rect 14232 11169 14266 11203
rect 15577 11169 15611 11203
rect 16624 11169 16658 11203
rect 19349 11169 19383 11203
rect 19717 11169 19751 11203
rect 20980 11169 21014 11203
rect 23372 11169 23406 11203
rect 24317 11169 24351 11203
rect 25456 11169 25490 11203
rect 26433 11169 26467 11203
rect 28457 11169 28491 11203
rect 28641 11169 28675 11203
rect 30941 11169 30975 11203
rect 32172 11169 32206 11203
rect 33241 11169 33275 11203
rect 2789 11101 2823 11135
rect 7941 11101 7975 11135
rect 6929 11033 6963 11067
rect 8493 11033 8527 11067
rect 10839 11033 10873 11067
rect 12909 11101 12943 11135
rect 18613 11101 18647 11135
rect 22109 11101 22143 11135
rect 28917 11101 28951 11135
rect 25559 11033 25593 11067
rect 3157 10965 3191 10999
rect 7205 10965 7239 10999
rect 9827 10965 9861 10999
rect 11805 10965 11839 10999
rect 12035 10965 12069 10999
rect 12633 10965 12667 10999
rect 14335 10965 14369 10999
rect 16037 10965 16071 10999
rect 17601 10965 17635 10999
rect 18245 10965 18279 10999
rect 20269 10965 20303 10999
rect 21051 10965 21085 10999
rect 23443 10965 23477 10999
rect 25881 10965 25915 10999
rect 26663 10965 26697 10999
rect 27721 10965 27755 10999
rect 29285 10965 29319 10999
rect 31171 10965 31205 10999
rect 32275 10965 32309 10999
rect 6285 10761 6319 10795
rect 9689 10761 9723 10795
rect 10977 10761 11011 10795
rect 21189 10761 21223 10795
rect 26617 10761 26651 10795
rect 32597 10761 32631 10795
rect 2881 10693 2915 10727
rect 13921 10693 13955 10727
rect 15761 10693 15795 10727
rect 19993 10693 20027 10727
rect 31125 10693 31159 10727
rect 3065 10625 3099 10659
rect 7113 10625 7147 10659
rect 7389 10625 7423 10659
rect 8677 10625 8711 10659
rect 8953 10625 8987 10659
rect 14565 10625 14599 10659
rect 20177 10625 20211 10659
rect 23857 10625 23891 10659
rect 29009 10625 29043 10659
rect 31677 10625 31711 10659
rect 33977 10625 34011 10659
rect 1593 10557 1627 10591
rect 1961 10557 1995 10591
rect 5089 10557 5123 10591
rect 5457 10557 5491 10591
rect 5641 10557 5675 10591
rect 6561 10557 6595 10591
rect 10216 10557 10250 10591
rect 11196 10557 11230 10591
rect 11897 10557 11931 10591
rect 12541 10557 12575 10591
rect 13001 10557 13035 10591
rect 14105 10557 14139 10591
rect 14657 10557 14691 10591
rect 15669 10557 15703 10591
rect 15945 10557 15979 10591
rect 18429 10557 18463 10591
rect 18797 10557 18831 10591
rect 19073 10557 19107 10591
rect 22604 10557 22638 10591
rect 23029 10557 23063 10591
rect 24869 10557 24903 10591
rect 25605 10557 25639 10591
rect 26065 10557 26099 10591
rect 27445 10557 27479 10591
rect 27629 10557 27663 10591
rect 28181 10557 28215 10591
rect 29285 10557 29319 10591
rect 29745 10557 29779 10591
rect 33216 10557 33250 10591
rect 33609 10557 33643 10591
rect 2145 10489 2179 10523
rect 3157 10489 3191 10523
rect 3709 10489 3743 10523
rect 7205 10489 7239 10523
rect 8769 10489 8803 10523
rect 13277 10489 13311 10523
rect 17049 10489 17083 10523
rect 19257 10489 19291 10523
rect 20269 10489 20303 10523
rect 20821 10489 20855 10523
rect 23949 10489 23983 10523
rect 24501 10489 24535 10523
rect 26341 10489 26375 10523
rect 28365 10489 28399 10523
rect 30021 10489 30055 10523
rect 31493 10489 31527 10523
rect 31769 10489 31803 10523
rect 32321 10489 32355 10523
rect 2421 10421 2455 10455
rect 4721 10421 4755 10455
rect 5273 10421 5307 10455
rect 8033 10421 8067 10455
rect 8401 10421 8435 10455
rect 10287 10421 10321 10455
rect 10701 10421 10735 10455
rect 11299 10421 11333 10455
rect 13645 10421 13679 10455
rect 15117 10421 15151 10455
rect 15577 10421 15611 10455
rect 16129 10421 16163 10455
rect 16681 10421 16715 10455
rect 17785 10421 17819 10455
rect 19533 10421 19567 10455
rect 22707 10421 22741 10455
rect 23489 10421 23523 10455
rect 25421 10421 25455 10455
rect 28733 10421 28767 10455
rect 33287 10421 33321 10455
rect 1961 10217 1995 10251
rect 2237 10217 2271 10251
rect 3157 10217 3191 10251
rect 5733 10217 5767 10251
rect 7113 10217 7147 10251
rect 8677 10217 8711 10251
rect 11161 10217 11195 10251
rect 13093 10217 13127 10251
rect 13737 10217 13771 10251
rect 17049 10217 17083 10251
rect 17969 10217 18003 10251
rect 22753 10217 22787 10251
rect 27077 10217 27111 10251
rect 31677 10217 31711 10251
rect 1685 10149 1719 10183
rect 4261 10149 4295 10183
rect 7389 10149 7423 10183
rect 7849 10149 7883 10183
rect 9781 10149 9815 10183
rect 9873 10149 9907 10183
rect 15117 10149 15151 10183
rect 15485 10149 15519 10183
rect 18245 10149 18279 10183
rect 21097 10149 21131 10183
rect 24501 10149 24535 10183
rect 27721 10149 27755 10183
rect 27813 10149 27847 10183
rect 32229 10149 32263 10183
rect 32321 10149 32355 10183
rect 33885 10149 33919 10183
rect 2421 10081 2455 10115
rect 2697 10081 2731 10115
rect 5641 10081 5675 10115
rect 6193 10081 6227 10115
rect 12357 10081 12391 10115
rect 12541 10081 12575 10115
rect 13277 10081 13311 10115
rect 13645 10081 13679 10115
rect 14197 10081 14231 10115
rect 16865 10081 16899 10115
rect 19717 10081 19751 10115
rect 22477 10081 22511 10115
rect 22937 10081 22971 10115
rect 24225 10081 24259 10115
rect 26617 10081 26651 10115
rect 29193 10081 29227 10115
rect 29653 10081 29687 10115
rect 30824 10081 30858 10115
rect 35265 10081 35299 10115
rect 4169 10013 4203 10047
rect 7757 10013 7791 10047
rect 8033 10013 8067 10047
rect 10057 10013 10091 10047
rect 12817 10013 12851 10047
rect 4721 9945 4755 9979
rect 15393 10013 15427 10047
rect 16037 10013 16071 10047
rect 18153 10013 18187 10047
rect 21005 10013 21039 10047
rect 24409 10013 24443 10047
rect 24685 10013 24719 10047
rect 28365 10013 28399 10047
rect 29929 10013 29963 10047
rect 32505 10013 32539 10047
rect 33793 10013 33827 10047
rect 34069 10013 34103 10047
rect 18705 9945 18739 9979
rect 21557 9945 21591 9979
rect 30895 9945 30929 9979
rect 33241 9945 33275 9979
rect 5181 9877 5215 9911
rect 13277 9877 13311 9911
rect 13461 9877 13495 9911
rect 14657 9877 14691 9911
rect 19901 9877 19935 9911
rect 20177 9877 20211 9911
rect 23765 9877 23799 9911
rect 25697 9877 25731 9911
rect 26801 9877 26835 9911
rect 28641 9877 28675 9911
rect 30665 9877 30699 9911
rect 35403 9877 35437 9911
rect 6101 9673 6135 9707
rect 8217 9673 8251 9707
rect 8585 9673 8619 9707
rect 10149 9673 10183 9707
rect 11253 9673 11287 9707
rect 15393 9673 15427 9707
rect 17233 9673 17267 9707
rect 20729 9673 20763 9707
rect 21097 9673 21131 9707
rect 27905 9673 27939 9707
rect 30481 9673 30515 9707
rect 32229 9673 32263 9707
rect 33793 9673 33827 9707
rect 35265 9673 35299 9707
rect 36001 9673 36035 9707
rect 7941 9605 7975 9639
rect 9873 9605 9907 9639
rect 13737 9605 13771 9639
rect 14381 9605 14415 9639
rect 21373 9605 21407 9639
rect 24685 9605 24719 9639
rect 34069 9605 34103 9639
rect 35633 9605 35667 9639
rect 2605 9537 2639 9571
rect 4721 9537 4755 9571
rect 7021 9537 7055 9571
rect 8861 9537 8895 9571
rect 10471 9537 10505 9571
rect 12541 9537 12575 9571
rect 12817 9537 12851 9571
rect 18061 9537 18095 9571
rect 19809 9537 19843 9571
rect 21649 9537 21683 9571
rect 21925 9537 21959 9571
rect 23765 9537 23799 9571
rect 24409 9537 24443 9571
rect 25605 9537 25639 9571
rect 26985 9537 27019 9571
rect 29699 9537 29733 9571
rect 30665 9537 30699 9571
rect 30941 9537 30975 9571
rect 32413 9537 32447 9571
rect 32689 9537 32723 9571
rect 1409 9469 1443 9503
rect 1961 9469 1995 9503
rect 3525 9469 3559 9503
rect 10384 9469 10418 9503
rect 11412 9469 11446 9503
rect 11805 9469 11839 9503
rect 14473 9469 14507 9503
rect 15761 9469 15795 9503
rect 16497 9469 16531 9503
rect 16681 9469 16715 9503
rect 18981 9469 19015 9503
rect 28089 9469 28123 9503
rect 28641 9469 28675 9503
rect 29612 9469 29646 9503
rect 35449 9469 35483 9503
rect 2926 9401 2960 9435
rect 4169 9401 4203 9435
rect 4445 9401 4479 9435
rect 4537 9401 4571 9435
rect 7342 9401 7376 9435
rect 8953 9401 8987 9435
rect 9505 9401 9539 9435
rect 12633 9401 12667 9435
rect 14835 9401 14869 9435
rect 16037 9401 16071 9435
rect 16957 9401 16991 9435
rect 17877 9401 17911 9435
rect 18423 9401 18457 9435
rect 19717 9401 19751 9435
rect 20130 9401 20164 9435
rect 21741 9401 21775 9435
rect 23857 9401 23891 9435
rect 25329 9401 25363 9435
rect 25421 9401 25455 9435
rect 26341 9401 26375 9435
rect 27077 9401 27111 9435
rect 27629 9401 27663 9435
rect 30757 9401 30791 9435
rect 32505 9401 32539 9435
rect 1593 9333 1627 9367
rect 2513 9333 2547 9367
rect 3801 9333 3835 9367
rect 5641 9333 5675 9367
rect 6561 9333 6595 9367
rect 10885 9333 10919 9367
rect 11483 9333 11517 9367
rect 12265 9333 12299 9367
rect 19257 9333 19291 9367
rect 22569 9333 22603 9367
rect 23029 9333 23063 9367
rect 23489 9333 23523 9367
rect 25053 9333 25087 9367
rect 26617 9333 26651 9367
rect 28089 9333 28123 9367
rect 28273 9333 28307 9367
rect 29009 9333 29043 9367
rect 30113 9333 30147 9367
rect 31677 9333 31711 9367
rect 33333 9333 33367 9367
rect 2053 9129 2087 9163
rect 2605 9129 2639 9163
rect 3157 9129 3191 9163
rect 3893 9129 3927 9163
rect 4997 9129 5031 9163
rect 6101 9129 6135 9163
rect 6837 9129 6871 9163
rect 7297 9129 7331 9163
rect 7849 9129 7883 9163
rect 8861 9129 8895 9163
rect 13829 9129 13863 9163
rect 15025 9129 15059 9163
rect 16957 9129 16991 9163
rect 18153 9129 18187 9163
rect 18429 9129 18463 9163
rect 20269 9129 20303 9163
rect 20729 9129 20763 9163
rect 21925 9129 21959 9163
rect 23489 9129 23523 9163
rect 24409 9129 24443 9163
rect 24961 9129 24995 9163
rect 25881 9129 25915 9163
rect 27445 9129 27479 9163
rect 29561 9129 29595 9163
rect 31861 9129 31895 9163
rect 32505 9129 32539 9163
rect 33057 9129 33091 9163
rect 3433 9061 3467 9095
rect 4629 9061 4663 9095
rect 5543 9061 5577 9095
rect 9873 9061 9907 9095
rect 11989 9061 12023 9095
rect 12081 9061 12115 9095
rect 14749 9061 14783 9095
rect 15485 9061 15519 9095
rect 16405 9061 16439 9095
rect 19435 9061 19469 9095
rect 21097 9061 21131 9095
rect 26887 9061 26921 9095
rect 28457 9061 28491 9095
rect 29009 9061 29043 9095
rect 30573 9061 30607 9095
rect 30665 9061 30699 9095
rect 34529 9061 34563 9095
rect 2237 8993 2271 9027
rect 4077 8993 4111 9027
rect 5181 8993 5215 9027
rect 13461 8993 13495 9027
rect 16865 8993 16899 9027
rect 17417 8993 17451 9027
rect 19073 8993 19107 9027
rect 19993 8993 20027 9027
rect 25145 8993 25179 9027
rect 25329 8993 25363 9027
rect 32137 8993 32171 9027
rect 35909 8993 35943 9027
rect 6929 8925 6963 8959
rect 9781 8925 9815 8959
rect 12633 8925 12667 8959
rect 15393 8925 15427 8959
rect 16037 8925 16071 8959
rect 21005 8925 21039 8959
rect 23121 8925 23155 8959
rect 24685 8925 24719 8959
rect 26525 8925 26559 8959
rect 28365 8925 28399 8959
rect 30849 8925 30883 8959
rect 34437 8925 34471 8959
rect 35081 8925 35115 8959
rect 4261 8857 4295 8891
rect 10333 8857 10367 8891
rect 14381 8857 14415 8891
rect 21557 8857 21591 8891
rect 24041 8857 24075 8891
rect 8309 8789 8343 8823
rect 13001 8789 13035 8823
rect 18981 8789 19015 8823
rect 36093 8789 36127 8823
rect 3157 8585 3191 8619
rect 3893 8585 3927 8619
rect 7343 8585 7377 8619
rect 7757 8585 7791 8619
rect 9137 8585 9171 8619
rect 9505 8585 9539 8619
rect 9873 8585 9907 8619
rect 11069 8585 11103 8619
rect 11529 8585 11563 8619
rect 11897 8585 11931 8619
rect 13369 8585 13403 8619
rect 15301 8585 15335 8619
rect 15577 8585 15611 8619
rect 17509 8585 17543 8619
rect 18613 8585 18647 8619
rect 18889 8585 18923 8619
rect 20269 8585 20303 8619
rect 22109 8585 22143 8619
rect 22845 8585 22879 8619
rect 25697 8585 25731 8619
rect 27445 8585 27479 8619
rect 28365 8585 28399 8619
rect 31125 8585 31159 8619
rect 33241 8585 33275 8619
rect 37611 8585 37645 8619
rect 3433 8517 3467 8551
rect 10609 8517 10643 8551
rect 2237 8449 2271 8483
rect 4353 8449 4387 8483
rect 8217 8449 8251 8483
rect 14381 8449 14415 8483
rect 16497 8449 16531 8483
rect 17141 8449 17175 8483
rect 20545 8517 20579 8551
rect 30849 8517 30883 8551
rect 35909 8517 35943 8551
rect 19349 8449 19383 8483
rect 26525 8449 26559 8483
rect 27721 8449 27755 8483
rect 28641 8449 28675 8483
rect 29561 8449 29595 8483
rect 31677 8449 31711 8483
rect 34621 8449 34655 8483
rect 34989 8449 35023 8483
rect 35265 8449 35299 8483
rect 36921 8449 36955 8483
rect 5616 8381 5650 8415
rect 6009 8381 6043 8415
rect 7272 8381 7306 8415
rect 12449 8381 12483 8415
rect 18388 8381 18422 8415
rect 18613 8381 18647 8415
rect 20913 8381 20947 8415
rect 21097 8381 21131 8415
rect 21557 8381 21591 8415
rect 23816 8381 23850 8415
rect 24317 8381 24351 8415
rect 24777 8381 24811 8415
rect 30481 8381 30515 8415
rect 32597 8381 32631 8415
rect 33609 8381 33643 8415
rect 33860 8381 33894 8415
rect 34253 8381 34287 8415
rect 36496 8381 36530 8415
rect 37540 8381 37574 8415
rect 4077 8313 4111 8347
rect 4169 8313 4203 8347
rect 5181 8313 5215 8347
rect 7021 8313 7055 8347
rect 8033 8313 8067 8347
rect 8538 8313 8572 8347
rect 10057 8313 10091 8347
rect 10149 8313 10183 8347
rect 12265 8313 12299 8347
rect 12770 8313 12804 8347
rect 13645 8313 13679 8347
rect 16589 8313 16623 8347
rect 18475 8313 18509 8347
rect 19711 8313 19745 8347
rect 21833 8313 21867 8347
rect 23903 8313 23937 8347
rect 25139 8313 25173 8347
rect 26065 8313 26099 8347
rect 26433 8313 26467 8347
rect 26887 8313 26921 8347
rect 32039 8313 32073 8347
rect 35081 8313 35115 8347
rect 1777 8245 1811 8279
rect 2145 8245 2179 8279
rect 2605 8245 2639 8279
rect 5687 8245 5721 8279
rect 6653 8245 6687 8279
rect 14289 8245 14323 8279
rect 14749 8245 14783 8279
rect 16221 8245 16255 8279
rect 19257 8245 19291 8279
rect 23213 8245 23247 8279
rect 24685 8245 24719 8279
rect 29929 8245 29963 8279
rect 31585 8245 31619 8279
rect 32873 8245 32907 8279
rect 33931 8245 33965 8279
rect 36599 8245 36633 8279
rect 38025 8245 38059 8279
rect 2145 8041 2179 8075
rect 3893 8041 3927 8075
rect 4261 8041 4295 8075
rect 4629 8041 4663 8075
rect 5181 8041 5215 8075
rect 5825 8041 5859 8075
rect 11345 8041 11379 8075
rect 13553 8041 13587 8075
rect 14657 8041 14691 8075
rect 15117 8041 15151 8075
rect 16497 8041 16531 8075
rect 17785 8041 17819 8075
rect 18153 8041 18187 8075
rect 19073 8041 19107 8075
rect 22569 8041 22603 8075
rect 23949 8041 23983 8075
rect 26341 8041 26375 8075
rect 26617 8041 26651 8075
rect 29653 8041 29687 8075
rect 30849 8041 30883 8075
rect 31677 8041 31711 8075
rect 32505 8041 32539 8075
rect 34253 8041 34287 8075
rect 35357 8041 35391 8075
rect 2421 7973 2455 8007
rect 8217 7973 8251 8007
rect 9781 7973 9815 8007
rect 9873 7973 9907 8007
rect 10425 7973 10459 8007
rect 13829 7973 13863 8007
rect 15485 7973 15519 8007
rect 16037 7973 16071 8007
rect 17227 7973 17261 8007
rect 20729 7973 20763 8007
rect 23115 7973 23149 8007
rect 24593 7973 24627 8007
rect 24685 7973 24719 8007
rect 30250 7973 30284 8007
rect 34437 7973 34471 8007
rect 34529 7973 34563 8007
rect 35081 7973 35115 8007
rect 36001 7973 36035 8007
rect 36093 7973 36127 8007
rect 4077 7905 4111 7939
rect 5457 7905 5491 7939
rect 6377 7905 6411 7939
rect 8769 7905 8803 7939
rect 11529 7905 11563 7939
rect 11805 7905 11839 7939
rect 16865 7905 16899 7939
rect 18981 7905 19015 7939
rect 19441 7905 19475 7939
rect 21189 7905 21223 7939
rect 21373 7905 21407 7939
rect 22753 7905 22787 7939
rect 23673 7905 23707 7939
rect 26525 7905 26559 7939
rect 26985 7905 27019 7939
rect 28365 7905 28399 7939
rect 28825 7905 28859 7939
rect 29101 7905 29135 7939
rect 2329 7837 2363 7871
rect 2973 7837 3007 7871
rect 8125 7837 8159 7871
rect 13737 7837 13771 7871
rect 14381 7837 14415 7871
rect 15393 7837 15427 7871
rect 18889 7837 18923 7871
rect 21649 7837 21683 7871
rect 21925 7837 21959 7871
rect 24869 7837 24903 7871
rect 29929 7837 29963 7871
rect 32137 7837 32171 7871
rect 36277 7837 36311 7871
rect 28181 7769 28215 7803
rect 1777 7701 1811 7735
rect 10701 7701 10735 7735
rect 12541 7701 12575 7735
rect 20085 7701 20119 7735
rect 24409 7701 24443 7735
rect 25513 7701 25547 7735
rect 27721 7701 27755 7735
rect 33057 7701 33091 7735
rect 2237 7497 2271 7531
rect 3709 7497 3743 7531
rect 4813 7497 4847 7531
rect 5181 7497 5215 7531
rect 8125 7497 8159 7531
rect 8677 7497 8711 7531
rect 11713 7497 11747 7531
rect 15301 7497 15335 7531
rect 17325 7497 17359 7531
rect 17785 7497 17819 7531
rect 19073 7497 19107 7531
rect 19441 7497 19475 7531
rect 19901 7497 19935 7531
rect 23213 7497 23247 7531
rect 24777 7497 24811 7531
rect 27445 7497 27479 7531
rect 29009 7497 29043 7531
rect 33701 7497 33735 7531
rect 34345 7497 34379 7531
rect 36277 7497 36311 7531
rect 36645 7497 36679 7531
rect 5779 7429 5813 7463
rect 13277 7429 13311 7463
rect 17049 7429 17083 7463
rect 18705 7429 18739 7463
rect 22845 7429 22879 7463
rect 38025 7429 38059 7463
rect 2421 7361 2455 7395
rect 8861 7361 8895 7395
rect 12909 7361 12943 7395
rect 15025 7361 15059 7395
rect 16037 7361 16071 7395
rect 18153 7361 18187 7395
rect 21189 7361 21223 7395
rect 21649 7361 21683 7395
rect 23765 7361 23799 7395
rect 25329 7361 25363 7395
rect 30021 7361 30055 7395
rect 31217 7361 31251 7395
rect 34621 7361 34655 7395
rect 35265 7361 35299 7395
rect 36001 7361 36035 7395
rect 3065 7293 3099 7327
rect 3893 7293 3927 7327
rect 5708 7293 5742 7327
rect 6101 7293 6135 7327
rect 6653 7293 6687 7327
rect 7113 7293 7147 7327
rect 7297 7293 7331 7327
rect 10609 7293 10643 7327
rect 11161 7293 11195 7327
rect 13369 7293 13403 7327
rect 14289 7293 14323 7327
rect 20085 7293 20119 7327
rect 20637 7293 20671 7327
rect 22569 7293 22603 7327
rect 24409 7293 24443 7327
rect 27629 7293 27663 7327
rect 28181 7293 28215 7327
rect 29285 7293 29319 7327
rect 29745 7293 29779 7327
rect 30665 7293 30699 7327
rect 31769 7293 31803 7327
rect 33828 7293 33862 7327
rect 36461 7293 36495 7327
rect 37013 7293 37047 7327
rect 37611 7293 37645 7327
rect 1869 7225 1903 7259
rect 2513 7225 2547 7259
rect 4255 7225 4289 7259
rect 9182 7225 9216 7259
rect 10517 7225 10551 7259
rect 13731 7225 13765 7259
rect 14565 7225 14599 7259
rect 16129 7225 16163 7259
rect 16681 7225 16715 7259
rect 18245 7225 18279 7259
rect 20821 7225 20855 7259
rect 21557 7225 21591 7259
rect 22011 7225 22045 7259
rect 23857 7225 23891 7259
rect 25421 7225 25455 7259
rect 25973 7225 26007 7259
rect 28365 7225 28399 7259
rect 32131 7225 32165 7259
rect 32965 7225 32999 7259
rect 33931 7225 33965 7259
rect 34989 7225 35023 7259
rect 35081 7225 35115 7259
rect 3341 7157 3375 7191
rect 5457 7157 5491 7191
rect 6929 7157 6963 7191
rect 9781 7157 9815 7191
rect 10057 7157 10091 7191
rect 10701 7157 10735 7191
rect 12081 7157 12115 7191
rect 15761 7157 15795 7191
rect 25145 7157 25179 7191
rect 26525 7157 26559 7191
rect 26893 7157 26927 7191
rect 28733 7157 28767 7191
rect 30389 7157 30423 7191
rect 31585 7157 31619 7191
rect 32689 7157 32723 7191
rect 37703 7157 37737 7191
rect 1961 6953 1995 6987
rect 3893 6953 3927 6987
rect 6837 6953 6871 6987
rect 9137 6953 9171 6987
rect 9505 6953 9539 6987
rect 9873 6953 9907 6987
rect 13369 6953 13403 6987
rect 15117 6953 15151 6987
rect 16773 6953 16807 6987
rect 20177 6953 20211 6987
rect 22109 6953 22143 6987
rect 23765 6953 23799 6987
rect 25237 6953 25271 6987
rect 25605 6953 25639 6987
rect 27629 6953 27663 6987
rect 28457 6953 28491 6987
rect 30665 6953 30699 6987
rect 31217 6953 31251 6987
rect 34161 6953 34195 6987
rect 35265 6953 35299 6987
rect 2329 6885 2363 6919
rect 2605 6885 2639 6919
rect 4261 6885 4295 6919
rect 4813 6885 4847 6919
rect 5825 6885 5859 6919
rect 8125 6885 8159 6919
rect 8217 6885 8251 6919
rect 10425 6885 10459 6919
rect 10517 6885 10551 6919
rect 12633 6885 12667 6919
rect 13823 6885 13857 6919
rect 15393 6885 15427 6919
rect 15485 6885 15519 6919
rect 17049 6885 17083 6919
rect 17141 6885 17175 6919
rect 18705 6885 18739 6919
rect 21097 6885 21131 6919
rect 22655 6885 22689 6919
rect 24225 6885 24259 6919
rect 26617 6885 26651 6919
rect 26709 6885 26743 6919
rect 28917 6885 28951 6919
rect 32499 6885 32533 6919
rect 34437 6885 34471 6919
rect 36001 6885 36035 6919
rect 36553 6885 36587 6919
rect 1476 6817 1510 6851
rect 11989 6817 12023 6851
rect 12449 6817 12483 6851
rect 13461 6817 13495 6851
rect 21281 6817 21315 6851
rect 21741 6817 21775 6851
rect 22293 6817 22327 6851
rect 23213 6817 23247 6851
rect 30297 6817 30331 6851
rect 32137 6817 32171 6851
rect 2513 6749 2547 6783
rect 4169 6749 4203 6783
rect 5733 6749 5767 6783
rect 6009 6749 6043 6783
rect 8401 6749 8435 6783
rect 10701 6749 10735 6783
rect 17325 6749 17359 6783
rect 18613 6749 18647 6783
rect 18889 6749 18923 6783
rect 24133 6749 24167 6783
rect 24777 6749 24811 6783
rect 26893 6749 26927 6783
rect 28825 6749 28859 6783
rect 29469 6749 29503 6783
rect 34345 6749 34379 6783
rect 34989 6749 35023 6783
rect 35909 6749 35943 6783
rect 1547 6681 1581 6715
rect 3065 6681 3099 6715
rect 7941 6681 7975 6715
rect 14381 6681 14415 6715
rect 15945 6681 15979 6715
rect 21419 6681 21453 6715
rect 3433 6613 3467 6647
rect 7297 6613 7331 6647
rect 12909 6613 12943 6647
rect 16313 6613 16347 6647
rect 18153 6613 18187 6647
rect 19533 6613 19567 6647
rect 30205 6613 30239 6647
rect 31769 6613 31803 6647
rect 33057 6613 33091 6647
rect 1869 6409 1903 6443
rect 5641 6409 5675 6443
rect 6285 6409 6319 6443
rect 8861 6409 8895 6443
rect 11621 6409 11655 6443
rect 13829 6409 13863 6443
rect 15393 6409 15427 6443
rect 17785 6409 17819 6443
rect 19073 6409 19107 6443
rect 19717 6409 19751 6443
rect 22661 6409 22695 6443
rect 24685 6409 24719 6443
rect 25053 6409 25087 6443
rect 26893 6409 26927 6443
rect 27353 6409 27387 6443
rect 28825 6409 28859 6443
rect 29469 6409 29503 6443
rect 33333 6409 33367 6443
rect 34253 6409 34287 6443
rect 34621 6409 34655 6443
rect 35909 6409 35943 6443
rect 36369 6409 36403 6443
rect 37013 6409 37047 6443
rect 2329 6341 2363 6375
rect 3065 6341 3099 6375
rect 15669 6341 15703 6375
rect 17141 6341 17175 6375
rect 22937 6341 22971 6375
rect 26525 6341 26559 6375
rect 36599 6341 36633 6375
rect 2513 6273 2547 6307
rect 5871 6273 5905 6307
rect 17417 6273 17451 6307
rect 18153 6273 18187 6307
rect 19993 6273 20027 6307
rect 21741 6273 21775 6307
rect 23765 6273 23799 6307
rect 25329 6273 25363 6307
rect 25973 6273 26007 6307
rect 28273 6273 28307 6307
rect 30665 6273 30699 6307
rect 30941 6273 30975 6307
rect 32137 6273 32171 6307
rect 33701 6273 33735 6307
rect 34989 6273 35023 6307
rect 35357 6273 35391 6307
rect 1460 6205 1494 6239
rect 3985 6205 4019 6239
rect 5784 6205 5818 6239
rect 7297 6205 7331 6239
rect 9781 6205 9815 6239
rect 12725 6205 12759 6239
rect 13001 6205 13035 6239
rect 14473 6205 14507 6239
rect 16221 6205 16255 6239
rect 20177 6205 20211 6239
rect 20637 6205 20671 6239
rect 23397 6205 23431 6239
rect 27537 6205 27571 6239
rect 28089 6205 28123 6239
rect 29285 6205 29319 6239
rect 29745 6205 29779 6239
rect 36528 6205 36562 6239
rect 1547 6137 1581 6171
rect 2605 6137 2639 6171
rect 3525 6137 3559 6171
rect 4347 6137 4381 6171
rect 7618 6137 7652 6171
rect 9689 6137 9723 6171
rect 10143 6137 10177 6171
rect 14381 6137 14415 6171
rect 14835 6137 14869 6171
rect 16129 6137 16163 6171
rect 16583 6137 16617 6171
rect 18245 6137 18279 6171
rect 18797 6137 18831 6171
rect 20913 6137 20947 6171
rect 22103 6137 22137 6171
rect 23857 6137 23891 6171
rect 24409 6137 24443 6171
rect 25421 6137 25455 6171
rect 30757 6137 30791 6171
rect 32458 6137 32492 6171
rect 35081 6137 35115 6171
rect 3893 6069 3927 6103
rect 4905 6069 4939 6103
rect 5273 6069 5307 6103
rect 7113 6069 7147 6103
rect 8217 6069 8251 6103
rect 8493 6069 8527 6103
rect 9229 6069 9263 6103
rect 10701 6069 10735 6103
rect 10977 6069 11011 6103
rect 11989 6069 12023 6103
rect 12541 6069 12575 6103
rect 13461 6069 13495 6103
rect 21373 6069 21407 6103
rect 30297 6069 30331 6103
rect 31585 6069 31619 6103
rect 31953 6069 31987 6103
rect 33057 6069 33091 6103
rect 3157 5865 3191 5899
rect 3525 5865 3559 5899
rect 5641 5865 5675 5899
rect 9965 5865 9999 5899
rect 11805 5865 11839 5899
rect 15025 5865 15059 5899
rect 15945 5865 15979 5899
rect 18061 5865 18095 5899
rect 18797 5865 18831 5899
rect 22385 5865 22419 5899
rect 22661 5865 22695 5899
rect 23121 5865 23155 5899
rect 24869 5865 24903 5899
rect 29929 5865 29963 5899
rect 31125 5865 31159 5899
rect 34897 5865 34931 5899
rect 35265 5865 35299 5899
rect 2558 5797 2592 5831
rect 4261 5797 4295 5831
rect 4813 5797 4847 5831
rect 6653 5797 6687 5831
rect 7205 5797 7239 5831
rect 8217 5797 8251 5831
rect 10609 5797 10643 5831
rect 12173 5797 12207 5831
rect 14381 5797 14415 5831
rect 16865 5797 16899 5831
rect 16957 5797 16991 5831
rect 18429 5797 18463 5831
rect 21827 5797 21861 5831
rect 23397 5797 23431 5831
rect 27261 5797 27295 5831
rect 30849 5797 30883 5831
rect 32321 5797 32355 5831
rect 33977 5797 34011 5831
rect 34529 5797 34563 5831
rect 13921 5729 13955 5763
rect 14197 5729 14231 5763
rect 15761 5729 15795 5763
rect 19257 5729 19291 5763
rect 19809 5729 19843 5763
rect 24777 5729 24811 5763
rect 25237 5729 25271 5763
rect 30481 5729 30515 5763
rect 2237 5661 2271 5695
rect 4169 5661 4203 5695
rect 6561 5661 6595 5695
rect 8114 5661 8148 5695
rect 8769 5661 8803 5695
rect 10333 5661 10367 5695
rect 10517 5661 10551 5695
rect 10793 5661 10827 5695
rect 12081 5661 12115 5695
rect 12357 5661 12391 5695
rect 14749 5661 14783 5695
rect 19993 5661 20027 5695
rect 21281 5661 21315 5695
rect 21465 5661 21499 5695
rect 23305 5661 23339 5695
rect 23949 5661 23983 5695
rect 27169 5661 27203 5695
rect 27813 5661 27847 5695
rect 29561 5661 29595 5695
rect 32229 5661 32263 5695
rect 33885 5661 33919 5695
rect 35357 5661 35391 5695
rect 17417 5593 17451 5627
rect 32781 5593 32815 5627
rect 1777 5525 1811 5559
rect 2145 5525 2179 5559
rect 3801 5525 3835 5559
rect 6285 5525 6319 5559
rect 13001 5525 13035 5559
rect 13369 5525 13403 5559
rect 15577 5525 15611 5559
rect 16497 5525 16531 5559
rect 24225 5525 24259 5559
rect 24685 5525 24719 5559
rect 28733 5525 28767 5559
rect 3341 5321 3375 5355
rect 3985 5321 4019 5355
rect 4721 5321 4755 5355
rect 6561 5321 6595 5355
rect 8125 5321 8159 5355
rect 8401 5321 8435 5355
rect 10149 5321 10183 5355
rect 11897 5321 11931 5355
rect 14105 5321 14139 5355
rect 14381 5321 14415 5355
rect 17049 5321 17083 5355
rect 19257 5321 19291 5355
rect 22201 5321 22235 5355
rect 23121 5321 23155 5355
rect 25237 5321 25271 5355
rect 28641 5321 28675 5355
rect 31953 5321 31987 5355
rect 33425 5321 33459 5355
rect 33885 5321 33919 5355
rect 34161 5321 34195 5355
rect 1547 5253 1581 5287
rect 8769 5253 8803 5287
rect 12265 5253 12299 5287
rect 13737 5253 13771 5287
rect 22477 5253 22511 5287
rect 26617 5253 26651 5287
rect 27445 5253 27479 5287
rect 29469 5253 29503 5287
rect 2421 5185 2455 5219
rect 4307 5185 4341 5219
rect 7205 5185 7239 5219
rect 9321 5185 9355 5219
rect 10609 5185 10643 5219
rect 12817 5185 12851 5219
rect 15301 5185 15335 5219
rect 16129 5185 16163 5219
rect 20729 5185 20763 5219
rect 21281 5185 21315 5219
rect 23397 5185 23431 5219
rect 23765 5185 23799 5219
rect 27169 5185 27203 5219
rect 28365 5185 28399 5219
rect 32781 5185 32815 5219
rect 1476 5117 1510 5151
rect 1869 5117 1903 5151
rect 4220 5117 4254 5151
rect 5089 5117 5123 5151
rect 5457 5117 5491 5151
rect 5733 5117 5767 5151
rect 14841 5117 14875 5151
rect 15025 5117 15059 5151
rect 17785 5117 17819 5151
rect 18061 5117 18095 5151
rect 18521 5117 18555 5151
rect 19717 5117 19751 5151
rect 20177 5117 20211 5151
rect 25697 5117 25731 5151
rect 27629 5117 27663 5151
rect 28089 5117 28123 5151
rect 29285 5117 29319 5151
rect 30113 5117 30147 5151
rect 30665 5117 30699 5151
rect 31585 5117 31619 5151
rect 32229 5117 32263 5151
rect 35484 5117 35518 5151
rect 35909 5117 35943 5151
rect 2329 5049 2363 5083
rect 2783 5049 2817 5083
rect 7526 5049 7560 5083
rect 9045 5049 9079 5083
rect 9137 5049 9171 5083
rect 10517 5049 10551 5083
rect 10971 5049 11005 5083
rect 16037 5049 16071 5083
rect 16450 5049 16484 5083
rect 20453 5049 20487 5083
rect 23857 5049 23891 5083
rect 24409 5049 24443 5083
rect 26018 5049 26052 5083
rect 30986 5049 31020 5083
rect 32505 5049 32539 5083
rect 32597 5049 32631 5083
rect 35587 5049 35621 5083
rect 3709 4981 3743 5015
rect 5457 4981 5491 5015
rect 7021 4981 7055 5015
rect 11529 4981 11563 5015
rect 12725 4981 12759 5015
rect 13185 4981 13219 5015
rect 15577 4981 15611 5015
rect 17325 4981 17359 5015
rect 18153 4981 18187 5015
rect 21189 4981 21223 5015
rect 21649 4981 21683 5015
rect 24869 4981 24903 5015
rect 25605 4981 25639 5015
rect 29009 4981 29043 5015
rect 29837 4981 29871 5015
rect 30481 4981 30515 5015
rect 2145 4777 2179 4811
rect 4169 4777 4203 4811
rect 7941 4777 7975 4811
rect 9873 4777 9907 4811
rect 10241 4777 10275 4811
rect 13921 4777 13955 4811
rect 14657 4777 14691 4811
rect 17141 4777 17175 4811
rect 19809 4777 19843 4811
rect 20177 4777 20211 4811
rect 21557 4777 21591 4811
rect 22017 4777 22051 4811
rect 22569 4777 22603 4811
rect 26709 4777 26743 4811
rect 29285 4777 29319 4811
rect 30757 4777 30791 4811
rect 33885 4777 33919 4811
rect 2513 4709 2547 4743
rect 3801 4709 3835 4743
rect 5962 4709 5996 4743
rect 8769 4709 8803 4743
rect 10977 4709 11011 4743
rect 11253 4709 11287 4743
rect 15301 4709 15335 4743
rect 23305 4709 23339 4743
rect 23581 4709 23615 4743
rect 25099 4709 25133 4743
rect 28175 4709 28209 4743
rect 29882 4709 29916 4743
rect 32321 4709 32355 4743
rect 2237 4641 2271 4675
rect 4077 4641 4111 4675
rect 4629 4641 4663 4675
rect 8309 4641 8343 4675
rect 8585 4641 8619 4675
rect 10057 4641 10091 4675
rect 13093 4641 13127 4675
rect 13277 4641 13311 4675
rect 15485 4641 15519 4675
rect 16957 4641 16991 4675
rect 17693 4641 17727 4675
rect 18797 4641 18831 4675
rect 19073 4641 19107 4675
rect 19533 4641 19567 4675
rect 24961 4641 24995 4675
rect 26525 4641 26559 4675
rect 33701 4641 33735 4675
rect 34780 4641 34814 4675
rect 5641 4573 5675 4607
rect 9045 4573 9079 4607
rect 11161 4573 11195 4607
rect 11437 4573 11471 4607
rect 13369 4573 13403 4607
rect 15853 4573 15887 4607
rect 16405 4573 16439 4607
rect 16589 4573 16623 4607
rect 18429 4573 18463 4607
rect 21649 4573 21683 4607
rect 23489 4573 23523 4607
rect 23949 4573 23983 4607
rect 27629 4573 27663 4607
rect 27813 4573 27847 4607
rect 29561 4573 29595 4607
rect 32229 4573 32263 4607
rect 12173 4505 12207 4539
rect 16773 4505 16807 4539
rect 18889 4505 18923 4539
rect 32781 4505 32815 4539
rect 1685 4437 1719 4471
rect 3157 4437 3191 4471
rect 5273 4437 5307 4471
rect 6561 4437 6595 4471
rect 6837 4437 6871 4471
rect 7297 4437 7331 4471
rect 10609 4437 10643 4471
rect 12541 4437 12575 4471
rect 15025 4437 15059 4471
rect 18153 4437 18187 4471
rect 25789 4437 25823 4471
rect 27261 4437 27295 4471
rect 28733 4437 28767 4471
rect 30481 4437 30515 4471
rect 33149 4437 33183 4471
rect 34851 4437 34885 4471
rect 2513 4233 2547 4267
rect 6101 4233 6135 4267
rect 8125 4233 8159 4267
rect 14013 4233 14047 4267
rect 21925 4233 21959 4267
rect 23029 4233 23063 4267
rect 26525 4233 26559 4267
rect 28457 4233 28491 4267
rect 29101 4233 29135 4267
rect 30297 4233 30331 4267
rect 32229 4233 32263 4267
rect 32873 4233 32907 4267
rect 4629 4165 4663 4199
rect 12541 4165 12575 4199
rect 13553 4165 13587 4199
rect 16681 4165 16715 4199
rect 17049 4165 17083 4199
rect 22569 4165 22603 4199
rect 26801 4165 26835 4199
rect 30665 4165 30699 4199
rect 33563 4165 33597 4199
rect 2145 4097 2179 4131
rect 2881 4097 2915 4131
rect 3065 4097 3099 4131
rect 3341 4097 3375 4131
rect 5273 4097 5307 4131
rect 7573 4097 7607 4131
rect 10609 4097 10643 4131
rect 14381 4097 14415 4131
rect 15577 4097 15611 4131
rect 16313 4097 16347 4131
rect 16773 4097 16807 4131
rect 20177 4097 20211 4131
rect 22201 4097 22235 4131
rect 23765 4097 23799 4131
rect 24041 4097 24075 4131
rect 28089 4097 28123 4131
rect 29377 4097 29411 4131
rect 1685 4029 1719 4063
rect 1961 4029 1995 4063
rect 4997 4029 5031 4063
rect 5181 4029 5215 4063
rect 8493 4029 8527 4063
rect 9045 4029 9079 4063
rect 10517 4029 10551 4063
rect 10793 4029 10827 4063
rect 12081 4029 12115 4063
rect 12449 4029 12483 4063
rect 12725 4029 12759 4063
rect 14841 4029 14875 4063
rect 14933 4029 14967 4063
rect 15117 4029 15151 4063
rect 16037 4029 16071 4063
rect 16405 4029 16439 4063
rect 16552 4029 16586 4063
rect 18061 4029 18095 4063
rect 18521 4029 18555 4063
rect 18889 4029 18923 4063
rect 19257 4029 19291 4063
rect 19533 4029 19567 4063
rect 21005 4029 21039 4063
rect 25145 4029 25179 4063
rect 25605 4029 25639 4063
rect 30021 4029 30055 4063
rect 30849 4029 30883 4063
rect 31309 4029 31343 4063
rect 33492 4029 33526 4063
rect 33885 4029 33919 4063
rect 3157 3961 3191 3995
rect 6929 3961 6963 3995
rect 7021 3961 7055 3995
rect 9689 3961 9723 3995
rect 11253 3961 11287 3995
rect 11805 3961 11839 3995
rect 17785 3961 17819 3995
rect 20913 3961 20947 3995
rect 21367 3961 21401 3995
rect 23397 3961 23431 3995
rect 23857 3961 23891 3995
rect 25513 3961 25547 3995
rect 25967 3961 26001 3995
rect 27445 3961 27479 3995
rect 27537 3961 27571 3995
rect 29469 3961 29503 3995
rect 32413 3961 32447 3995
rect 4169 3893 4203 3927
rect 5733 3893 5767 3927
rect 6561 3893 6595 3927
rect 8769 3893 8803 3927
rect 10057 3893 10091 3927
rect 10333 3893 10367 3927
rect 12081 3893 12115 3927
rect 12173 3893 12207 3927
rect 12909 3893 12943 3927
rect 14749 3893 14783 3927
rect 15945 3893 15979 3927
rect 16037 3893 16071 3927
rect 17417 3893 17451 3927
rect 19809 3893 19843 3927
rect 24777 3893 24811 3927
rect 27261 3893 27295 3927
rect 30941 3893 30975 3927
rect 34253 3893 34287 3927
rect 35173 3893 35207 3927
rect 1685 3689 1719 3723
rect 2053 3689 2087 3723
rect 2237 3689 2271 3723
rect 3157 3689 3191 3723
rect 4353 3689 4387 3723
rect 4813 3689 4847 3723
rect 5917 3689 5951 3723
rect 7205 3689 7239 3723
rect 8677 3689 8711 3723
rect 9965 3689 9999 3723
rect 11805 3689 11839 3723
rect 14105 3689 14139 3723
rect 20361 3689 20395 3723
rect 21097 3689 21131 3723
rect 23489 3689 23523 3723
rect 24961 3689 24995 3723
rect 25559 3689 25593 3723
rect 26341 3689 26375 3723
rect 27905 3689 27939 3723
rect 29377 3689 29411 3723
rect 33287 3689 33321 3723
rect 10609 3621 10643 3655
rect 15301 3621 15335 3655
rect 16405 3621 16439 3655
rect 22154 3621 22188 3655
rect 23121 3621 23155 3655
rect 23949 3621 23983 3655
rect 24041 3621 24075 3655
rect 27261 3621 27295 3655
rect 29745 3621 29779 3655
rect 30941 3621 30975 3655
rect 2421 3553 2455 3587
rect 2697 3553 2731 3587
rect 4972 3553 5006 3587
rect 7205 3553 7239 3587
rect 7389 3553 7423 3587
rect 8493 3553 8527 3587
rect 9505 3553 9539 3587
rect 9781 3553 9815 3587
rect 10885 3553 10919 3587
rect 11529 3553 11563 3587
rect 12357 3553 12391 3587
rect 12633 3553 12667 3587
rect 13921 3553 13955 3587
rect 14381 3553 14415 3587
rect 16865 3553 16899 3587
rect 17969 3553 18003 3587
rect 18153 3553 18187 3587
rect 18521 3553 18555 3587
rect 18889 3553 18923 3587
rect 25421 3553 25455 3587
rect 26801 3553 26835 3587
rect 27077 3553 27111 3587
rect 28140 3553 28174 3587
rect 30297 3553 30331 3587
rect 32204 3553 32238 3587
rect 33216 3553 33250 3587
rect 6837 3485 6871 3519
rect 12817 3485 12851 3519
rect 15669 3485 15703 3519
rect 17233 3485 17267 3519
rect 19165 3485 19199 3519
rect 21649 3485 21683 3519
rect 21833 3485 21867 3519
rect 24593 3485 24627 3519
rect 28227 3485 28261 3519
rect 29653 3485 29687 3519
rect 6469 3417 6503 3451
rect 12449 3417 12483 3451
rect 13829 3417 13863 3451
rect 15577 3417 15611 3451
rect 19809 3417 19843 3451
rect 22753 3417 22787 3451
rect 32275 3417 32309 3451
rect 5043 3349 5077 3383
rect 12265 3349 12299 3383
rect 13369 3349 13403 3383
rect 15025 3349 15059 3383
rect 15439 3349 15473 3383
rect 15761 3349 15795 3383
rect 17509 3349 17543 3383
rect 19533 3349 19567 3383
rect 25973 3349 26007 3383
rect 2513 3145 2547 3179
rect 2881 3145 2915 3179
rect 4077 3145 4111 3179
rect 4721 3145 4755 3179
rect 8125 3145 8159 3179
rect 8309 3145 8343 3179
rect 2191 3077 2225 3111
rect 3065 3009 3099 3043
rect 5917 3009 5951 3043
rect 7481 3009 7515 3043
rect 1961 2941 1995 2975
rect 2120 2941 2154 2975
rect 4220 2941 4254 2975
rect 5089 2941 5123 2975
rect 5825 2941 5859 2975
rect 6285 2941 6319 2975
rect 6653 2941 6687 2975
rect 7205 2941 7239 2975
rect 7389 2941 7423 2975
rect 4307 2873 4341 2907
rect 9413 3145 9447 3179
rect 10793 3145 10827 3179
rect 11345 3145 11379 3179
rect 13921 3145 13955 3179
rect 14013 3145 14047 3179
rect 19809 3145 19843 3179
rect 21925 3145 21959 3179
rect 23121 3145 23155 3179
rect 28733 3145 28767 3179
rect 30389 3145 30423 3179
rect 31999 3145 32033 3179
rect 32689 3145 32723 3179
rect 33241 3145 33275 3179
rect 9229 3009 9263 3043
rect 8585 2941 8619 2975
rect 9689 3009 9723 3043
rect 10057 3009 10091 3043
rect 11805 3009 11839 3043
rect 12173 3009 12207 3043
rect 13185 3009 13219 3043
rect 9321 2941 9355 2975
rect 9597 2941 9631 2975
rect 9873 2941 9907 2975
rect 11161 2941 11195 2975
rect 12449 2941 12483 2975
rect 12541 2941 12575 2975
rect 12725 2941 12759 2975
rect 13461 2873 13495 2907
rect 8309 2805 8343 2839
rect 8493 2805 8527 2839
rect 8769 2805 8803 2839
rect 9045 2805 9079 2839
rect 9229 2805 9263 2839
rect 14841 3077 14875 3111
rect 15761 3077 15795 3111
rect 16865 3077 16899 3111
rect 18245 3077 18279 3111
rect 20085 3077 20119 3111
rect 20177 3077 20211 3111
rect 20453 3077 20487 3111
rect 24777 3077 24811 3111
rect 32413 3077 32447 3111
rect 17693 3009 17727 3043
rect 18613 3009 18647 3043
rect 19533 3009 19567 3043
rect 14289 2941 14323 2975
rect 14473 2941 14507 2975
rect 16497 2941 16531 2975
rect 18797 2941 18831 2975
rect 18889 2941 18923 2975
rect 19073 2941 19107 2975
rect 20821 3009 20855 3043
rect 22753 3009 22787 3043
rect 23489 3009 23523 3043
rect 24225 3009 24259 3043
rect 26801 3009 26835 3043
rect 26893 3009 26927 3043
rect 27169 3009 27203 3043
rect 27997 3009 28031 3043
rect 29101 3009 29135 3043
rect 30021 3009 30055 3043
rect 20361 2941 20395 2975
rect 20637 2941 20671 2975
rect 22661 2941 22695 2975
rect 25973 2941 26007 2975
rect 26157 2941 26191 2975
rect 16221 2873 16255 2907
rect 20085 2873 20119 2907
rect 24317 2873 24351 2907
rect 27261 2941 27295 2975
rect 27813 2941 27847 2975
rect 29285 2941 29319 2975
rect 29837 2941 29871 2975
rect 31928 2941 31962 2975
rect 30849 2873 30883 2907
rect 14013 2805 14047 2839
rect 15393 2805 15427 2839
rect 21373 2805 21407 2839
rect 24041 2805 24075 2839
rect 25421 2805 25455 2839
rect 25789 2805 25823 2839
rect 26893 2805 26927 2839
rect 28365 2805 28399 2839
rect 2145 2601 2179 2635
rect 3111 2601 3145 2635
rect 4399 2601 4433 2635
rect 7021 2601 7055 2635
rect 9597 2601 9631 2635
rect 12817 2601 12851 2635
rect 14473 2601 14507 2635
rect 14933 2601 14967 2635
rect 20085 2601 20119 2635
rect 20545 2601 20579 2635
rect 22201 2601 22235 2635
rect 22891 2601 22925 2635
rect 25421 2601 25455 2635
rect 26617 2601 26651 2635
rect 27353 2601 27387 2635
rect 28917 2601 28951 2635
rect 29285 2601 29319 2635
rect 29929 2601 29963 2635
rect 3525 2533 3559 2567
rect 1961 2465 1995 2499
rect 3040 2465 3074 2499
rect 4296 2465 4330 2499
rect 4721 2465 4755 2499
rect 5917 2465 5951 2499
rect 6009 2465 6043 2499
rect 5181 2397 5215 2431
rect 7849 2533 7883 2567
rect 11713 2533 11747 2567
rect 13369 2533 13403 2567
rect 13829 2533 13863 2567
rect 17233 2533 17267 2567
rect 17785 2533 17819 2567
rect 20913 2533 20947 2567
rect 24041 2533 24075 2567
rect 28641 2533 28675 2567
rect 7113 2465 7147 2499
rect 7205 2465 7239 2499
rect 7389 2465 7423 2499
rect 8217 2465 8251 2499
rect 8677 2465 8711 2499
rect 9965 2465 9999 2499
rect 10425 2465 10459 2499
rect 10701 2465 10735 2499
rect 11069 2465 11103 2499
rect 12357 2465 12391 2499
rect 12633 2465 12667 2499
rect 16037 2465 16071 2499
rect 16405 2465 16439 2499
rect 16773 2465 16807 2499
rect 16865 2465 16899 2499
rect 18153 2465 18187 2499
rect 18337 2465 18371 2499
rect 18429 2465 18463 2499
rect 18613 2465 18647 2499
rect 19717 2465 19751 2499
rect 19901 2465 19935 2499
rect 21097 2465 21131 2499
rect 21281 2465 21315 2499
rect 21465 2465 21499 2499
rect 22788 2465 22822 2499
rect 23213 2465 23247 2499
rect 23857 2465 23891 2499
rect 24685 2465 24719 2499
rect 25053 2465 25087 2499
rect 25605 2465 25639 2499
rect 26157 2465 26191 2499
rect 26709 2465 26743 2499
rect 26928 2465 26962 2499
rect 27905 2465 27939 2499
rect 28457 2465 28491 2499
rect 29745 2465 29779 2499
rect 30824 2465 30858 2499
rect 7021 2329 7055 2363
rect 8861 2329 8895 2363
rect 11989 2397 12023 2431
rect 14197 2397 14231 2431
rect 18797 2397 18831 2431
rect 21925 2397 21959 2431
rect 25789 2329 25823 2363
rect 30205 2397 30239 2431
rect 27813 2329 27847 2363
rect 30895 2329 30929 2363
rect 2513 2261 2547 2295
rect 6285 2261 6319 2295
rect 6653 2261 6687 2295
rect 9229 2261 9263 2295
rect 10149 2261 10183 2295
rect 10701 2261 10735 2295
rect 10793 2261 10827 2295
rect 13645 2261 13679 2295
rect 13967 2261 14001 2295
rect 14105 2261 14139 2295
rect 15209 2261 15243 2295
rect 19349 2261 19383 2295
rect 22569 2261 22603 2295
rect 26709 2261 26743 2295
rect 27031 2261 27065 2295
rect 31217 2261 31251 2295
<< metal1 >>
rect 1104 13626 38824 13648
rect 1104 13574 14315 13626
rect 14367 13574 14379 13626
rect 14431 13574 14443 13626
rect 14495 13574 14507 13626
rect 14559 13574 27648 13626
rect 27700 13574 27712 13626
rect 27764 13574 27776 13626
rect 27828 13574 27840 13626
rect 27892 13574 38824 13626
rect 1104 13552 38824 13574
rect 106 13132 112 13184
rect 164 13172 170 13184
rect 28258 13172 28264 13184
rect 164 13144 28264 13172
rect 164 13132 170 13144
rect 28258 13132 28264 13144
rect 28316 13132 28322 13184
rect 1104 13082 38824 13104
rect 1104 13030 7648 13082
rect 7700 13030 7712 13082
rect 7764 13030 7776 13082
rect 7828 13030 7840 13082
rect 7892 13030 20982 13082
rect 21034 13030 21046 13082
rect 21098 13030 21110 13082
rect 21162 13030 21174 13082
rect 21226 13030 34315 13082
rect 34367 13030 34379 13082
rect 34431 13030 34443 13082
rect 34495 13030 34507 13082
rect 34559 13030 38824 13082
rect 1104 13008 38824 13030
rect 18509 12971 18567 12977
rect 18509 12937 18521 12971
rect 18555 12968 18567 12971
rect 19610 12968 19616 12980
rect 18555 12940 19616 12968
rect 18555 12937 18567 12940
rect 18509 12931 18567 12937
rect 19610 12928 19616 12940
rect 19668 12928 19674 12980
rect 28258 12968 28264 12980
rect 28219 12940 28264 12968
rect 28258 12928 28264 12940
rect 28316 12928 28322 12980
rect 31941 12971 31999 12977
rect 31941 12937 31953 12971
rect 31987 12968 31999 12971
rect 34054 12968 34060 12980
rect 31987 12940 34060 12968
rect 31987 12937 31999 12940
rect 31941 12931 31999 12937
rect 34054 12928 34060 12940
rect 34112 12928 34118 12980
rect 35618 12968 35624 12980
rect 35579 12940 35624 12968
rect 35618 12928 35624 12940
rect 35676 12928 35682 12980
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12764 1455 12767
rect 7285 12767 7343 12773
rect 1443 12736 1808 12764
rect 1443 12733 1455 12736
rect 1397 12727 1455 12733
rect 1780 12640 1808 12736
rect 7285 12733 7297 12767
rect 7331 12764 7343 12767
rect 7331 12736 7880 12764
rect 7331 12733 7343 12736
rect 7285 12727 7343 12733
rect 7852 12705 7880 12736
rect 8202 12724 8208 12776
rect 8260 12764 8266 12776
rect 8386 12773 8392 12776
rect 8332 12767 8392 12773
rect 8332 12764 8344 12767
rect 8260 12736 8344 12764
rect 8260 12724 8266 12736
rect 8332 12733 8344 12736
rect 8378 12733 8392 12767
rect 8332 12727 8392 12733
rect 8386 12724 8392 12727
rect 8444 12764 8450 12776
rect 8757 12767 8815 12773
rect 8757 12764 8769 12767
rect 8444 12736 8769 12764
rect 8444 12724 8450 12736
rect 8757 12733 8769 12736
rect 8803 12733 8815 12767
rect 8757 12727 8815 12733
rect 18325 12767 18383 12773
rect 18325 12733 18337 12767
rect 18371 12764 18383 12767
rect 18693 12767 18751 12773
rect 18693 12764 18705 12767
rect 18371 12736 18705 12764
rect 18371 12733 18383 12736
rect 18325 12727 18383 12733
rect 18693 12733 18705 12736
rect 18739 12733 18751 12767
rect 18693 12727 18751 12733
rect 28077 12767 28135 12773
rect 28077 12733 28089 12767
rect 28123 12764 28135 12767
rect 28718 12764 28724 12776
rect 28123 12736 28724 12764
rect 28123 12733 28135 12736
rect 28077 12727 28135 12733
rect 28718 12724 28724 12736
rect 28776 12724 28782 12776
rect 31386 12724 31392 12776
rect 31444 12764 31450 12776
rect 31757 12767 31815 12773
rect 31757 12764 31769 12767
rect 31444 12736 31769 12764
rect 31444 12724 31450 12736
rect 31757 12733 31769 12736
rect 31803 12764 31815 12767
rect 32309 12767 32367 12773
rect 32309 12764 32321 12767
rect 31803 12736 32321 12764
rect 31803 12733 31815 12736
rect 31757 12727 31815 12733
rect 32309 12733 32321 12736
rect 32355 12733 32367 12767
rect 32309 12727 32367 12733
rect 34790 12724 34796 12776
rect 34848 12764 34854 12776
rect 35437 12767 35495 12773
rect 35437 12764 35449 12767
rect 34848 12736 35449 12764
rect 34848 12724 34854 12736
rect 35437 12733 35449 12736
rect 35483 12764 35495 12767
rect 35989 12767 36047 12773
rect 35989 12764 36001 12767
rect 35483 12736 36001 12764
rect 35483 12733 35495 12736
rect 35437 12727 35495 12733
rect 35989 12733 36001 12736
rect 36035 12733 36047 12767
rect 35989 12727 36047 12733
rect 7837 12699 7895 12705
rect 7837 12665 7849 12699
rect 7883 12696 7895 12699
rect 12894 12696 12900 12708
rect 7883 12668 12900 12696
rect 7883 12665 7895 12668
rect 7837 12659 7895 12665
rect 12894 12656 12900 12668
rect 12952 12656 12958 12708
rect 16850 12656 16856 12708
rect 16908 12696 16914 12708
rect 39574 12696 39580 12708
rect 16908 12668 39580 12696
rect 16908 12656 16914 12668
rect 39574 12656 39580 12668
rect 39632 12656 39638 12708
rect 106 12588 112 12640
rect 164 12628 170 12640
rect 1581 12631 1639 12637
rect 1581 12628 1593 12631
rect 164 12600 1593 12628
rect 164 12588 170 12600
rect 1581 12597 1593 12600
rect 1627 12597 1639 12631
rect 1581 12591 1639 12597
rect 1762 12588 1768 12640
rect 1820 12628 1826 12640
rect 1949 12631 2007 12637
rect 1949 12628 1961 12631
rect 1820 12600 1961 12628
rect 1820 12588 1826 12600
rect 1949 12597 1961 12600
rect 1995 12597 2007 12631
rect 7466 12628 7472 12640
rect 7427 12600 7472 12628
rect 1949 12591 2007 12597
rect 7466 12588 7472 12600
rect 7524 12588 7530 12640
rect 8018 12588 8024 12640
rect 8076 12628 8082 12640
rect 8435 12631 8493 12637
rect 8435 12628 8447 12631
rect 8076 12600 8447 12628
rect 8076 12588 8082 12600
rect 8435 12597 8447 12600
rect 8481 12597 8493 12631
rect 8435 12591 8493 12597
rect 18693 12631 18751 12637
rect 18693 12597 18705 12631
rect 18739 12628 18751 12631
rect 18969 12631 19027 12637
rect 18969 12628 18981 12631
rect 18739 12600 18981 12628
rect 18739 12597 18751 12600
rect 18693 12591 18751 12597
rect 18969 12597 18981 12600
rect 19015 12628 19027 12631
rect 19242 12628 19248 12640
rect 19015 12600 19248 12628
rect 19015 12597 19027 12600
rect 18969 12591 19027 12597
rect 19242 12588 19248 12600
rect 19300 12588 19306 12640
rect 28718 12628 28724 12640
rect 28679 12600 28724 12628
rect 28718 12588 28724 12600
rect 28776 12588 28782 12640
rect 1104 12538 38824 12560
rect 1104 12486 14315 12538
rect 14367 12486 14379 12538
rect 14431 12486 14443 12538
rect 14495 12486 14507 12538
rect 14559 12486 27648 12538
rect 27700 12486 27712 12538
rect 27764 12486 27776 12538
rect 27828 12486 27840 12538
rect 27892 12486 38824 12538
rect 1104 12464 38824 12486
rect 1397 12291 1455 12297
rect 1397 12257 1409 12291
rect 1443 12288 1455 12291
rect 2038 12288 2044 12300
rect 1443 12260 2044 12288
rect 1443 12257 1455 12260
rect 1397 12251 1455 12257
rect 2038 12248 2044 12260
rect 2096 12248 2102 12300
rect 6546 12248 6552 12300
rect 6604 12288 6610 12300
rect 6676 12291 6734 12297
rect 6676 12288 6688 12291
rect 6604 12260 6688 12288
rect 6604 12248 6610 12260
rect 6676 12257 6688 12260
rect 6722 12257 6734 12291
rect 6676 12251 6734 12257
rect 7720 12291 7778 12297
rect 7720 12257 7732 12291
rect 7766 12288 7778 12291
rect 8110 12288 8116 12300
rect 7766 12260 8116 12288
rect 7766 12257 7778 12260
rect 7720 12251 7778 12257
rect 8110 12248 8116 12260
rect 8168 12248 8174 12300
rect 9582 12288 9588 12300
rect 9543 12260 9588 12288
rect 9582 12248 9588 12260
rect 9640 12248 9646 12300
rect 10689 12291 10747 12297
rect 10689 12257 10701 12291
rect 10735 12288 10747 12291
rect 10778 12288 10784 12300
rect 10735 12260 10784 12288
rect 10735 12257 10747 12260
rect 10689 12251 10747 12257
rect 10778 12248 10784 12260
rect 10836 12248 10842 12300
rect 15654 12288 15660 12300
rect 15615 12260 15660 12288
rect 15654 12248 15660 12260
rect 15712 12248 15718 12300
rect 16828 12291 16886 12297
rect 16828 12257 16840 12291
rect 16874 12288 16886 12291
rect 17034 12288 17040 12300
rect 16874 12260 17040 12288
rect 16874 12257 16886 12260
rect 16828 12251 16886 12257
rect 17034 12248 17040 12260
rect 17092 12248 17098 12300
rect 18852 12291 18910 12297
rect 18852 12257 18864 12291
rect 18898 12288 18910 12291
rect 19242 12288 19248 12300
rect 18898 12260 19248 12288
rect 18898 12257 18910 12260
rect 18852 12251 18910 12257
rect 19242 12248 19248 12260
rect 19300 12248 19306 12300
rect 19702 12248 19708 12300
rect 19760 12288 19766 12300
rect 19797 12291 19855 12297
rect 19797 12288 19809 12291
rect 19760 12260 19809 12288
rect 19760 12248 19766 12260
rect 19797 12257 19809 12260
rect 19843 12257 19855 12291
rect 19797 12251 19855 12257
rect 23474 12248 23480 12300
rect 23532 12288 23538 12300
rect 24489 12291 24547 12297
rect 23532 12260 23577 12288
rect 23532 12248 23538 12260
rect 24489 12257 24501 12291
rect 24535 12288 24547 12291
rect 25130 12288 25136 12300
rect 24535 12260 25136 12288
rect 24535 12257 24547 12260
rect 24489 12251 24547 12257
rect 25130 12248 25136 12260
rect 25188 12248 25194 12300
rect 27341 12291 27399 12297
rect 27341 12257 27353 12291
rect 27387 12288 27399 12291
rect 28074 12288 28080 12300
rect 27387 12260 28080 12288
rect 27387 12257 27399 12260
rect 27341 12251 27399 12257
rect 28074 12248 28080 12260
rect 28132 12248 28138 12300
rect 2682 12220 2688 12232
rect 2643 12192 2688 12220
rect 2682 12180 2688 12192
rect 2740 12180 2746 12232
rect 17773 12223 17831 12229
rect 17773 12189 17785 12223
rect 17819 12220 17831 12223
rect 18138 12220 18144 12232
rect 17819 12192 18144 12220
rect 17819 12189 17831 12192
rect 17773 12183 17831 12189
rect 18138 12180 18144 12192
rect 18196 12180 18202 12232
rect 1578 12152 1584 12164
rect 1539 12124 1584 12152
rect 1578 12112 1584 12124
rect 1636 12112 1642 12164
rect 15887 12155 15945 12161
rect 15887 12121 15899 12155
rect 15933 12152 15945 12155
rect 18598 12152 18604 12164
rect 15933 12124 18604 12152
rect 15933 12121 15945 12124
rect 15887 12115 15945 12121
rect 18598 12112 18604 12124
rect 18656 12112 18662 12164
rect 6779 12087 6837 12093
rect 6779 12053 6791 12087
rect 6825 12084 6837 12087
rect 6914 12084 6920 12096
rect 6825 12056 6920 12084
rect 6825 12053 6837 12056
rect 6779 12047 6837 12053
rect 6914 12044 6920 12056
rect 6972 12044 6978 12096
rect 7791 12087 7849 12093
rect 7791 12053 7803 12087
rect 7837 12084 7849 12087
rect 8846 12084 8852 12096
rect 7837 12056 8852 12084
rect 7837 12053 7849 12056
rect 7791 12047 7849 12053
rect 8846 12044 8852 12056
rect 8904 12044 8910 12096
rect 9030 12044 9036 12096
rect 9088 12084 9094 12096
rect 9815 12087 9873 12093
rect 9815 12084 9827 12087
rect 9088 12056 9827 12084
rect 9088 12044 9094 12056
rect 9815 12053 9827 12056
rect 9861 12053 9873 12087
rect 9815 12047 9873 12053
rect 10502 12044 10508 12096
rect 10560 12084 10566 12096
rect 10827 12087 10885 12093
rect 10827 12084 10839 12087
rect 10560 12056 10839 12084
rect 10560 12044 10566 12056
rect 10827 12053 10839 12056
rect 10873 12053 10885 12087
rect 10827 12047 10885 12053
rect 16758 12044 16764 12096
rect 16816 12084 16822 12096
rect 16899 12087 16957 12093
rect 16899 12084 16911 12087
rect 16816 12056 16911 12084
rect 16816 12044 16822 12056
rect 16899 12053 16911 12056
rect 16945 12053 16957 12087
rect 16899 12047 16957 12053
rect 18414 12044 18420 12096
rect 18472 12084 18478 12096
rect 18923 12087 18981 12093
rect 18923 12084 18935 12087
rect 18472 12056 18935 12084
rect 18472 12044 18478 12056
rect 18923 12053 18935 12056
rect 18969 12053 18981 12087
rect 18923 12047 18981 12053
rect 19794 12044 19800 12096
rect 19852 12084 19858 12096
rect 19981 12087 20039 12093
rect 19981 12084 19993 12087
rect 19852 12056 19993 12084
rect 19852 12044 19858 12056
rect 19981 12053 19993 12056
rect 20027 12053 20039 12087
rect 19981 12047 20039 12053
rect 23615 12087 23673 12093
rect 23615 12053 23627 12087
rect 23661 12084 23673 12087
rect 24118 12084 24124 12096
rect 23661 12056 24124 12084
rect 23661 12053 23673 12056
rect 23615 12047 23673 12053
rect 24118 12044 24124 12056
rect 24176 12044 24182 12096
rect 24670 12084 24676 12096
rect 24631 12056 24676 12084
rect 24670 12044 24676 12056
rect 24728 12044 24734 12096
rect 27522 12084 27528 12096
rect 27483 12056 27528 12084
rect 27522 12044 27528 12056
rect 27580 12044 27586 12096
rect 1104 11994 38824 12016
rect 1104 11942 7648 11994
rect 7700 11942 7712 11994
rect 7764 11942 7776 11994
rect 7828 11942 7840 11994
rect 7892 11942 20982 11994
rect 21034 11942 21046 11994
rect 21098 11942 21110 11994
rect 21162 11942 21174 11994
rect 21226 11942 34315 11994
rect 34367 11942 34379 11994
rect 34431 11942 34443 11994
rect 34495 11942 34507 11994
rect 34559 11942 38824 11994
rect 1104 11920 38824 11942
rect 1118 11840 1124 11892
rect 1176 11880 1182 11892
rect 1581 11883 1639 11889
rect 1581 11880 1593 11883
rect 1176 11852 1593 11880
rect 1176 11840 1182 11852
rect 1581 11849 1593 11852
rect 1627 11849 1639 11883
rect 1581 11843 1639 11849
rect 1946 11840 1952 11892
rect 2004 11880 2010 11892
rect 2685 11883 2743 11889
rect 2685 11880 2697 11883
rect 2004 11852 2697 11880
rect 2004 11840 2010 11852
rect 2685 11849 2697 11852
rect 2731 11849 2743 11883
rect 2685 11843 2743 11849
rect 4798 11840 4804 11892
rect 4856 11880 4862 11892
rect 8665 11883 8723 11889
rect 8665 11880 8677 11883
rect 4856 11852 8677 11880
rect 4856 11840 4862 11852
rect 8665 11849 8677 11852
rect 8711 11880 8723 11883
rect 8849 11883 8907 11889
rect 8849 11880 8861 11883
rect 8711 11852 8861 11880
rect 8711 11849 8723 11852
rect 8665 11843 8723 11849
rect 8849 11849 8861 11852
rect 8895 11849 8907 11883
rect 17034 11880 17040 11892
rect 16995 11852 17040 11880
rect 8849 11843 8907 11849
rect 17034 11840 17040 11852
rect 17092 11880 17098 11892
rect 23014 11880 23020 11892
rect 17092 11852 23020 11880
rect 17092 11840 17098 11852
rect 1670 11812 1676 11824
rect 1412 11784 1676 11812
rect 1412 11685 1440 11784
rect 1670 11772 1676 11784
rect 1728 11812 1734 11824
rect 6546 11812 6552 11824
rect 1728 11784 6552 11812
rect 1728 11772 1734 11784
rect 6546 11772 6552 11784
rect 6604 11772 6610 11824
rect 19702 11772 19708 11824
rect 19760 11812 19766 11824
rect 20533 11815 20591 11821
rect 20533 11812 20545 11815
rect 19760 11784 20545 11812
rect 19760 11772 19766 11784
rect 20533 11781 20545 11784
rect 20579 11781 20591 11815
rect 20533 11775 20591 11781
rect 2038 11744 2044 11756
rect 1999 11716 2044 11744
rect 2038 11704 2044 11716
rect 2096 11704 2102 11756
rect 4522 11704 4528 11756
rect 4580 11744 4586 11756
rect 9582 11744 9588 11756
rect 4580 11716 9588 11744
rect 4580 11704 4586 11716
rect 9582 11704 9588 11716
rect 9640 11744 9646 11756
rect 9858 11744 9864 11756
rect 9640 11716 9864 11744
rect 9640 11704 9646 11716
rect 9858 11704 9864 11716
rect 9916 11704 9922 11756
rect 14093 11747 14151 11753
rect 14093 11713 14105 11747
rect 14139 11744 14151 11747
rect 15654 11744 15660 11756
rect 14139 11716 15660 11744
rect 14139 11713 14151 11716
rect 14093 11707 14151 11713
rect 15654 11704 15660 11716
rect 15712 11744 15718 11756
rect 15841 11747 15899 11753
rect 15841 11744 15853 11747
rect 15712 11716 15853 11744
rect 15712 11704 15718 11716
rect 15841 11713 15853 11716
rect 15887 11744 15899 11747
rect 20346 11744 20352 11756
rect 15887 11716 20352 11744
rect 15887 11713 15899 11716
rect 15841 11707 15899 11713
rect 20346 11704 20352 11716
rect 20404 11704 20410 11756
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11645 1455 11679
rect 1397 11639 1455 11645
rect 2501 11679 2559 11685
rect 2501 11645 2513 11679
rect 2547 11676 2559 11679
rect 7006 11676 7012 11688
rect 2547 11648 3004 11676
rect 6967 11648 7012 11676
rect 2547 11645 2559 11648
rect 2501 11639 2559 11645
rect 2976 11552 3004 11648
rect 7006 11636 7012 11648
rect 7064 11636 7070 11688
rect 7377 11679 7435 11685
rect 7377 11645 7389 11679
rect 7423 11676 7435 11679
rect 7466 11676 7472 11688
rect 7423 11648 7472 11676
rect 7423 11645 7435 11648
rect 7377 11639 7435 11645
rect 6270 11608 6276 11620
rect 6183 11580 6276 11608
rect 6270 11568 6276 11580
rect 6328 11608 6334 11620
rect 7392 11608 7420 11639
rect 7466 11636 7472 11648
rect 7524 11636 7530 11688
rect 8456 11679 8514 11685
rect 8456 11645 8468 11679
rect 8502 11676 8514 11679
rect 8665 11679 8723 11685
rect 8665 11676 8677 11679
rect 8502 11648 8677 11676
rect 8502 11645 8514 11648
rect 8456 11639 8514 11645
rect 8665 11645 8677 11648
rect 8711 11676 8723 11679
rect 9122 11676 9128 11688
rect 8711 11648 9128 11676
rect 8711 11645 8723 11648
rect 8665 11639 8723 11645
rect 9122 11636 9128 11648
rect 9180 11636 9186 11688
rect 9306 11636 9312 11688
rect 9364 11676 9370 11688
rect 9436 11679 9494 11685
rect 9436 11676 9448 11679
rect 9364 11648 9448 11676
rect 9364 11636 9370 11648
rect 9436 11645 9448 11648
rect 9482 11676 9494 11679
rect 10229 11679 10287 11685
rect 10229 11676 10241 11679
rect 9482 11648 10241 11676
rect 9482 11645 9494 11648
rect 9436 11639 9494 11645
rect 10229 11645 10241 11648
rect 10275 11645 10287 11679
rect 10229 11639 10287 11645
rect 10480 11679 10538 11685
rect 10480 11645 10492 11679
rect 10526 11676 10538 11679
rect 11057 11679 11115 11685
rect 11057 11676 11069 11679
rect 10526 11648 11069 11676
rect 10526 11645 10538 11648
rect 10480 11639 10538 11645
rect 11057 11645 11069 11648
rect 11103 11645 11115 11679
rect 11057 11639 11115 11645
rect 6328 11580 7420 11608
rect 10244 11608 10272 11639
rect 11790 11636 11796 11688
rect 11848 11676 11854 11688
rect 13884 11679 13942 11685
rect 13884 11676 13896 11679
rect 11848 11648 13896 11676
rect 11848 11636 11854 11648
rect 13884 11645 13896 11648
rect 13930 11676 13942 11679
rect 18230 11676 18236 11688
rect 13930 11648 14412 11676
rect 18191 11648 18236 11676
rect 13930 11645 13942 11648
rect 13884 11639 13942 11645
rect 14384 11617 14412 11648
rect 18230 11636 18236 11648
rect 18288 11636 18294 11688
rect 18690 11676 18696 11688
rect 18651 11648 18696 11676
rect 18690 11636 18696 11648
rect 18748 11636 18754 11688
rect 19740 11679 19798 11685
rect 19740 11676 19752 11679
rect 19076 11648 19752 11676
rect 14093 11611 14151 11617
rect 14093 11608 14105 11611
rect 10244 11580 14105 11608
rect 6328 11568 6334 11580
rect 14093 11577 14105 11580
rect 14139 11577 14151 11611
rect 14093 11571 14151 11577
rect 14369 11611 14427 11617
rect 14369 11577 14381 11611
rect 14415 11608 14427 11611
rect 17218 11608 17224 11620
rect 14415 11580 17224 11608
rect 14415 11577 14427 11580
rect 14369 11571 14427 11577
rect 17218 11568 17224 11580
rect 17276 11568 17282 11620
rect 17865 11611 17923 11617
rect 17865 11577 17877 11611
rect 17911 11608 17923 11611
rect 18708 11608 18736 11636
rect 17911 11580 18736 11608
rect 17911 11577 17923 11580
rect 17865 11571 17923 11577
rect 19076 11552 19104 11648
rect 19740 11645 19752 11648
rect 19786 11676 19798 11679
rect 20165 11679 20223 11685
rect 20165 11676 20177 11679
rect 19786 11648 20177 11676
rect 19786 11645 19798 11648
rect 19740 11639 19798 11645
rect 20165 11645 20177 11648
rect 20211 11676 20223 11679
rect 22370 11676 22376 11688
rect 20211 11648 22376 11676
rect 20211 11645 20223 11648
rect 20165 11639 20223 11645
rect 22370 11636 22376 11648
rect 22428 11636 22434 11688
rect 22639 11685 22667 11852
rect 23014 11840 23020 11852
rect 23072 11840 23078 11892
rect 35618 11880 35624 11892
rect 35579 11852 35624 11880
rect 35618 11840 35624 11852
rect 35676 11840 35682 11892
rect 24394 11772 24400 11824
rect 24452 11812 24458 11824
rect 25547 11815 25605 11821
rect 25547 11812 25559 11815
rect 24452 11784 25559 11812
rect 24452 11772 24458 11784
rect 25547 11781 25559 11784
rect 25593 11781 25605 11815
rect 25547 11775 25605 11781
rect 25317 11747 25375 11753
rect 25317 11744 25329 11747
rect 24412 11716 25329 11744
rect 24412 11685 24440 11716
rect 25317 11713 25329 11716
rect 25363 11744 25375 11747
rect 26326 11744 26332 11756
rect 25363 11716 26332 11744
rect 25363 11713 25375 11716
rect 25317 11707 25375 11713
rect 26326 11704 26332 11716
rect 26384 11704 26390 11756
rect 22624 11679 22682 11685
rect 22624 11645 22636 11679
rect 22670 11645 22682 11679
rect 22624 11639 22682 11645
rect 24397 11679 24455 11685
rect 24397 11645 24409 11679
rect 24443 11645 24455 11679
rect 24397 11639 24455 11645
rect 25476 11679 25534 11685
rect 25476 11645 25488 11679
rect 25522 11676 25534 11679
rect 35434 11676 35440 11688
rect 25522 11648 26004 11676
rect 35395 11648 35440 11676
rect 25522 11645 25534 11648
rect 25476 11639 25534 11645
rect 19843 11611 19901 11617
rect 19843 11577 19855 11611
rect 19889 11608 19901 11611
rect 21634 11608 21640 11620
rect 19889 11580 21640 11608
rect 19889 11577 19901 11580
rect 19843 11571 19901 11577
rect 21634 11568 21640 11580
rect 21692 11568 21698 11620
rect 25976 11617 26004 11648
rect 35434 11636 35440 11648
rect 35492 11676 35498 11688
rect 35989 11679 36047 11685
rect 35989 11676 36001 11679
rect 35492 11648 36001 11676
rect 35492 11636 35498 11648
rect 35989 11645 36001 11648
rect 36035 11645 36047 11679
rect 35989 11639 36047 11645
rect 25961 11611 26019 11617
rect 25961 11577 25973 11611
rect 26007 11608 26019 11611
rect 30926 11608 30932 11620
rect 26007 11580 30932 11608
rect 26007 11577 26019 11580
rect 25961 11571 26019 11577
rect 30926 11568 30932 11580
rect 30984 11568 30990 11620
rect 2958 11500 2964 11552
rect 3016 11540 3022 11552
rect 3053 11543 3111 11549
rect 3053 11540 3065 11543
rect 3016 11512 3065 11540
rect 3016 11500 3022 11512
rect 3053 11509 3065 11512
rect 3099 11509 3111 11543
rect 7098 11540 7104 11552
rect 7059 11512 7104 11540
rect 3053 11503 3111 11509
rect 7098 11500 7104 11512
rect 7156 11500 7162 11552
rect 7929 11543 7987 11549
rect 7929 11509 7941 11543
rect 7975 11540 7987 11543
rect 8110 11540 8116 11552
rect 7975 11512 8116 11540
rect 7975 11509 7987 11512
rect 7929 11503 7987 11509
rect 8110 11500 8116 11512
rect 8168 11500 8174 11552
rect 8527 11543 8585 11549
rect 8527 11509 8539 11543
rect 8573 11540 8585 11543
rect 8662 11540 8668 11552
rect 8573 11512 8668 11540
rect 8573 11509 8585 11512
rect 8527 11503 8585 11509
rect 8662 11500 8668 11512
rect 8720 11500 8726 11552
rect 8938 11500 8944 11552
rect 8996 11540 9002 11552
rect 9539 11543 9597 11549
rect 9539 11540 9551 11543
rect 8996 11512 9551 11540
rect 8996 11500 9002 11512
rect 9539 11509 9551 11512
rect 9585 11509 9597 11543
rect 9539 11503 9597 11509
rect 10318 11500 10324 11552
rect 10376 11540 10382 11552
rect 10551 11543 10609 11549
rect 10551 11540 10563 11543
rect 10376 11512 10563 11540
rect 10376 11500 10382 11512
rect 10551 11509 10563 11512
rect 10597 11509 10609 11543
rect 10551 11503 10609 11509
rect 10778 11500 10784 11552
rect 10836 11540 10842 11552
rect 10873 11543 10931 11549
rect 10873 11540 10885 11543
rect 10836 11512 10885 11540
rect 10836 11500 10842 11512
rect 10873 11509 10885 11512
rect 10919 11509 10931 11543
rect 10873 11503 10931 11509
rect 11057 11543 11115 11549
rect 11057 11509 11069 11543
rect 11103 11540 11115 11543
rect 11333 11543 11391 11549
rect 11333 11540 11345 11543
rect 11103 11512 11345 11540
rect 11103 11509 11115 11512
rect 11057 11503 11115 11509
rect 11333 11509 11345 11512
rect 11379 11540 11391 11543
rect 11790 11540 11796 11552
rect 11379 11512 11796 11540
rect 11379 11509 11391 11512
rect 11333 11503 11391 11509
rect 11790 11500 11796 11512
rect 11848 11500 11854 11552
rect 13955 11543 14013 11549
rect 13955 11509 13967 11543
rect 14001 11540 14013 11543
rect 14182 11540 14188 11552
rect 14001 11512 14188 11540
rect 14001 11509 14013 11512
rect 13955 11503 14013 11509
rect 14182 11500 14188 11512
rect 14240 11500 14246 11552
rect 14826 11540 14832 11552
rect 14787 11512 14832 11540
rect 14826 11500 14832 11512
rect 14884 11500 14890 11552
rect 16577 11543 16635 11549
rect 16577 11509 16589 11543
rect 16623 11540 16635 11543
rect 17402 11540 17408 11552
rect 16623 11512 17408 11540
rect 16623 11509 16635 11512
rect 16577 11503 16635 11509
rect 17402 11500 17408 11512
rect 17460 11500 17466 11552
rect 17954 11500 17960 11552
rect 18012 11540 18018 11552
rect 18233 11543 18291 11549
rect 18233 11540 18245 11543
rect 18012 11512 18245 11540
rect 18012 11500 18018 11512
rect 18233 11509 18245 11512
rect 18279 11509 18291 11543
rect 18233 11503 18291 11509
rect 19058 11500 19064 11552
rect 19116 11500 19122 11552
rect 19242 11540 19248 11552
rect 19155 11512 19248 11540
rect 19242 11500 19248 11512
rect 19300 11540 19306 11552
rect 19978 11540 19984 11552
rect 19300 11512 19984 11540
rect 19300 11500 19306 11512
rect 19978 11500 19984 11512
rect 20036 11500 20042 11552
rect 22695 11543 22753 11549
rect 22695 11509 22707 11543
rect 22741 11540 22753 11543
rect 22922 11540 22928 11552
rect 22741 11512 22928 11540
rect 22741 11509 22753 11512
rect 22695 11503 22753 11509
rect 22922 11500 22928 11512
rect 22980 11500 22986 11552
rect 23474 11500 23480 11552
rect 23532 11540 23538 11552
rect 23845 11543 23903 11549
rect 23845 11540 23857 11543
rect 23532 11512 23857 11540
rect 23532 11500 23538 11512
rect 23845 11509 23857 11512
rect 23891 11509 23903 11543
rect 23845 11503 23903 11509
rect 24302 11500 24308 11552
rect 24360 11540 24366 11552
rect 24581 11543 24639 11549
rect 24581 11540 24593 11543
rect 24360 11512 24593 11540
rect 24360 11500 24366 11512
rect 24581 11509 24593 11512
rect 24627 11509 24639 11543
rect 24581 11503 24639 11509
rect 24949 11543 25007 11549
rect 24949 11509 24961 11543
rect 24995 11540 25007 11543
rect 25130 11540 25136 11552
rect 24995 11512 25136 11540
rect 24995 11509 25007 11512
rect 24949 11503 25007 11509
rect 25130 11500 25136 11512
rect 25188 11500 25194 11552
rect 27338 11540 27344 11552
rect 27299 11512 27344 11540
rect 27338 11500 27344 11512
rect 27396 11500 27402 11552
rect 27893 11543 27951 11549
rect 27893 11509 27905 11543
rect 27939 11540 27951 11543
rect 28074 11540 28080 11552
rect 27939 11512 28080 11540
rect 27939 11509 27951 11512
rect 27893 11503 27951 11509
rect 28074 11500 28080 11512
rect 28132 11500 28138 11552
rect 1104 11450 38824 11472
rect 1104 11398 14315 11450
rect 14367 11398 14379 11450
rect 14431 11398 14443 11450
rect 14495 11398 14507 11450
rect 14559 11398 27648 11450
rect 27700 11398 27712 11450
rect 27764 11398 27776 11450
rect 27828 11398 27840 11450
rect 27892 11398 38824 11450
rect 1104 11376 38824 11398
rect 1670 11336 1676 11348
rect 1631 11308 1676 11336
rect 1670 11296 1676 11308
rect 1728 11296 1734 11348
rect 4755 11339 4813 11345
rect 4755 11305 4767 11339
rect 4801 11305 4813 11339
rect 4755 11299 4813 11305
rect 4770 11268 4798 11299
rect 5442 11296 5448 11348
rect 5500 11336 5506 11348
rect 5721 11339 5779 11345
rect 5721 11336 5733 11339
rect 5500 11308 5733 11336
rect 5500 11296 5506 11308
rect 5721 11305 5733 11308
rect 5767 11305 5779 11339
rect 8570 11336 8576 11348
rect 5721 11299 5779 11305
rect 5828 11308 8576 11336
rect 5828 11268 5856 11308
rect 8570 11296 8576 11308
rect 8628 11296 8634 11348
rect 8846 11336 8852 11348
rect 8807 11308 8852 11336
rect 8846 11296 8852 11308
rect 8904 11296 8910 11348
rect 15749 11339 15807 11345
rect 15749 11305 15761 11339
rect 15795 11305 15807 11339
rect 15749 11299 15807 11305
rect 16715 11339 16773 11345
rect 16715 11305 16727 11339
rect 16761 11336 16773 11339
rect 16850 11336 16856 11348
rect 16761 11308 16856 11336
rect 16761 11305 16773 11308
rect 16715 11299 16773 11305
rect 4770 11240 5856 11268
rect 7190 11228 7196 11280
rect 7248 11268 7254 11280
rect 8021 11271 8079 11277
rect 8021 11268 8033 11271
rect 7248 11240 8033 11268
rect 7248 11228 7254 11240
rect 8021 11237 8033 11240
rect 8067 11237 8079 11271
rect 8021 11231 8079 11237
rect 14642 11228 14648 11280
rect 14700 11268 14706 11280
rect 15764 11268 15792 11299
rect 16850 11296 16856 11308
rect 16908 11296 16914 11348
rect 19058 11296 19064 11348
rect 19116 11336 19122 11348
rect 19245 11339 19303 11345
rect 19245 11336 19257 11339
rect 19116 11308 19257 11336
rect 19116 11296 19122 11308
rect 19245 11305 19257 11308
rect 19291 11305 19303 11339
rect 19245 11299 19303 11305
rect 22922 11296 22928 11348
rect 22980 11336 22986 11348
rect 23753 11339 23811 11345
rect 23753 11336 23765 11339
rect 22980 11308 23765 11336
rect 22980 11296 22986 11308
rect 23753 11305 23765 11308
rect 23799 11336 23811 11339
rect 23842 11336 23848 11348
rect 23799 11308 23848 11336
rect 23799 11305 23811 11308
rect 23753 11299 23811 11305
rect 23842 11296 23848 11308
rect 23900 11296 23906 11348
rect 24486 11336 24492 11348
rect 24447 11308 24492 11336
rect 24486 11296 24492 11308
rect 24544 11296 24550 11348
rect 33459 11339 33517 11345
rect 33459 11305 33471 11339
rect 33505 11336 33517 11339
rect 37734 11336 37740 11348
rect 33505 11308 37740 11336
rect 33505 11305 33517 11308
rect 33459 11299 33517 11305
rect 37734 11296 37740 11308
rect 37792 11296 37798 11348
rect 17494 11268 17500 11280
rect 14700 11240 17500 11268
rect 14700 11228 14706 11240
rect 17494 11228 17500 11240
rect 17552 11228 17558 11280
rect 17586 11228 17592 11280
rect 17644 11268 17650 11280
rect 17819 11271 17877 11277
rect 17819 11268 17831 11271
rect 17644 11240 17831 11268
rect 17644 11228 17650 11240
rect 17819 11237 17831 11240
rect 17865 11237 17877 11271
rect 17819 11231 17877 11237
rect 23014 11228 23020 11280
rect 23072 11268 23078 11280
rect 23072 11240 24348 11268
rect 23072 11228 23078 11240
rect 2406 11200 2412 11212
rect 2367 11172 2412 11200
rect 2406 11160 2412 11172
rect 2464 11160 2470 11212
rect 2685 11203 2743 11209
rect 2685 11169 2697 11203
rect 2731 11200 2743 11203
rect 2866 11200 2872 11212
rect 2731 11172 2872 11200
rect 2731 11169 2743 11172
rect 2685 11163 2743 11169
rect 2866 11160 2872 11172
rect 2924 11160 2930 11212
rect 4617 11203 4675 11209
rect 4617 11169 4629 11203
rect 4663 11200 4675 11203
rect 4706 11200 4712 11212
rect 4663 11172 4712 11200
rect 4663 11169 4675 11172
rect 4617 11163 4675 11169
rect 4706 11160 4712 11172
rect 4764 11160 4770 11212
rect 5905 11203 5963 11209
rect 5905 11169 5917 11203
rect 5951 11169 5963 11203
rect 6178 11200 6184 11212
rect 6139 11172 6184 11200
rect 5905 11163 5963 11169
rect 2774 11132 2780 11144
rect 2735 11104 2780 11132
rect 2774 11092 2780 11104
rect 2832 11092 2838 11144
rect 5920 11132 5948 11163
rect 6178 11160 6184 11172
rect 6236 11160 6242 11212
rect 9582 11160 9588 11212
rect 9640 11200 9646 11212
rect 9712 11203 9770 11209
rect 9712 11200 9724 11203
rect 9640 11172 9724 11200
rect 9640 11160 9646 11172
rect 9712 11169 9724 11172
rect 9758 11169 9770 11203
rect 9712 11163 9770 11169
rect 9858 11160 9864 11212
rect 9916 11200 9922 11212
rect 10724 11203 10782 11209
rect 10724 11200 10736 11203
rect 9916 11172 10736 11200
rect 9916 11160 9922 11172
rect 10724 11169 10736 11172
rect 10770 11200 10782 11203
rect 10962 11200 10968 11212
rect 10770 11172 10968 11200
rect 10770 11169 10782 11172
rect 10724 11163 10782 11169
rect 10962 11160 10968 11172
rect 11020 11160 11026 11212
rect 13906 11160 13912 11212
rect 13964 11200 13970 11212
rect 14220 11203 14278 11209
rect 14220 11200 14232 11203
rect 13964 11172 14232 11200
rect 13964 11160 13970 11172
rect 14220 11169 14232 11172
rect 14266 11169 14278 11203
rect 14220 11163 14278 11169
rect 15565 11203 15623 11209
rect 15565 11169 15577 11203
rect 15611 11200 15623 11203
rect 15838 11200 15844 11212
rect 15611 11172 15844 11200
rect 15611 11169 15623 11172
rect 15565 11163 15623 11169
rect 15838 11160 15844 11172
rect 15896 11160 15902 11212
rect 16482 11160 16488 11212
rect 16540 11200 16546 11212
rect 16612 11203 16670 11209
rect 16612 11200 16624 11203
rect 16540 11172 16624 11200
rect 16540 11160 16546 11172
rect 16612 11169 16624 11172
rect 16658 11169 16670 11203
rect 19334 11200 19340 11212
rect 19295 11172 19340 11200
rect 16612 11163 16670 11169
rect 19334 11160 19340 11172
rect 19392 11160 19398 11212
rect 19705 11203 19763 11209
rect 19705 11169 19717 11203
rect 19751 11200 19763 11203
rect 19794 11200 19800 11212
rect 19751 11172 19800 11200
rect 19751 11169 19763 11172
rect 19705 11163 19763 11169
rect 7929 11135 7987 11141
rect 5920 11104 6408 11132
rect 6380 11076 6408 11104
rect 7929 11101 7941 11135
rect 7975 11132 7987 11135
rect 8662 11132 8668 11144
rect 7975 11104 8668 11132
rect 7975 11101 7987 11104
rect 7929 11095 7987 11101
rect 8662 11092 8668 11104
rect 8720 11092 8726 11144
rect 12250 11092 12256 11144
rect 12308 11132 12314 11144
rect 12897 11135 12955 11141
rect 12897 11132 12909 11135
rect 12308 11104 12909 11132
rect 12308 11092 12314 11104
rect 12897 11101 12909 11104
rect 12943 11101 12955 11135
rect 12897 11095 12955 11101
rect 18601 11135 18659 11141
rect 18601 11101 18613 11135
rect 18647 11132 18659 11135
rect 18690 11132 18696 11144
rect 18647 11104 18696 11132
rect 18647 11101 18659 11104
rect 18601 11095 18659 11101
rect 18690 11092 18696 11104
rect 18748 11132 18754 11144
rect 19720 11132 19748 11163
rect 19794 11160 19800 11172
rect 19852 11160 19858 11212
rect 19978 11160 19984 11212
rect 20036 11200 20042 11212
rect 20968 11203 21026 11209
rect 20968 11200 20980 11203
rect 20036 11172 20980 11200
rect 20036 11160 20042 11172
rect 20968 11169 20980 11172
rect 21014 11200 21026 11203
rect 23360 11203 23418 11209
rect 21014 11172 21312 11200
rect 21014 11169 21026 11172
rect 20968 11163 21026 11169
rect 18748 11104 19748 11132
rect 18748 11092 18754 11104
rect 21284 11076 21312 11172
rect 23360 11169 23372 11203
rect 23406 11200 23418 11203
rect 23474 11200 23480 11212
rect 23406 11172 23480 11200
rect 23406 11169 23418 11172
rect 23360 11163 23418 11169
rect 23474 11160 23480 11172
rect 23532 11160 23538 11212
rect 24320 11209 24348 11240
rect 26252 11240 32203 11268
rect 24305 11203 24363 11209
rect 24305 11169 24317 11203
rect 24351 11200 24363 11203
rect 24854 11200 24860 11212
rect 24351 11172 24860 11200
rect 24351 11169 24363 11172
rect 24305 11163 24363 11169
rect 24854 11160 24860 11172
rect 24912 11160 24918 11212
rect 25222 11160 25228 11212
rect 25280 11200 25286 11212
rect 25444 11203 25502 11209
rect 25444 11200 25456 11203
rect 25280 11172 25456 11200
rect 25280 11160 25286 11172
rect 25444 11169 25456 11172
rect 25490 11200 25502 11203
rect 26252 11200 26280 11240
rect 26418 11200 26424 11212
rect 25490 11172 26280 11200
rect 26379 11172 26424 11200
rect 25490 11169 25502 11172
rect 25444 11163 25502 11169
rect 26418 11160 26424 11172
rect 26476 11160 26482 11212
rect 28445 11203 28503 11209
rect 28445 11169 28457 11203
rect 28491 11169 28503 11203
rect 28626 11200 28632 11212
rect 28587 11172 28632 11200
rect 28445 11163 28503 11169
rect 22097 11135 22155 11141
rect 22097 11101 22109 11135
rect 22143 11132 22155 11135
rect 23014 11132 23020 11144
rect 22143 11104 23020 11132
rect 22143 11101 22155 11104
rect 22097 11095 22155 11101
rect 23014 11092 23020 11104
rect 23072 11092 23078 11144
rect 26970 11132 26976 11144
rect 23446 11104 26976 11132
rect 6362 11024 6368 11076
rect 6420 11064 6426 11076
rect 6917 11067 6975 11073
rect 6917 11064 6929 11067
rect 6420 11036 6929 11064
rect 6420 11024 6426 11036
rect 6917 11033 6929 11036
rect 6963 11064 6975 11067
rect 7006 11064 7012 11076
rect 6963 11036 7012 11064
rect 6963 11033 6975 11036
rect 6917 11027 6975 11033
rect 7006 11024 7012 11036
rect 7064 11064 7070 11076
rect 8478 11064 8484 11076
rect 7064 11036 8340 11064
rect 8439 11036 8484 11064
rect 7064 11024 7070 11036
rect 3142 10996 3148 11008
rect 3103 10968 3148 10996
rect 3142 10956 3148 10968
rect 3200 10956 3206 11008
rect 7190 10996 7196 11008
rect 7151 10968 7196 10996
rect 7190 10956 7196 10968
rect 7248 10956 7254 11008
rect 8312 10996 8340 11036
rect 8478 11024 8484 11036
rect 8536 11024 8542 11076
rect 10226 11064 10232 11076
rect 8588 11036 10232 11064
rect 8588 10996 8616 11036
rect 10226 11024 10232 11036
rect 10284 11024 10290 11076
rect 10827 11067 10885 11073
rect 10827 11033 10839 11067
rect 10873 11064 10885 11067
rect 16390 11064 16396 11076
rect 10873 11036 16396 11064
rect 10873 11033 10885 11036
rect 10827 11027 10885 11033
rect 16390 11024 16396 11036
rect 16448 11024 16454 11076
rect 21266 11024 21272 11076
rect 21324 11064 21330 11076
rect 23446 11064 23474 11104
rect 26970 11092 26976 11104
rect 27028 11092 27034 11144
rect 28460 11132 28488 11163
rect 28626 11160 28632 11172
rect 28684 11160 28690 11212
rect 30926 11200 30932 11212
rect 30887 11172 30932 11200
rect 30926 11160 30932 11172
rect 30984 11160 30990 11212
rect 32175 11209 32203 11240
rect 32160 11203 32218 11209
rect 32160 11169 32172 11203
rect 32206 11200 32218 11203
rect 32582 11200 32588 11212
rect 32206 11172 32588 11200
rect 32206 11169 32218 11172
rect 32160 11163 32218 11169
rect 32582 11160 32588 11172
rect 32640 11160 32646 11212
rect 32674 11160 32680 11212
rect 32732 11200 32738 11212
rect 33229 11203 33287 11209
rect 33229 11200 33241 11203
rect 32732 11172 33241 11200
rect 32732 11160 32738 11172
rect 33229 11169 33241 11172
rect 33275 11169 33287 11203
rect 33229 11163 33287 11169
rect 28534 11132 28540 11144
rect 28460 11104 28540 11132
rect 28534 11092 28540 11104
rect 28592 11092 28598 11144
rect 28902 11132 28908 11144
rect 28863 11104 28908 11132
rect 28902 11092 28908 11104
rect 28960 11092 28966 11144
rect 21324 11036 23474 11064
rect 21324 11024 21330 11036
rect 24210 11024 24216 11076
rect 24268 11064 24274 11076
rect 25547 11067 25605 11073
rect 25547 11064 25559 11067
rect 24268 11036 25559 11064
rect 24268 11024 24274 11036
rect 25547 11033 25559 11036
rect 25593 11033 25605 11067
rect 25547 11027 25605 11033
rect 8312 10968 8616 10996
rect 9674 10956 9680 11008
rect 9732 10996 9738 11008
rect 9815 10999 9873 11005
rect 9815 10996 9827 10999
rect 9732 10968 9827 10996
rect 9732 10956 9738 10968
rect 9815 10965 9827 10968
rect 9861 10965 9873 10999
rect 9815 10959 9873 10965
rect 11793 10999 11851 11005
rect 11793 10965 11805 10999
rect 11839 10996 11851 10999
rect 11882 10996 11888 11008
rect 11839 10968 11888 10996
rect 11839 10965 11851 10968
rect 11793 10959 11851 10965
rect 11882 10956 11888 10968
rect 11940 10956 11946 11008
rect 12023 10999 12081 11005
rect 12023 10965 12035 10999
rect 12069 10996 12081 10999
rect 12434 10996 12440 11008
rect 12069 10968 12440 10996
rect 12069 10965 12081 10968
rect 12023 10959 12081 10965
rect 12434 10956 12440 10968
rect 12492 10956 12498 11008
rect 12618 10996 12624 11008
rect 12579 10968 12624 10996
rect 12618 10956 12624 10968
rect 12676 10956 12682 11008
rect 13538 10956 13544 11008
rect 13596 10996 13602 11008
rect 14323 10999 14381 11005
rect 14323 10996 14335 10999
rect 13596 10968 14335 10996
rect 13596 10956 13602 10968
rect 14323 10965 14335 10968
rect 14369 10965 14381 10999
rect 16022 10996 16028 11008
rect 15983 10968 16028 10996
rect 14323 10959 14381 10965
rect 16022 10956 16028 10968
rect 16080 10956 16086 11008
rect 17589 10999 17647 11005
rect 17589 10965 17601 10999
rect 17635 10996 17647 10999
rect 17770 10996 17776 11008
rect 17635 10968 17776 10996
rect 17635 10965 17647 10968
rect 17589 10959 17647 10965
rect 17770 10956 17776 10968
rect 17828 10956 17834 11008
rect 18230 10996 18236 11008
rect 18191 10968 18236 10996
rect 18230 10956 18236 10968
rect 18288 10956 18294 11008
rect 20162 10956 20168 11008
rect 20220 10996 20226 11008
rect 20257 10999 20315 11005
rect 20257 10996 20269 10999
rect 20220 10968 20269 10996
rect 20220 10956 20226 10968
rect 20257 10965 20269 10968
rect 20303 10996 20315 10999
rect 21039 10999 21097 11005
rect 21039 10996 21051 10999
rect 20303 10968 21051 10996
rect 20303 10965 20315 10968
rect 20257 10959 20315 10965
rect 21039 10965 21051 10968
rect 21085 10965 21097 10999
rect 21039 10959 21097 10965
rect 23290 10956 23296 11008
rect 23348 10996 23354 11008
rect 23431 10999 23489 11005
rect 23431 10996 23443 10999
rect 23348 10968 23443 10996
rect 23348 10956 23354 10968
rect 23431 10965 23443 10968
rect 23477 10965 23489 10999
rect 25866 10996 25872 11008
rect 25827 10968 25872 10996
rect 23431 10959 23489 10965
rect 25866 10956 25872 10968
rect 25924 10956 25930 11008
rect 26651 10999 26709 11005
rect 26651 10965 26663 10999
rect 26697 10996 26709 10999
rect 27062 10996 27068 11008
rect 26697 10968 27068 10996
rect 26697 10965 26709 10968
rect 26651 10959 26709 10965
rect 27062 10956 27068 10968
rect 27120 10956 27126 11008
rect 27706 10996 27712 11008
rect 27667 10968 27712 10996
rect 27706 10956 27712 10968
rect 27764 10956 27770 11008
rect 29270 10996 29276 11008
rect 29231 10968 29276 10996
rect 29270 10956 29276 10968
rect 29328 10956 29334 11008
rect 31159 10999 31217 11005
rect 31159 10965 31171 10999
rect 31205 10996 31217 10999
rect 31570 10996 31576 11008
rect 31205 10968 31576 10996
rect 31205 10965 31217 10968
rect 31159 10959 31217 10965
rect 31570 10956 31576 10968
rect 31628 10956 31634 11008
rect 31662 10956 31668 11008
rect 31720 10996 31726 11008
rect 32263 10999 32321 11005
rect 32263 10996 32275 10999
rect 31720 10968 32275 10996
rect 31720 10956 31726 10968
rect 32263 10965 32275 10968
rect 32309 10965 32321 10999
rect 32263 10959 32321 10965
rect 1104 10906 38824 10928
rect 1104 10854 7648 10906
rect 7700 10854 7712 10906
rect 7764 10854 7776 10906
rect 7828 10854 7840 10906
rect 7892 10854 20982 10906
rect 21034 10854 21046 10906
rect 21098 10854 21110 10906
rect 21162 10854 21174 10906
rect 21226 10854 34315 10906
rect 34367 10854 34379 10906
rect 34431 10854 34443 10906
rect 34495 10854 34507 10906
rect 34559 10854 38824 10906
rect 1104 10832 38824 10854
rect 6273 10795 6331 10801
rect 6273 10761 6285 10795
rect 6319 10792 6331 10795
rect 6362 10792 6368 10804
rect 6319 10764 6368 10792
rect 6319 10761 6331 10764
rect 6273 10755 6331 10761
rect 6362 10752 6368 10764
rect 6420 10752 6426 10804
rect 6546 10752 6552 10804
rect 6604 10792 6610 10804
rect 9582 10792 9588 10804
rect 6604 10764 9588 10792
rect 6604 10752 6610 10764
rect 9582 10752 9588 10764
rect 9640 10792 9646 10804
rect 9677 10795 9735 10801
rect 9677 10792 9689 10795
rect 9640 10764 9689 10792
rect 9640 10752 9646 10764
rect 9677 10761 9689 10764
rect 9723 10761 9735 10795
rect 10962 10792 10968 10804
rect 10923 10764 10968 10792
rect 9677 10755 9735 10761
rect 10962 10752 10968 10764
rect 11020 10752 11026 10804
rect 21177 10795 21235 10801
rect 21177 10761 21189 10795
rect 21223 10792 21235 10795
rect 21266 10792 21272 10804
rect 21223 10764 21272 10792
rect 21223 10761 21235 10764
rect 21177 10755 21235 10761
rect 21266 10752 21272 10764
rect 21324 10752 21330 10804
rect 26418 10792 26424 10804
rect 23032 10764 26424 10792
rect 2866 10724 2872 10736
rect 2779 10696 2872 10724
rect 2866 10684 2872 10696
rect 2924 10724 2930 10736
rect 2924 10696 3924 10724
rect 2924 10684 2930 10696
rect 2682 10616 2688 10668
rect 2740 10656 2746 10668
rect 3050 10656 3056 10668
rect 2740 10628 3056 10656
rect 2740 10616 2746 10628
rect 3050 10616 3056 10628
rect 3108 10616 3114 10668
rect 3896 10656 3924 10696
rect 4154 10684 4160 10736
rect 4212 10724 4218 10736
rect 4212 10696 7420 10724
rect 4212 10684 4218 10696
rect 6270 10656 6276 10668
rect 3896 10628 6276 10656
rect 6270 10616 6276 10628
rect 6328 10616 6334 10668
rect 6914 10616 6920 10668
rect 6972 10656 6978 10668
rect 7392 10665 7420 10696
rect 7944 10696 8984 10724
rect 7944 10668 7972 10696
rect 7101 10659 7159 10665
rect 7101 10656 7113 10659
rect 6972 10628 7113 10656
rect 6972 10616 6978 10628
rect 7101 10625 7113 10628
rect 7147 10625 7159 10659
rect 7101 10619 7159 10625
rect 7377 10659 7435 10665
rect 7377 10625 7389 10659
rect 7423 10656 7435 10659
rect 7926 10656 7932 10668
rect 7423 10628 7932 10656
rect 7423 10625 7435 10628
rect 7377 10619 7435 10625
rect 7926 10616 7932 10628
rect 7984 10616 7990 10668
rect 8665 10659 8723 10665
rect 8665 10625 8677 10659
rect 8711 10656 8723 10659
rect 8846 10656 8852 10668
rect 8711 10628 8852 10656
rect 8711 10625 8723 10628
rect 8665 10619 8723 10625
rect 8846 10616 8852 10628
rect 8904 10616 8910 10668
rect 8956 10665 8984 10696
rect 11882 10684 11888 10736
rect 11940 10724 11946 10736
rect 13906 10724 13912 10736
rect 11940 10696 13912 10724
rect 11940 10684 11946 10696
rect 13906 10684 13912 10696
rect 13964 10684 13970 10736
rect 15749 10727 15807 10733
rect 15749 10693 15761 10727
rect 15795 10724 15807 10727
rect 16022 10724 16028 10736
rect 15795 10696 16028 10724
rect 15795 10693 15807 10696
rect 15749 10687 15807 10693
rect 16022 10684 16028 10696
rect 16080 10724 16086 10736
rect 16298 10724 16304 10736
rect 16080 10696 16304 10724
rect 16080 10684 16086 10696
rect 16298 10684 16304 10696
rect 16356 10684 16362 10736
rect 19794 10684 19800 10736
rect 19852 10724 19858 10736
rect 19981 10727 20039 10733
rect 19981 10724 19993 10727
rect 19852 10696 19993 10724
rect 19852 10684 19858 10696
rect 19981 10693 19993 10696
rect 20027 10724 20039 10727
rect 22830 10724 22836 10736
rect 20027 10696 22836 10724
rect 20027 10693 20039 10696
rect 19981 10687 20039 10693
rect 22830 10684 22836 10696
rect 22888 10684 22894 10736
rect 8941 10659 8999 10665
rect 8941 10625 8953 10659
rect 8987 10625 8999 10659
rect 8941 10619 8999 10625
rect 13630 10616 13636 10668
rect 13688 10656 13694 10668
rect 14553 10659 14611 10665
rect 14553 10656 14565 10659
rect 13688 10628 14565 10656
rect 13688 10616 13694 10628
rect 14553 10625 14565 10628
rect 14599 10625 14611 10659
rect 16666 10656 16672 10668
rect 14553 10619 14611 10625
rect 15672 10628 16672 10656
rect 1578 10588 1584 10600
rect 1539 10560 1584 10588
rect 1578 10548 1584 10560
rect 1636 10548 1642 10600
rect 1949 10591 2007 10597
rect 1949 10557 1961 10591
rect 1995 10588 2007 10591
rect 2866 10588 2872 10600
rect 1995 10560 2872 10588
rect 1995 10557 2007 10560
rect 1949 10551 2007 10557
rect 2866 10548 2872 10560
rect 2924 10548 2930 10600
rect 5077 10591 5135 10597
rect 5077 10557 5089 10591
rect 5123 10588 5135 10591
rect 5445 10591 5503 10597
rect 5445 10588 5457 10591
rect 5123 10560 5457 10588
rect 5123 10557 5135 10560
rect 5077 10551 5135 10557
rect 5445 10557 5457 10560
rect 5491 10557 5503 10591
rect 5626 10588 5632 10600
rect 5587 10560 5632 10588
rect 5445 10551 5503 10557
rect 2130 10520 2136 10532
rect 2091 10492 2136 10520
rect 2130 10480 2136 10492
rect 2188 10480 2194 10532
rect 3142 10480 3148 10532
rect 3200 10520 3206 10532
rect 3697 10523 3755 10529
rect 3200 10492 3245 10520
rect 3200 10480 3206 10492
rect 3697 10489 3709 10523
rect 3743 10520 3755 10523
rect 5460 10520 5488 10551
rect 5626 10548 5632 10560
rect 5684 10588 5690 10600
rect 6178 10588 6184 10600
rect 5684 10560 6184 10588
rect 5684 10548 5690 10560
rect 6178 10548 6184 10560
rect 6236 10588 6242 10600
rect 6549 10591 6607 10597
rect 6549 10588 6561 10591
rect 6236 10560 6561 10588
rect 6236 10548 6242 10560
rect 6549 10557 6561 10560
rect 6595 10557 6607 10591
rect 6549 10551 6607 10557
rect 10204 10591 10262 10597
rect 10204 10557 10216 10591
rect 10250 10588 10262 10591
rect 10250 10560 10732 10588
rect 10250 10557 10262 10560
rect 10204 10551 10262 10557
rect 3743 10492 4154 10520
rect 5460 10492 5810 10520
rect 3743 10489 3755 10492
rect 3697 10483 3755 10489
rect 1670 10412 1676 10464
rect 1728 10452 1734 10464
rect 2406 10452 2412 10464
rect 1728 10424 2412 10452
rect 1728 10412 1734 10424
rect 2406 10412 2412 10424
rect 2464 10412 2470 10464
rect 4126 10452 4154 10492
rect 4706 10452 4712 10464
rect 4126 10424 4712 10452
rect 4706 10412 4712 10424
rect 4764 10412 4770 10464
rect 5074 10412 5080 10464
rect 5132 10452 5138 10464
rect 5261 10455 5319 10461
rect 5261 10452 5273 10455
rect 5132 10424 5273 10452
rect 5132 10412 5138 10424
rect 5261 10421 5273 10424
rect 5307 10421 5319 10455
rect 5782 10452 5810 10492
rect 6086 10480 6092 10532
rect 6144 10520 6150 10532
rect 7190 10520 7196 10532
rect 6144 10492 7196 10520
rect 6144 10480 6150 10492
rect 7190 10480 7196 10492
rect 7248 10480 7254 10532
rect 8757 10523 8815 10529
rect 8757 10489 8769 10523
rect 8803 10489 8815 10523
rect 8757 10483 8815 10489
rect 7006 10452 7012 10464
rect 5782 10424 7012 10452
rect 5261 10415 5319 10421
rect 7006 10412 7012 10424
rect 7064 10412 7070 10464
rect 7208 10452 7236 10480
rect 8021 10455 8079 10461
rect 8021 10452 8033 10455
rect 7208 10424 8033 10452
rect 8021 10421 8033 10424
rect 8067 10421 8079 10455
rect 8386 10452 8392 10464
rect 8347 10424 8392 10452
rect 8021 10415 8079 10421
rect 8386 10412 8392 10424
rect 8444 10452 8450 10464
rect 8772 10452 8800 10483
rect 8444 10424 8800 10452
rect 8444 10412 8450 10424
rect 9766 10412 9772 10464
rect 9824 10452 9830 10464
rect 10704 10461 10732 10560
rect 10962 10548 10968 10600
rect 11020 10588 11026 10600
rect 11184 10591 11242 10597
rect 11184 10588 11196 10591
rect 11020 10560 11196 10588
rect 11020 10548 11026 10560
rect 11184 10557 11196 10560
rect 11230 10557 11242 10591
rect 11882 10588 11888 10600
rect 11843 10560 11888 10588
rect 11184 10551 11242 10557
rect 11882 10548 11888 10560
rect 11940 10548 11946 10600
rect 12250 10548 12256 10600
rect 12308 10588 12314 10600
rect 12529 10591 12587 10597
rect 12529 10588 12541 10591
rect 12308 10560 12541 10588
rect 12308 10548 12314 10560
rect 12529 10557 12541 10560
rect 12575 10557 12587 10591
rect 12529 10551 12587 10557
rect 12618 10548 12624 10600
rect 12676 10588 12682 10600
rect 12989 10591 13047 10597
rect 12989 10588 13001 10591
rect 12676 10560 13001 10588
rect 12676 10548 12682 10560
rect 12989 10557 13001 10560
rect 13035 10557 13047 10591
rect 12989 10551 13047 10557
rect 14090 10548 14096 10600
rect 14148 10588 14154 10600
rect 14642 10588 14648 10600
rect 14148 10560 14193 10588
rect 14603 10560 14648 10588
rect 14148 10548 14154 10560
rect 14642 10548 14648 10560
rect 14700 10548 14706 10600
rect 15672 10597 15700 10628
rect 16666 10616 16672 10628
rect 16724 10616 16730 10668
rect 15657 10591 15715 10597
rect 15657 10557 15669 10591
rect 15703 10557 15715 10591
rect 15657 10551 15715 10557
rect 15933 10591 15991 10597
rect 15933 10557 15945 10591
rect 15979 10557 15991 10591
rect 15933 10551 15991 10557
rect 18417 10591 18475 10597
rect 18417 10557 18429 10591
rect 18463 10588 18475 10591
rect 18785 10591 18843 10597
rect 18785 10588 18797 10591
rect 18463 10560 18797 10588
rect 18463 10557 18475 10560
rect 18417 10551 18475 10557
rect 18785 10557 18797 10560
rect 18831 10588 18843 10591
rect 18874 10588 18880 10600
rect 18831 10560 18880 10588
rect 18831 10557 18843 10560
rect 18785 10551 18843 10557
rect 13262 10520 13268 10532
rect 13223 10492 13268 10520
rect 13262 10480 13268 10492
rect 13320 10480 13326 10532
rect 15948 10520 15976 10551
rect 18874 10548 18880 10560
rect 18932 10548 18938 10600
rect 19061 10591 19119 10597
rect 19061 10557 19073 10591
rect 19107 10588 19119 10591
rect 19426 10588 19432 10600
rect 19107 10560 19432 10588
rect 19107 10557 19119 10560
rect 19061 10551 19119 10557
rect 19426 10548 19432 10560
rect 19484 10588 19490 10600
rect 19812 10588 19840 10684
rect 20162 10656 20168 10668
rect 20123 10628 20168 10656
rect 20162 10616 20168 10628
rect 20220 10616 20226 10668
rect 19484 10560 19840 10588
rect 19484 10548 19490 10560
rect 22370 10548 22376 10600
rect 22428 10588 22434 10600
rect 22554 10588 22560 10600
rect 22612 10597 22618 10600
rect 23032 10597 23060 10764
rect 26418 10752 26424 10764
rect 26476 10792 26482 10804
rect 26605 10795 26663 10801
rect 26605 10792 26617 10795
rect 26476 10764 26617 10792
rect 26476 10752 26482 10764
rect 26605 10761 26617 10764
rect 26651 10761 26663 10795
rect 32582 10792 32588 10804
rect 32543 10764 32588 10792
rect 26605 10755 26663 10761
rect 32582 10752 32588 10764
rect 32640 10792 32646 10804
rect 35434 10792 35440 10804
rect 32640 10764 35440 10792
rect 32640 10752 32646 10764
rect 35434 10752 35440 10764
rect 35492 10752 35498 10804
rect 28810 10684 28816 10736
rect 28868 10724 28874 10736
rect 29270 10724 29276 10736
rect 28868 10696 29276 10724
rect 28868 10684 28874 10696
rect 29270 10684 29276 10696
rect 29328 10724 29334 10736
rect 29328 10696 29408 10724
rect 29328 10684 29334 10696
rect 23842 10656 23848 10668
rect 23803 10628 23848 10656
rect 23842 10616 23848 10628
rect 23900 10616 23906 10668
rect 24670 10616 24676 10668
rect 24728 10656 24734 10668
rect 28997 10659 29055 10665
rect 28997 10656 29009 10659
rect 24728 10628 29009 10656
rect 24728 10616 24734 10628
rect 28997 10625 29009 10628
rect 29043 10656 29055 10659
rect 29043 10628 29316 10656
rect 29043 10625 29055 10628
rect 28997 10619 29055 10625
rect 22612 10591 22650 10597
rect 22428 10560 22560 10588
rect 22428 10548 22434 10560
rect 22554 10548 22560 10560
rect 22638 10588 22650 10591
rect 23017 10591 23075 10597
rect 23017 10588 23029 10591
rect 22638 10560 23029 10588
rect 22638 10557 22650 10560
rect 22612 10551 22650 10557
rect 23017 10557 23029 10560
rect 23063 10557 23075 10591
rect 24854 10588 24860 10600
rect 24767 10560 24860 10588
rect 23017 10551 23075 10557
rect 22612 10548 22618 10551
rect 24854 10548 24860 10560
rect 24912 10588 24918 10600
rect 25406 10588 25412 10600
rect 24912 10560 25412 10588
rect 24912 10548 24918 10560
rect 25406 10548 25412 10560
rect 25464 10548 25470 10600
rect 25498 10548 25504 10600
rect 25556 10588 25562 10600
rect 25593 10591 25651 10597
rect 25593 10588 25605 10591
rect 25556 10560 25605 10588
rect 25556 10548 25562 10560
rect 25593 10557 25605 10560
rect 25639 10588 25651 10591
rect 25866 10588 25872 10600
rect 25639 10560 25872 10588
rect 25639 10557 25651 10560
rect 25593 10551 25651 10557
rect 25866 10548 25872 10560
rect 25924 10548 25930 10600
rect 26050 10588 26056 10600
rect 26011 10560 26056 10588
rect 26050 10548 26056 10560
rect 26108 10548 26114 10600
rect 27433 10591 27491 10597
rect 27433 10588 27445 10591
rect 26160 10560 27445 10588
rect 15120 10492 15976 10520
rect 10275 10455 10333 10461
rect 10275 10452 10287 10455
rect 9824 10424 10287 10452
rect 9824 10412 9830 10424
rect 10275 10421 10287 10424
rect 10321 10421 10333 10455
rect 10275 10415 10333 10421
rect 10689 10455 10747 10461
rect 10689 10421 10701 10455
rect 10735 10452 10747 10455
rect 10778 10452 10784 10464
rect 10735 10424 10784 10452
rect 10735 10421 10747 10424
rect 10689 10415 10747 10421
rect 10778 10412 10784 10424
rect 10836 10412 10842 10464
rect 11054 10412 11060 10464
rect 11112 10452 11118 10464
rect 11287 10455 11345 10461
rect 11287 10452 11299 10455
rect 11112 10424 11299 10452
rect 11112 10412 11118 10424
rect 11287 10421 11299 10424
rect 11333 10421 11345 10455
rect 11287 10415 11345 10421
rect 13633 10455 13691 10461
rect 13633 10421 13645 10455
rect 13679 10452 13691 10455
rect 13814 10452 13820 10464
rect 13679 10424 13820 10452
rect 13679 10421 13691 10424
rect 13633 10415 13691 10421
rect 13814 10412 13820 10424
rect 13872 10412 13878 10464
rect 14918 10412 14924 10464
rect 14976 10452 14982 10464
rect 15120 10461 15148 10492
rect 16022 10480 16028 10532
rect 16080 10520 16086 10532
rect 16482 10520 16488 10532
rect 16080 10492 16488 10520
rect 16080 10480 16086 10492
rect 16482 10480 16488 10492
rect 16540 10520 16546 10532
rect 17037 10523 17095 10529
rect 17037 10520 17049 10523
rect 16540 10492 17049 10520
rect 16540 10480 16546 10492
rect 17037 10489 17049 10492
rect 17083 10489 17095 10523
rect 19242 10520 19248 10532
rect 19203 10492 19248 10520
rect 17037 10483 17095 10489
rect 19242 10480 19248 10492
rect 19300 10480 19306 10532
rect 20162 10480 20168 10532
rect 20220 10520 20226 10532
rect 20257 10523 20315 10529
rect 20257 10520 20269 10523
rect 20220 10492 20269 10520
rect 20220 10480 20226 10492
rect 20257 10489 20269 10492
rect 20303 10489 20315 10523
rect 20806 10520 20812 10532
rect 20767 10492 20812 10520
rect 20257 10483 20315 10489
rect 20806 10480 20812 10492
rect 20864 10480 20870 10532
rect 22462 10480 22468 10532
rect 22520 10520 22526 10532
rect 23934 10520 23940 10532
rect 22520 10492 23831 10520
rect 23895 10492 23940 10520
rect 22520 10480 22526 10492
rect 15105 10455 15163 10461
rect 15105 10452 15117 10455
rect 14976 10424 15117 10452
rect 14976 10412 14982 10424
rect 15105 10421 15117 10424
rect 15151 10421 15163 10455
rect 15105 10415 15163 10421
rect 15565 10455 15623 10461
rect 15565 10421 15577 10455
rect 15611 10452 15623 10455
rect 15838 10452 15844 10464
rect 15611 10424 15844 10452
rect 15611 10421 15623 10424
rect 15565 10415 15623 10421
rect 15838 10412 15844 10424
rect 15896 10412 15902 10464
rect 16114 10452 16120 10464
rect 16075 10424 16120 10452
rect 16114 10412 16120 10424
rect 16172 10412 16178 10464
rect 16666 10452 16672 10464
rect 16627 10424 16672 10452
rect 16666 10412 16672 10424
rect 16724 10412 16730 10464
rect 17770 10452 17776 10464
rect 17731 10424 17776 10452
rect 17770 10412 17776 10424
rect 17828 10412 17834 10464
rect 19334 10412 19340 10464
rect 19392 10452 19398 10464
rect 19521 10455 19579 10461
rect 19521 10452 19533 10455
rect 19392 10424 19533 10452
rect 19392 10412 19398 10424
rect 19521 10421 19533 10424
rect 19567 10421 19579 10455
rect 19521 10415 19579 10421
rect 22695 10455 22753 10461
rect 22695 10421 22707 10455
rect 22741 10452 22753 10455
rect 22922 10452 22928 10464
rect 22741 10424 22928 10452
rect 22741 10421 22753 10424
rect 22695 10415 22753 10421
rect 22922 10412 22928 10424
rect 22980 10412 22986 10464
rect 23474 10412 23480 10464
rect 23532 10452 23538 10464
rect 23803 10452 23831 10492
rect 23934 10480 23940 10492
rect 23992 10480 23998 10532
rect 24489 10523 24547 10529
rect 24489 10489 24501 10523
rect 24535 10520 24547 10523
rect 24578 10520 24584 10532
rect 24535 10492 24584 10520
rect 24535 10489 24547 10492
rect 24489 10483 24547 10489
rect 24578 10480 24584 10492
rect 24636 10480 24642 10532
rect 26160 10520 26188 10560
rect 27433 10557 27445 10560
rect 27479 10588 27491 10591
rect 27522 10588 27528 10600
rect 27479 10560 27528 10588
rect 27479 10557 27491 10560
rect 27433 10551 27491 10557
rect 27522 10548 27528 10560
rect 27580 10588 27586 10600
rect 27617 10591 27675 10597
rect 27617 10588 27629 10591
rect 27580 10560 27629 10588
rect 27580 10548 27586 10560
rect 27617 10557 27629 10560
rect 27663 10557 27675 10591
rect 27617 10551 27675 10557
rect 27706 10548 27712 10600
rect 27764 10588 27770 10600
rect 28169 10591 28227 10597
rect 28169 10588 28181 10591
rect 27764 10560 28181 10588
rect 27764 10548 27770 10560
rect 28169 10557 28181 10560
rect 28215 10588 28227 10591
rect 28810 10588 28816 10600
rect 28215 10560 28816 10588
rect 28215 10557 28227 10560
rect 28169 10551 28227 10557
rect 28810 10548 28816 10560
rect 28868 10548 28874 10600
rect 29288 10597 29316 10628
rect 29273 10591 29331 10597
rect 29273 10557 29285 10591
rect 29319 10557 29331 10591
rect 29380 10588 29408 10696
rect 30926 10684 30932 10736
rect 30984 10724 30990 10736
rect 31113 10727 31171 10733
rect 31113 10724 31125 10727
rect 30984 10696 31125 10724
rect 30984 10684 30990 10696
rect 31113 10693 31125 10696
rect 31159 10724 31171 10727
rect 35250 10724 35256 10736
rect 31159 10696 35256 10724
rect 31159 10693 31171 10696
rect 31113 10687 31171 10693
rect 35250 10684 35256 10696
rect 35308 10684 35314 10736
rect 31662 10656 31668 10668
rect 31623 10628 31668 10656
rect 31662 10616 31668 10628
rect 31720 10616 31726 10668
rect 32674 10616 32680 10668
rect 32732 10656 32738 10668
rect 33965 10659 34023 10665
rect 33965 10656 33977 10659
rect 32732 10628 33977 10656
rect 32732 10616 32738 10628
rect 33965 10625 33977 10628
rect 34011 10625 34023 10659
rect 33965 10619 34023 10625
rect 29733 10591 29791 10597
rect 29733 10588 29745 10591
rect 29380 10560 29745 10588
rect 29273 10551 29331 10557
rect 29733 10557 29745 10560
rect 29779 10557 29791 10591
rect 29733 10551 29791 10557
rect 33204 10591 33262 10597
rect 33204 10557 33216 10591
rect 33250 10588 33262 10591
rect 33597 10591 33655 10597
rect 33597 10588 33609 10591
rect 33250 10560 33609 10588
rect 33250 10557 33262 10560
rect 33204 10551 33262 10557
rect 33597 10557 33609 10560
rect 33643 10588 33655 10591
rect 35894 10588 35900 10600
rect 33643 10560 35900 10588
rect 33643 10557 33655 10560
rect 33597 10551 33655 10557
rect 35894 10548 35900 10560
rect 35952 10548 35958 10600
rect 26326 10520 26332 10532
rect 24688 10492 26188 10520
rect 26287 10492 26332 10520
rect 24688 10452 24716 10492
rect 26326 10480 26332 10492
rect 26384 10480 26390 10532
rect 28353 10523 28411 10529
rect 28353 10489 28365 10523
rect 28399 10520 28411 10523
rect 29822 10520 29828 10532
rect 28399 10492 29828 10520
rect 28399 10489 28411 10492
rect 28353 10483 28411 10489
rect 29822 10480 29828 10492
rect 29880 10480 29886 10532
rect 30006 10520 30012 10532
rect 29967 10492 30012 10520
rect 30006 10480 30012 10492
rect 30064 10480 30070 10532
rect 31478 10520 31484 10532
rect 31391 10492 31484 10520
rect 31478 10480 31484 10492
rect 31536 10520 31542 10532
rect 31757 10523 31815 10529
rect 31757 10520 31769 10523
rect 31536 10492 31769 10520
rect 31536 10480 31542 10492
rect 31757 10489 31769 10492
rect 31803 10489 31815 10523
rect 31757 10483 31815 10489
rect 32309 10523 32367 10529
rect 32309 10489 32321 10523
rect 32355 10520 32367 10523
rect 32490 10520 32496 10532
rect 32355 10492 32496 10520
rect 32355 10489 32367 10492
rect 32309 10483 32367 10489
rect 32490 10480 32496 10492
rect 32548 10480 32554 10532
rect 23532 10424 23577 10452
rect 23803 10424 24716 10452
rect 23532 10412 23538 10424
rect 24762 10412 24768 10464
rect 24820 10452 24826 10464
rect 25222 10452 25228 10464
rect 24820 10424 25228 10452
rect 24820 10412 24826 10424
rect 25222 10412 25228 10424
rect 25280 10452 25286 10464
rect 25409 10455 25467 10461
rect 25409 10452 25421 10455
rect 25280 10424 25421 10452
rect 25280 10412 25286 10424
rect 25409 10421 25421 10424
rect 25455 10421 25467 10455
rect 25409 10415 25467 10421
rect 28626 10412 28632 10464
rect 28684 10452 28690 10464
rect 28721 10455 28779 10461
rect 28721 10452 28733 10455
rect 28684 10424 28733 10452
rect 28684 10412 28690 10424
rect 28721 10421 28733 10424
rect 28767 10452 28779 10455
rect 29638 10452 29644 10464
rect 28767 10424 29644 10452
rect 28767 10421 28779 10424
rect 28721 10415 28779 10421
rect 29638 10412 29644 10424
rect 29696 10412 29702 10464
rect 33275 10455 33333 10461
rect 33275 10421 33287 10455
rect 33321 10452 33333 10455
rect 33502 10452 33508 10464
rect 33321 10424 33508 10452
rect 33321 10421 33333 10424
rect 33275 10415 33333 10421
rect 33502 10412 33508 10424
rect 33560 10412 33566 10464
rect 1104 10362 38824 10384
rect 1104 10310 14315 10362
rect 14367 10310 14379 10362
rect 14431 10310 14443 10362
rect 14495 10310 14507 10362
rect 14559 10310 27648 10362
rect 27700 10310 27712 10362
rect 27764 10310 27776 10362
rect 27828 10310 27840 10362
rect 27892 10310 38824 10362
rect 1104 10288 38824 10310
rect 1578 10208 1584 10260
rect 1636 10248 1642 10260
rect 1949 10251 2007 10257
rect 1949 10248 1961 10251
rect 1636 10220 1961 10248
rect 1636 10208 1642 10220
rect 1949 10217 1961 10220
rect 1995 10217 2007 10251
rect 2222 10248 2228 10260
rect 2183 10220 2228 10248
rect 1949 10211 2007 10217
rect 2222 10208 2228 10220
rect 2280 10208 2286 10260
rect 3050 10208 3056 10260
rect 3108 10248 3114 10260
rect 3145 10251 3203 10257
rect 3145 10248 3157 10251
rect 3108 10220 3157 10248
rect 3108 10208 3114 10220
rect 3145 10217 3157 10220
rect 3191 10217 3203 10251
rect 5718 10248 5724 10260
rect 5679 10220 5724 10248
rect 3145 10211 3203 10217
rect 5718 10208 5724 10220
rect 5776 10208 5782 10260
rect 7098 10248 7104 10260
rect 7059 10220 7104 10248
rect 7098 10208 7104 10220
rect 7156 10208 7162 10260
rect 8662 10248 8668 10260
rect 8623 10220 8668 10248
rect 8662 10208 8668 10220
rect 8720 10208 8726 10260
rect 10962 10208 10968 10260
rect 11020 10248 11026 10260
rect 11149 10251 11207 10257
rect 11149 10248 11161 10251
rect 11020 10220 11161 10248
rect 11020 10208 11026 10220
rect 11149 10217 11161 10220
rect 11195 10217 11207 10251
rect 11149 10211 11207 10217
rect 12434 10208 12440 10260
rect 12492 10248 12498 10260
rect 13081 10251 13139 10257
rect 13081 10248 13093 10251
rect 12492 10220 13093 10248
rect 12492 10208 12498 10220
rect 13081 10217 13093 10220
rect 13127 10217 13139 10251
rect 13722 10248 13728 10260
rect 13683 10220 13728 10248
rect 13081 10211 13139 10217
rect 13722 10208 13728 10220
rect 13780 10208 13786 10260
rect 16574 10208 16580 10260
rect 16632 10248 16638 10260
rect 17037 10251 17095 10257
rect 17037 10248 17049 10251
rect 16632 10220 17049 10248
rect 16632 10208 16638 10220
rect 17037 10217 17049 10220
rect 17083 10217 17095 10251
rect 17954 10248 17960 10260
rect 17915 10220 17960 10248
rect 17037 10211 17095 10217
rect 17954 10208 17960 10220
rect 18012 10208 18018 10260
rect 22738 10248 22744 10260
rect 22699 10220 22744 10248
rect 22738 10208 22744 10220
rect 22796 10208 22802 10260
rect 27062 10248 27068 10260
rect 27023 10220 27068 10248
rect 27062 10208 27068 10220
rect 27120 10208 27126 10260
rect 31662 10248 31668 10260
rect 31623 10220 31668 10248
rect 31662 10208 31668 10220
rect 31720 10208 31726 10260
rect 1673 10183 1731 10189
rect 1673 10149 1685 10183
rect 1719 10180 1731 10183
rect 2038 10180 2044 10192
rect 1719 10152 2044 10180
rect 1719 10149 1731 10152
rect 1673 10143 1731 10149
rect 2038 10140 2044 10152
rect 2096 10180 2102 10192
rect 2096 10152 2728 10180
rect 2096 10140 2102 10152
rect 2700 10121 2728 10152
rect 3970 10140 3976 10192
rect 4028 10180 4034 10192
rect 4249 10183 4307 10189
rect 4249 10180 4261 10183
rect 4028 10152 4261 10180
rect 4028 10140 4034 10152
rect 4249 10149 4261 10152
rect 4295 10149 4307 10183
rect 4249 10143 4307 10149
rect 6914 10140 6920 10192
rect 6972 10180 6978 10192
rect 7377 10183 7435 10189
rect 7377 10180 7389 10183
rect 6972 10152 7389 10180
rect 6972 10140 6978 10152
rect 7377 10149 7389 10152
rect 7423 10149 7435 10183
rect 7377 10143 7435 10149
rect 7837 10183 7895 10189
rect 7837 10149 7849 10183
rect 7883 10180 7895 10183
rect 8202 10180 8208 10192
rect 7883 10152 8208 10180
rect 7883 10149 7895 10152
rect 7837 10143 7895 10149
rect 8202 10140 8208 10152
rect 8260 10140 8266 10192
rect 9766 10180 9772 10192
rect 9727 10152 9772 10180
rect 9766 10140 9772 10152
rect 9824 10140 9830 10192
rect 9858 10140 9864 10192
rect 9916 10180 9922 10192
rect 15105 10183 15163 10189
rect 9916 10152 9961 10180
rect 9916 10140 9922 10152
rect 15105 10149 15117 10183
rect 15151 10180 15163 10183
rect 15378 10180 15384 10192
rect 15151 10152 15384 10180
rect 15151 10149 15163 10152
rect 15105 10143 15163 10149
rect 15378 10140 15384 10152
rect 15436 10180 15442 10192
rect 15473 10183 15531 10189
rect 15473 10180 15485 10183
rect 15436 10152 15485 10180
rect 15436 10140 15442 10152
rect 15473 10149 15485 10152
rect 15519 10149 15531 10183
rect 18230 10180 18236 10192
rect 18191 10152 18236 10180
rect 15473 10143 15531 10149
rect 18230 10140 18236 10152
rect 18288 10140 18294 10192
rect 21085 10183 21143 10189
rect 21085 10149 21097 10183
rect 21131 10180 21143 10183
rect 21266 10180 21272 10192
rect 21131 10152 21272 10180
rect 21131 10149 21143 10152
rect 21085 10143 21143 10149
rect 21266 10140 21272 10152
rect 21324 10140 21330 10192
rect 23934 10140 23940 10192
rect 23992 10180 23998 10192
rect 24489 10183 24547 10189
rect 24489 10180 24501 10183
rect 23992 10152 24501 10180
rect 23992 10140 23998 10152
rect 24489 10149 24501 10152
rect 24535 10149 24547 10183
rect 24489 10143 24547 10149
rect 27338 10140 27344 10192
rect 27396 10180 27402 10192
rect 27706 10180 27712 10192
rect 27396 10152 27712 10180
rect 27396 10140 27402 10152
rect 27706 10140 27712 10152
rect 27764 10140 27770 10192
rect 27801 10183 27859 10189
rect 27801 10149 27813 10183
rect 27847 10180 27859 10183
rect 28166 10180 28172 10192
rect 27847 10152 28172 10180
rect 27847 10149 27859 10152
rect 27801 10143 27859 10149
rect 28166 10140 28172 10152
rect 28224 10140 28230 10192
rect 31570 10140 31576 10192
rect 31628 10180 31634 10192
rect 32217 10183 32275 10189
rect 32217 10180 32229 10183
rect 31628 10152 32229 10180
rect 31628 10140 31634 10152
rect 32217 10149 32229 10152
rect 32263 10149 32275 10183
rect 32217 10143 32275 10149
rect 32306 10140 32312 10192
rect 32364 10180 32370 10192
rect 33870 10180 33876 10192
rect 32364 10152 32409 10180
rect 33831 10152 33876 10180
rect 32364 10140 32370 10152
rect 33870 10140 33876 10152
rect 33928 10140 33934 10192
rect 2409 10115 2467 10121
rect 2409 10081 2421 10115
rect 2455 10081 2467 10115
rect 2409 10075 2467 10081
rect 2685 10115 2743 10121
rect 2685 10081 2697 10115
rect 2731 10112 2743 10115
rect 2866 10112 2872 10124
rect 2731 10084 2872 10112
rect 2731 10081 2743 10084
rect 2685 10075 2743 10081
rect 2424 10044 2452 10075
rect 2866 10072 2872 10084
rect 2924 10072 2930 10124
rect 5534 10072 5540 10124
rect 5592 10112 5598 10124
rect 5629 10115 5687 10121
rect 5629 10112 5641 10115
rect 5592 10084 5641 10112
rect 5592 10072 5598 10084
rect 5629 10081 5641 10084
rect 5675 10081 5687 10115
rect 5629 10075 5687 10081
rect 6181 10115 6239 10121
rect 6181 10081 6193 10115
rect 6227 10112 6239 10115
rect 6270 10112 6276 10124
rect 6227 10084 6276 10112
rect 6227 10081 6239 10084
rect 6181 10075 6239 10081
rect 3602 10044 3608 10056
rect 2424 10016 3608 10044
rect 3602 10004 3608 10016
rect 3660 10004 3666 10056
rect 4154 10004 4160 10056
rect 4212 10044 4218 10056
rect 4212 10016 4257 10044
rect 4212 10004 4218 10016
rect 4706 9976 4712 9988
rect 4667 9948 4712 9976
rect 4706 9936 4712 9948
rect 4764 9936 4770 9988
rect 5644 9976 5672 10075
rect 6270 10072 6276 10084
rect 6328 10072 6334 10124
rect 12342 10112 12348 10124
rect 12303 10084 12348 10112
rect 12342 10072 12348 10084
rect 12400 10072 12406 10124
rect 12526 10112 12532 10124
rect 12487 10084 12532 10112
rect 12526 10072 12532 10084
rect 12584 10072 12590 10124
rect 13265 10115 13323 10121
rect 13265 10081 13277 10115
rect 13311 10112 13323 10115
rect 13633 10115 13691 10121
rect 13633 10112 13645 10115
rect 13311 10084 13645 10112
rect 13311 10081 13323 10084
rect 13265 10075 13323 10081
rect 13633 10081 13645 10084
rect 13679 10081 13691 10115
rect 13633 10075 13691 10081
rect 6822 10004 6828 10056
rect 6880 10044 6886 10056
rect 7745 10047 7803 10053
rect 7745 10044 7757 10047
rect 6880 10016 7757 10044
rect 6880 10004 6886 10016
rect 7745 10013 7757 10016
rect 7791 10013 7803 10047
rect 7745 10007 7803 10013
rect 7926 10004 7932 10056
rect 7984 10044 7990 10056
rect 8021 10047 8079 10053
rect 8021 10044 8033 10047
rect 7984 10016 8033 10044
rect 7984 10004 7990 10016
rect 8021 10013 8033 10016
rect 8067 10013 8079 10047
rect 10042 10044 10048 10056
rect 10003 10016 10048 10044
rect 8021 10007 8079 10013
rect 10042 10004 10048 10016
rect 10100 10004 10106 10056
rect 12805 10047 12863 10053
rect 12805 10013 12817 10047
rect 12851 10044 12863 10047
rect 13354 10044 13360 10056
rect 12851 10016 13360 10044
rect 12851 10013 12863 10016
rect 12805 10007 12863 10013
rect 13354 10004 13360 10016
rect 13412 10004 13418 10056
rect 13446 10004 13452 10056
rect 13504 10044 13510 10056
rect 13648 10044 13676 10075
rect 13814 10072 13820 10124
rect 13872 10112 13878 10124
rect 14090 10112 14096 10124
rect 13872 10084 14096 10112
rect 13872 10072 13878 10084
rect 14090 10072 14096 10084
rect 14148 10112 14154 10124
rect 14185 10115 14243 10121
rect 14185 10112 14197 10115
rect 14148 10084 14197 10112
rect 14148 10072 14154 10084
rect 14185 10081 14197 10084
rect 14231 10112 14243 10115
rect 14642 10112 14648 10124
rect 14231 10084 14648 10112
rect 14231 10081 14243 10084
rect 14185 10075 14243 10081
rect 14642 10072 14648 10084
rect 14700 10072 14706 10124
rect 16853 10115 16911 10121
rect 16853 10081 16865 10115
rect 16899 10112 16911 10115
rect 17218 10112 17224 10124
rect 16899 10084 17224 10112
rect 16899 10081 16911 10084
rect 16853 10075 16911 10081
rect 17218 10072 17224 10084
rect 17276 10072 17282 10124
rect 19518 10072 19524 10124
rect 19576 10112 19582 10124
rect 19705 10115 19763 10121
rect 19705 10112 19717 10115
rect 19576 10084 19717 10112
rect 19576 10072 19582 10084
rect 19705 10081 19717 10084
rect 19751 10081 19763 10115
rect 22462 10112 22468 10124
rect 22423 10084 22468 10112
rect 19705 10075 19763 10081
rect 22462 10072 22468 10084
rect 22520 10072 22526 10124
rect 22830 10072 22836 10124
rect 22888 10112 22894 10124
rect 22925 10115 22983 10121
rect 22925 10112 22937 10115
rect 22888 10084 22937 10112
rect 22888 10072 22894 10084
rect 22925 10081 22937 10084
rect 22971 10081 22983 10115
rect 24210 10112 24216 10124
rect 24171 10084 24216 10112
rect 22925 10075 22983 10081
rect 24210 10072 24216 10084
rect 24268 10072 24274 10124
rect 26234 10072 26240 10124
rect 26292 10112 26298 10124
rect 26605 10115 26663 10121
rect 26605 10112 26617 10115
rect 26292 10084 26617 10112
rect 26292 10072 26298 10084
rect 26605 10081 26617 10084
rect 26651 10081 26663 10115
rect 26605 10075 26663 10081
rect 28626 10072 28632 10124
rect 28684 10112 28690 10124
rect 29181 10115 29239 10121
rect 29181 10112 29193 10115
rect 28684 10084 29193 10112
rect 28684 10072 28690 10084
rect 29181 10081 29193 10084
rect 29227 10081 29239 10115
rect 29638 10112 29644 10124
rect 29599 10084 29644 10112
rect 29181 10075 29239 10081
rect 29638 10072 29644 10084
rect 29696 10072 29702 10124
rect 30812 10115 30870 10121
rect 30812 10112 30824 10115
rect 29748 10084 30824 10112
rect 14734 10044 14740 10056
rect 13504 10016 13584 10044
rect 13648 10016 14740 10044
rect 13504 10004 13510 10016
rect 12250 9976 12256 9988
rect 5644 9948 12256 9976
rect 12250 9936 12256 9948
rect 12308 9936 12314 9988
rect 4982 9868 4988 9920
rect 5040 9908 5046 9920
rect 5169 9911 5227 9917
rect 5169 9908 5181 9911
rect 5040 9880 5181 9908
rect 5040 9868 5046 9880
rect 5169 9877 5181 9880
rect 5215 9908 5227 9911
rect 5626 9908 5632 9920
rect 5215 9880 5632 9908
rect 5215 9877 5227 9880
rect 5169 9871 5227 9877
rect 5626 9868 5632 9880
rect 5684 9868 5690 9920
rect 13078 9868 13084 9920
rect 13136 9908 13142 9920
rect 13265 9911 13323 9917
rect 13265 9908 13277 9911
rect 13136 9880 13277 9908
rect 13136 9868 13142 9880
rect 13265 9877 13277 9880
rect 13311 9908 13323 9911
rect 13449 9911 13507 9917
rect 13449 9908 13461 9911
rect 13311 9880 13461 9908
rect 13311 9877 13323 9880
rect 13265 9871 13323 9877
rect 13449 9877 13461 9880
rect 13495 9877 13507 9911
rect 13556 9908 13584 10016
rect 14734 10004 14740 10016
rect 14792 10004 14798 10056
rect 14826 10004 14832 10056
rect 14884 10044 14890 10056
rect 15381 10047 15439 10053
rect 15381 10044 15393 10047
rect 14884 10016 15393 10044
rect 14884 10004 14890 10016
rect 15381 10013 15393 10016
rect 15427 10013 15439 10047
rect 16022 10044 16028 10056
rect 15983 10016 16028 10044
rect 15381 10007 15439 10013
rect 16022 10004 16028 10016
rect 16080 10004 16086 10056
rect 18138 10044 18144 10056
rect 18099 10016 18144 10044
rect 18138 10004 18144 10016
rect 18196 10004 18202 10056
rect 20806 10004 20812 10056
rect 20864 10044 20870 10056
rect 20993 10047 21051 10053
rect 20993 10044 21005 10047
rect 20864 10016 21005 10044
rect 20864 10004 20870 10016
rect 20993 10013 21005 10016
rect 21039 10044 21051 10047
rect 23198 10044 23204 10056
rect 21039 10016 23204 10044
rect 21039 10013 21051 10016
rect 20993 10007 21051 10013
rect 23198 10004 23204 10016
rect 23256 10004 23262 10056
rect 24394 10044 24400 10056
rect 24355 10016 24400 10044
rect 24394 10004 24400 10016
rect 24452 10004 24458 10056
rect 24486 10004 24492 10056
rect 24544 10044 24550 10056
rect 24673 10047 24731 10053
rect 24673 10044 24685 10047
rect 24544 10016 24685 10044
rect 24544 10004 24550 10016
rect 24673 10013 24685 10016
rect 24719 10013 24731 10047
rect 24673 10007 24731 10013
rect 28353 10047 28411 10053
rect 28353 10013 28365 10047
rect 28399 10044 28411 10047
rect 28994 10044 29000 10056
rect 28399 10016 29000 10044
rect 28399 10013 28411 10016
rect 28353 10007 28411 10013
rect 28994 10004 29000 10016
rect 29052 10004 29058 10056
rect 17770 9936 17776 9988
rect 17828 9976 17834 9988
rect 18693 9979 18751 9985
rect 18693 9976 18705 9979
rect 17828 9948 18705 9976
rect 17828 9936 17834 9948
rect 18693 9945 18705 9948
rect 18739 9976 18751 9979
rect 21542 9976 21548 9988
rect 18739 9948 21548 9976
rect 18739 9945 18751 9948
rect 18693 9939 18751 9945
rect 21542 9936 21548 9948
rect 21600 9936 21606 9988
rect 23474 9936 23480 9988
rect 23532 9976 23538 9988
rect 29748 9976 29776 10084
rect 30812 10081 30824 10084
rect 30858 10112 30870 10115
rect 31754 10112 31760 10124
rect 30858 10084 31760 10112
rect 30858 10081 30870 10084
rect 30812 10075 30870 10081
rect 31754 10072 31760 10084
rect 31812 10072 31818 10124
rect 35250 10112 35256 10124
rect 35211 10084 35256 10112
rect 35250 10072 35256 10084
rect 35308 10072 35314 10124
rect 29917 10047 29975 10053
rect 29917 10013 29929 10047
rect 29963 10044 29975 10047
rect 32030 10044 32036 10056
rect 29963 10016 32036 10044
rect 29963 10013 29975 10016
rect 29917 10007 29975 10013
rect 32030 10004 32036 10016
rect 32088 10004 32094 10056
rect 32490 10044 32496 10056
rect 32451 10016 32496 10044
rect 32490 10004 32496 10016
rect 32548 10044 32554 10056
rect 32548 10016 33134 10044
rect 32548 10004 32554 10016
rect 23532 9948 24072 9976
rect 23532 9936 23538 9948
rect 13998 9908 14004 9920
rect 13556 9880 14004 9908
rect 13449 9871 13507 9877
rect 13998 9868 14004 9880
rect 14056 9908 14062 9920
rect 14645 9911 14703 9917
rect 14645 9908 14657 9911
rect 14056 9880 14657 9908
rect 14056 9868 14062 9880
rect 14645 9877 14657 9880
rect 14691 9877 14703 9911
rect 19886 9908 19892 9920
rect 19847 9880 19892 9908
rect 14645 9871 14703 9877
rect 19886 9868 19892 9880
rect 19944 9868 19950 9920
rect 20162 9908 20168 9920
rect 20123 9880 20168 9908
rect 20162 9868 20168 9880
rect 20220 9868 20226 9920
rect 23382 9868 23388 9920
rect 23440 9908 23446 9920
rect 23753 9911 23811 9917
rect 23753 9908 23765 9911
rect 23440 9880 23765 9908
rect 23440 9868 23446 9880
rect 23753 9877 23765 9880
rect 23799 9908 23811 9911
rect 23934 9908 23940 9920
rect 23799 9880 23940 9908
rect 23799 9877 23811 9880
rect 23753 9871 23811 9877
rect 23934 9868 23940 9880
rect 23992 9868 23998 9920
rect 24044 9908 24072 9948
rect 25424 9948 29776 9976
rect 25424 9908 25452 9948
rect 30558 9936 30564 9988
rect 30616 9976 30622 9988
rect 30883 9979 30941 9985
rect 30883 9976 30895 9979
rect 30616 9948 30895 9976
rect 30616 9936 30622 9948
rect 30883 9945 30895 9948
rect 30929 9945 30941 9979
rect 33106 9976 33134 10016
rect 33502 10004 33508 10056
rect 33560 10044 33566 10056
rect 33781 10047 33839 10053
rect 33781 10044 33793 10047
rect 33560 10016 33793 10044
rect 33560 10004 33566 10016
rect 33781 10013 33793 10016
rect 33827 10013 33839 10047
rect 34057 10047 34115 10053
rect 34057 10044 34069 10047
rect 33781 10007 33839 10013
rect 33888 10016 34069 10044
rect 33229 9979 33287 9985
rect 33229 9976 33241 9979
rect 33106 9948 33241 9976
rect 30883 9939 30941 9945
rect 33229 9945 33241 9948
rect 33275 9976 33287 9979
rect 33888 9976 33916 10016
rect 34057 10013 34069 10016
rect 34103 10013 34115 10047
rect 34057 10007 34115 10013
rect 33275 9948 33916 9976
rect 33275 9945 33287 9948
rect 33229 9939 33287 9945
rect 24044 9880 25452 9908
rect 25685 9911 25743 9917
rect 25685 9877 25697 9911
rect 25731 9908 25743 9911
rect 26050 9908 26056 9920
rect 25731 9880 26056 9908
rect 25731 9877 25743 9880
rect 25685 9871 25743 9877
rect 26050 9868 26056 9880
rect 26108 9908 26114 9920
rect 26602 9908 26608 9920
rect 26108 9880 26608 9908
rect 26108 9868 26114 9880
rect 26602 9868 26608 9880
rect 26660 9868 26666 9920
rect 26786 9908 26792 9920
rect 26747 9880 26792 9908
rect 26786 9868 26792 9880
rect 26844 9868 26850 9920
rect 28534 9868 28540 9920
rect 28592 9908 28598 9920
rect 28629 9911 28687 9917
rect 28629 9908 28641 9911
rect 28592 9880 28641 9908
rect 28592 9868 28598 9880
rect 28629 9877 28641 9880
rect 28675 9877 28687 9911
rect 30650 9908 30656 9920
rect 30611 9880 30656 9908
rect 28629 9871 28687 9877
rect 30650 9868 30656 9880
rect 30708 9868 30714 9920
rect 34974 9868 34980 9920
rect 35032 9908 35038 9920
rect 35391 9911 35449 9917
rect 35391 9908 35403 9911
rect 35032 9880 35403 9908
rect 35032 9868 35038 9880
rect 35391 9877 35403 9880
rect 35437 9877 35449 9911
rect 35391 9871 35449 9877
rect 1104 9818 38824 9840
rect 1104 9766 7648 9818
rect 7700 9766 7712 9818
rect 7764 9766 7776 9818
rect 7828 9766 7840 9818
rect 7892 9766 20982 9818
rect 21034 9766 21046 9818
rect 21098 9766 21110 9818
rect 21162 9766 21174 9818
rect 21226 9766 34315 9818
rect 34367 9766 34379 9818
rect 34431 9766 34443 9818
rect 34495 9766 34507 9818
rect 34559 9766 38824 9818
rect 1104 9744 38824 9766
rect 106 9664 112 9716
rect 164 9704 170 9716
rect 5994 9704 6000 9716
rect 164 9676 6000 9704
rect 164 9664 170 9676
rect 5994 9664 6000 9676
rect 6052 9664 6058 9716
rect 6089 9707 6147 9713
rect 6089 9673 6101 9707
rect 6135 9704 6147 9707
rect 6270 9704 6276 9716
rect 6135 9676 6276 9704
rect 6135 9673 6147 9676
rect 6089 9667 6147 9673
rect 6270 9664 6276 9676
rect 6328 9664 6334 9716
rect 8202 9704 8208 9716
rect 8163 9676 8208 9704
rect 8202 9664 8208 9676
rect 8260 9704 8266 9716
rect 8573 9707 8631 9713
rect 8573 9704 8585 9707
rect 8260 9676 8585 9704
rect 8260 9664 8266 9676
rect 8573 9673 8585 9676
rect 8619 9673 8631 9707
rect 8573 9667 8631 9673
rect 9766 9664 9772 9716
rect 9824 9704 9830 9716
rect 10137 9707 10195 9713
rect 10137 9704 10149 9707
rect 9824 9676 10149 9704
rect 9824 9664 9830 9676
rect 10137 9673 10149 9676
rect 10183 9673 10195 9707
rect 10137 9667 10195 9673
rect 10226 9664 10232 9716
rect 10284 9704 10290 9716
rect 11241 9707 11299 9713
rect 11241 9704 11253 9707
rect 10284 9676 11253 9704
rect 10284 9664 10290 9676
rect 11241 9673 11253 9676
rect 11287 9704 11299 9707
rect 12342 9704 12348 9716
rect 11287 9676 12348 9704
rect 11287 9673 11299 9676
rect 11241 9667 11299 9673
rect 12342 9664 12348 9676
rect 12400 9664 12406 9716
rect 15378 9704 15384 9716
rect 15339 9676 15384 9704
rect 15378 9664 15384 9676
rect 15436 9664 15442 9716
rect 17218 9704 17224 9716
rect 17179 9676 17224 9704
rect 17218 9664 17224 9676
rect 17276 9664 17282 9716
rect 20717 9707 20775 9713
rect 20717 9673 20729 9707
rect 20763 9704 20775 9707
rect 21085 9707 21143 9713
rect 21085 9704 21097 9707
rect 20763 9676 21097 9704
rect 20763 9673 20775 9676
rect 20717 9667 20775 9673
rect 21085 9673 21097 9676
rect 21131 9704 21143 9707
rect 21266 9704 21272 9716
rect 21131 9676 21272 9704
rect 21131 9673 21143 9676
rect 21085 9667 21143 9673
rect 21266 9664 21272 9676
rect 21324 9664 21330 9716
rect 27706 9664 27712 9716
rect 27764 9704 27770 9716
rect 27893 9707 27951 9713
rect 27893 9704 27905 9707
rect 27764 9676 27905 9704
rect 27764 9664 27770 9676
rect 27893 9673 27905 9676
rect 27939 9673 27951 9707
rect 27893 9667 27951 9673
rect 30469 9707 30527 9713
rect 30469 9673 30481 9707
rect 30515 9704 30527 9707
rect 30742 9704 30748 9716
rect 30515 9676 30748 9704
rect 30515 9673 30527 9676
rect 30469 9667 30527 9673
rect 30742 9664 30748 9676
rect 30800 9704 30806 9716
rect 32217 9707 32275 9713
rect 32217 9704 32229 9707
rect 30800 9676 32229 9704
rect 30800 9664 30806 9676
rect 32217 9673 32229 9676
rect 32263 9704 32275 9707
rect 32306 9704 32312 9716
rect 32263 9676 32312 9704
rect 32263 9673 32275 9676
rect 32217 9667 32275 9673
rect 32306 9664 32312 9676
rect 32364 9664 32370 9716
rect 33781 9707 33839 9713
rect 33781 9704 33793 9707
rect 33106 9676 33793 9704
rect 7929 9639 7987 9645
rect 7929 9605 7941 9639
rect 7975 9636 7987 9639
rect 8386 9636 8392 9648
rect 7975 9608 8392 9636
rect 7975 9605 7987 9608
rect 7929 9599 7987 9605
rect 8386 9596 8392 9608
rect 8444 9636 8450 9648
rect 9858 9636 9864 9648
rect 8444 9608 9864 9636
rect 8444 9596 8450 9608
rect 9858 9596 9864 9608
rect 9916 9596 9922 9648
rect 12434 9596 12440 9648
rect 12492 9636 12498 9648
rect 12492 9608 12572 9636
rect 12492 9596 12498 9608
rect 2593 9571 2651 9577
rect 2593 9537 2605 9571
rect 2639 9568 2651 9571
rect 2774 9568 2780 9580
rect 2639 9540 2780 9568
rect 2639 9537 2651 9540
rect 2593 9531 2651 9537
rect 2774 9528 2780 9540
rect 2832 9528 2838 9580
rect 4706 9568 4712 9580
rect 4667 9540 4712 9568
rect 4706 9528 4712 9540
rect 4764 9528 4770 9580
rect 7009 9571 7067 9577
rect 7009 9537 7021 9571
rect 7055 9568 7067 9571
rect 7098 9568 7104 9580
rect 7055 9540 7104 9568
rect 7055 9537 7067 9540
rect 7009 9531 7067 9537
rect 7098 9528 7104 9540
rect 7156 9528 7162 9580
rect 8846 9568 8852 9580
rect 8759 9540 8852 9568
rect 8846 9528 8852 9540
rect 8904 9568 8910 9580
rect 12544 9577 12572 9608
rect 12710 9596 12716 9648
rect 12768 9636 12774 9648
rect 13725 9639 13783 9645
rect 13725 9636 13737 9639
rect 12768 9608 13737 9636
rect 12768 9596 12774 9608
rect 13725 9605 13737 9608
rect 13771 9636 13783 9639
rect 14090 9636 14096 9648
rect 13771 9608 14096 9636
rect 13771 9605 13783 9608
rect 13725 9599 13783 9605
rect 14090 9596 14096 9608
rect 14148 9596 14154 9648
rect 14369 9639 14427 9645
rect 14369 9605 14381 9639
rect 14415 9636 14427 9639
rect 14734 9636 14740 9648
rect 14415 9608 14740 9636
rect 14415 9605 14427 9608
rect 14369 9599 14427 9605
rect 14734 9596 14740 9608
rect 14792 9636 14798 9648
rect 15010 9636 15016 9648
rect 14792 9608 15016 9636
rect 14792 9596 14798 9608
rect 15010 9596 15016 9608
rect 15068 9636 15074 9648
rect 17862 9636 17868 9648
rect 15068 9608 17868 9636
rect 15068 9596 15074 9608
rect 17862 9596 17868 9608
rect 17920 9596 17926 9648
rect 20162 9596 20168 9648
rect 20220 9636 20226 9648
rect 21361 9639 21419 9645
rect 21361 9636 21373 9639
rect 20220 9608 21373 9636
rect 20220 9596 20226 9608
rect 21361 9605 21373 9608
rect 21407 9636 21419 9639
rect 21726 9636 21732 9648
rect 21407 9608 21732 9636
rect 21407 9605 21419 9608
rect 21361 9599 21419 9605
rect 21726 9596 21732 9608
rect 21784 9596 21790 9648
rect 23382 9596 23388 9648
rect 23440 9636 23446 9648
rect 24673 9639 24731 9645
rect 24673 9636 24685 9639
rect 23440 9608 24685 9636
rect 23440 9596 23446 9608
rect 24673 9605 24685 9608
rect 24719 9605 24731 9639
rect 24673 9599 24731 9605
rect 27154 9596 27160 9648
rect 27212 9636 27218 9648
rect 33106 9636 33134 9676
rect 33781 9673 33793 9676
rect 33827 9704 33839 9707
rect 33870 9704 33876 9716
rect 33827 9676 33876 9704
rect 33827 9673 33839 9676
rect 33781 9667 33839 9673
rect 33870 9664 33876 9676
rect 33928 9664 33934 9716
rect 35250 9704 35256 9716
rect 35211 9676 35256 9704
rect 35250 9664 35256 9676
rect 35308 9704 35314 9716
rect 35989 9707 36047 9713
rect 35989 9704 36001 9707
rect 35308 9676 36001 9704
rect 35308 9664 35314 9676
rect 35989 9673 36001 9676
rect 36035 9673 36047 9707
rect 35989 9667 36047 9673
rect 27212 9608 33134 9636
rect 27212 9596 27218 9608
rect 33502 9596 33508 9648
rect 33560 9636 33566 9648
rect 34057 9639 34115 9645
rect 34057 9636 34069 9639
rect 33560 9608 34069 9636
rect 33560 9596 33566 9608
rect 34057 9605 34069 9608
rect 34103 9605 34115 9639
rect 35618 9636 35624 9648
rect 35579 9608 35624 9636
rect 34057 9599 34115 9605
rect 35618 9596 35624 9608
rect 35676 9596 35682 9648
rect 10459 9571 10517 9577
rect 10459 9568 10471 9571
rect 8904 9540 10471 9568
rect 8904 9528 8910 9540
rect 10459 9537 10471 9540
rect 10505 9537 10517 9571
rect 10459 9531 10517 9537
rect 12529 9571 12587 9577
rect 12529 9537 12541 9571
rect 12575 9537 12587 9571
rect 12802 9568 12808 9580
rect 12763 9540 12808 9568
rect 12529 9531 12587 9537
rect 12802 9528 12808 9540
rect 12860 9568 12866 9580
rect 15378 9568 15384 9580
rect 12860 9540 15384 9568
rect 12860 9528 12866 9540
rect 15378 9528 15384 9540
rect 15436 9528 15442 9580
rect 17954 9528 17960 9580
rect 18012 9568 18018 9580
rect 18049 9571 18107 9577
rect 18049 9568 18061 9571
rect 18012 9540 18061 9568
rect 18012 9528 18018 9540
rect 18049 9537 18061 9540
rect 18095 9537 18107 9571
rect 18049 9531 18107 9537
rect 19242 9528 19248 9580
rect 19300 9568 19306 9580
rect 19797 9571 19855 9577
rect 19797 9568 19809 9571
rect 19300 9540 19809 9568
rect 19300 9528 19306 9540
rect 19797 9537 19809 9540
rect 19843 9568 19855 9571
rect 20254 9568 20260 9580
rect 19843 9540 20260 9568
rect 19843 9537 19855 9540
rect 19797 9531 19855 9537
rect 20254 9528 20260 9540
rect 20312 9528 20318 9580
rect 21634 9568 21640 9580
rect 21595 9540 21640 9568
rect 21634 9528 21640 9540
rect 21692 9528 21698 9580
rect 21910 9568 21916 9580
rect 21871 9540 21916 9568
rect 21910 9528 21916 9540
rect 21968 9528 21974 9580
rect 23753 9571 23811 9577
rect 23753 9537 23765 9571
rect 23799 9568 23811 9571
rect 24210 9568 24216 9580
rect 23799 9540 24216 9568
rect 23799 9537 23811 9540
rect 23753 9531 23811 9537
rect 24210 9528 24216 9540
rect 24268 9528 24274 9580
rect 24397 9571 24455 9577
rect 24397 9537 24409 9571
rect 24443 9568 24455 9571
rect 24486 9568 24492 9580
rect 24443 9540 24492 9568
rect 24443 9537 24455 9540
rect 24397 9531 24455 9537
rect 24486 9528 24492 9540
rect 24544 9528 24550 9580
rect 24578 9528 24584 9580
rect 24636 9568 24642 9580
rect 25593 9571 25651 9577
rect 25593 9568 25605 9571
rect 24636 9540 25605 9568
rect 24636 9528 24642 9540
rect 25593 9537 25605 9540
rect 25639 9537 25651 9571
rect 25593 9531 25651 9537
rect 26973 9571 27031 9577
rect 26973 9537 26985 9571
rect 27019 9568 27031 9571
rect 27062 9568 27068 9580
rect 27019 9540 27068 9568
rect 27019 9537 27031 9540
rect 26973 9531 27031 9537
rect 27062 9528 27068 9540
rect 27120 9528 27126 9580
rect 29687 9571 29745 9577
rect 29687 9537 29699 9571
rect 29733 9568 29745 9571
rect 30650 9568 30656 9580
rect 29733 9540 30656 9568
rect 29733 9537 29745 9540
rect 29687 9531 29745 9537
rect 30650 9528 30656 9540
rect 30708 9528 30714 9580
rect 30926 9568 30932 9580
rect 30887 9540 30932 9568
rect 30926 9528 30932 9540
rect 30984 9528 30990 9580
rect 32401 9571 32459 9577
rect 32401 9537 32413 9571
rect 32447 9568 32459 9571
rect 32490 9568 32496 9580
rect 32447 9540 32496 9568
rect 32447 9537 32459 9540
rect 32401 9531 32459 9537
rect 32490 9528 32496 9540
rect 32548 9528 32554 9580
rect 32674 9568 32680 9580
rect 32635 9540 32680 9568
rect 32674 9528 32680 9540
rect 32732 9528 32738 9580
rect 1394 9500 1400 9512
rect 1355 9472 1400 9500
rect 1394 9460 1400 9472
rect 1452 9500 1458 9512
rect 1946 9500 1952 9512
rect 1452 9472 1952 9500
rect 1452 9460 1458 9472
rect 1946 9460 1952 9472
rect 2004 9460 2010 9512
rect 3513 9503 3571 9509
rect 3513 9469 3525 9503
rect 3559 9500 3571 9503
rect 3970 9500 3976 9512
rect 3559 9472 3976 9500
rect 3559 9469 3571 9472
rect 3513 9463 3571 9469
rect 3970 9460 3976 9472
rect 4028 9460 4034 9512
rect 10372 9503 10430 9509
rect 10372 9469 10384 9503
rect 10418 9500 10430 9503
rect 11400 9503 11458 9509
rect 10418 9472 10916 9500
rect 10418 9469 10430 9472
rect 10372 9463 10430 9469
rect 2914 9435 2972 9441
rect 2914 9432 2926 9435
rect 2516 9404 2926 9432
rect 2516 9376 2544 9404
rect 2914 9401 2926 9404
rect 2960 9401 2972 9435
rect 2914 9395 2972 9401
rect 3234 9392 3240 9444
rect 3292 9432 3298 9444
rect 4157 9435 4215 9441
rect 4157 9432 4169 9435
rect 3292 9404 4169 9432
rect 3292 9392 3298 9404
rect 4157 9401 4169 9404
rect 4203 9401 4215 9435
rect 4430 9432 4436 9444
rect 4391 9404 4436 9432
rect 4157 9395 4215 9401
rect 106 9324 112 9376
rect 164 9364 170 9376
rect 1581 9367 1639 9373
rect 1581 9364 1593 9367
rect 164 9336 1593 9364
rect 164 9324 170 9336
rect 1581 9333 1593 9336
rect 1627 9333 1639 9367
rect 2498 9364 2504 9376
rect 2459 9336 2504 9364
rect 1581 9327 1639 9333
rect 2498 9324 2504 9336
rect 2556 9324 2562 9376
rect 3602 9324 3608 9376
rect 3660 9364 3666 9376
rect 3789 9367 3847 9373
rect 3789 9364 3801 9367
rect 3660 9336 3801 9364
rect 3660 9324 3666 9336
rect 3789 9333 3801 9336
rect 3835 9333 3847 9367
rect 4172 9364 4200 9395
rect 4430 9392 4436 9404
rect 4488 9392 4494 9444
rect 4525 9435 4583 9441
rect 4525 9401 4537 9435
rect 4571 9401 4583 9435
rect 7282 9432 7288 9444
rect 4525 9395 4583 9401
rect 6564 9404 7288 9432
rect 4540 9364 4568 9395
rect 4172 9336 4568 9364
rect 3789 9327 3847 9333
rect 5534 9324 5540 9376
rect 5592 9364 5598 9376
rect 5629 9367 5687 9373
rect 5629 9364 5641 9367
rect 5592 9336 5641 9364
rect 5592 9324 5598 9336
rect 5629 9333 5641 9336
rect 5675 9333 5687 9367
rect 5629 9327 5687 9333
rect 5810 9324 5816 9376
rect 5868 9364 5874 9376
rect 6564 9373 6592 9404
rect 7282 9392 7288 9404
rect 7340 9441 7346 9444
rect 7340 9435 7388 9441
rect 7340 9401 7342 9435
rect 7376 9401 7388 9435
rect 7340 9395 7388 9401
rect 7340 9392 7346 9395
rect 8202 9392 8208 9444
rect 8260 9432 8266 9444
rect 8941 9435 8999 9441
rect 8941 9432 8953 9435
rect 8260 9404 8953 9432
rect 8260 9392 8266 9404
rect 8941 9401 8953 9404
rect 8987 9401 8999 9435
rect 8941 9395 8999 9401
rect 9493 9435 9551 9441
rect 9493 9401 9505 9435
rect 9539 9432 9551 9435
rect 10042 9432 10048 9444
rect 9539 9404 10048 9432
rect 9539 9401 9551 9404
rect 9493 9395 9551 9401
rect 6549 9367 6607 9373
rect 6549 9364 6561 9367
rect 5868 9336 6561 9364
rect 5868 9324 5874 9336
rect 6549 9333 6561 9336
rect 6595 9333 6607 9367
rect 6549 9327 6607 9333
rect 7098 9324 7104 9376
rect 7156 9364 7162 9376
rect 8478 9364 8484 9376
rect 7156 9336 8484 9364
rect 7156 9324 7162 9336
rect 8478 9324 8484 9336
rect 8536 9364 8542 9376
rect 9508 9364 9536 9395
rect 10042 9392 10048 9404
rect 10100 9392 10106 9444
rect 10888 9376 10916 9472
rect 11400 9469 11412 9503
rect 11446 9500 11458 9503
rect 11790 9500 11796 9512
rect 11446 9472 11796 9500
rect 11446 9469 11458 9472
rect 11400 9463 11458 9469
rect 11790 9460 11796 9472
rect 11848 9460 11854 9512
rect 14461 9503 14519 9509
rect 14461 9469 14473 9503
rect 14507 9500 14519 9503
rect 14642 9500 14648 9512
rect 14507 9472 14648 9500
rect 14507 9469 14519 9472
rect 14461 9463 14519 9469
rect 14642 9460 14648 9472
rect 14700 9460 14706 9512
rect 15749 9503 15807 9509
rect 15749 9469 15761 9503
rect 15795 9500 15807 9503
rect 16482 9500 16488 9512
rect 15795 9472 16488 9500
rect 15795 9469 15807 9472
rect 15749 9463 15807 9469
rect 16482 9460 16488 9472
rect 16540 9460 16546 9512
rect 16669 9503 16727 9509
rect 16669 9469 16681 9503
rect 16715 9469 16727 9503
rect 16669 9463 16727 9469
rect 12621 9435 12679 9441
rect 12621 9401 12633 9435
rect 12667 9432 12679 9435
rect 12986 9432 12992 9444
rect 12667 9404 12992 9432
rect 12667 9401 12679 9404
rect 12621 9395 12679 9401
rect 12986 9392 12992 9404
rect 13044 9392 13050 9444
rect 14823 9435 14881 9441
rect 13280 9404 14733 9432
rect 10870 9364 10876 9376
rect 8536 9336 9536 9364
rect 10831 9336 10876 9364
rect 8536 9324 8542 9336
rect 10870 9324 10876 9336
rect 10928 9324 10934 9376
rect 11471 9367 11529 9373
rect 11471 9333 11483 9367
rect 11517 9364 11529 9367
rect 11698 9364 11704 9376
rect 11517 9336 11704 9364
rect 11517 9333 11529 9336
rect 11471 9327 11529 9333
rect 11698 9324 11704 9336
rect 11756 9324 11762 9376
rect 12253 9367 12311 9373
rect 12253 9333 12265 9367
rect 12299 9364 12311 9367
rect 12526 9364 12532 9376
rect 12299 9336 12532 9364
rect 12299 9333 12311 9336
rect 12253 9327 12311 9333
rect 12526 9324 12532 9336
rect 12584 9364 12590 9376
rect 13280 9364 13308 9404
rect 12584 9336 13308 9364
rect 14705 9364 14733 9404
rect 14823 9401 14835 9435
rect 14869 9432 14881 9435
rect 15010 9432 15016 9444
rect 14869 9404 15016 9432
rect 14869 9401 14881 9404
rect 14823 9395 14881 9401
rect 15010 9392 15016 9404
rect 15068 9392 15074 9444
rect 16025 9435 16083 9441
rect 16025 9432 16037 9435
rect 15580 9404 16037 9432
rect 15580 9376 15608 9404
rect 16025 9401 16037 9404
rect 16071 9432 16083 9435
rect 16684 9432 16712 9463
rect 18230 9460 18236 9512
rect 18288 9500 18294 9512
rect 18969 9503 19027 9509
rect 18969 9500 18981 9503
rect 18288 9472 18981 9500
rect 18288 9460 18294 9472
rect 18969 9469 18981 9472
rect 19015 9469 19027 9503
rect 18969 9463 19027 9469
rect 28077 9503 28135 9509
rect 28077 9469 28089 9503
rect 28123 9500 28135 9503
rect 28626 9500 28632 9512
rect 28123 9472 28632 9500
rect 28123 9469 28135 9472
rect 28077 9463 28135 9469
rect 28626 9460 28632 9472
rect 28684 9460 28690 9512
rect 28718 9460 28724 9512
rect 28776 9500 28782 9512
rect 29600 9503 29658 9509
rect 29600 9500 29612 9503
rect 28776 9472 29612 9500
rect 28776 9460 28782 9472
rect 29600 9469 29612 9472
rect 29646 9500 29658 9503
rect 29646 9472 30144 9500
rect 29646 9469 29658 9472
rect 29600 9463 29658 9469
rect 16942 9432 16948 9444
rect 16071 9404 16712 9432
rect 16903 9404 16948 9432
rect 16071 9401 16083 9404
rect 16025 9395 16083 9401
rect 16942 9392 16948 9404
rect 17000 9392 17006 9444
rect 17862 9432 17868 9444
rect 17775 9404 17868 9432
rect 17862 9392 17868 9404
rect 17920 9432 17926 9444
rect 18411 9435 18469 9441
rect 18411 9432 18423 9435
rect 17920 9404 18423 9432
rect 17920 9392 17926 9404
rect 18411 9401 18423 9404
rect 18457 9432 18469 9435
rect 19705 9435 19763 9441
rect 19705 9432 19717 9435
rect 18457 9404 19717 9432
rect 18457 9401 18469 9404
rect 18411 9395 18469 9401
rect 19705 9401 19717 9404
rect 19751 9432 19763 9435
rect 20070 9432 20076 9444
rect 19751 9404 20076 9432
rect 19751 9401 19763 9404
rect 19705 9395 19763 9401
rect 20070 9392 20076 9404
rect 20128 9441 20134 9444
rect 20128 9435 20176 9441
rect 20128 9401 20130 9435
rect 20164 9401 20176 9435
rect 20128 9395 20176 9401
rect 20128 9392 20134 9395
rect 21726 9392 21732 9444
rect 21784 9432 21790 9444
rect 23845 9435 23903 9441
rect 21784 9404 21829 9432
rect 21784 9392 21790 9404
rect 23845 9401 23857 9435
rect 23891 9401 23903 9435
rect 23845 9395 23903 9401
rect 15562 9364 15568 9376
rect 14705 9336 15568 9364
rect 12584 9324 12590 9336
rect 15562 9324 15568 9336
rect 15620 9324 15626 9376
rect 18782 9324 18788 9376
rect 18840 9364 18846 9376
rect 19245 9367 19303 9373
rect 19245 9364 19257 9367
rect 18840 9336 19257 9364
rect 18840 9324 18846 9336
rect 19245 9333 19257 9336
rect 19291 9364 19303 9367
rect 19518 9364 19524 9376
rect 19291 9336 19524 9364
rect 19291 9333 19303 9336
rect 19245 9327 19303 9333
rect 19518 9324 19524 9336
rect 19576 9324 19582 9376
rect 19978 9324 19984 9376
rect 20036 9364 20042 9376
rect 22462 9364 22468 9376
rect 20036 9336 22468 9364
rect 20036 9324 20042 9336
rect 22462 9324 22468 9336
rect 22520 9364 22526 9376
rect 22557 9367 22615 9373
rect 22557 9364 22569 9367
rect 22520 9336 22569 9364
rect 22520 9324 22526 9336
rect 22557 9333 22569 9336
rect 22603 9333 22615 9367
rect 22557 9327 22615 9333
rect 22830 9324 22836 9376
rect 22888 9364 22894 9376
rect 23017 9367 23075 9373
rect 23017 9364 23029 9367
rect 22888 9336 23029 9364
rect 22888 9324 22894 9336
rect 23017 9333 23029 9336
rect 23063 9364 23075 9367
rect 23198 9364 23204 9376
rect 23063 9336 23204 9364
rect 23063 9333 23075 9336
rect 23017 9327 23075 9333
rect 23198 9324 23204 9336
rect 23256 9324 23262 9376
rect 23477 9367 23535 9373
rect 23477 9333 23489 9367
rect 23523 9364 23535 9367
rect 23658 9364 23664 9376
rect 23523 9336 23664 9364
rect 23523 9333 23535 9336
rect 23477 9327 23535 9333
rect 23658 9324 23664 9336
rect 23716 9364 23722 9376
rect 23860 9364 23888 9395
rect 24118 9392 24124 9444
rect 24176 9432 24182 9444
rect 25314 9432 25320 9444
rect 24176 9404 25320 9432
rect 24176 9392 24182 9404
rect 25314 9392 25320 9404
rect 25372 9392 25378 9444
rect 25409 9435 25467 9441
rect 25409 9401 25421 9435
rect 25455 9401 25467 9435
rect 25409 9395 25467 9401
rect 25041 9367 25099 9373
rect 25041 9364 25053 9367
rect 23716 9336 25053 9364
rect 23716 9324 23722 9336
rect 25041 9333 25053 9336
rect 25087 9364 25099 9367
rect 25424 9364 25452 9395
rect 25682 9392 25688 9444
rect 25740 9432 25746 9444
rect 26329 9435 26387 9441
rect 26329 9432 26341 9435
rect 25740 9404 26341 9432
rect 25740 9392 25746 9404
rect 26329 9401 26341 9404
rect 26375 9432 26387 9435
rect 27065 9435 27123 9441
rect 27065 9432 27077 9435
rect 26375 9404 27077 9432
rect 26375 9401 26387 9404
rect 26329 9395 26387 9401
rect 27065 9401 27077 9404
rect 27111 9432 27123 9435
rect 27154 9432 27160 9444
rect 27111 9404 27160 9432
rect 27111 9401 27123 9404
rect 27065 9395 27123 9401
rect 27154 9392 27160 9404
rect 27212 9392 27218 9444
rect 27617 9435 27675 9441
rect 27617 9401 27629 9435
rect 27663 9432 27675 9435
rect 28350 9432 28356 9444
rect 27663 9404 28356 9432
rect 27663 9401 27675 9404
rect 27617 9395 27675 9401
rect 28350 9392 28356 9404
rect 28408 9392 28414 9444
rect 30116 9376 30144 9472
rect 35250 9460 35256 9512
rect 35308 9500 35314 9512
rect 35437 9503 35495 9509
rect 35437 9500 35449 9503
rect 35308 9472 35449 9500
rect 35308 9460 35314 9472
rect 35437 9469 35449 9472
rect 35483 9469 35495 9503
rect 35437 9463 35495 9469
rect 30742 9432 30748 9444
rect 30703 9404 30748 9432
rect 30742 9392 30748 9404
rect 30800 9392 30806 9444
rect 32493 9435 32551 9441
rect 32493 9401 32505 9435
rect 32539 9432 32551 9435
rect 32539 9404 32628 9432
rect 32539 9401 32551 9404
rect 32493 9395 32551 9401
rect 25087 9336 25452 9364
rect 25087 9333 25099 9336
rect 25041 9327 25099 9333
rect 26234 9324 26240 9376
rect 26292 9364 26298 9376
rect 26605 9367 26663 9373
rect 26605 9364 26617 9367
rect 26292 9336 26617 9364
rect 26292 9324 26298 9336
rect 26605 9333 26617 9336
rect 26651 9364 26663 9367
rect 28077 9367 28135 9373
rect 28077 9364 28089 9367
rect 26651 9336 28089 9364
rect 26651 9333 26663 9336
rect 26605 9327 26663 9333
rect 28077 9333 28089 9336
rect 28123 9333 28135 9367
rect 28258 9364 28264 9376
rect 28219 9336 28264 9364
rect 28077 9327 28135 9333
rect 28258 9324 28264 9336
rect 28316 9324 28322 9376
rect 28718 9324 28724 9376
rect 28776 9364 28782 9376
rect 28997 9367 29055 9373
rect 28997 9364 29009 9367
rect 28776 9336 29009 9364
rect 28776 9324 28782 9336
rect 28997 9333 29009 9336
rect 29043 9364 29055 9367
rect 29638 9364 29644 9376
rect 29043 9336 29644 9364
rect 29043 9333 29055 9336
rect 28997 9327 29055 9333
rect 29638 9324 29644 9336
rect 29696 9324 29702 9376
rect 30098 9364 30104 9376
rect 30059 9336 30104 9364
rect 30098 9324 30104 9336
rect 30156 9324 30162 9376
rect 31665 9367 31723 9373
rect 31665 9333 31677 9367
rect 31711 9364 31723 9367
rect 31754 9364 31760 9376
rect 31711 9336 31760 9364
rect 31711 9333 31723 9336
rect 31665 9327 31723 9333
rect 31754 9324 31760 9336
rect 31812 9324 31818 9376
rect 32600 9364 32628 9404
rect 33134 9364 33140 9376
rect 32600 9336 33140 9364
rect 33134 9324 33140 9336
rect 33192 9364 33198 9376
rect 33321 9367 33379 9373
rect 33321 9364 33333 9367
rect 33192 9336 33333 9364
rect 33192 9324 33198 9336
rect 33321 9333 33333 9336
rect 33367 9333 33379 9367
rect 33321 9327 33379 9333
rect 1104 9274 38824 9296
rect 1104 9222 14315 9274
rect 14367 9222 14379 9274
rect 14431 9222 14443 9274
rect 14495 9222 14507 9274
rect 14559 9222 27648 9274
rect 27700 9222 27712 9274
rect 27764 9222 27776 9274
rect 27828 9222 27840 9274
rect 27892 9222 38824 9274
rect 1104 9200 38824 9222
rect 2038 9160 2044 9172
rect 1999 9132 2044 9160
rect 2038 9120 2044 9132
rect 2096 9120 2102 9172
rect 2498 9120 2504 9172
rect 2556 9160 2562 9172
rect 2593 9163 2651 9169
rect 2593 9160 2605 9163
rect 2556 9132 2605 9160
rect 2556 9120 2562 9132
rect 2593 9129 2605 9132
rect 2639 9129 2651 9163
rect 2593 9123 2651 9129
rect 3145 9163 3203 9169
rect 3145 9129 3157 9163
rect 3191 9160 3203 9163
rect 3234 9160 3240 9172
rect 3191 9132 3240 9160
rect 3191 9129 3203 9132
rect 3145 9123 3203 9129
rect 3234 9120 3240 9132
rect 3292 9120 3298 9172
rect 3881 9163 3939 9169
rect 3881 9129 3893 9163
rect 3927 9160 3939 9163
rect 4154 9160 4160 9172
rect 3927 9132 4160 9160
rect 3927 9129 3939 9132
rect 3881 9123 3939 9129
rect 4154 9120 4160 9132
rect 4212 9120 4218 9172
rect 4430 9120 4436 9172
rect 4488 9160 4494 9172
rect 4985 9163 5043 9169
rect 4985 9160 4997 9163
rect 4488 9132 4997 9160
rect 4488 9120 4494 9132
rect 4985 9129 4997 9132
rect 5031 9160 5043 9163
rect 6086 9160 6092 9172
rect 5031 9132 5993 9160
rect 6047 9132 6092 9160
rect 5031 9129 5043 9132
rect 4985 9123 5043 9129
rect 2774 9052 2780 9104
rect 2832 9092 2838 9104
rect 3421 9095 3479 9101
rect 3421 9092 3433 9095
rect 2832 9064 3433 9092
rect 2832 9052 2838 9064
rect 3421 9061 3433 9064
rect 3467 9061 3479 9095
rect 3421 9055 3479 9061
rect 3970 9052 3976 9104
rect 4028 9092 4034 9104
rect 4617 9095 4675 9101
rect 4617 9092 4629 9095
rect 4028 9064 4629 9092
rect 4028 9052 4034 9064
rect 4617 9061 4629 9064
rect 4663 9061 4675 9095
rect 4617 9055 4675 9061
rect 5531 9095 5589 9101
rect 5531 9061 5543 9095
rect 5577 9092 5589 9095
rect 5810 9092 5816 9104
rect 5577 9064 5816 9092
rect 5577 9061 5589 9064
rect 5531 9055 5589 9061
rect 5810 9052 5816 9064
rect 5868 9052 5874 9104
rect 5965 9092 5993 9132
rect 6086 9120 6092 9132
rect 6144 9120 6150 9172
rect 6822 9160 6828 9172
rect 6783 9132 6828 9160
rect 6822 9120 6828 9132
rect 6880 9120 6886 9172
rect 7282 9160 7288 9172
rect 7243 9132 7288 9160
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 7837 9163 7895 9169
rect 7837 9129 7849 9163
rect 7883 9160 7895 9163
rect 8202 9160 8208 9172
rect 7883 9132 8208 9160
rect 7883 9129 7895 9132
rect 7837 9123 7895 9129
rect 8202 9120 8208 9132
rect 8260 9120 8266 9172
rect 8846 9160 8852 9172
rect 8807 9132 8852 9160
rect 8846 9120 8852 9132
rect 8904 9120 8910 9172
rect 13814 9120 13820 9172
rect 13872 9160 13878 9172
rect 13872 9132 13917 9160
rect 13872 9120 13878 9132
rect 14826 9120 14832 9172
rect 14884 9160 14890 9172
rect 15013 9163 15071 9169
rect 15013 9160 15025 9163
rect 14884 9132 15025 9160
rect 14884 9120 14890 9132
rect 15013 9129 15025 9132
rect 15059 9129 15071 9163
rect 16945 9163 17003 9169
rect 16945 9160 16957 9163
rect 15013 9123 15071 9129
rect 15304 9132 16957 9160
rect 7098 9092 7104 9104
rect 5965 9064 7104 9092
rect 7098 9052 7104 9064
rect 7156 9052 7162 9104
rect 9858 9092 9864 9104
rect 9819 9064 9864 9092
rect 9858 9052 9864 9064
rect 9916 9052 9922 9104
rect 11698 9052 11704 9104
rect 11756 9092 11762 9104
rect 11977 9095 12035 9101
rect 11977 9092 11989 9095
rect 11756 9064 11989 9092
rect 11756 9052 11762 9064
rect 11977 9061 11989 9064
rect 12023 9061 12035 9095
rect 11977 9055 12035 9061
rect 12069 9095 12127 9101
rect 12069 9061 12081 9095
rect 12115 9092 12127 9095
rect 12986 9092 12992 9104
rect 12115 9064 12992 9092
rect 12115 9061 12127 9064
rect 12069 9055 12127 9061
rect 12986 9052 12992 9064
rect 13044 9052 13050 9104
rect 14642 9052 14648 9104
rect 14700 9092 14706 9104
rect 14737 9095 14795 9101
rect 14737 9092 14749 9095
rect 14700 9064 14749 9092
rect 14700 9052 14706 9064
rect 14737 9061 14749 9064
rect 14783 9092 14795 9095
rect 15304 9092 15332 9132
rect 16945 9129 16957 9132
rect 16991 9129 17003 9163
rect 18138 9160 18144 9172
rect 18099 9132 18144 9160
rect 16945 9123 17003 9129
rect 18138 9120 18144 9132
rect 18196 9120 18202 9172
rect 18230 9120 18236 9172
rect 18288 9160 18294 9172
rect 18417 9163 18475 9169
rect 18417 9160 18429 9163
rect 18288 9132 18429 9160
rect 18288 9120 18294 9132
rect 18417 9129 18429 9132
rect 18463 9129 18475 9163
rect 20070 9160 20076 9172
rect 18417 9123 18475 9129
rect 19438 9132 20076 9160
rect 15470 9092 15476 9104
rect 14783 9064 15332 9092
rect 15431 9064 15476 9092
rect 14783 9061 14795 9064
rect 14737 9055 14795 9061
rect 15470 9052 15476 9064
rect 15528 9052 15534 9104
rect 16390 9092 16396 9104
rect 16351 9064 16396 9092
rect 16390 9052 16396 9064
rect 16448 9052 16454 9104
rect 19438 9101 19466 9132
rect 20070 9120 20076 9132
rect 20128 9120 20134 9172
rect 20254 9160 20260 9172
rect 20215 9132 20260 9160
rect 20254 9120 20260 9132
rect 20312 9120 20318 9172
rect 20717 9163 20775 9169
rect 20717 9129 20729 9163
rect 20763 9160 20775 9163
rect 20806 9160 20812 9172
rect 20763 9132 20812 9160
rect 20763 9129 20775 9132
rect 20717 9123 20775 9129
rect 20806 9120 20812 9132
rect 20864 9120 20870 9172
rect 21634 9120 21640 9172
rect 21692 9160 21698 9172
rect 21913 9163 21971 9169
rect 21913 9160 21925 9163
rect 21692 9132 21925 9160
rect 21692 9120 21698 9132
rect 21913 9129 21925 9132
rect 21959 9129 21971 9163
rect 23474 9160 23480 9172
rect 23435 9132 23480 9160
rect 21913 9123 21971 9129
rect 23474 9120 23480 9132
rect 23532 9120 23538 9172
rect 24394 9160 24400 9172
rect 24355 9132 24400 9160
rect 24394 9120 24400 9132
rect 24452 9120 24458 9172
rect 24949 9163 25007 9169
rect 24949 9160 24961 9163
rect 24780 9132 24961 9160
rect 19423 9095 19481 9101
rect 19423 9061 19435 9095
rect 19469 9061 19481 9095
rect 21085 9095 21143 9101
rect 21085 9092 21097 9095
rect 19423 9055 19481 9061
rect 19996 9064 21097 9092
rect 2222 9024 2228 9036
rect 2183 8996 2228 9024
rect 2222 8984 2228 8996
rect 2280 8984 2286 9036
rect 4062 9024 4068 9036
rect 4023 8996 4068 9024
rect 4062 8984 4068 8996
rect 4120 9024 4126 9036
rect 5166 9024 5172 9036
rect 4120 8984 4154 9024
rect 5079 8996 5172 9024
rect 5166 8984 5172 8996
rect 5224 9024 5230 9036
rect 5718 9024 5724 9036
rect 5224 8996 5724 9024
rect 5224 8984 5230 8996
rect 5718 8984 5724 8996
rect 5776 8984 5782 9036
rect 8110 9024 8116 9036
rect 5828 8996 8116 9024
rect 4126 8956 4154 8984
rect 5828 8956 5856 8996
rect 8110 8984 8116 8996
rect 8168 8984 8174 9036
rect 13449 9027 13507 9033
rect 13449 8993 13461 9027
rect 13495 9024 13507 9027
rect 13722 9024 13728 9036
rect 13495 8996 13728 9024
rect 13495 8993 13507 8996
rect 13449 8987 13507 8993
rect 13722 8984 13728 8996
rect 13780 8984 13786 9036
rect 16850 9024 16856 9036
rect 16811 8996 16856 9024
rect 16850 8984 16856 8996
rect 16908 8984 16914 9036
rect 17405 9027 17463 9033
rect 17405 8993 17417 9027
rect 17451 9024 17463 9027
rect 17494 9024 17500 9036
rect 17451 8996 17500 9024
rect 17451 8993 17463 8996
rect 17405 8987 17463 8993
rect 17494 8984 17500 8996
rect 17552 8984 17558 9036
rect 19058 9024 19064 9036
rect 19019 8996 19064 9024
rect 19058 8984 19064 8996
rect 19116 8984 19122 9036
rect 19996 9033 20024 9064
rect 21085 9061 21097 9064
rect 21131 9092 21143 9095
rect 22094 9092 22100 9104
rect 21131 9064 22100 9092
rect 21131 9061 21143 9064
rect 21085 9055 21143 9061
rect 22094 9052 22100 9064
rect 22152 9052 22158 9104
rect 19981 9027 20039 9033
rect 19981 8993 19993 9027
rect 20027 8993 20039 9027
rect 24780 9024 24808 9132
rect 24949 9129 24961 9132
rect 24995 9129 25007 9163
rect 24949 9123 25007 9129
rect 25314 9120 25320 9172
rect 25372 9160 25378 9172
rect 25869 9163 25927 9169
rect 25869 9160 25881 9163
rect 25372 9132 25881 9160
rect 25372 9120 25378 9132
rect 25869 9129 25881 9132
rect 25915 9129 25927 9163
rect 25869 9123 25927 9129
rect 27433 9163 27491 9169
rect 27433 9129 27445 9163
rect 27479 9160 27491 9163
rect 28258 9160 28264 9172
rect 27479 9132 28264 9160
rect 27479 9129 27491 9132
rect 27433 9123 27491 9129
rect 28258 9120 28264 9132
rect 28316 9120 28322 9172
rect 28902 9120 28908 9172
rect 28960 9160 28966 9172
rect 29546 9160 29552 9172
rect 28960 9132 29552 9160
rect 28960 9120 28966 9132
rect 29546 9120 29552 9132
rect 29604 9120 29610 9172
rect 31570 9120 31576 9172
rect 31628 9160 31634 9172
rect 31849 9163 31907 9169
rect 31849 9160 31861 9163
rect 31628 9132 31861 9160
rect 31628 9120 31634 9132
rect 31849 9129 31861 9132
rect 31895 9129 31907 9163
rect 32490 9160 32496 9172
rect 32451 9132 32496 9160
rect 31849 9123 31907 9129
rect 32490 9120 32496 9132
rect 32548 9120 32554 9172
rect 33045 9163 33103 9169
rect 33045 9129 33057 9163
rect 33091 9160 33103 9163
rect 33134 9160 33140 9172
rect 33091 9132 33140 9160
rect 33091 9129 33103 9132
rect 33045 9123 33103 9129
rect 33134 9120 33140 9132
rect 33192 9120 33198 9172
rect 25498 9092 25504 9104
rect 25148 9064 25504 9092
rect 25148 9033 25176 9064
rect 25498 9052 25504 9064
rect 25556 9052 25562 9104
rect 26875 9095 26933 9101
rect 26875 9061 26887 9095
rect 26921 9092 26933 9095
rect 26970 9092 26976 9104
rect 26921 9064 26976 9092
rect 26921 9061 26933 9064
rect 26875 9055 26933 9061
rect 26970 9052 26976 9064
rect 27028 9052 27034 9104
rect 28442 9092 28448 9104
rect 28403 9064 28448 9092
rect 28442 9052 28448 9064
rect 28500 9052 28506 9104
rect 28994 9092 29000 9104
rect 28955 9064 29000 9092
rect 28994 9052 29000 9064
rect 29052 9052 29058 9104
rect 30558 9092 30564 9104
rect 30519 9064 30564 9092
rect 30558 9052 30564 9064
rect 30616 9052 30622 9104
rect 30653 9095 30711 9101
rect 30653 9061 30665 9095
rect 30699 9092 30711 9095
rect 30834 9092 30840 9104
rect 30699 9064 30840 9092
rect 30699 9061 30711 9064
rect 30653 9055 30711 9061
rect 30834 9052 30840 9064
rect 30892 9092 30898 9104
rect 31478 9092 31484 9104
rect 30892 9064 31484 9092
rect 30892 9052 30898 9064
rect 31478 9052 31484 9064
rect 31536 9052 31542 9104
rect 34517 9095 34575 9101
rect 34517 9061 34529 9095
rect 34563 9092 34575 9095
rect 34606 9092 34612 9104
rect 34563 9064 34612 9092
rect 34563 9061 34575 9064
rect 34517 9055 34575 9061
rect 34606 9052 34612 9064
rect 34664 9052 34670 9104
rect 19981 8987 20039 8993
rect 23124 8996 24808 9024
rect 25133 9027 25191 9033
rect 23124 8968 23152 8996
rect 25133 8993 25145 9027
rect 25179 8993 25191 9027
rect 25133 8987 25191 8993
rect 25317 9027 25375 9033
rect 25317 8993 25329 9027
rect 25363 8993 25375 9027
rect 25317 8987 25375 8993
rect 6914 8956 6920 8968
rect 4126 8928 5856 8956
rect 6875 8928 6920 8956
rect 6914 8916 6920 8928
rect 6972 8916 6978 8968
rect 9769 8959 9827 8965
rect 9769 8925 9781 8959
rect 9815 8956 9827 8959
rect 11054 8956 11060 8968
rect 9815 8928 11060 8956
rect 9815 8925 9827 8928
rect 9769 8919 9827 8925
rect 11054 8916 11060 8928
rect 11112 8916 11118 8968
rect 11146 8916 11152 8968
rect 11204 8956 11210 8968
rect 12621 8959 12679 8965
rect 12621 8956 12633 8959
rect 11204 8928 12633 8956
rect 11204 8916 11210 8928
rect 12621 8925 12633 8928
rect 12667 8956 12679 8959
rect 15102 8956 15108 8968
rect 12667 8928 15108 8956
rect 12667 8925 12679 8928
rect 12621 8919 12679 8925
rect 15102 8916 15108 8928
rect 15160 8956 15166 8968
rect 15381 8959 15439 8965
rect 15381 8956 15393 8959
rect 15160 8928 15393 8956
rect 15160 8916 15166 8928
rect 15381 8925 15393 8928
rect 15427 8925 15439 8959
rect 16022 8956 16028 8968
rect 15983 8928 16028 8956
rect 15381 8919 15439 8925
rect 16022 8916 16028 8928
rect 16080 8916 16086 8968
rect 20714 8916 20720 8968
rect 20772 8956 20778 8968
rect 20993 8959 21051 8965
rect 20993 8956 21005 8959
rect 20772 8928 21005 8956
rect 20772 8916 20778 8928
rect 20993 8925 21005 8928
rect 21039 8956 21051 8959
rect 21910 8956 21916 8968
rect 21039 8928 21916 8956
rect 21039 8925 21051 8928
rect 20993 8919 21051 8925
rect 21910 8916 21916 8928
rect 21968 8916 21974 8968
rect 23106 8956 23112 8968
rect 23067 8928 23112 8956
rect 23106 8916 23112 8928
rect 23164 8916 23170 8968
rect 23198 8916 23204 8968
rect 23256 8956 23262 8968
rect 24673 8959 24731 8965
rect 24673 8956 24685 8959
rect 23256 8928 24685 8956
rect 23256 8916 23262 8928
rect 24673 8925 24685 8928
rect 24719 8956 24731 8959
rect 25332 8956 25360 8987
rect 32030 8984 32036 9036
rect 32088 9024 32094 9036
rect 32125 9027 32183 9033
rect 32125 9024 32137 9027
rect 32088 8996 32137 9024
rect 32088 8984 32094 8996
rect 32125 8993 32137 8996
rect 32171 9024 32183 9027
rect 33226 9024 33232 9036
rect 32171 8996 33232 9024
rect 32171 8993 32183 8996
rect 32125 8987 32183 8993
rect 33226 8984 33232 8996
rect 33284 8984 33290 9036
rect 35894 9024 35900 9036
rect 35855 8996 35900 9024
rect 35894 8984 35900 8996
rect 35952 8984 35958 9036
rect 26510 8956 26516 8968
rect 24719 8928 25360 8956
rect 26471 8928 26516 8956
rect 24719 8925 24731 8928
rect 24673 8919 24731 8925
rect 26510 8916 26516 8928
rect 26568 8916 26574 8968
rect 28350 8956 28356 8968
rect 28311 8928 28356 8956
rect 28350 8916 28356 8928
rect 28408 8956 28414 8968
rect 30837 8959 30895 8965
rect 30837 8956 30849 8959
rect 28408 8928 30849 8956
rect 28408 8916 28414 8928
rect 30837 8925 30849 8928
rect 30883 8956 30895 8959
rect 30926 8956 30932 8968
rect 30883 8928 30932 8956
rect 30883 8925 30895 8928
rect 30837 8919 30895 8925
rect 30926 8916 30932 8928
rect 30984 8916 30990 8968
rect 34425 8959 34483 8965
rect 34425 8925 34437 8959
rect 34471 8956 34483 8959
rect 34698 8956 34704 8968
rect 34471 8928 34704 8956
rect 34471 8925 34483 8928
rect 34425 8919 34483 8925
rect 34698 8916 34704 8928
rect 34756 8916 34762 8968
rect 35069 8959 35127 8965
rect 35069 8925 35081 8959
rect 35115 8956 35127 8959
rect 36262 8956 36268 8968
rect 35115 8928 36268 8956
rect 35115 8925 35127 8928
rect 35069 8919 35127 8925
rect 36262 8916 36268 8928
rect 36320 8916 36326 8968
rect 14 8848 20 8900
rect 72 8888 78 8900
rect 4249 8891 4307 8897
rect 4249 8888 4261 8891
rect 72 8860 4261 8888
rect 72 8848 78 8860
rect 4249 8857 4261 8860
rect 4295 8857 4307 8891
rect 4249 8851 4307 8857
rect 8754 8848 8760 8900
rect 8812 8888 8818 8900
rect 10321 8891 10379 8897
rect 10321 8888 10333 8891
rect 8812 8860 10333 8888
rect 8812 8848 8818 8860
rect 10321 8857 10333 8860
rect 10367 8888 10379 8891
rect 12802 8888 12808 8900
rect 10367 8860 12808 8888
rect 10367 8857 10379 8860
rect 10321 8851 10379 8857
rect 12802 8848 12808 8860
rect 12860 8848 12866 8900
rect 14369 8891 14427 8897
rect 14369 8857 14381 8891
rect 14415 8888 14427 8891
rect 15010 8888 15016 8900
rect 14415 8860 15016 8888
rect 14415 8857 14427 8860
rect 14369 8851 14427 8857
rect 15010 8848 15016 8860
rect 15068 8848 15074 8900
rect 21542 8888 21548 8900
rect 21503 8860 21548 8888
rect 21542 8848 21548 8860
rect 21600 8848 21606 8900
rect 23382 8848 23388 8900
rect 23440 8888 23446 8900
rect 24029 8891 24087 8897
rect 24029 8888 24041 8891
rect 23440 8860 24041 8888
rect 23440 8848 23446 8860
rect 24029 8857 24041 8860
rect 24075 8857 24087 8891
rect 24029 8851 24087 8857
rect 30098 8848 30104 8900
rect 30156 8888 30162 8900
rect 36630 8888 36636 8900
rect 30156 8860 36636 8888
rect 30156 8848 30162 8860
rect 36630 8848 36636 8860
rect 36688 8848 36694 8900
rect 8294 8820 8300 8832
rect 8255 8792 8300 8820
rect 8294 8780 8300 8792
rect 8352 8780 8358 8832
rect 12986 8820 12992 8832
rect 12947 8792 12992 8820
rect 12986 8780 12992 8792
rect 13044 8780 13050 8832
rect 18966 8820 18972 8832
rect 18927 8792 18972 8820
rect 18966 8780 18972 8792
rect 19024 8780 19030 8832
rect 21266 8780 21272 8832
rect 21324 8820 21330 8832
rect 24670 8820 24676 8832
rect 21324 8792 24676 8820
rect 21324 8780 21330 8792
rect 24670 8780 24676 8792
rect 24728 8780 24734 8832
rect 36081 8823 36139 8829
rect 36081 8789 36093 8823
rect 36127 8820 36139 8823
rect 39574 8820 39580 8832
rect 36127 8792 39580 8820
rect 36127 8789 36139 8792
rect 36081 8783 36139 8789
rect 39574 8780 39580 8792
rect 39632 8780 39638 8832
rect 1104 8730 38824 8752
rect 1104 8678 7648 8730
rect 7700 8678 7712 8730
rect 7764 8678 7776 8730
rect 7828 8678 7840 8730
rect 7892 8678 20982 8730
rect 21034 8678 21046 8730
rect 21098 8678 21110 8730
rect 21162 8678 21174 8730
rect 21226 8678 34315 8730
rect 34367 8678 34379 8730
rect 34431 8678 34443 8730
rect 34495 8678 34507 8730
rect 34559 8678 38824 8730
rect 1104 8656 38824 8678
rect 2222 8576 2228 8628
rect 2280 8616 2286 8628
rect 3142 8616 3148 8628
rect 2280 8588 2957 8616
rect 3103 8588 3148 8616
rect 2280 8576 2286 8588
rect 1854 8508 1860 8560
rect 1912 8548 1918 8560
rect 2929 8548 2957 8588
rect 3142 8576 3148 8588
rect 3200 8576 3206 8628
rect 3881 8619 3939 8625
rect 3881 8585 3893 8619
rect 3927 8616 3939 8619
rect 4062 8616 4068 8628
rect 3927 8588 4068 8616
rect 3927 8585 3939 8588
rect 3881 8579 3939 8585
rect 4062 8576 4068 8588
rect 4120 8576 4126 8628
rect 6822 8576 6828 8628
rect 6880 8616 6886 8628
rect 7331 8619 7389 8625
rect 7331 8616 7343 8619
rect 6880 8588 7343 8616
rect 6880 8576 6886 8588
rect 7331 8585 7343 8588
rect 7377 8585 7389 8619
rect 7331 8579 7389 8585
rect 7745 8619 7803 8625
rect 7745 8585 7757 8619
rect 7791 8616 7803 8619
rect 8202 8616 8208 8628
rect 7791 8588 8208 8616
rect 7791 8585 7803 8588
rect 7745 8579 7803 8585
rect 3421 8551 3479 8557
rect 3421 8548 3433 8551
rect 1912 8520 2360 8548
rect 2929 8520 3433 8548
rect 1912 8508 1918 8520
rect 2130 8440 2136 8492
rect 2188 8480 2194 8492
rect 2225 8483 2283 8489
rect 2225 8480 2237 8483
rect 2188 8452 2237 8480
rect 2188 8440 2194 8452
rect 2225 8449 2237 8452
rect 2271 8449 2283 8483
rect 2332 8480 2360 8520
rect 3421 8517 3433 8520
rect 3467 8517 3479 8551
rect 7190 8548 7196 8560
rect 3421 8511 3479 8517
rect 3528 8520 7196 8548
rect 3528 8480 3556 8520
rect 7190 8508 7196 8520
rect 7248 8508 7254 8560
rect 2332 8452 3556 8480
rect 2225 8443 2283 8449
rect 3786 8440 3792 8492
rect 3844 8480 3850 8492
rect 4341 8483 4399 8489
rect 4341 8480 4353 8483
rect 3844 8452 4353 8480
rect 3844 8440 3850 8452
rect 4341 8449 4353 8452
rect 4387 8449 4399 8483
rect 4341 8443 4399 8449
rect 5604 8415 5662 8421
rect 5604 8381 5616 8415
rect 5650 8412 5662 8415
rect 5994 8412 6000 8424
rect 5650 8384 6000 8412
rect 5650 8381 5662 8384
rect 5604 8375 5662 8381
rect 5994 8372 6000 8384
rect 6052 8372 6058 8424
rect 6362 8372 6368 8424
rect 6420 8412 6426 8424
rect 7260 8415 7318 8421
rect 7260 8412 7272 8415
rect 6420 8384 7272 8412
rect 6420 8372 6426 8384
rect 7260 8381 7272 8384
rect 7306 8412 7318 8415
rect 7760 8412 7788 8579
rect 8202 8576 8208 8588
rect 8260 8576 8266 8628
rect 9125 8619 9183 8625
rect 9125 8585 9137 8619
rect 9171 8616 9183 8619
rect 9493 8619 9551 8625
rect 9493 8616 9505 8619
rect 9171 8588 9505 8616
rect 9171 8585 9183 8588
rect 9125 8579 9183 8585
rect 9493 8585 9505 8588
rect 9539 8616 9551 8619
rect 9858 8616 9864 8628
rect 9539 8588 9864 8616
rect 9539 8585 9551 8588
rect 9493 8579 9551 8585
rect 9858 8576 9864 8588
rect 9916 8576 9922 8628
rect 11054 8616 11060 8628
rect 11015 8588 11060 8616
rect 11054 8576 11060 8588
rect 11112 8576 11118 8628
rect 11517 8619 11575 8625
rect 11517 8585 11529 8619
rect 11563 8616 11575 8619
rect 11698 8616 11704 8628
rect 11563 8588 11704 8616
rect 11563 8585 11575 8588
rect 11517 8579 11575 8585
rect 11698 8576 11704 8588
rect 11756 8576 11762 8628
rect 11885 8619 11943 8625
rect 11885 8585 11897 8619
rect 11931 8616 11943 8619
rect 12986 8616 12992 8628
rect 11931 8588 12992 8616
rect 11931 8585 11943 8588
rect 11885 8579 11943 8585
rect 12986 8576 12992 8588
rect 13044 8616 13050 8628
rect 13357 8619 13415 8625
rect 13357 8616 13369 8619
rect 13044 8588 13369 8616
rect 13044 8576 13050 8588
rect 13357 8585 13369 8588
rect 13403 8585 13415 8619
rect 13357 8579 13415 8585
rect 15289 8619 15347 8625
rect 15289 8585 15301 8619
rect 15335 8616 15347 8619
rect 15470 8616 15476 8628
rect 15335 8588 15476 8616
rect 15335 8585 15347 8588
rect 15289 8579 15347 8585
rect 15470 8576 15476 8588
rect 15528 8616 15534 8628
rect 15565 8619 15623 8625
rect 15565 8616 15577 8619
rect 15528 8588 15577 8616
rect 15528 8576 15534 8588
rect 15565 8585 15577 8588
rect 15611 8585 15623 8619
rect 17494 8616 17500 8628
rect 17455 8588 17500 8616
rect 15565 8579 15623 8585
rect 17494 8576 17500 8588
rect 17552 8576 17558 8628
rect 18601 8619 18659 8625
rect 18601 8585 18613 8619
rect 18647 8616 18659 8619
rect 18877 8619 18935 8625
rect 18877 8616 18889 8619
rect 18647 8588 18889 8616
rect 18647 8585 18659 8588
rect 18601 8579 18659 8585
rect 18877 8585 18889 8588
rect 18923 8616 18935 8619
rect 19150 8616 19156 8628
rect 18923 8588 19156 8616
rect 18923 8585 18935 8588
rect 18877 8579 18935 8585
rect 19150 8576 19156 8588
rect 19208 8576 19214 8628
rect 20162 8576 20168 8628
rect 20220 8616 20226 8628
rect 20257 8619 20315 8625
rect 20257 8616 20269 8619
rect 20220 8588 20269 8616
rect 20220 8576 20226 8588
rect 20257 8585 20269 8588
rect 20303 8585 20315 8619
rect 22094 8616 22100 8628
rect 22055 8588 22100 8616
rect 20257 8579 20315 8585
rect 22094 8576 22100 8588
rect 22152 8576 22158 8628
rect 22833 8619 22891 8625
rect 22833 8585 22845 8619
rect 22879 8616 22891 8619
rect 23106 8616 23112 8628
rect 22879 8588 23112 8616
rect 22879 8585 22891 8588
rect 22833 8579 22891 8585
rect 23106 8576 23112 8588
rect 23164 8576 23170 8628
rect 25682 8616 25688 8628
rect 25643 8588 25688 8616
rect 25682 8576 25688 8588
rect 25740 8576 25746 8628
rect 27433 8619 27491 8625
rect 27433 8585 27445 8619
rect 27479 8616 27491 8619
rect 28353 8619 28411 8625
rect 28353 8616 28365 8619
rect 27479 8588 28365 8616
rect 27479 8585 27491 8588
rect 27433 8579 27491 8585
rect 28353 8585 28365 8588
rect 28399 8616 28411 8619
rect 28442 8616 28448 8628
rect 28399 8588 28448 8616
rect 28399 8585 28411 8588
rect 28353 8579 28411 8585
rect 28442 8576 28448 8588
rect 28500 8576 28506 8628
rect 30558 8576 30564 8628
rect 30616 8616 30622 8628
rect 31113 8619 31171 8625
rect 31113 8616 31125 8619
rect 30616 8588 31125 8616
rect 30616 8576 30622 8588
rect 31113 8585 31125 8588
rect 31159 8585 31171 8619
rect 33226 8616 33232 8628
rect 33187 8588 33232 8616
rect 31113 8579 31171 8585
rect 33226 8576 33232 8588
rect 33284 8576 33290 8628
rect 34698 8576 34704 8628
rect 34756 8616 34762 8628
rect 37599 8619 37657 8625
rect 37599 8616 37611 8619
rect 34756 8588 37611 8616
rect 34756 8576 34762 8588
rect 37599 8585 37611 8588
rect 37645 8585 37657 8619
rect 37599 8579 37657 8585
rect 10410 8508 10416 8560
rect 10468 8548 10474 8560
rect 10597 8551 10655 8557
rect 10597 8548 10609 8551
rect 10468 8520 10609 8548
rect 10468 8508 10474 8520
rect 10597 8517 10609 8520
rect 10643 8548 10655 8551
rect 11146 8548 11152 8560
rect 10643 8520 11152 8548
rect 10643 8517 10655 8520
rect 10597 8511 10655 8517
rect 11146 8508 11152 8520
rect 11204 8508 11210 8560
rect 16390 8508 16396 8560
rect 16448 8548 16454 8560
rect 16448 8520 16528 8548
rect 16448 8508 16454 8520
rect 8205 8483 8263 8489
rect 8205 8449 8217 8483
rect 8251 8480 8263 8483
rect 8294 8480 8300 8492
rect 8251 8452 8300 8480
rect 8251 8449 8263 8452
rect 8205 8443 8263 8449
rect 8294 8440 8300 8452
rect 8352 8480 8358 8492
rect 10686 8480 10692 8492
rect 8352 8452 10692 8480
rect 8352 8440 8358 8452
rect 10686 8440 10692 8452
rect 10744 8440 10750 8492
rect 13630 8440 13636 8492
rect 13688 8480 13694 8492
rect 14369 8483 14427 8489
rect 14369 8480 14381 8483
rect 13688 8452 14381 8480
rect 13688 8440 13694 8452
rect 14369 8449 14381 8452
rect 14415 8480 14427 8483
rect 14642 8480 14648 8492
rect 14415 8452 14648 8480
rect 14415 8449 14427 8452
rect 14369 8443 14427 8449
rect 14642 8440 14648 8452
rect 14700 8440 14706 8492
rect 16500 8489 16528 8520
rect 19886 8508 19892 8560
rect 19944 8548 19950 8560
rect 20533 8551 20591 8557
rect 20533 8548 20545 8551
rect 19944 8520 20545 8548
rect 19944 8508 19950 8520
rect 20533 8517 20545 8520
rect 20579 8517 20591 8551
rect 30834 8548 30840 8560
rect 30795 8520 30840 8548
rect 20533 8511 20591 8517
rect 16485 8483 16543 8489
rect 16485 8449 16497 8483
rect 16531 8449 16543 8483
rect 17126 8480 17132 8492
rect 17039 8452 17132 8480
rect 16485 8443 16543 8449
rect 17126 8440 17132 8452
rect 17184 8480 17190 8492
rect 18874 8480 18880 8492
rect 17184 8452 18880 8480
rect 17184 8440 17190 8452
rect 18874 8440 18880 8452
rect 18932 8440 18938 8492
rect 18966 8440 18972 8492
rect 19024 8480 19030 8492
rect 19337 8483 19395 8489
rect 19337 8480 19349 8483
rect 19024 8452 19349 8480
rect 19024 8440 19030 8452
rect 19337 8449 19349 8452
rect 19383 8449 19395 8483
rect 20548 8480 20576 8511
rect 30834 8508 30840 8520
rect 30892 8508 30898 8560
rect 35894 8548 35900 8560
rect 35855 8520 35900 8548
rect 35894 8508 35900 8520
rect 35952 8508 35958 8560
rect 21358 8480 21364 8492
rect 20548 8452 21364 8480
rect 19337 8443 19395 8449
rect 21358 8440 21364 8452
rect 21416 8480 21422 8492
rect 21416 8452 21588 8480
rect 21416 8440 21422 8452
rect 7306 8384 7788 8412
rect 12437 8415 12495 8421
rect 7306 8381 7318 8384
rect 7260 8375 7318 8381
rect 12437 8381 12449 8415
rect 12483 8412 12495 8415
rect 12618 8412 12624 8424
rect 12483 8384 12624 8412
rect 12483 8381 12495 8384
rect 12437 8375 12495 8381
rect 12618 8372 12624 8384
rect 12676 8372 12682 8424
rect 18376 8415 18434 8421
rect 18376 8381 18388 8415
rect 18422 8412 18434 8415
rect 18601 8415 18659 8421
rect 18601 8412 18613 8415
rect 18422 8384 18613 8412
rect 18422 8381 18434 8384
rect 18376 8375 18434 8381
rect 18601 8381 18613 8384
rect 18647 8381 18659 8415
rect 18601 8375 18659 8381
rect 18690 8372 18696 8424
rect 18748 8412 18754 8424
rect 20901 8415 20959 8421
rect 20901 8412 20913 8415
rect 18748 8384 20913 8412
rect 18748 8372 18754 8384
rect 20901 8381 20913 8384
rect 20947 8412 20959 8415
rect 21085 8415 21143 8421
rect 21085 8412 21097 8415
rect 20947 8384 21097 8412
rect 20947 8381 20959 8384
rect 20901 8375 20959 8381
rect 21085 8381 21097 8384
rect 21131 8412 21143 8415
rect 21266 8412 21272 8424
rect 21131 8384 21272 8412
rect 21131 8381 21143 8384
rect 21085 8375 21143 8381
rect 21266 8372 21272 8384
rect 21324 8372 21330 8424
rect 21560 8421 21588 8452
rect 26326 8440 26332 8492
rect 26384 8480 26390 8492
rect 26513 8483 26571 8489
rect 26513 8480 26525 8483
rect 26384 8452 26525 8480
rect 26384 8440 26390 8452
rect 26513 8449 26525 8452
rect 26559 8480 26571 8483
rect 27709 8483 27767 8489
rect 27709 8480 27721 8483
rect 26559 8452 27721 8480
rect 26559 8449 26571 8452
rect 26513 8443 26571 8449
rect 27709 8449 27721 8452
rect 27755 8449 27767 8483
rect 27709 8443 27767 8449
rect 28350 8440 28356 8492
rect 28408 8480 28414 8492
rect 28629 8483 28687 8489
rect 28629 8480 28641 8483
rect 28408 8452 28641 8480
rect 28408 8440 28414 8452
rect 28629 8449 28641 8452
rect 28675 8449 28687 8483
rect 29546 8480 29552 8492
rect 29507 8452 29552 8480
rect 28629 8443 28687 8449
rect 29546 8440 29552 8452
rect 29604 8440 29610 8492
rect 30006 8440 30012 8492
rect 30064 8480 30070 8492
rect 31662 8480 31668 8492
rect 30064 8452 31668 8480
rect 30064 8440 30070 8452
rect 31662 8440 31668 8452
rect 31720 8440 31726 8492
rect 34606 8480 34612 8492
rect 33612 8452 34612 8480
rect 21545 8415 21603 8421
rect 21545 8381 21557 8415
rect 21591 8381 21603 8415
rect 23750 8412 23756 8424
rect 23714 8384 23756 8412
rect 21545 8375 21603 8381
rect 23750 8372 23756 8384
rect 23808 8421 23814 8424
rect 23808 8415 23862 8421
rect 23808 8381 23816 8415
rect 23850 8412 23862 8415
rect 24305 8415 24363 8421
rect 24305 8412 24317 8415
rect 23850 8384 24317 8412
rect 23850 8381 23862 8384
rect 23808 8375 23862 8381
rect 24305 8381 24317 8384
rect 24351 8412 24363 8415
rect 24578 8412 24584 8424
rect 24351 8384 24584 8412
rect 24351 8381 24363 8384
rect 24305 8375 24363 8381
rect 23808 8372 23814 8375
rect 24578 8372 24584 8384
rect 24636 8372 24642 8424
rect 24765 8415 24823 8421
rect 24765 8381 24777 8415
rect 24811 8412 24823 8415
rect 24854 8412 24860 8424
rect 24811 8384 24860 8412
rect 24811 8381 24823 8384
rect 24765 8375 24823 8381
rect 24854 8372 24860 8384
rect 24912 8372 24918 8424
rect 30469 8415 30527 8421
rect 30469 8381 30481 8415
rect 30515 8412 30527 8415
rect 30742 8412 30748 8424
rect 30515 8384 30748 8412
rect 30515 8381 30527 8384
rect 30469 8375 30527 8381
rect 30742 8372 30748 8384
rect 30800 8372 30806 8424
rect 33612 8421 33640 8452
rect 34606 8440 34612 8452
rect 34664 8440 34670 8492
rect 34974 8480 34980 8492
rect 34935 8452 34980 8480
rect 34974 8440 34980 8452
rect 35032 8440 35038 8492
rect 35250 8480 35256 8492
rect 35211 8452 35256 8480
rect 35250 8440 35256 8452
rect 35308 8440 35314 8492
rect 35434 8440 35440 8492
rect 35492 8480 35498 8492
rect 36909 8483 36967 8489
rect 36909 8480 36921 8483
rect 35492 8452 36921 8480
rect 35492 8440 35498 8452
rect 32585 8415 32643 8421
rect 32585 8381 32597 8415
rect 32631 8412 32643 8415
rect 33597 8415 33655 8421
rect 33597 8412 33609 8415
rect 32631 8384 33609 8412
rect 32631 8381 32643 8384
rect 32585 8375 32643 8381
rect 33597 8381 33609 8384
rect 33643 8381 33655 8415
rect 33597 8375 33655 8381
rect 33848 8415 33906 8421
rect 33848 8381 33860 8415
rect 33894 8412 33906 8415
rect 34146 8412 34152 8424
rect 33894 8384 34152 8412
rect 33894 8381 33906 8384
rect 33848 8375 33906 8381
rect 34146 8372 34152 8384
rect 34204 8412 34210 8424
rect 34241 8415 34299 8421
rect 34241 8412 34253 8415
rect 34204 8384 34253 8412
rect 34204 8372 34210 8384
rect 34241 8381 34253 8384
rect 34287 8381 34299 8415
rect 34241 8375 34299 8381
rect 3878 8304 3884 8356
rect 3936 8344 3942 8356
rect 4065 8347 4123 8353
rect 4065 8344 4077 8347
rect 3936 8316 4077 8344
rect 3936 8304 3942 8316
rect 4065 8313 4077 8316
rect 4111 8313 4123 8347
rect 4065 8307 4123 8313
rect 4157 8347 4215 8353
rect 4157 8313 4169 8347
rect 4203 8344 4215 8347
rect 4522 8344 4528 8356
rect 4203 8316 4528 8344
rect 4203 8313 4215 8316
rect 4157 8307 4215 8313
rect 4522 8304 4528 8316
rect 4580 8304 4586 8356
rect 5169 8347 5227 8353
rect 5169 8313 5181 8347
rect 5215 8344 5227 8347
rect 5810 8344 5816 8356
rect 5215 8316 5816 8344
rect 5215 8313 5227 8316
rect 5169 8307 5227 8313
rect 5810 8304 5816 8316
rect 5868 8344 5874 8356
rect 7009 8347 7067 8353
rect 7009 8344 7021 8347
rect 5868 8316 7021 8344
rect 5868 8304 5874 8316
rect 7009 8313 7021 8316
rect 7055 8344 7067 8347
rect 8021 8347 8079 8353
rect 8021 8344 8033 8347
rect 7055 8316 8033 8344
rect 7055 8313 7067 8316
rect 7009 8307 7067 8313
rect 8021 8313 8033 8316
rect 8067 8344 8079 8347
rect 8526 8347 8584 8353
rect 8526 8344 8538 8347
rect 8067 8316 8538 8344
rect 8067 8313 8079 8316
rect 8021 8307 8079 8313
rect 8526 8313 8538 8316
rect 8572 8344 8584 8347
rect 8662 8344 8668 8356
rect 8572 8316 8668 8344
rect 8572 8313 8584 8316
rect 8526 8307 8584 8313
rect 8662 8304 8668 8316
rect 8720 8304 8726 8356
rect 10042 8344 10048 8356
rect 10003 8316 10048 8344
rect 10042 8304 10048 8316
rect 10100 8304 10106 8356
rect 10137 8347 10195 8353
rect 10137 8313 10149 8347
rect 10183 8313 10195 8347
rect 10137 8307 10195 8313
rect 12253 8347 12311 8353
rect 12253 8313 12265 8347
rect 12299 8344 12311 8347
rect 12758 8347 12816 8353
rect 12758 8344 12770 8347
rect 12299 8316 12770 8344
rect 12299 8313 12311 8316
rect 12253 8307 12311 8313
rect 12758 8313 12770 8316
rect 12804 8344 12816 8347
rect 13633 8347 13691 8353
rect 13633 8344 13645 8347
rect 12804 8316 13645 8344
rect 12804 8313 12816 8316
rect 12758 8307 12816 8313
rect 13633 8313 13645 8316
rect 13679 8344 13691 8347
rect 13679 8316 13814 8344
rect 13679 8313 13691 8316
rect 13633 8307 13691 8313
rect 1765 8279 1823 8285
rect 1765 8245 1777 8279
rect 1811 8276 1823 8279
rect 2133 8279 2191 8285
rect 2133 8276 2145 8279
rect 1811 8248 2145 8276
rect 1811 8245 1823 8248
rect 1765 8239 1823 8245
rect 2133 8245 2145 8248
rect 2179 8276 2191 8279
rect 2498 8276 2504 8288
rect 2179 8248 2504 8276
rect 2179 8245 2191 8248
rect 2133 8239 2191 8245
rect 2498 8236 2504 8248
rect 2556 8276 2562 8288
rect 2593 8279 2651 8285
rect 2593 8276 2605 8279
rect 2556 8248 2605 8276
rect 2556 8236 2562 8248
rect 2593 8245 2605 8248
rect 2639 8276 2651 8279
rect 3326 8276 3332 8288
rect 2639 8248 3332 8276
rect 2639 8245 2651 8248
rect 2593 8239 2651 8245
rect 3326 8236 3332 8248
rect 3384 8236 3390 8288
rect 5258 8236 5264 8288
rect 5316 8276 5322 8288
rect 5675 8279 5733 8285
rect 5675 8276 5687 8279
rect 5316 8248 5687 8276
rect 5316 8236 5322 8248
rect 5675 8245 5687 8248
rect 5721 8245 5733 8279
rect 5675 8239 5733 8245
rect 6641 8279 6699 8285
rect 6641 8245 6653 8279
rect 6687 8276 6699 8279
rect 6914 8276 6920 8288
rect 6687 8248 6920 8276
rect 6687 8245 6699 8248
rect 6641 8239 6699 8245
rect 6914 8236 6920 8248
rect 6972 8236 6978 8288
rect 9858 8236 9864 8288
rect 9916 8276 9922 8288
rect 10152 8276 10180 8307
rect 9916 8248 10180 8276
rect 13786 8276 13814 8316
rect 16574 8304 16580 8356
rect 16632 8344 16638 8356
rect 18463 8347 18521 8353
rect 16632 8316 16677 8344
rect 16632 8304 16638 8316
rect 18463 8313 18475 8347
rect 18509 8344 18521 8347
rect 19518 8344 19524 8356
rect 18509 8316 19524 8344
rect 18509 8313 18521 8316
rect 18463 8307 18521 8313
rect 19518 8304 19524 8316
rect 19576 8304 19582 8356
rect 19699 8347 19757 8353
rect 19699 8313 19711 8347
rect 19745 8344 19757 8347
rect 20070 8344 20076 8356
rect 19745 8316 20076 8344
rect 19745 8313 19757 8316
rect 19699 8307 19757 8313
rect 13906 8276 13912 8288
rect 13786 8248 13912 8276
rect 9916 8236 9922 8248
rect 13906 8236 13912 8248
rect 13964 8276 13970 8288
rect 14277 8279 14335 8285
rect 14277 8276 14289 8279
rect 13964 8248 14289 8276
rect 13964 8236 13970 8248
rect 14277 8245 14289 8248
rect 14323 8276 14335 8279
rect 14734 8276 14740 8288
rect 14323 8248 14740 8276
rect 14323 8245 14335 8248
rect 14277 8239 14335 8245
rect 14734 8236 14740 8248
rect 14792 8236 14798 8288
rect 15930 8236 15936 8288
rect 15988 8276 15994 8288
rect 16209 8279 16267 8285
rect 16209 8276 16221 8279
rect 15988 8248 16221 8276
rect 15988 8236 15994 8248
rect 16209 8245 16221 8248
rect 16255 8276 16267 8279
rect 16850 8276 16856 8288
rect 16255 8248 16856 8276
rect 16255 8245 16267 8248
rect 16209 8239 16267 8245
rect 16850 8236 16856 8248
rect 16908 8236 16914 8288
rect 19245 8279 19303 8285
rect 19245 8245 19257 8279
rect 19291 8276 19303 8279
rect 19714 8276 19742 8307
rect 20070 8304 20076 8316
rect 20128 8304 20134 8356
rect 21818 8344 21824 8356
rect 21779 8316 21824 8344
rect 21818 8304 21824 8316
rect 21876 8304 21882 8356
rect 23891 8347 23949 8353
rect 23891 8313 23903 8347
rect 23937 8344 23949 8347
rect 24946 8344 24952 8356
rect 23937 8316 24952 8344
rect 23937 8313 23949 8316
rect 23891 8307 23949 8313
rect 24946 8304 24952 8316
rect 25004 8304 25010 8356
rect 25127 8347 25185 8353
rect 25127 8344 25139 8347
rect 25102 8313 25139 8344
rect 25173 8344 25185 8347
rect 26053 8347 26111 8353
rect 26053 8344 26065 8347
rect 25173 8316 26065 8344
rect 25173 8313 25185 8316
rect 25102 8307 25185 8313
rect 26053 8313 26065 8316
rect 26099 8344 26111 8347
rect 26421 8347 26479 8353
rect 26421 8344 26433 8347
rect 26099 8316 26433 8344
rect 26099 8313 26111 8316
rect 26053 8307 26111 8313
rect 26421 8313 26433 8316
rect 26467 8344 26479 8347
rect 26875 8347 26933 8353
rect 26875 8344 26887 8347
rect 26467 8316 26887 8344
rect 26467 8313 26479 8316
rect 26421 8307 26479 8313
rect 26875 8313 26887 8316
rect 26921 8344 26933 8347
rect 26970 8344 26976 8356
rect 26921 8316 26976 8344
rect 26921 8313 26933 8316
rect 26875 8307 26933 8313
rect 19291 8248 19742 8276
rect 23201 8279 23259 8285
rect 19291 8245 19303 8248
rect 19245 8239 19303 8245
rect 23201 8245 23213 8279
rect 23247 8276 23259 8279
rect 23474 8276 23480 8288
rect 23247 8248 23480 8276
rect 23247 8245 23259 8248
rect 23201 8239 23259 8245
rect 23474 8236 23480 8248
rect 23532 8276 23538 8288
rect 24673 8279 24731 8285
rect 24673 8276 24685 8279
rect 23532 8248 24685 8276
rect 23532 8236 23538 8248
rect 24673 8245 24685 8248
rect 24719 8276 24731 8279
rect 25102 8276 25130 8307
rect 26970 8304 26976 8316
rect 27028 8304 27034 8356
rect 32027 8347 32085 8353
rect 32027 8313 32039 8347
rect 32073 8313 32085 8347
rect 34624 8344 34652 8440
rect 36499 8421 36527 8452
rect 36909 8449 36921 8452
rect 36955 8449 36967 8483
rect 36909 8443 36967 8449
rect 36484 8415 36542 8421
rect 36484 8381 36496 8415
rect 36530 8381 36542 8415
rect 36484 8375 36542 8381
rect 36630 8372 36636 8424
rect 36688 8412 36694 8424
rect 37528 8415 37586 8421
rect 37528 8412 37540 8415
rect 36688 8384 37540 8412
rect 36688 8372 36694 8384
rect 37528 8381 37540 8384
rect 37574 8412 37586 8415
rect 37574 8384 38056 8412
rect 37574 8381 37586 8384
rect 37528 8375 37586 8381
rect 35069 8347 35127 8353
rect 35069 8344 35081 8347
rect 34624 8316 35081 8344
rect 32027 8307 32085 8313
rect 35069 8313 35081 8316
rect 35115 8313 35127 8347
rect 35069 8307 35127 8313
rect 29914 8276 29920 8288
rect 24719 8248 25130 8276
rect 29875 8248 29920 8276
rect 24719 8245 24731 8248
rect 24673 8239 24731 8245
rect 29914 8236 29920 8248
rect 29972 8236 29978 8288
rect 31573 8279 31631 8285
rect 31573 8245 31585 8279
rect 31619 8276 31631 8279
rect 32048 8276 32076 8307
rect 32490 8276 32496 8288
rect 31619 8248 32496 8276
rect 31619 8245 31631 8248
rect 31573 8239 31631 8245
rect 32490 8236 32496 8248
rect 32548 8276 32554 8288
rect 32861 8279 32919 8285
rect 32861 8276 32873 8279
rect 32548 8248 32873 8276
rect 32548 8236 32554 8248
rect 32861 8245 32873 8248
rect 32907 8245 32919 8279
rect 32861 8239 32919 8245
rect 33919 8279 33977 8285
rect 33919 8245 33931 8279
rect 33965 8276 33977 8279
rect 34146 8276 34152 8288
rect 33965 8248 34152 8276
rect 33965 8245 33977 8248
rect 33919 8239 33977 8245
rect 34146 8236 34152 8248
rect 34204 8236 34210 8288
rect 35986 8236 35992 8288
rect 36044 8276 36050 8288
rect 38028 8285 38056 8384
rect 36587 8279 36645 8285
rect 36587 8276 36599 8279
rect 36044 8248 36599 8276
rect 36044 8236 36050 8248
rect 36587 8245 36599 8248
rect 36633 8245 36645 8279
rect 36587 8239 36645 8245
rect 38013 8279 38071 8285
rect 38013 8245 38025 8279
rect 38059 8276 38071 8279
rect 38102 8276 38108 8288
rect 38059 8248 38108 8276
rect 38059 8245 38071 8248
rect 38013 8239 38071 8245
rect 38102 8236 38108 8248
rect 38160 8236 38166 8288
rect 1104 8186 38824 8208
rect 1104 8134 14315 8186
rect 14367 8134 14379 8186
rect 14431 8134 14443 8186
rect 14495 8134 14507 8186
rect 14559 8134 27648 8186
rect 27700 8134 27712 8186
rect 27764 8134 27776 8186
rect 27828 8134 27840 8186
rect 27892 8134 38824 8186
rect 1104 8112 38824 8134
rect 2130 8072 2136 8084
rect 2091 8044 2136 8072
rect 2130 8032 2136 8044
rect 2188 8032 2194 8084
rect 3878 8072 3884 8084
rect 3839 8044 3884 8072
rect 3878 8032 3884 8044
rect 3936 8032 3942 8084
rect 3970 8032 3976 8084
rect 4028 8072 4034 8084
rect 4249 8075 4307 8081
rect 4249 8072 4261 8075
rect 4028 8044 4261 8072
rect 4028 8032 4034 8044
rect 4249 8041 4261 8044
rect 4295 8041 4307 8075
rect 4249 8035 4307 8041
rect 4522 8032 4528 8084
rect 4580 8072 4586 8084
rect 4617 8075 4675 8081
rect 4617 8072 4629 8075
rect 4580 8044 4629 8072
rect 4580 8032 4586 8044
rect 4617 8041 4629 8044
rect 4663 8041 4675 8075
rect 5166 8072 5172 8084
rect 5127 8044 5172 8072
rect 4617 8035 4675 8041
rect 5166 8032 5172 8044
rect 5224 8032 5230 8084
rect 5810 8072 5816 8084
rect 5771 8044 5816 8072
rect 5810 8032 5816 8044
rect 5868 8032 5874 8084
rect 9674 8032 9680 8084
rect 9732 8072 9738 8084
rect 11330 8072 11336 8084
rect 9732 8044 9812 8072
rect 11291 8044 11336 8072
rect 9732 8032 9738 8044
rect 2406 8004 2412 8016
rect 2319 7976 2412 8004
rect 2406 7964 2412 7976
rect 2464 8004 2470 8016
rect 2464 7976 5574 8004
rect 2464 7964 2470 7976
rect 3694 7896 3700 7948
rect 3752 7936 3758 7948
rect 4065 7939 4123 7945
rect 4065 7936 4077 7939
rect 3752 7908 4077 7936
rect 3752 7896 3758 7908
rect 4065 7905 4077 7908
rect 4111 7905 4123 7939
rect 5442 7936 5448 7948
rect 5403 7908 5448 7936
rect 4065 7899 4123 7905
rect 5442 7896 5448 7908
rect 5500 7896 5506 7948
rect 5546 7936 5574 7976
rect 8110 7964 8116 8016
rect 8168 8004 8174 8016
rect 9784 8013 9812 8044
rect 11330 8032 11336 8044
rect 11388 8032 11394 8084
rect 13541 8075 13599 8081
rect 13541 8041 13553 8075
rect 13587 8072 13599 8075
rect 13722 8072 13728 8084
rect 13587 8044 13728 8072
rect 13587 8041 13599 8044
rect 13541 8035 13599 8041
rect 13722 8032 13728 8044
rect 13780 8032 13786 8084
rect 14642 8072 14648 8084
rect 14603 8044 14648 8072
rect 14642 8032 14648 8044
rect 14700 8032 14706 8084
rect 15102 8072 15108 8084
rect 15063 8044 15108 8072
rect 15102 8032 15108 8044
rect 15160 8032 15166 8084
rect 16485 8075 16543 8081
rect 16485 8041 16497 8075
rect 16531 8072 16543 8075
rect 16574 8072 16580 8084
rect 16531 8044 16580 8072
rect 16531 8041 16543 8044
rect 16485 8035 16543 8041
rect 16574 8032 16580 8044
rect 16632 8072 16638 8084
rect 17770 8072 17776 8084
rect 16632 8044 17776 8072
rect 16632 8032 16638 8044
rect 17770 8032 17776 8044
rect 17828 8032 17834 8084
rect 18141 8075 18199 8081
rect 18141 8041 18153 8075
rect 18187 8072 18199 8075
rect 18414 8072 18420 8084
rect 18187 8044 18420 8072
rect 18187 8041 18199 8044
rect 18141 8035 18199 8041
rect 18414 8032 18420 8044
rect 18472 8032 18478 8084
rect 18966 8032 18972 8084
rect 19024 8072 19030 8084
rect 19061 8075 19119 8081
rect 19061 8072 19073 8075
rect 19024 8044 19073 8072
rect 19024 8032 19030 8044
rect 19061 8041 19073 8044
rect 19107 8041 19119 8075
rect 19061 8035 19119 8041
rect 19518 8032 19524 8084
rect 19576 8072 19582 8084
rect 22557 8075 22615 8081
rect 22557 8072 22569 8075
rect 19576 8044 22569 8072
rect 19576 8032 19582 8044
rect 22557 8041 22569 8044
rect 22603 8072 22615 8075
rect 22646 8072 22652 8084
rect 22603 8044 22652 8072
rect 22603 8041 22615 8044
rect 22557 8035 22615 8041
rect 22646 8032 22652 8044
rect 22704 8032 22710 8084
rect 23290 8032 23296 8084
rect 23348 8072 23354 8084
rect 23937 8075 23995 8081
rect 23937 8072 23949 8075
rect 23348 8044 23949 8072
rect 23348 8032 23354 8044
rect 23937 8041 23949 8044
rect 23983 8072 23995 8075
rect 26329 8075 26387 8081
rect 23983 8044 24624 8072
rect 23983 8041 23995 8044
rect 23937 8035 23995 8041
rect 8205 8007 8263 8013
rect 8205 8004 8217 8007
rect 8168 7976 8217 8004
rect 8168 7964 8174 7976
rect 8205 7973 8217 7976
rect 8251 8004 8263 8007
rect 9769 8007 9827 8013
rect 8251 7976 9168 8004
rect 8251 7973 8263 7976
rect 8205 7967 8263 7973
rect 5902 7936 5908 7948
rect 5546 7908 5908 7936
rect 5902 7896 5908 7908
rect 5960 7936 5966 7948
rect 6365 7939 6423 7945
rect 6365 7936 6377 7939
rect 5960 7908 6377 7936
rect 5960 7896 5966 7908
rect 6365 7905 6377 7908
rect 6411 7905 6423 7939
rect 6365 7899 6423 7905
rect 8754 7896 8760 7948
rect 8812 7936 8818 7948
rect 8812 7908 8857 7936
rect 8812 7896 8818 7908
rect 2317 7871 2375 7877
rect 2317 7837 2329 7871
rect 2363 7837 2375 7871
rect 2317 7831 2375 7837
rect 2961 7871 3019 7877
rect 2961 7837 2973 7871
rect 3007 7868 3019 7871
rect 3418 7868 3424 7880
rect 3007 7840 3424 7868
rect 3007 7837 3019 7840
rect 2961 7831 3019 7837
rect 1946 7760 1952 7812
rect 2004 7800 2010 7812
rect 2332 7800 2360 7831
rect 3418 7828 3424 7840
rect 3476 7828 3482 7880
rect 8113 7871 8171 7877
rect 8113 7837 8125 7871
rect 8159 7868 8171 7871
rect 8202 7868 8208 7880
rect 8159 7840 8208 7868
rect 8159 7837 8171 7840
rect 8113 7831 8171 7837
rect 8202 7828 8208 7840
rect 8260 7868 8266 7880
rect 8938 7868 8944 7880
rect 8260 7840 8944 7868
rect 8260 7828 8266 7840
rect 8938 7828 8944 7840
rect 8996 7828 9002 7880
rect 9140 7868 9168 7976
rect 9769 7973 9781 8007
rect 9815 7973 9827 8007
rect 9769 7967 9827 7973
rect 9858 7964 9864 8016
rect 9916 8004 9922 8016
rect 10410 8004 10416 8016
rect 9916 7976 9961 8004
rect 10371 7976 10416 8004
rect 9916 7964 9922 7976
rect 10410 7964 10416 7976
rect 10468 7964 10474 8016
rect 13814 7964 13820 8016
rect 13872 8004 13878 8016
rect 13872 7976 13917 8004
rect 13872 7964 13878 7976
rect 15010 7964 15016 8016
rect 15068 8004 15074 8016
rect 15473 8007 15531 8013
rect 15473 8004 15485 8007
rect 15068 7976 15485 8004
rect 15068 7964 15074 7976
rect 15473 7973 15485 7976
rect 15519 7973 15531 8007
rect 16022 8004 16028 8016
rect 15983 7976 16028 8004
rect 15473 7967 15531 7973
rect 16022 7964 16028 7976
rect 16080 7964 16086 8016
rect 17034 7964 17040 8016
rect 17092 8004 17098 8016
rect 17215 8007 17273 8013
rect 17215 8004 17227 8007
rect 17092 7976 17227 8004
rect 17092 7964 17098 7976
rect 17215 7973 17227 7976
rect 17261 8004 17273 8007
rect 17862 8004 17868 8016
rect 17261 7976 17868 8004
rect 17261 7973 17273 7976
rect 17215 7967 17273 7973
rect 17862 7964 17868 7976
rect 17920 7964 17926 8016
rect 20714 8004 20720 8016
rect 20675 7976 20720 8004
rect 20714 7964 20720 7976
rect 20772 7964 20778 8016
rect 22830 7964 22836 8016
rect 22888 8004 22894 8016
rect 23103 8007 23161 8013
rect 23103 8004 23115 8007
rect 22888 7976 23115 8004
rect 22888 7964 22894 7976
rect 23103 7973 23115 7976
rect 23149 8004 23161 8007
rect 23474 8004 23480 8016
rect 23149 7976 23480 8004
rect 23149 7973 23161 7976
rect 23103 7967 23161 7973
rect 23474 7964 23480 7976
rect 23532 7964 23538 8016
rect 24596 8013 24624 8044
rect 26329 8041 26341 8075
rect 26375 8072 26387 8075
rect 26510 8072 26516 8084
rect 26375 8044 26516 8072
rect 26375 8041 26387 8044
rect 26329 8035 26387 8041
rect 26510 8032 26516 8044
rect 26568 8072 26574 8084
rect 26605 8075 26663 8081
rect 26605 8072 26617 8075
rect 26568 8044 26617 8072
rect 26568 8032 26574 8044
rect 26605 8041 26617 8044
rect 26651 8041 26663 8075
rect 26605 8035 26663 8041
rect 26970 8032 26976 8084
rect 27028 8072 27034 8084
rect 29641 8075 29699 8081
rect 29641 8072 29653 8075
rect 27028 8044 29653 8072
rect 27028 8032 27034 8044
rect 29641 8041 29653 8044
rect 29687 8072 29699 8075
rect 29914 8072 29920 8084
rect 29687 8044 29920 8072
rect 29687 8041 29699 8044
rect 29641 8035 29699 8041
rect 29914 8032 29920 8044
rect 29972 8072 29978 8084
rect 30650 8072 30656 8084
rect 29972 8044 30656 8072
rect 29972 8032 29978 8044
rect 24581 8007 24639 8013
rect 24581 7973 24593 8007
rect 24627 7973 24639 8007
rect 24581 7967 24639 7973
rect 24673 8007 24731 8013
rect 24673 7973 24685 8007
rect 24719 8004 24731 8007
rect 24762 8004 24768 8016
rect 24719 7976 24768 8004
rect 24719 7973 24731 7976
rect 24673 7967 24731 7973
rect 24762 7964 24768 7976
rect 24820 7964 24826 8016
rect 28718 8004 28724 8016
rect 26988 7976 28724 8004
rect 11517 7939 11575 7945
rect 11517 7905 11529 7939
rect 11563 7905 11575 7939
rect 11517 7899 11575 7905
rect 9858 7868 9864 7880
rect 9140 7840 9864 7868
rect 9858 7828 9864 7840
rect 9916 7828 9922 7880
rect 11532 7868 11560 7899
rect 11698 7896 11704 7948
rect 11756 7936 11762 7948
rect 11793 7939 11851 7945
rect 11793 7936 11805 7939
rect 11756 7908 11805 7936
rect 11756 7896 11762 7908
rect 11793 7905 11805 7908
rect 11839 7936 11851 7939
rect 12710 7936 12716 7948
rect 11839 7908 12716 7936
rect 11839 7905 11851 7908
rect 11793 7899 11851 7905
rect 12710 7896 12716 7908
rect 12768 7896 12774 7948
rect 16853 7939 16911 7945
rect 16853 7905 16865 7939
rect 16899 7936 16911 7939
rect 16942 7936 16948 7948
rect 16899 7908 16948 7936
rect 16899 7905 16911 7908
rect 16853 7899 16911 7905
rect 16942 7896 16948 7908
rect 17000 7896 17006 7948
rect 18690 7896 18696 7948
rect 18748 7936 18754 7948
rect 18966 7936 18972 7948
rect 18748 7908 18972 7936
rect 18748 7896 18754 7908
rect 18966 7896 18972 7908
rect 19024 7896 19030 7948
rect 19426 7936 19432 7948
rect 19387 7908 19432 7936
rect 19426 7896 19432 7908
rect 19484 7896 19490 7948
rect 21177 7939 21235 7945
rect 21177 7905 21189 7939
rect 21223 7905 21235 7939
rect 21358 7936 21364 7948
rect 21319 7908 21364 7936
rect 21177 7899 21235 7905
rect 12066 7868 12072 7880
rect 11532 7840 12072 7868
rect 12066 7828 12072 7840
rect 12124 7828 12130 7880
rect 13538 7828 13544 7880
rect 13596 7868 13602 7880
rect 13725 7871 13783 7877
rect 13725 7868 13737 7871
rect 13596 7840 13737 7868
rect 13596 7828 13602 7840
rect 13725 7837 13737 7840
rect 13771 7837 13783 7871
rect 13725 7831 13783 7837
rect 14369 7871 14427 7877
rect 14369 7837 14381 7871
rect 14415 7868 14427 7871
rect 14642 7868 14648 7880
rect 14415 7840 14648 7868
rect 14415 7837 14427 7840
rect 14369 7831 14427 7837
rect 14642 7828 14648 7840
rect 14700 7828 14706 7880
rect 15378 7868 15384 7880
rect 15339 7840 15384 7868
rect 15378 7828 15384 7840
rect 15436 7828 15442 7880
rect 18877 7871 18935 7877
rect 18877 7837 18889 7871
rect 18923 7868 18935 7871
rect 19058 7868 19064 7880
rect 18923 7840 19064 7868
rect 18923 7837 18935 7840
rect 18877 7831 18935 7837
rect 19058 7828 19064 7840
rect 19116 7828 19122 7880
rect 21192 7868 21220 7899
rect 21358 7896 21364 7908
rect 21416 7896 21422 7948
rect 22738 7936 22744 7948
rect 22699 7908 22744 7936
rect 22738 7896 22744 7908
rect 22796 7896 22802 7948
rect 23658 7936 23664 7948
rect 23619 7908 23664 7936
rect 23658 7896 23664 7908
rect 23716 7896 23722 7948
rect 26418 7896 26424 7948
rect 26476 7936 26482 7948
rect 26513 7939 26571 7945
rect 26513 7936 26525 7939
rect 26476 7908 26525 7936
rect 26476 7896 26482 7908
rect 26513 7905 26525 7908
rect 26559 7905 26571 7939
rect 26513 7899 26571 7905
rect 26602 7896 26608 7948
rect 26660 7936 26666 7948
rect 26988 7945 27016 7976
rect 28718 7964 28724 7976
rect 28776 7964 28782 8016
rect 30253 8013 30281 8044
rect 30650 8032 30656 8044
rect 30708 8032 30714 8084
rect 30834 8072 30840 8084
rect 30795 8044 30840 8072
rect 30834 8032 30840 8044
rect 30892 8032 30898 8084
rect 31662 8072 31668 8084
rect 31623 8044 31668 8072
rect 31662 8032 31668 8044
rect 31720 8032 31726 8084
rect 32490 8072 32496 8084
rect 32451 8044 32496 8072
rect 32490 8032 32496 8044
rect 32548 8032 32554 8084
rect 34241 8075 34299 8081
rect 34241 8041 34253 8075
rect 34287 8072 34299 8075
rect 34698 8072 34704 8084
rect 34287 8044 34704 8072
rect 34287 8041 34299 8044
rect 34241 8035 34299 8041
rect 34698 8032 34704 8044
rect 34756 8032 34762 8084
rect 34974 8032 34980 8084
rect 35032 8072 35038 8084
rect 35345 8075 35403 8081
rect 35345 8072 35357 8075
rect 35032 8044 35357 8072
rect 35032 8032 35038 8044
rect 35345 8041 35357 8044
rect 35391 8041 35403 8075
rect 35345 8035 35403 8041
rect 30238 8007 30296 8013
rect 30238 8004 30250 8007
rect 30216 7976 30250 8004
rect 30238 7973 30250 7976
rect 30284 7973 30296 8007
rect 30238 7967 30296 7973
rect 34146 7964 34152 8016
rect 34204 8004 34210 8016
rect 34425 8007 34483 8013
rect 34425 8004 34437 8007
rect 34204 7976 34437 8004
rect 34204 7964 34210 7976
rect 34425 7973 34437 7976
rect 34471 7973 34483 8007
rect 34425 7967 34483 7973
rect 34514 7964 34520 8016
rect 34572 8004 34578 8016
rect 35069 8007 35127 8013
rect 34572 7976 34617 8004
rect 34572 7964 34578 7976
rect 35069 7973 35081 8007
rect 35115 8004 35127 8007
rect 35250 8004 35256 8016
rect 35115 7976 35256 8004
rect 35115 7973 35127 7976
rect 35069 7967 35127 7973
rect 35250 7964 35256 7976
rect 35308 7964 35314 8016
rect 35986 8004 35992 8016
rect 35947 7976 35992 8004
rect 35986 7964 35992 7976
rect 36044 7964 36050 8016
rect 36078 7964 36084 8016
rect 36136 8004 36142 8016
rect 36136 7976 36181 8004
rect 36136 7964 36142 7976
rect 26973 7939 27031 7945
rect 26973 7936 26985 7939
rect 26660 7908 26985 7936
rect 26660 7896 26666 7908
rect 26973 7905 26985 7908
rect 27019 7905 27031 7939
rect 28353 7939 28411 7945
rect 28353 7936 28365 7939
rect 26973 7899 27031 7905
rect 28184 7908 28365 7936
rect 21266 7868 21272 7880
rect 21192 7840 21272 7868
rect 5258 7800 5264 7812
rect 2004 7772 5264 7800
rect 2004 7760 2010 7772
rect 5258 7760 5264 7772
rect 5316 7760 5322 7812
rect 16482 7760 16488 7812
rect 16540 7800 16546 7812
rect 21192 7800 21220 7840
rect 21266 7828 21272 7840
rect 21324 7828 21330 7880
rect 21634 7868 21640 7880
rect 21547 7840 21640 7868
rect 21634 7828 21640 7840
rect 21692 7868 21698 7880
rect 21913 7871 21971 7877
rect 21913 7868 21925 7871
rect 21692 7840 21925 7868
rect 21692 7828 21698 7840
rect 21913 7837 21925 7840
rect 21959 7837 21971 7871
rect 21913 7831 21971 7837
rect 24670 7828 24676 7880
rect 24728 7868 24734 7880
rect 24857 7871 24915 7877
rect 24857 7868 24869 7871
rect 24728 7840 24869 7868
rect 24728 7828 24734 7840
rect 24857 7837 24869 7840
rect 24903 7837 24915 7871
rect 24857 7831 24915 7837
rect 16540 7772 21220 7800
rect 16540 7760 16546 7772
rect 24302 7760 24308 7812
rect 24360 7800 24366 7812
rect 28184 7809 28212 7908
rect 28353 7905 28365 7908
rect 28399 7905 28411 7939
rect 28810 7936 28816 7948
rect 28771 7908 28816 7936
rect 28353 7899 28411 7905
rect 28810 7896 28816 7908
rect 28868 7896 28874 7948
rect 29089 7939 29147 7945
rect 29089 7905 29101 7939
rect 29135 7936 29147 7939
rect 31846 7936 31852 7948
rect 29135 7908 31852 7936
rect 29135 7905 29147 7908
rect 29089 7899 29147 7905
rect 31846 7896 31852 7908
rect 31904 7896 31910 7948
rect 29914 7868 29920 7880
rect 29875 7840 29920 7868
rect 29914 7828 29920 7840
rect 29972 7828 29978 7880
rect 32122 7868 32128 7880
rect 32083 7840 32128 7868
rect 32122 7828 32128 7840
rect 32180 7828 32186 7880
rect 33686 7828 33692 7880
rect 33744 7868 33750 7880
rect 34514 7868 34520 7880
rect 33744 7840 34520 7868
rect 33744 7828 33750 7840
rect 34514 7828 34520 7840
rect 34572 7868 34578 7880
rect 36078 7868 36084 7880
rect 34572 7840 36084 7868
rect 34572 7828 34578 7840
rect 36078 7828 36084 7840
rect 36136 7828 36142 7880
rect 36262 7868 36268 7880
rect 36223 7840 36268 7868
rect 36262 7828 36268 7840
rect 36320 7828 36326 7880
rect 28169 7803 28227 7809
rect 28169 7800 28181 7803
rect 24360 7772 28181 7800
rect 24360 7760 24366 7772
rect 28169 7769 28181 7772
rect 28215 7769 28227 7803
rect 28169 7763 28227 7769
rect 30374 7760 30380 7812
rect 30432 7800 30438 7812
rect 31754 7800 31760 7812
rect 30432 7772 31760 7800
rect 30432 7760 30438 7772
rect 31754 7760 31760 7772
rect 31812 7800 31818 7812
rect 36446 7800 36452 7812
rect 31812 7772 36452 7800
rect 31812 7760 31818 7772
rect 36446 7760 36452 7772
rect 36504 7760 36510 7812
rect 1765 7735 1823 7741
rect 1765 7701 1777 7735
rect 1811 7732 1823 7735
rect 2682 7732 2688 7744
rect 1811 7704 2688 7732
rect 1811 7701 1823 7704
rect 1765 7695 1823 7701
rect 2682 7692 2688 7704
rect 2740 7692 2746 7744
rect 10042 7692 10048 7744
rect 10100 7732 10106 7744
rect 10689 7735 10747 7741
rect 10689 7732 10701 7735
rect 10100 7704 10701 7732
rect 10100 7692 10106 7704
rect 10689 7701 10701 7704
rect 10735 7701 10747 7735
rect 10689 7695 10747 7701
rect 12529 7735 12587 7741
rect 12529 7701 12541 7735
rect 12575 7732 12587 7735
rect 12618 7732 12624 7744
rect 12575 7704 12624 7732
rect 12575 7701 12587 7704
rect 12529 7695 12587 7701
rect 12618 7692 12624 7704
rect 12676 7692 12682 7744
rect 20070 7732 20076 7744
rect 19983 7704 20076 7732
rect 20070 7692 20076 7704
rect 20128 7732 20134 7744
rect 21542 7732 21548 7744
rect 20128 7704 21548 7732
rect 20128 7692 20134 7704
rect 21542 7692 21548 7704
rect 21600 7692 21606 7744
rect 24397 7735 24455 7741
rect 24397 7701 24409 7735
rect 24443 7732 24455 7735
rect 24854 7732 24860 7744
rect 24443 7704 24860 7732
rect 24443 7701 24455 7704
rect 24397 7695 24455 7701
rect 24854 7692 24860 7704
rect 24912 7692 24918 7744
rect 25498 7732 25504 7744
rect 25459 7704 25504 7732
rect 25498 7692 25504 7704
rect 25556 7732 25562 7744
rect 27522 7732 27528 7744
rect 25556 7704 27528 7732
rect 25556 7692 25562 7704
rect 27522 7692 27528 7704
rect 27580 7692 27586 7744
rect 27706 7732 27712 7744
rect 27667 7704 27712 7732
rect 27706 7692 27712 7704
rect 27764 7692 27770 7744
rect 33045 7735 33103 7741
rect 33045 7701 33057 7735
rect 33091 7732 33103 7735
rect 33686 7732 33692 7744
rect 33091 7704 33692 7732
rect 33091 7701 33103 7704
rect 33045 7695 33103 7701
rect 33686 7692 33692 7704
rect 33744 7692 33750 7744
rect 1104 7642 38824 7664
rect 1104 7590 7648 7642
rect 7700 7590 7712 7642
rect 7764 7590 7776 7642
rect 7828 7590 7840 7642
rect 7892 7590 20982 7642
rect 21034 7590 21046 7642
rect 21098 7590 21110 7642
rect 21162 7590 21174 7642
rect 21226 7590 34315 7642
rect 34367 7590 34379 7642
rect 34431 7590 34443 7642
rect 34495 7590 34507 7642
rect 34559 7590 38824 7642
rect 1104 7568 38824 7590
rect 2225 7531 2283 7537
rect 2225 7497 2237 7531
rect 2271 7528 2283 7531
rect 2406 7528 2412 7540
rect 2271 7500 2412 7528
rect 2271 7497 2283 7500
rect 2225 7491 2283 7497
rect 2406 7488 2412 7500
rect 2464 7488 2470 7540
rect 2590 7488 2596 7540
rect 2648 7528 2654 7540
rect 3694 7528 3700 7540
rect 2648 7500 3700 7528
rect 2648 7488 2654 7500
rect 3694 7488 3700 7500
rect 3752 7488 3758 7540
rect 4522 7488 4528 7540
rect 4580 7528 4586 7540
rect 4801 7531 4859 7537
rect 4801 7528 4813 7531
rect 4580 7500 4813 7528
rect 4580 7488 4586 7500
rect 4801 7497 4813 7500
rect 4847 7497 4859 7531
rect 4801 7491 4859 7497
rect 5169 7531 5227 7537
rect 5169 7497 5181 7531
rect 5215 7528 5227 7531
rect 5442 7528 5448 7540
rect 5215 7500 5448 7528
rect 5215 7497 5227 7500
rect 5169 7491 5227 7497
rect 5442 7488 5448 7500
rect 5500 7488 5506 7540
rect 8110 7528 8116 7540
rect 8071 7500 8116 7528
rect 8110 7488 8116 7500
rect 8168 7488 8174 7540
rect 8662 7528 8668 7540
rect 8623 7500 8668 7528
rect 8662 7488 8668 7500
rect 8720 7488 8726 7540
rect 11698 7528 11704 7540
rect 11659 7500 11704 7528
rect 11698 7488 11704 7500
rect 11756 7488 11762 7540
rect 15010 7488 15016 7540
rect 15068 7528 15074 7540
rect 15289 7531 15347 7537
rect 15289 7528 15301 7531
rect 15068 7500 15301 7528
rect 15068 7488 15074 7500
rect 15289 7497 15301 7500
rect 15335 7497 15347 7531
rect 15289 7491 15347 7497
rect 16942 7488 16948 7540
rect 17000 7528 17006 7540
rect 17313 7531 17371 7537
rect 17313 7528 17325 7531
rect 17000 7500 17325 7528
rect 17000 7488 17006 7500
rect 17313 7497 17325 7500
rect 17359 7497 17371 7531
rect 17770 7528 17776 7540
rect 17731 7500 17776 7528
rect 17313 7491 17371 7497
rect 17770 7488 17776 7500
rect 17828 7488 17834 7540
rect 18966 7488 18972 7540
rect 19024 7528 19030 7540
rect 19061 7531 19119 7537
rect 19061 7528 19073 7531
rect 19024 7500 19073 7528
rect 19024 7488 19030 7500
rect 19061 7497 19073 7500
rect 19107 7497 19119 7531
rect 19426 7528 19432 7540
rect 19387 7500 19432 7528
rect 19061 7491 19119 7497
rect 19426 7488 19432 7500
rect 19484 7488 19490 7540
rect 19886 7528 19892 7540
rect 19847 7500 19892 7528
rect 19886 7488 19892 7500
rect 19944 7488 19950 7540
rect 22738 7488 22744 7540
rect 22796 7528 22802 7540
rect 23201 7531 23259 7537
rect 23201 7528 23213 7531
rect 22796 7500 23213 7528
rect 22796 7488 22802 7500
rect 23201 7497 23213 7500
rect 23247 7497 23259 7531
rect 24762 7528 24768 7540
rect 24675 7500 24768 7528
rect 23201 7491 23259 7497
rect 24762 7488 24768 7500
rect 24820 7528 24826 7540
rect 26786 7528 26792 7540
rect 24820 7500 26792 7528
rect 24820 7488 24826 7500
rect 26786 7488 26792 7500
rect 26844 7488 26850 7540
rect 26878 7488 26884 7540
rect 26936 7528 26942 7540
rect 27433 7531 27491 7537
rect 27433 7528 27445 7531
rect 26936 7500 27445 7528
rect 26936 7488 26942 7500
rect 27433 7497 27445 7500
rect 27479 7497 27491 7531
rect 27433 7491 27491 7497
rect 3878 7420 3884 7472
rect 3936 7460 3942 7472
rect 5767 7463 5825 7469
rect 5767 7460 5779 7463
rect 3936 7432 5779 7460
rect 3936 7420 3942 7432
rect 5767 7429 5779 7432
rect 5813 7429 5825 7463
rect 5767 7423 5825 7429
rect 13265 7463 13323 7469
rect 13265 7429 13277 7463
rect 13311 7460 13323 7463
rect 13906 7460 13912 7472
rect 13311 7432 13912 7460
rect 13311 7429 13323 7432
rect 13265 7423 13323 7429
rect 13906 7420 13912 7432
rect 13964 7420 13970 7472
rect 17034 7460 17040 7472
rect 16995 7432 17040 7460
rect 17034 7420 17040 7432
rect 17092 7420 17098 7472
rect 17954 7420 17960 7472
rect 18012 7460 18018 7472
rect 18693 7463 18751 7469
rect 18693 7460 18705 7463
rect 18012 7432 18705 7460
rect 18012 7420 18018 7432
rect 18693 7429 18705 7432
rect 18739 7429 18751 7463
rect 22830 7460 22836 7472
rect 22791 7432 22836 7460
rect 18693 7423 18751 7429
rect 22830 7420 22836 7432
rect 22888 7420 22894 7472
rect 22922 7420 22928 7472
rect 22980 7460 22986 7472
rect 22980 7432 25360 7460
rect 22980 7420 22986 7432
rect 2409 7395 2467 7401
rect 2409 7361 2421 7395
rect 2455 7392 2467 7395
rect 2682 7392 2688 7404
rect 2455 7364 2688 7392
rect 2455 7361 2467 7364
rect 2409 7355 2467 7361
rect 2682 7352 2688 7364
rect 2740 7352 2746 7404
rect 5074 7392 5080 7404
rect 3896 7364 5080 7392
rect 3896 7336 3924 7364
rect 5074 7352 5080 7364
rect 5132 7352 5138 7404
rect 6270 7352 6276 7404
rect 6328 7392 6334 7404
rect 6730 7392 6736 7404
rect 6328 7364 6736 7392
rect 6328 7352 6334 7364
rect 6730 7352 6736 7364
rect 6788 7392 6794 7404
rect 8849 7395 8907 7401
rect 6788 7364 7328 7392
rect 6788 7352 6794 7364
rect 3053 7327 3111 7333
rect 3053 7293 3065 7327
rect 3099 7324 3111 7327
rect 3418 7324 3424 7336
rect 3099 7296 3424 7324
rect 3099 7293 3111 7296
rect 3053 7287 3111 7293
rect 3418 7284 3424 7296
rect 3476 7284 3482 7336
rect 3878 7324 3884 7336
rect 3839 7296 3884 7324
rect 3878 7284 3884 7296
rect 3936 7284 3942 7336
rect 4522 7324 4528 7336
rect 4126 7296 4528 7324
rect 1857 7259 1915 7265
rect 1857 7225 1869 7259
rect 1903 7256 1915 7259
rect 2501 7259 2559 7265
rect 1903 7228 2360 7256
rect 1903 7225 1915 7228
rect 1857 7219 1915 7225
rect 2332 7188 2360 7228
rect 2501 7225 2513 7259
rect 2547 7225 2559 7259
rect 4126 7256 4154 7296
rect 4522 7284 4528 7296
rect 4580 7284 4586 7336
rect 4614 7284 4620 7336
rect 4672 7324 4678 7336
rect 5696 7327 5754 7333
rect 5696 7324 5708 7327
rect 4672 7296 5708 7324
rect 4672 7284 4678 7296
rect 5696 7293 5708 7296
rect 5742 7324 5754 7327
rect 6089 7327 6147 7333
rect 6089 7324 6101 7327
rect 5742 7296 6101 7324
rect 5742 7293 5754 7296
rect 5696 7287 5754 7293
rect 6089 7293 6101 7296
rect 6135 7293 6147 7327
rect 6089 7287 6147 7293
rect 6641 7327 6699 7333
rect 6641 7293 6653 7327
rect 6687 7324 6699 7327
rect 7098 7324 7104 7336
rect 6687 7296 7104 7324
rect 6687 7293 6699 7296
rect 6641 7287 6699 7293
rect 7098 7284 7104 7296
rect 7156 7284 7162 7336
rect 7300 7333 7328 7364
rect 8849 7361 8861 7395
rect 8895 7392 8907 7395
rect 9122 7392 9128 7404
rect 8895 7364 9128 7392
rect 8895 7361 8907 7364
rect 8849 7355 8907 7361
rect 9122 7352 9128 7364
rect 9180 7392 9186 7404
rect 11330 7392 11336 7404
rect 9180 7364 11336 7392
rect 9180 7352 9186 7364
rect 11330 7352 11336 7364
rect 11388 7352 11394 7404
rect 12897 7395 12955 7401
rect 12897 7361 12909 7395
rect 12943 7392 12955 7395
rect 13814 7392 13820 7404
rect 12943 7364 13820 7392
rect 12943 7361 12955 7364
rect 12897 7355 12955 7361
rect 13786 7352 13820 7364
rect 13872 7352 13878 7404
rect 15013 7395 15071 7401
rect 15013 7361 15025 7395
rect 15059 7392 15071 7395
rect 15378 7392 15384 7404
rect 15059 7364 15384 7392
rect 15059 7361 15071 7364
rect 15013 7355 15071 7361
rect 15378 7352 15384 7364
rect 15436 7352 15442 7404
rect 16022 7392 16028 7404
rect 15935 7364 16028 7392
rect 16022 7352 16028 7364
rect 16080 7392 16086 7404
rect 17126 7392 17132 7404
rect 16080 7364 17132 7392
rect 16080 7352 16086 7364
rect 17126 7352 17132 7364
rect 17184 7352 17190 7404
rect 18141 7395 18199 7401
rect 18141 7361 18153 7395
rect 18187 7392 18199 7395
rect 18414 7392 18420 7404
rect 18187 7364 18420 7392
rect 18187 7361 18199 7364
rect 18141 7355 18199 7361
rect 18414 7352 18420 7364
rect 18472 7352 18478 7404
rect 21174 7392 21180 7404
rect 21135 7364 21180 7392
rect 21174 7352 21180 7364
rect 21232 7352 21238 7404
rect 21634 7392 21640 7404
rect 21595 7364 21640 7392
rect 21634 7352 21640 7364
rect 21692 7352 21698 7404
rect 22646 7352 22652 7404
rect 22704 7392 22710 7404
rect 25332 7401 25360 7432
rect 23753 7395 23811 7401
rect 23753 7392 23765 7395
rect 22704 7364 23765 7392
rect 22704 7352 22710 7364
rect 23753 7361 23765 7364
rect 23799 7361 23811 7395
rect 23753 7355 23811 7361
rect 25317 7395 25375 7401
rect 25317 7361 25329 7395
rect 25363 7392 25375 7395
rect 25590 7392 25596 7404
rect 25363 7364 25596 7392
rect 25363 7361 25375 7364
rect 25317 7355 25375 7361
rect 25590 7352 25596 7364
rect 25648 7352 25654 7404
rect 7285 7327 7343 7333
rect 7285 7293 7297 7327
rect 7331 7293 7343 7327
rect 10597 7327 10655 7333
rect 10597 7324 10609 7327
rect 7285 7287 7343 7293
rect 10060 7296 10609 7324
rect 2501 7219 2559 7225
rect 3160 7228 4154 7256
rect 4243 7259 4301 7265
rect 2516 7188 2544 7219
rect 3160 7188 3188 7228
rect 4243 7225 4255 7259
rect 4289 7225 4301 7259
rect 4243 7219 4301 7225
rect 3326 7188 3332 7200
rect 2332 7160 3188 7188
rect 3287 7160 3332 7188
rect 3326 7148 3332 7160
rect 3384 7188 3390 7200
rect 4258 7188 4286 7219
rect 8662 7216 8668 7268
rect 8720 7256 8726 7268
rect 9170 7259 9228 7265
rect 9170 7256 9182 7259
rect 8720 7228 9182 7256
rect 8720 7216 8726 7228
rect 9170 7225 9182 7228
rect 9216 7256 9228 7259
rect 9306 7256 9312 7268
rect 9216 7228 9312 7256
rect 9216 7225 9228 7228
rect 9170 7219 9228 7225
rect 9306 7216 9312 7228
rect 9364 7216 9370 7268
rect 5445 7191 5503 7197
rect 5445 7188 5457 7191
rect 3384 7160 5457 7188
rect 3384 7148 3390 7160
rect 5445 7157 5457 7160
rect 5491 7188 5503 7191
rect 5810 7188 5816 7200
rect 5491 7160 5816 7188
rect 5491 7157 5503 7160
rect 5445 7151 5503 7157
rect 5810 7148 5816 7160
rect 5868 7148 5874 7200
rect 6914 7188 6920 7200
rect 6875 7160 6920 7188
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 9769 7191 9827 7197
rect 9769 7157 9781 7191
rect 9815 7188 9827 7191
rect 9858 7188 9864 7200
rect 9815 7160 9864 7188
rect 9815 7157 9827 7160
rect 9769 7151 9827 7157
rect 9858 7148 9864 7160
rect 9916 7148 9922 7200
rect 9950 7148 9956 7200
rect 10008 7188 10014 7200
rect 10060 7197 10088 7296
rect 10597 7293 10609 7296
rect 10643 7293 10655 7327
rect 10597 7287 10655 7293
rect 11149 7327 11207 7333
rect 11149 7293 11161 7327
rect 11195 7324 11207 7327
rect 11698 7324 11704 7336
rect 11195 7296 11704 7324
rect 11195 7293 11207 7296
rect 11149 7287 11207 7293
rect 10505 7259 10563 7265
rect 10505 7225 10517 7259
rect 10551 7256 10563 7259
rect 11164 7256 11192 7287
rect 11698 7284 11704 7296
rect 11756 7284 11762 7336
rect 13354 7324 13360 7336
rect 13315 7296 13360 7324
rect 13354 7284 13360 7296
rect 13412 7284 13418 7336
rect 13786 7324 13814 7352
rect 14277 7327 14335 7333
rect 14277 7324 14289 7327
rect 13786 7296 14289 7324
rect 14277 7293 14289 7296
rect 14323 7324 14335 7327
rect 15654 7324 15660 7336
rect 14323 7296 15660 7324
rect 14323 7293 14335 7296
rect 14277 7287 14335 7293
rect 15654 7284 15660 7296
rect 15712 7284 15718 7336
rect 19886 7284 19892 7336
rect 19944 7324 19950 7336
rect 20073 7327 20131 7333
rect 20073 7324 20085 7327
rect 19944 7296 20085 7324
rect 19944 7284 19950 7296
rect 20073 7293 20085 7296
rect 20119 7293 20131 7327
rect 20073 7287 20131 7293
rect 20162 7284 20168 7336
rect 20220 7324 20226 7336
rect 20625 7327 20683 7333
rect 20625 7324 20637 7327
rect 20220 7296 20637 7324
rect 20220 7284 20226 7296
rect 20625 7293 20637 7296
rect 20671 7324 20683 7327
rect 21358 7324 21364 7336
rect 20671 7296 21364 7324
rect 20671 7293 20683 7296
rect 20625 7287 20683 7293
rect 21358 7284 21364 7296
rect 21416 7284 21422 7336
rect 22557 7327 22615 7333
rect 22557 7293 22569 7327
rect 22603 7324 22615 7327
rect 24397 7327 24455 7333
rect 22603 7296 23474 7324
rect 22603 7293 22615 7296
rect 22557 7287 22615 7293
rect 10551 7228 11192 7256
rect 10551 7225 10563 7228
rect 10505 7219 10563 7225
rect 10045 7191 10103 7197
rect 10045 7188 10057 7191
rect 10008 7160 10057 7188
rect 10008 7148 10014 7160
rect 10045 7157 10057 7160
rect 10091 7157 10103 7191
rect 10686 7188 10692 7200
rect 10647 7160 10692 7188
rect 10045 7151 10103 7157
rect 10686 7148 10692 7160
rect 10744 7148 10750 7200
rect 12066 7188 12072 7200
rect 12027 7160 12072 7188
rect 12066 7148 12072 7160
rect 12124 7148 12130 7200
rect 13372 7188 13400 7284
rect 13768 7265 13774 7268
rect 13719 7259 13774 7265
rect 13719 7225 13731 7259
rect 13765 7225 13774 7259
rect 13719 7219 13774 7225
rect 13768 7216 13774 7219
rect 13826 7256 13832 7268
rect 14553 7259 14611 7265
rect 14553 7256 14565 7259
rect 13826 7228 13867 7256
rect 13899 7228 14565 7256
rect 13826 7216 13832 7228
rect 13899 7188 13927 7228
rect 14553 7225 14565 7228
rect 14599 7225 14611 7259
rect 14553 7219 14611 7225
rect 16117 7259 16175 7265
rect 16117 7225 16129 7259
rect 16163 7225 16175 7259
rect 16117 7219 16175 7225
rect 16669 7259 16727 7265
rect 16669 7225 16681 7259
rect 16715 7256 16727 7259
rect 17310 7256 17316 7268
rect 16715 7228 17316 7256
rect 16715 7225 16727 7228
rect 16669 7219 16727 7225
rect 15746 7188 15752 7200
rect 13372 7160 13927 7188
rect 15707 7160 15752 7188
rect 15746 7148 15752 7160
rect 15804 7188 15810 7200
rect 16132 7188 16160 7219
rect 17310 7216 17316 7228
rect 17368 7216 17374 7268
rect 18233 7259 18291 7265
rect 18233 7225 18245 7259
rect 18279 7225 18291 7259
rect 20806 7256 20812 7268
rect 20767 7228 20812 7256
rect 18233 7219 18291 7225
rect 15804 7160 16160 7188
rect 15804 7148 15810 7160
rect 17770 7148 17776 7200
rect 17828 7188 17834 7200
rect 18248 7188 18276 7219
rect 20806 7216 20812 7228
rect 20864 7216 20870 7268
rect 21542 7256 21548 7268
rect 21455 7228 21548 7256
rect 21542 7216 21548 7228
rect 21600 7256 21606 7268
rect 21999 7259 22057 7265
rect 21999 7256 22011 7259
rect 21600 7228 22011 7256
rect 21600 7216 21606 7228
rect 21999 7225 22011 7228
rect 22045 7256 22057 7259
rect 22830 7256 22836 7268
rect 22045 7228 22836 7256
rect 22045 7225 22057 7228
rect 21999 7219 22057 7225
rect 22830 7216 22836 7228
rect 22888 7216 22894 7268
rect 23446 7256 23474 7296
rect 24397 7293 24409 7327
rect 24443 7324 24455 7327
rect 24670 7324 24676 7336
rect 24443 7296 24676 7324
rect 24443 7293 24455 7296
rect 24397 7287 24455 7293
rect 24670 7284 24676 7296
rect 24728 7284 24734 7336
rect 26418 7284 26424 7336
rect 26476 7324 26482 7336
rect 27448 7324 27476 7491
rect 27522 7488 27528 7540
rect 27580 7528 27586 7540
rect 28997 7531 29055 7537
rect 28997 7528 29009 7531
rect 27580 7500 29009 7528
rect 27580 7488 27586 7500
rect 28997 7497 29009 7500
rect 29043 7497 29055 7531
rect 33686 7528 33692 7540
rect 33647 7500 33692 7528
rect 28997 7491 29055 7497
rect 27617 7327 27675 7333
rect 27617 7324 27629 7327
rect 26476 7296 26924 7324
rect 27448 7296 27629 7324
rect 26476 7284 26482 7296
rect 23845 7259 23903 7265
rect 23845 7256 23857 7259
rect 23446 7228 23857 7256
rect 23845 7225 23857 7228
rect 23891 7225 23903 7259
rect 25409 7259 25467 7265
rect 23845 7219 23903 7225
rect 24504 7228 25176 7256
rect 17828 7160 18276 7188
rect 17828 7148 17834 7160
rect 23750 7148 23756 7200
rect 23808 7188 23814 7200
rect 23860 7188 23888 7219
rect 24504 7188 24532 7228
rect 25148 7197 25176 7228
rect 25409 7225 25421 7259
rect 25455 7225 25467 7259
rect 25409 7219 25467 7225
rect 25961 7259 26019 7265
rect 25961 7225 25973 7259
rect 26007 7256 26019 7259
rect 26694 7256 26700 7268
rect 26007 7228 26700 7256
rect 26007 7225 26019 7228
rect 25961 7219 26019 7225
rect 23808 7160 24532 7188
rect 25133 7191 25191 7197
rect 23808 7148 23814 7160
rect 25133 7157 25145 7191
rect 25179 7188 25191 7191
rect 25424 7188 25452 7219
rect 26694 7216 26700 7228
rect 26752 7216 26758 7268
rect 26896 7200 26924 7296
rect 27617 7293 27629 7296
rect 27663 7293 27675 7327
rect 27617 7287 27675 7293
rect 27706 7284 27712 7336
rect 27764 7324 27770 7336
rect 28169 7327 28227 7333
rect 28169 7324 28181 7327
rect 27764 7296 28181 7324
rect 27764 7284 27770 7296
rect 28169 7293 28181 7296
rect 28215 7293 28227 7327
rect 29012 7324 29040 7491
rect 33686 7488 33692 7500
rect 33744 7488 33750 7540
rect 34333 7531 34391 7537
rect 34333 7528 34345 7531
rect 33796 7500 34345 7528
rect 30009 7395 30067 7401
rect 30009 7361 30021 7395
rect 30055 7392 30067 7395
rect 31205 7395 31263 7401
rect 31205 7392 31217 7395
rect 30055 7364 31217 7392
rect 30055 7361 30067 7364
rect 30009 7355 30067 7361
rect 31205 7361 31217 7364
rect 31251 7392 31263 7395
rect 32122 7392 32128 7404
rect 31251 7364 32128 7392
rect 31251 7361 31263 7364
rect 31205 7355 31263 7361
rect 32122 7352 32128 7364
rect 32180 7352 32186 7404
rect 29273 7327 29331 7333
rect 29273 7324 29285 7327
rect 29012 7296 29285 7324
rect 28169 7287 28227 7293
rect 29273 7293 29285 7296
rect 29319 7324 29331 7327
rect 29454 7324 29460 7336
rect 29319 7296 29460 7324
rect 29319 7293 29331 7296
rect 29273 7287 29331 7293
rect 25179 7160 25452 7188
rect 25179 7157 25191 7160
rect 25133 7151 25191 7157
rect 25498 7148 25504 7200
rect 25556 7188 25562 7200
rect 26234 7188 26240 7200
rect 25556 7160 26240 7188
rect 25556 7148 25562 7160
rect 26234 7148 26240 7160
rect 26292 7148 26298 7200
rect 26510 7188 26516 7200
rect 26471 7160 26516 7188
rect 26510 7148 26516 7160
rect 26568 7148 26574 7200
rect 26878 7188 26884 7200
rect 26839 7160 26884 7188
rect 26878 7148 26884 7160
rect 26936 7148 26942 7200
rect 28184 7188 28212 7287
rect 29454 7284 29460 7296
rect 29512 7284 29518 7336
rect 29730 7324 29736 7336
rect 29691 7296 29736 7324
rect 29730 7284 29736 7296
rect 29788 7284 29794 7336
rect 29914 7284 29920 7336
rect 29972 7324 29978 7336
rect 30653 7327 30711 7333
rect 30653 7324 30665 7327
rect 29972 7296 30665 7324
rect 29972 7284 29978 7296
rect 30653 7293 30665 7296
rect 30699 7293 30711 7327
rect 31754 7324 31760 7336
rect 31715 7296 31760 7324
rect 30653 7287 30711 7293
rect 31754 7284 31760 7296
rect 31812 7284 31818 7336
rect 32398 7284 32404 7336
rect 32456 7324 32462 7336
rect 33796 7333 33824 7500
rect 34333 7497 34345 7500
rect 34379 7528 34391 7531
rect 34790 7528 34796 7540
rect 34379 7500 34796 7528
rect 34379 7497 34391 7500
rect 34333 7491 34391 7497
rect 34790 7488 34796 7500
rect 34848 7488 34854 7540
rect 35986 7488 35992 7540
rect 36044 7528 36050 7540
rect 36265 7531 36323 7537
rect 36265 7528 36277 7531
rect 36044 7500 36277 7528
rect 36044 7488 36050 7500
rect 36265 7497 36277 7500
rect 36311 7497 36323 7531
rect 36630 7528 36636 7540
rect 36591 7500 36636 7528
rect 36265 7491 36323 7497
rect 36630 7488 36636 7500
rect 36688 7488 36694 7540
rect 35894 7420 35900 7472
rect 35952 7460 35958 7472
rect 38013 7463 38071 7469
rect 38013 7460 38025 7463
rect 35952 7432 38025 7460
rect 35952 7420 35958 7432
rect 33962 7352 33968 7404
rect 34020 7392 34026 7404
rect 34609 7395 34667 7401
rect 34609 7392 34621 7395
rect 34020 7364 34621 7392
rect 34020 7352 34026 7364
rect 34609 7361 34621 7364
rect 34655 7392 34667 7395
rect 35066 7392 35072 7404
rect 34655 7364 35072 7392
rect 34655 7361 34667 7364
rect 34609 7355 34667 7361
rect 35066 7352 35072 7364
rect 35124 7352 35130 7404
rect 35250 7392 35256 7404
rect 35211 7364 35256 7392
rect 35250 7352 35256 7364
rect 35308 7352 35314 7404
rect 35989 7395 36047 7401
rect 35989 7361 36001 7395
rect 36035 7392 36047 7395
rect 36078 7392 36084 7404
rect 36035 7364 36084 7392
rect 36035 7361 36047 7364
rect 35989 7355 36047 7361
rect 36078 7352 36084 7364
rect 36136 7352 36142 7404
rect 33796 7327 33874 7333
rect 33796 7324 33828 7327
rect 32456 7296 33828 7324
rect 32456 7284 32462 7296
rect 33816 7293 33828 7296
rect 33862 7293 33874 7327
rect 36446 7324 36452 7336
rect 36407 7296 36452 7324
rect 33816 7287 33874 7293
rect 36446 7284 36452 7296
rect 36504 7324 36510 7336
rect 37614 7333 37642 7432
rect 38013 7429 38025 7432
rect 38059 7429 38071 7463
rect 38013 7423 38071 7429
rect 37001 7327 37059 7333
rect 37001 7324 37013 7327
rect 36504 7296 37013 7324
rect 36504 7284 36510 7296
rect 37001 7293 37013 7296
rect 37047 7293 37059 7327
rect 37001 7287 37059 7293
rect 37599 7327 37657 7333
rect 37599 7293 37611 7327
rect 37645 7293 37657 7327
rect 37599 7287 37657 7293
rect 28353 7259 28411 7265
rect 28353 7225 28365 7259
rect 28399 7256 28411 7259
rect 31938 7256 31944 7268
rect 28399 7228 31944 7256
rect 28399 7225 28411 7228
rect 28353 7219 28411 7225
rect 31938 7216 31944 7228
rect 31996 7216 32002 7268
rect 32119 7259 32177 7265
rect 32119 7225 32131 7259
rect 32165 7256 32177 7259
rect 32490 7256 32496 7268
rect 32165 7228 32496 7256
rect 32165 7225 32177 7228
rect 32119 7219 32177 7225
rect 28442 7188 28448 7200
rect 28184 7160 28448 7188
rect 28442 7148 28448 7160
rect 28500 7188 28506 7200
rect 28721 7191 28779 7197
rect 28721 7188 28733 7191
rect 28500 7160 28733 7188
rect 28500 7148 28506 7160
rect 28721 7157 28733 7160
rect 28767 7188 28779 7191
rect 28810 7188 28816 7200
rect 28767 7160 28816 7188
rect 28767 7157 28779 7160
rect 28721 7151 28779 7157
rect 28810 7148 28816 7160
rect 28868 7188 28874 7200
rect 29730 7188 29736 7200
rect 28868 7160 29736 7188
rect 28868 7148 28874 7160
rect 29730 7148 29736 7160
rect 29788 7148 29794 7200
rect 30377 7191 30435 7197
rect 30377 7157 30389 7191
rect 30423 7188 30435 7191
rect 30650 7188 30656 7200
rect 30423 7160 30656 7188
rect 30423 7157 30435 7160
rect 30377 7151 30435 7157
rect 30650 7148 30656 7160
rect 30708 7188 30714 7200
rect 31573 7191 31631 7197
rect 31573 7188 31585 7191
rect 30708 7160 31585 7188
rect 30708 7148 30714 7160
rect 31573 7157 31585 7160
rect 31619 7188 31631 7191
rect 32134 7188 32162 7219
rect 32490 7216 32496 7228
rect 32548 7256 32554 7268
rect 32953 7259 33011 7265
rect 32953 7256 32965 7259
rect 32548 7228 32965 7256
rect 32548 7216 32554 7228
rect 32953 7225 32965 7228
rect 32999 7225 33011 7259
rect 32953 7219 33011 7225
rect 33919 7259 33977 7265
rect 33919 7225 33931 7259
rect 33965 7256 33977 7259
rect 34974 7256 34980 7268
rect 33965 7228 34980 7256
rect 33965 7225 33977 7228
rect 33919 7219 33977 7225
rect 34974 7216 34980 7228
rect 35032 7216 35038 7268
rect 35066 7216 35072 7268
rect 35124 7256 35130 7268
rect 35124 7228 35169 7256
rect 35124 7216 35130 7228
rect 32674 7188 32680 7200
rect 31619 7160 32162 7188
rect 32635 7160 32680 7188
rect 31619 7157 31631 7160
rect 31573 7151 31631 7157
rect 32674 7148 32680 7160
rect 32732 7148 32738 7200
rect 37090 7148 37096 7200
rect 37148 7188 37154 7200
rect 37691 7191 37749 7197
rect 37691 7188 37703 7191
rect 37148 7160 37703 7188
rect 37148 7148 37154 7160
rect 37691 7157 37703 7160
rect 37737 7157 37749 7191
rect 37691 7151 37749 7157
rect 1104 7098 38824 7120
rect 1104 7046 14315 7098
rect 14367 7046 14379 7098
rect 14431 7046 14443 7098
rect 14495 7046 14507 7098
rect 14559 7046 27648 7098
rect 27700 7046 27712 7098
rect 27764 7046 27776 7098
rect 27828 7046 27840 7098
rect 27892 7046 38824 7098
rect 1104 7024 38824 7046
rect 1946 6984 1952 6996
rect 1907 6956 1952 6984
rect 1946 6944 1952 6956
rect 2004 6944 2010 6996
rect 3878 6984 3884 6996
rect 3839 6956 3884 6984
rect 3878 6944 3884 6956
rect 3936 6944 3942 6996
rect 4062 6944 4068 6996
rect 4120 6984 4126 6996
rect 4120 6956 4384 6984
rect 4120 6944 4126 6956
rect 2317 6919 2375 6925
rect 2317 6885 2329 6919
rect 2363 6916 2375 6919
rect 2593 6919 2651 6925
rect 2593 6916 2605 6919
rect 2363 6888 2605 6916
rect 2363 6885 2375 6888
rect 2317 6879 2375 6885
rect 2593 6885 2605 6888
rect 2639 6916 2651 6919
rect 3142 6916 3148 6928
rect 2639 6888 3148 6916
rect 2639 6885 2651 6888
rect 2593 6879 2651 6885
rect 3142 6876 3148 6888
rect 3200 6876 3206 6928
rect 3970 6876 3976 6928
rect 4028 6916 4034 6928
rect 4249 6919 4307 6925
rect 4249 6916 4261 6919
rect 4028 6888 4261 6916
rect 4028 6876 4034 6888
rect 4249 6885 4261 6888
rect 4295 6885 4307 6919
rect 4356 6916 4384 6956
rect 6730 6944 6736 6996
rect 6788 6984 6794 6996
rect 6825 6987 6883 6993
rect 6825 6984 6837 6987
rect 6788 6956 6837 6984
rect 6788 6944 6794 6956
rect 6825 6953 6837 6956
rect 6871 6953 6883 6987
rect 6825 6947 6883 6953
rect 8018 6944 8024 6996
rect 8076 6984 8082 6996
rect 9122 6984 9128 6996
rect 8076 6956 8156 6984
rect 9083 6956 9128 6984
rect 8076 6944 8082 6956
rect 4801 6919 4859 6925
rect 4801 6916 4813 6919
rect 4356 6888 4813 6916
rect 4249 6879 4307 6885
rect 4801 6885 4813 6888
rect 4847 6885 4859 6919
rect 4801 6879 4859 6885
rect 5813 6919 5871 6925
rect 5813 6885 5825 6919
rect 5859 6916 5871 6919
rect 5902 6916 5908 6928
rect 5859 6888 5908 6916
rect 5859 6885 5871 6888
rect 5813 6879 5871 6885
rect 5902 6876 5908 6888
rect 5960 6876 5966 6928
rect 8128 6925 8156 6956
rect 9122 6944 9128 6956
rect 9180 6944 9186 6996
rect 9493 6987 9551 6993
rect 9493 6953 9505 6987
rect 9539 6984 9551 6987
rect 9674 6984 9680 6996
rect 9539 6956 9680 6984
rect 9539 6953 9551 6956
rect 9493 6947 9551 6953
rect 9674 6944 9680 6956
rect 9732 6944 9738 6996
rect 9858 6984 9864 6996
rect 9819 6956 9864 6984
rect 9858 6944 9864 6956
rect 9916 6944 9922 6996
rect 10318 6944 10324 6996
rect 10376 6984 10382 6996
rect 13357 6987 13415 6993
rect 10376 6956 10456 6984
rect 10376 6944 10382 6956
rect 8113 6919 8171 6925
rect 8113 6885 8125 6919
rect 8159 6885 8171 6919
rect 8113 6879 8171 6885
rect 8205 6919 8263 6925
rect 8205 6885 8217 6919
rect 8251 6916 8263 6919
rect 8386 6916 8392 6928
rect 8251 6888 8392 6916
rect 8251 6885 8263 6888
rect 8205 6879 8263 6885
rect 8386 6876 8392 6888
rect 8444 6876 8450 6928
rect 10428 6925 10456 6956
rect 13357 6953 13369 6987
rect 13403 6984 13415 6987
rect 13538 6984 13544 6996
rect 13403 6956 13544 6984
rect 13403 6953 13415 6956
rect 13357 6947 13415 6953
rect 13538 6944 13544 6956
rect 13596 6944 13602 6996
rect 14642 6944 14648 6996
rect 14700 6984 14706 6996
rect 15105 6987 15163 6993
rect 15105 6984 15117 6987
rect 14700 6956 15117 6984
rect 14700 6944 14706 6956
rect 15105 6953 15117 6956
rect 15151 6984 15163 6987
rect 16022 6984 16028 6996
rect 15151 6956 16028 6984
rect 15151 6953 15163 6956
rect 15105 6947 15163 6953
rect 16022 6944 16028 6956
rect 16080 6944 16086 6996
rect 16758 6984 16764 6996
rect 16719 6956 16764 6984
rect 16758 6944 16764 6956
rect 16816 6944 16822 6996
rect 20162 6984 20168 6996
rect 20123 6956 20168 6984
rect 20162 6944 20168 6956
rect 20220 6944 20226 6996
rect 20806 6944 20812 6996
rect 20864 6984 20870 6996
rect 21726 6984 21732 6996
rect 20864 6956 21732 6984
rect 20864 6944 20870 6956
rect 21726 6944 21732 6956
rect 21784 6984 21790 6996
rect 22097 6987 22155 6993
rect 22097 6984 22109 6987
rect 21784 6956 22109 6984
rect 21784 6944 21790 6956
rect 22097 6953 22109 6956
rect 22143 6953 22155 6987
rect 23750 6984 23756 6996
rect 23711 6956 23756 6984
rect 22097 6947 22155 6953
rect 23750 6944 23756 6956
rect 23808 6944 23814 6996
rect 24762 6984 24768 6996
rect 23952 6956 24768 6984
rect 10413 6919 10471 6925
rect 10413 6885 10425 6919
rect 10459 6885 10471 6919
rect 10413 6879 10471 6885
rect 10505 6919 10563 6925
rect 10505 6885 10517 6919
rect 10551 6916 10563 6919
rect 10686 6916 10692 6928
rect 10551 6888 10692 6916
rect 10551 6885 10563 6888
rect 10505 6879 10563 6885
rect 10686 6876 10692 6888
rect 10744 6876 10750 6928
rect 12618 6916 12624 6928
rect 12579 6888 12624 6916
rect 12618 6876 12624 6888
rect 12676 6876 12682 6928
rect 13811 6919 13869 6925
rect 13811 6885 13823 6919
rect 13857 6916 13869 6919
rect 13906 6916 13912 6928
rect 13857 6888 13912 6916
rect 13857 6885 13869 6888
rect 13811 6879 13869 6885
rect 13906 6876 13912 6888
rect 13964 6876 13970 6928
rect 14182 6876 14188 6928
rect 14240 6916 14246 6928
rect 15010 6916 15016 6928
rect 14240 6888 15016 6916
rect 14240 6876 14246 6888
rect 15010 6876 15016 6888
rect 15068 6916 15074 6928
rect 15381 6919 15439 6925
rect 15381 6916 15393 6919
rect 15068 6888 15393 6916
rect 15068 6876 15074 6888
rect 15381 6885 15393 6888
rect 15427 6885 15439 6919
rect 15381 6879 15439 6885
rect 15473 6919 15531 6925
rect 15473 6885 15485 6919
rect 15519 6916 15531 6919
rect 15654 6916 15660 6928
rect 15519 6888 15660 6916
rect 15519 6885 15531 6888
rect 15473 6879 15531 6885
rect 15654 6876 15660 6888
rect 15712 6876 15718 6928
rect 16776 6916 16804 6944
rect 17037 6919 17095 6925
rect 17037 6916 17049 6919
rect 16776 6888 17049 6916
rect 17037 6885 17049 6888
rect 17083 6885 17095 6919
rect 17037 6879 17095 6885
rect 17126 6876 17132 6928
rect 17184 6916 17190 6928
rect 18693 6919 18751 6925
rect 18693 6916 18705 6919
rect 17184 6888 18705 6916
rect 17184 6876 17190 6888
rect 18693 6885 18705 6888
rect 18739 6885 18751 6919
rect 20180 6916 20208 6944
rect 21085 6919 21143 6925
rect 21085 6916 21097 6919
rect 20180 6888 21097 6916
rect 18693 6879 18751 6885
rect 21085 6885 21097 6888
rect 21131 6885 21143 6919
rect 22643 6919 22701 6925
rect 22643 6916 22655 6919
rect 21085 6879 21143 6885
rect 21744 6888 22655 6916
rect 1464 6851 1522 6857
rect 1464 6817 1476 6851
rect 1510 6848 1522 6851
rect 1854 6848 1860 6860
rect 1510 6820 1860 6848
rect 1510 6817 1522 6820
rect 1464 6811 1522 6817
rect 1854 6808 1860 6820
rect 1912 6808 1918 6860
rect 3694 6808 3700 6860
rect 3752 6848 3758 6860
rect 11974 6848 11980 6860
rect 3752 6820 4016 6848
rect 11935 6820 11980 6848
rect 3752 6808 3758 6820
rect 2498 6780 2504 6792
rect 2459 6752 2504 6780
rect 2498 6740 2504 6752
rect 2556 6740 2562 6792
rect 2929 6752 3924 6780
rect 1535 6715 1593 6721
rect 1535 6681 1547 6715
rect 1581 6712 1593 6715
rect 2929 6712 2957 6752
rect 3050 6712 3056 6724
rect 1581 6684 2957 6712
rect 3011 6684 3056 6712
rect 1581 6681 1593 6684
rect 1535 6675 1593 6681
rect 3050 6672 3056 6684
rect 3108 6672 3114 6724
rect 3418 6644 3424 6656
rect 3379 6616 3424 6644
rect 3418 6604 3424 6616
rect 3476 6604 3482 6656
rect 3896 6644 3924 6752
rect 3988 6712 4016 6820
rect 11974 6808 11980 6820
rect 12032 6808 12038 6860
rect 12437 6851 12495 6857
rect 12437 6817 12449 6851
rect 12483 6848 12495 6851
rect 12710 6848 12716 6860
rect 12483 6820 12716 6848
rect 12483 6817 12495 6820
rect 12437 6811 12495 6817
rect 12710 6808 12716 6820
rect 12768 6808 12774 6860
rect 13262 6808 13268 6860
rect 13320 6848 13326 6860
rect 13449 6851 13507 6857
rect 13449 6848 13461 6851
rect 13320 6820 13461 6848
rect 13320 6808 13326 6820
rect 13449 6817 13461 6820
rect 13495 6817 13507 6851
rect 13449 6811 13507 6817
rect 20346 6808 20352 6860
rect 20404 6848 20410 6860
rect 21269 6851 21327 6857
rect 21269 6848 21281 6851
rect 20404 6820 21281 6848
rect 20404 6808 20410 6820
rect 21269 6817 21281 6820
rect 21315 6848 21327 6851
rect 21358 6848 21364 6860
rect 21315 6820 21364 6848
rect 21315 6817 21327 6820
rect 21269 6811 21327 6817
rect 21358 6808 21364 6820
rect 21416 6808 21422 6860
rect 21744 6857 21772 6888
rect 22643 6885 22655 6888
rect 22689 6916 22701 6919
rect 22830 6916 22836 6928
rect 22689 6888 22836 6916
rect 22689 6885 22701 6888
rect 22643 6879 22701 6885
rect 22830 6876 22836 6888
rect 22888 6876 22894 6928
rect 21729 6851 21787 6857
rect 21729 6817 21741 6851
rect 21775 6817 21787 6851
rect 21729 6811 21787 6817
rect 21818 6808 21824 6860
rect 21876 6848 21882 6860
rect 22281 6851 22339 6857
rect 22281 6848 22293 6851
rect 21876 6820 22293 6848
rect 21876 6808 21882 6820
rect 22281 6817 22293 6820
rect 22327 6848 22339 6851
rect 22462 6848 22468 6860
rect 22327 6820 22468 6848
rect 22327 6817 22339 6820
rect 22281 6811 22339 6817
rect 22462 6808 22468 6820
rect 22520 6808 22526 6860
rect 23201 6851 23259 6857
rect 23201 6817 23213 6851
rect 23247 6848 23259 6851
rect 23952 6848 23980 6956
rect 24762 6944 24768 6956
rect 24820 6944 24826 6996
rect 25225 6987 25283 6993
rect 25225 6984 25237 6987
rect 24872 6956 25237 6984
rect 24210 6916 24216 6928
rect 24171 6888 24216 6916
rect 24210 6876 24216 6888
rect 24268 6876 24274 6928
rect 24394 6876 24400 6928
rect 24452 6916 24458 6928
rect 24872 6916 24900 6956
rect 25225 6953 25237 6956
rect 25271 6984 25283 6987
rect 25314 6984 25320 6996
rect 25271 6956 25320 6984
rect 25271 6953 25283 6956
rect 25225 6947 25283 6953
rect 25314 6944 25320 6956
rect 25372 6944 25378 6996
rect 25590 6984 25596 6996
rect 25551 6956 25596 6984
rect 25590 6944 25596 6956
rect 25648 6944 25654 6996
rect 27617 6987 27675 6993
rect 27617 6953 27629 6987
rect 27663 6984 27675 6987
rect 28442 6984 28448 6996
rect 27663 6956 28448 6984
rect 27663 6953 27675 6956
rect 27617 6947 27675 6953
rect 28442 6944 28448 6956
rect 28500 6944 28506 6996
rect 30650 6984 30656 6996
rect 30611 6956 30656 6984
rect 30650 6944 30656 6956
rect 30708 6944 30714 6996
rect 31205 6987 31263 6993
rect 31205 6953 31217 6987
rect 31251 6984 31263 6987
rect 33962 6984 33968 6996
rect 31251 6956 33968 6984
rect 31251 6953 31263 6956
rect 31205 6947 31263 6953
rect 33962 6944 33968 6956
rect 34020 6944 34026 6996
rect 34146 6984 34152 6996
rect 34107 6956 34152 6984
rect 34146 6944 34152 6956
rect 34204 6944 34210 6996
rect 34974 6944 34980 6996
rect 35032 6984 35038 6996
rect 35253 6987 35311 6993
rect 35253 6984 35265 6987
rect 35032 6956 35265 6984
rect 35032 6944 35038 6956
rect 35253 6953 35265 6956
rect 35299 6953 35311 6987
rect 35253 6947 35311 6953
rect 24452 6888 24900 6916
rect 24452 6876 24458 6888
rect 24946 6876 24952 6928
rect 25004 6916 25010 6928
rect 26602 6916 26608 6928
rect 25004 6888 26608 6916
rect 25004 6876 25010 6888
rect 26602 6876 26608 6888
rect 26660 6876 26666 6928
rect 26697 6919 26755 6925
rect 26697 6885 26709 6919
rect 26743 6916 26755 6919
rect 26786 6916 26792 6928
rect 26743 6888 26792 6916
rect 26743 6885 26755 6888
rect 26697 6879 26755 6885
rect 26786 6876 26792 6888
rect 26844 6876 26850 6928
rect 28902 6916 28908 6928
rect 28863 6888 28908 6916
rect 28902 6876 28908 6888
rect 28960 6876 28966 6928
rect 32490 6925 32496 6928
rect 32487 6916 32496 6925
rect 32451 6888 32496 6916
rect 32487 6879 32496 6888
rect 32490 6876 32496 6879
rect 32548 6876 32554 6928
rect 32674 6876 32680 6928
rect 32732 6916 32738 6928
rect 34054 6916 34060 6928
rect 32732 6888 34060 6916
rect 32732 6876 32738 6888
rect 34054 6876 34060 6888
rect 34112 6916 34118 6928
rect 34425 6919 34483 6925
rect 34425 6916 34437 6919
rect 34112 6888 34437 6916
rect 34112 6876 34118 6888
rect 34425 6885 34437 6888
rect 34471 6885 34483 6919
rect 34425 6879 34483 6885
rect 35066 6876 35072 6928
rect 35124 6916 35130 6928
rect 35894 6916 35900 6928
rect 35124 6888 35900 6916
rect 35124 6876 35130 6888
rect 35894 6876 35900 6888
rect 35952 6916 35958 6928
rect 35989 6919 36047 6925
rect 35989 6916 36001 6919
rect 35952 6888 36001 6916
rect 35952 6876 35958 6888
rect 35989 6885 36001 6888
rect 36035 6885 36047 6919
rect 35989 6879 36047 6885
rect 36262 6876 36268 6928
rect 36320 6916 36326 6928
rect 36541 6919 36599 6925
rect 36541 6916 36553 6919
rect 36320 6888 36553 6916
rect 36320 6876 36326 6888
rect 36541 6885 36553 6888
rect 36587 6885 36599 6919
rect 36541 6879 36599 6885
rect 23247 6820 23980 6848
rect 23247 6817 23259 6820
rect 23201 6811 23259 6817
rect 29822 6808 29828 6860
rect 29880 6848 29886 6860
rect 30285 6851 30343 6857
rect 30285 6848 30297 6851
rect 29880 6820 30297 6848
rect 29880 6808 29886 6820
rect 30285 6817 30297 6820
rect 30331 6848 30343 6851
rect 31110 6848 31116 6860
rect 30331 6820 31116 6848
rect 30331 6817 30343 6820
rect 30285 6811 30343 6817
rect 31110 6808 31116 6820
rect 31168 6808 31174 6860
rect 31938 6808 31944 6860
rect 31996 6848 32002 6860
rect 32125 6851 32183 6857
rect 32125 6848 32137 6851
rect 31996 6820 32137 6848
rect 31996 6808 32002 6820
rect 32125 6817 32137 6820
rect 32171 6817 32183 6851
rect 32125 6811 32183 6817
rect 4157 6783 4215 6789
rect 4157 6749 4169 6783
rect 4203 6749 4215 6783
rect 4157 6743 4215 6749
rect 5721 6783 5779 6789
rect 5721 6749 5733 6783
rect 5767 6749 5779 6783
rect 5994 6780 6000 6792
rect 5955 6752 6000 6780
rect 5721 6743 5779 6749
rect 4172 6712 4200 6743
rect 3988 6684 4200 6712
rect 5626 6644 5632 6656
rect 3896 6616 5632 6644
rect 5626 6604 5632 6616
rect 5684 6644 5690 6656
rect 5736 6644 5764 6743
rect 5994 6740 6000 6752
rect 6052 6740 6058 6792
rect 8110 6740 8116 6792
rect 8168 6780 8174 6792
rect 8389 6783 8447 6789
rect 8389 6780 8401 6783
rect 8168 6752 8401 6780
rect 8168 6740 8174 6752
rect 8389 6749 8401 6752
rect 8435 6780 8447 6783
rect 10689 6783 10747 6789
rect 10689 6780 10701 6783
rect 8435 6752 10701 6780
rect 8435 6749 8447 6752
rect 8389 6743 8447 6749
rect 10689 6749 10701 6752
rect 10735 6780 10747 6783
rect 11790 6780 11796 6792
rect 10735 6752 11796 6780
rect 10735 6749 10747 6752
rect 10689 6743 10747 6749
rect 11790 6740 11796 6752
rect 11848 6740 11854 6792
rect 14182 6740 14188 6792
rect 14240 6780 14246 6792
rect 14918 6780 14924 6792
rect 14240 6752 14924 6780
rect 14240 6740 14246 6752
rect 14918 6740 14924 6752
rect 14976 6740 14982 6792
rect 17126 6780 17132 6792
rect 15488 6752 17132 6780
rect 7929 6715 7987 6721
rect 7929 6681 7941 6715
rect 7975 6712 7987 6715
rect 8202 6712 8208 6724
rect 7975 6684 8208 6712
rect 7975 6681 7987 6684
rect 7929 6675 7987 6681
rect 8202 6672 8208 6684
rect 8260 6672 8266 6724
rect 14369 6715 14427 6721
rect 14369 6681 14381 6715
rect 14415 6712 14427 6715
rect 15488 6712 15516 6752
rect 17126 6740 17132 6752
rect 17184 6740 17190 6792
rect 17313 6783 17371 6789
rect 17313 6749 17325 6783
rect 17359 6749 17371 6783
rect 18598 6780 18604 6792
rect 18559 6752 18604 6780
rect 17313 6743 17371 6749
rect 14415 6684 15516 6712
rect 15933 6715 15991 6721
rect 14415 6681 14427 6684
rect 14369 6675 14427 6681
rect 15933 6681 15945 6715
rect 15979 6712 15991 6715
rect 17328 6712 17356 6743
rect 18598 6740 18604 6752
rect 18656 6740 18662 6792
rect 18874 6780 18880 6792
rect 18835 6752 18880 6780
rect 18874 6740 18880 6752
rect 18932 6740 18938 6792
rect 24121 6783 24179 6789
rect 24121 6749 24133 6783
rect 24167 6780 24179 6783
rect 24302 6780 24308 6792
rect 24167 6752 24308 6780
rect 24167 6749 24179 6752
rect 24121 6743 24179 6749
rect 24302 6740 24308 6752
rect 24360 6740 24366 6792
rect 24762 6780 24768 6792
rect 24723 6752 24768 6780
rect 24762 6740 24768 6752
rect 24820 6740 24826 6792
rect 26694 6740 26700 6792
rect 26752 6780 26758 6792
rect 26881 6783 26939 6789
rect 26881 6780 26893 6783
rect 26752 6752 26893 6780
rect 26752 6740 26758 6752
rect 26881 6749 26893 6752
rect 26927 6749 26939 6783
rect 26881 6743 26939 6749
rect 28626 6740 28632 6792
rect 28684 6780 28690 6792
rect 28813 6783 28871 6789
rect 28813 6780 28825 6783
rect 28684 6752 28825 6780
rect 28684 6740 28690 6752
rect 28813 6749 28825 6752
rect 28859 6749 28871 6783
rect 28813 6743 28871 6749
rect 29457 6783 29515 6789
rect 29457 6749 29469 6783
rect 29503 6780 29515 6783
rect 29638 6780 29644 6792
rect 29503 6752 29644 6780
rect 29503 6749 29515 6752
rect 29457 6743 29515 6749
rect 29638 6740 29644 6752
rect 29696 6740 29702 6792
rect 34333 6783 34391 6789
rect 34333 6749 34345 6783
rect 34379 6749 34391 6783
rect 34333 6743 34391 6749
rect 34977 6783 35035 6789
rect 34977 6749 34989 6783
rect 35023 6780 35035 6783
rect 35342 6780 35348 6792
rect 35023 6752 35348 6780
rect 35023 6749 35035 6752
rect 34977 6743 35035 6749
rect 17954 6712 17960 6724
rect 15979 6684 17960 6712
rect 15979 6681 15991 6684
rect 15933 6675 15991 6681
rect 17954 6672 17960 6684
rect 18012 6712 18018 6724
rect 21407 6715 21465 6721
rect 18012 6684 18368 6712
rect 18012 6672 18018 6684
rect 5684 6616 5764 6644
rect 5684 6604 5690 6616
rect 7190 6604 7196 6656
rect 7248 6644 7254 6656
rect 7285 6647 7343 6653
rect 7285 6644 7297 6647
rect 7248 6616 7297 6644
rect 7248 6604 7254 6616
rect 7285 6613 7297 6616
rect 7331 6613 7343 6647
rect 7285 6607 7343 6613
rect 12802 6604 12808 6656
rect 12860 6644 12866 6656
rect 12897 6647 12955 6653
rect 12897 6644 12909 6647
rect 12860 6616 12909 6644
rect 12860 6604 12866 6616
rect 12897 6613 12909 6616
rect 12943 6613 12955 6647
rect 12897 6607 12955 6613
rect 16206 6604 16212 6656
rect 16264 6644 16270 6656
rect 16301 6647 16359 6653
rect 16301 6644 16313 6647
rect 16264 6616 16313 6644
rect 16264 6604 16270 6616
rect 16301 6613 16313 6616
rect 16347 6613 16359 6647
rect 16301 6607 16359 6613
rect 18141 6647 18199 6653
rect 18141 6613 18153 6647
rect 18187 6644 18199 6647
rect 18230 6644 18236 6656
rect 18187 6616 18236 6644
rect 18187 6613 18199 6616
rect 18141 6607 18199 6613
rect 18230 6604 18236 6616
rect 18288 6604 18294 6656
rect 18340 6644 18368 6684
rect 21407 6681 21419 6715
rect 21453 6712 21465 6715
rect 24394 6712 24400 6724
rect 21453 6684 24400 6712
rect 21453 6681 21465 6684
rect 21407 6675 21465 6681
rect 24394 6672 24400 6684
rect 24452 6672 24458 6724
rect 34348 6712 34376 6743
rect 35342 6740 35348 6752
rect 35400 6740 35406 6792
rect 35897 6783 35955 6789
rect 35897 6749 35909 6783
rect 35943 6780 35955 6783
rect 36354 6780 36360 6792
rect 35943 6752 36360 6780
rect 35943 6749 35955 6752
rect 35897 6743 35955 6749
rect 36354 6740 36360 6752
rect 36412 6780 36418 6792
rect 37090 6780 37096 6792
rect 36412 6752 37096 6780
rect 36412 6740 36418 6752
rect 37090 6740 37096 6752
rect 37148 6740 37154 6792
rect 34882 6712 34888 6724
rect 34348 6684 34888 6712
rect 34882 6672 34888 6684
rect 34940 6712 34946 6724
rect 36262 6712 36268 6724
rect 34940 6684 36268 6712
rect 34940 6672 34946 6684
rect 36262 6672 36268 6684
rect 36320 6672 36326 6724
rect 19521 6647 19579 6653
rect 19521 6644 19533 6647
rect 18340 6616 19533 6644
rect 19521 6613 19533 6616
rect 19567 6613 19579 6647
rect 30190 6644 30196 6656
rect 30151 6616 30196 6644
rect 19521 6607 19579 6613
rect 30190 6604 30196 6616
rect 30248 6604 30254 6656
rect 30466 6604 30472 6656
rect 30524 6644 30530 6656
rect 31754 6644 31760 6656
rect 30524 6616 31760 6644
rect 30524 6604 30530 6616
rect 31754 6604 31760 6616
rect 31812 6604 31818 6656
rect 33045 6647 33103 6653
rect 33045 6613 33057 6647
rect 33091 6644 33103 6647
rect 34606 6644 34612 6656
rect 33091 6616 34612 6644
rect 33091 6613 33103 6616
rect 33045 6607 33103 6613
rect 34606 6604 34612 6616
rect 34664 6604 34670 6656
rect 1104 6554 38824 6576
rect 1104 6502 7648 6554
rect 7700 6502 7712 6554
rect 7764 6502 7776 6554
rect 7828 6502 7840 6554
rect 7892 6502 20982 6554
rect 21034 6502 21046 6554
rect 21098 6502 21110 6554
rect 21162 6502 21174 6554
rect 21226 6502 34315 6554
rect 34367 6502 34379 6554
rect 34431 6502 34443 6554
rect 34495 6502 34507 6554
rect 34559 6502 38824 6554
rect 1104 6480 38824 6502
rect 1854 6440 1860 6452
rect 1815 6412 1860 6440
rect 1854 6400 1860 6412
rect 1912 6400 1918 6452
rect 2498 6400 2504 6452
rect 2556 6440 2562 6452
rect 3786 6440 3792 6452
rect 2556 6412 3792 6440
rect 2556 6400 2562 6412
rect 3786 6400 3792 6412
rect 3844 6400 3850 6452
rect 5629 6443 5687 6449
rect 5629 6409 5641 6443
rect 5675 6440 5687 6443
rect 5902 6440 5908 6452
rect 5675 6412 5908 6440
rect 5675 6409 5687 6412
rect 5629 6403 5687 6409
rect 5902 6400 5908 6412
rect 5960 6400 5966 6452
rect 6273 6443 6331 6449
rect 6273 6409 6285 6443
rect 6319 6440 6331 6443
rect 6362 6440 6368 6452
rect 6319 6412 6368 6440
rect 6319 6409 6331 6412
rect 6273 6403 6331 6409
rect 2317 6375 2375 6381
rect 2317 6341 2329 6375
rect 2363 6372 2375 6375
rect 2590 6372 2596 6384
rect 2363 6344 2596 6372
rect 2363 6341 2375 6344
rect 2317 6335 2375 6341
rect 1448 6239 1506 6245
rect 1448 6205 1460 6239
rect 1494 6236 1506 6239
rect 2332 6236 2360 6335
rect 2590 6332 2596 6344
rect 2648 6332 2654 6384
rect 3050 6372 3056 6384
rect 3011 6344 3056 6372
rect 3050 6332 3056 6344
rect 3108 6332 3114 6384
rect 6288 6372 6316 6403
rect 6362 6400 6368 6412
rect 6420 6400 6426 6452
rect 8018 6400 8024 6452
rect 8076 6440 8082 6452
rect 8849 6443 8907 6449
rect 8849 6440 8861 6443
rect 8076 6412 8861 6440
rect 8076 6400 8082 6412
rect 8849 6409 8861 6412
rect 8895 6409 8907 6443
rect 8849 6403 8907 6409
rect 11609 6443 11667 6449
rect 11609 6409 11621 6443
rect 11655 6440 11667 6443
rect 11698 6440 11704 6452
rect 11655 6412 11704 6440
rect 11655 6409 11667 6412
rect 11609 6403 11667 6409
rect 11698 6400 11704 6412
rect 11756 6400 11762 6452
rect 13262 6400 13268 6452
rect 13320 6440 13326 6452
rect 13817 6443 13875 6449
rect 13817 6440 13829 6443
rect 13320 6412 13829 6440
rect 13320 6400 13326 6412
rect 13817 6409 13829 6412
rect 13863 6409 13875 6443
rect 13817 6403 13875 6409
rect 15381 6443 15439 6449
rect 15381 6409 15393 6443
rect 15427 6440 15439 6443
rect 15746 6440 15752 6452
rect 15427 6412 15752 6440
rect 15427 6409 15439 6412
rect 15381 6403 15439 6409
rect 15746 6400 15752 6412
rect 15804 6400 15810 6452
rect 17218 6400 17224 6452
rect 17276 6440 17282 6452
rect 17773 6443 17831 6449
rect 17773 6440 17785 6443
rect 17276 6412 17785 6440
rect 17276 6400 17282 6412
rect 17773 6409 17785 6412
rect 17819 6440 17831 6443
rect 19061 6443 19119 6449
rect 19061 6440 19073 6443
rect 17819 6412 19073 6440
rect 17819 6409 17831 6412
rect 17773 6403 17831 6409
rect 19061 6409 19073 6412
rect 19107 6409 19119 6443
rect 19061 6403 19119 6409
rect 19705 6443 19763 6449
rect 19705 6409 19717 6443
rect 19751 6440 19763 6443
rect 19794 6440 19800 6452
rect 19751 6412 19800 6440
rect 19751 6409 19763 6412
rect 19705 6403 19763 6409
rect 19794 6400 19800 6412
rect 19852 6440 19858 6452
rect 20162 6440 20168 6452
rect 19852 6412 20168 6440
rect 19852 6400 19858 6412
rect 20162 6400 20168 6412
rect 20220 6400 20226 6452
rect 22649 6443 22707 6449
rect 22649 6409 22661 6443
rect 22695 6440 22707 6443
rect 24210 6440 24216 6452
rect 22695 6412 24216 6440
rect 22695 6409 22707 6412
rect 22649 6403 22707 6409
rect 24210 6400 24216 6412
rect 24268 6440 24274 6452
rect 24673 6443 24731 6449
rect 24673 6440 24685 6443
rect 24268 6412 24685 6440
rect 24268 6400 24274 6412
rect 24673 6409 24685 6412
rect 24719 6440 24731 6443
rect 25041 6443 25099 6449
rect 25041 6440 25053 6443
rect 24719 6412 25053 6440
rect 24719 6409 24731 6412
rect 24673 6403 24731 6409
rect 25041 6409 25053 6412
rect 25087 6440 25099 6443
rect 25087 6412 25176 6440
rect 25087 6409 25099 6412
rect 25041 6403 25099 6409
rect 15654 6372 15660 6384
rect 5803 6344 6316 6372
rect 15615 6344 15660 6372
rect 2501 6307 2559 6313
rect 2501 6273 2513 6307
rect 2547 6304 2559 6307
rect 3418 6304 3424 6316
rect 2547 6276 3424 6304
rect 2547 6273 2559 6276
rect 2501 6267 2559 6273
rect 3418 6264 3424 6276
rect 3476 6304 3482 6316
rect 4062 6304 4068 6316
rect 3476 6276 4068 6304
rect 3476 6264 3482 6276
rect 4062 6264 4068 6276
rect 4120 6264 4126 6316
rect 5258 6304 5264 6316
rect 4258 6276 5264 6304
rect 1494 6208 2360 6236
rect 3973 6239 4031 6245
rect 1494 6205 1506 6208
rect 1448 6199 1506 6205
rect 3973 6205 3985 6239
rect 4019 6236 4031 6239
rect 4258 6236 4286 6276
rect 5258 6264 5264 6276
rect 5316 6264 5322 6316
rect 4019 6208 4286 6236
rect 4019 6205 4031 6208
rect 3973 6199 4031 6205
rect 4706 6196 4712 6248
rect 4764 6236 4770 6248
rect 5803 6245 5831 6344
rect 15654 6332 15660 6344
rect 15712 6332 15718 6384
rect 17129 6375 17187 6381
rect 17129 6341 17141 6375
rect 17175 6372 17187 6375
rect 18230 6372 18236 6384
rect 17175 6344 18236 6372
rect 17175 6341 17187 6344
rect 17129 6335 17187 6341
rect 18230 6332 18236 6344
rect 18288 6332 18294 6384
rect 5859 6307 5917 6313
rect 5859 6273 5871 6307
rect 5905 6304 5917 6307
rect 10042 6304 10048 6316
rect 5905 6276 10048 6304
rect 5905 6273 5917 6276
rect 5859 6267 5917 6273
rect 10042 6264 10048 6276
rect 10100 6264 10106 6316
rect 17402 6304 17408 6316
rect 17363 6276 17408 6304
rect 17402 6264 17408 6276
rect 17460 6264 17466 6316
rect 17954 6264 17960 6316
rect 18012 6304 18018 6316
rect 18141 6307 18199 6313
rect 18141 6304 18153 6307
rect 18012 6276 18153 6304
rect 18012 6264 18018 6276
rect 18141 6273 18153 6276
rect 18187 6273 18199 6307
rect 18141 6267 18199 6273
rect 18506 6264 18512 6316
rect 18564 6304 18570 6316
rect 19334 6304 19340 6316
rect 18564 6276 19340 6304
rect 18564 6264 18570 6276
rect 19334 6264 19340 6276
rect 19392 6304 19398 6316
rect 19981 6307 20039 6313
rect 19981 6304 19993 6307
rect 19392 6276 19993 6304
rect 19392 6264 19398 6276
rect 19981 6273 19993 6276
rect 20027 6273 20039 6307
rect 20180 6304 20208 6400
rect 22830 6332 22836 6384
rect 22888 6372 22894 6384
rect 22925 6375 22983 6381
rect 22925 6372 22937 6375
rect 22888 6344 22937 6372
rect 22888 6332 22894 6344
rect 22925 6341 22937 6344
rect 22971 6341 22983 6375
rect 22925 6335 22983 6341
rect 23290 6332 23296 6384
rect 23348 6372 23354 6384
rect 24762 6372 24768 6384
rect 23348 6344 24768 6372
rect 23348 6332 23354 6344
rect 24762 6332 24768 6344
rect 24820 6332 24826 6384
rect 21726 6304 21732 6316
rect 20180 6276 20668 6304
rect 21687 6276 21732 6304
rect 19981 6267 20039 6273
rect 5772 6239 5831 6245
rect 5772 6236 5784 6239
rect 4764 6208 5784 6236
rect 4764 6196 4770 6208
rect 5772 6205 5784 6208
rect 5818 6208 5831 6239
rect 5818 6205 5830 6208
rect 5772 6199 5830 6205
rect 7190 6196 7196 6248
rect 7248 6236 7254 6248
rect 7285 6239 7343 6245
rect 7285 6236 7297 6239
rect 7248 6208 7297 6236
rect 7248 6196 7254 6208
rect 7285 6205 7297 6208
rect 7331 6205 7343 6239
rect 9769 6239 9827 6245
rect 9769 6236 9781 6239
rect 7285 6199 7343 6205
rect 9232 6208 9781 6236
rect 1535 6171 1593 6177
rect 1535 6137 1547 6171
rect 1581 6168 1593 6171
rect 2498 6168 2504 6180
rect 1581 6140 2504 6168
rect 1581 6137 1593 6140
rect 1535 6131 1593 6137
rect 2498 6128 2504 6140
rect 2556 6128 2562 6180
rect 2590 6128 2596 6180
rect 2648 6168 2654 6180
rect 3513 6171 3571 6177
rect 2648 6140 2693 6168
rect 2648 6128 2654 6140
rect 3513 6137 3525 6171
rect 3559 6168 3571 6171
rect 4335 6171 4393 6177
rect 3559 6140 4016 6168
rect 3559 6137 3571 6140
rect 3513 6131 3571 6137
rect 3988 6112 4016 6140
rect 4335 6137 4347 6171
rect 4381 6168 4393 6171
rect 4430 6168 4436 6180
rect 4381 6140 4436 6168
rect 4381 6137 4393 6140
rect 4335 6131 4393 6137
rect 4430 6128 4436 6140
rect 4488 6128 4494 6180
rect 7606 6171 7664 6177
rect 7606 6168 7618 6171
rect 7116 6140 7618 6168
rect 7116 6112 7144 6140
rect 7606 6137 7618 6140
rect 7652 6137 7664 6171
rect 7606 6131 7664 6137
rect 9232 6112 9260 6208
rect 9769 6205 9781 6208
rect 9815 6205 9827 6239
rect 9769 6199 9827 6205
rect 12713 6239 12771 6245
rect 12713 6205 12725 6239
rect 12759 6236 12771 6239
rect 12802 6236 12808 6248
rect 12759 6208 12808 6236
rect 12759 6205 12771 6208
rect 12713 6199 12771 6205
rect 9306 6128 9312 6180
rect 9364 6168 9370 6180
rect 9677 6171 9735 6177
rect 9677 6168 9689 6171
rect 9364 6140 9689 6168
rect 9364 6128 9370 6140
rect 9677 6137 9689 6140
rect 9723 6168 9735 6171
rect 10131 6171 10189 6177
rect 10131 6168 10143 6171
rect 9723 6140 10143 6168
rect 9723 6137 9735 6140
rect 9677 6131 9735 6137
rect 10131 6137 10143 6140
rect 10177 6168 10189 6171
rect 10226 6168 10232 6180
rect 10177 6140 10232 6168
rect 10177 6137 10189 6140
rect 10131 6131 10189 6137
rect 10226 6128 10232 6140
rect 10284 6128 10290 6180
rect 3326 6060 3332 6112
rect 3384 6100 3390 6112
rect 3878 6100 3884 6112
rect 3384 6072 3884 6100
rect 3384 6060 3390 6072
rect 3878 6060 3884 6072
rect 3936 6060 3942 6112
rect 3970 6060 3976 6112
rect 4028 6100 4034 6112
rect 4893 6103 4951 6109
rect 4893 6100 4905 6103
rect 4028 6072 4905 6100
rect 4028 6060 4034 6072
rect 4893 6069 4905 6072
rect 4939 6069 4951 6103
rect 5258 6100 5264 6112
rect 5219 6072 5264 6100
rect 4893 6063 4951 6069
rect 5258 6060 5264 6072
rect 5316 6060 5322 6112
rect 7098 6100 7104 6112
rect 7059 6072 7104 6100
rect 7098 6060 7104 6072
rect 7156 6060 7162 6112
rect 8205 6103 8263 6109
rect 8205 6069 8217 6103
rect 8251 6100 8263 6103
rect 8386 6100 8392 6112
rect 8251 6072 8392 6100
rect 8251 6069 8263 6072
rect 8205 6063 8263 6069
rect 8386 6060 8392 6072
rect 8444 6100 8450 6112
rect 8481 6103 8539 6109
rect 8481 6100 8493 6103
rect 8444 6072 8493 6100
rect 8444 6060 8450 6072
rect 8481 6069 8493 6072
rect 8527 6069 8539 6103
rect 9214 6100 9220 6112
rect 9175 6072 9220 6100
rect 8481 6063 8539 6069
rect 9214 6060 9220 6072
rect 9272 6060 9278 6112
rect 10686 6100 10692 6112
rect 10647 6072 10692 6100
rect 10686 6060 10692 6072
rect 10744 6100 10750 6112
rect 10965 6103 11023 6109
rect 10965 6100 10977 6103
rect 10744 6072 10977 6100
rect 10744 6060 10750 6072
rect 10965 6069 10977 6072
rect 11011 6069 11023 6103
rect 11974 6100 11980 6112
rect 11935 6072 11980 6100
rect 10965 6063 11023 6069
rect 11974 6060 11980 6072
rect 12032 6060 12038 6112
rect 12526 6100 12532 6112
rect 12487 6072 12532 6100
rect 12526 6060 12532 6072
rect 12584 6060 12590 6112
rect 12728 6100 12756 6199
rect 12802 6196 12808 6208
rect 12860 6196 12866 6248
rect 12986 6236 12992 6248
rect 12947 6208 12992 6236
rect 12986 6196 12992 6208
rect 13044 6196 13050 6248
rect 14461 6239 14519 6245
rect 14461 6205 14473 6239
rect 14507 6236 14519 6239
rect 14642 6236 14648 6248
rect 14507 6208 14648 6236
rect 14507 6205 14519 6208
rect 14461 6199 14519 6205
rect 14642 6196 14648 6208
rect 14700 6196 14706 6248
rect 16206 6236 16212 6248
rect 16167 6208 16212 6236
rect 16206 6196 16212 6208
rect 16264 6196 16270 6248
rect 19996 6236 20024 6267
rect 20162 6236 20168 6248
rect 19996 6208 20168 6236
rect 20162 6196 20168 6208
rect 20220 6196 20226 6248
rect 20640 6245 20668 6276
rect 21726 6264 21732 6276
rect 21784 6264 21790 6316
rect 23753 6307 23811 6313
rect 23753 6304 23765 6307
rect 23584 6276 23765 6304
rect 20625 6239 20683 6245
rect 20625 6205 20637 6239
rect 20671 6205 20683 6239
rect 20625 6199 20683 6205
rect 22370 6196 22376 6248
rect 22428 6236 22434 6248
rect 23385 6239 23443 6245
rect 23385 6236 23397 6239
rect 22428 6208 23397 6236
rect 22428 6196 22434 6208
rect 14369 6171 14427 6177
rect 14369 6168 14381 6171
rect 13786 6140 14381 6168
rect 13078 6100 13084 6112
rect 12728 6072 13084 6100
rect 13078 6060 13084 6072
rect 13136 6060 13142 6112
rect 13170 6060 13176 6112
rect 13228 6100 13234 6112
rect 13449 6103 13507 6109
rect 13449 6100 13461 6103
rect 13228 6072 13461 6100
rect 13228 6060 13234 6072
rect 13449 6069 13461 6072
rect 13495 6100 13507 6103
rect 13786 6100 13814 6140
rect 14369 6137 14381 6140
rect 14415 6168 14427 6171
rect 14823 6171 14881 6177
rect 14823 6168 14835 6171
rect 14415 6140 14835 6168
rect 14415 6137 14427 6140
rect 14369 6131 14427 6137
rect 14823 6137 14835 6140
rect 14869 6168 14881 6171
rect 16022 6168 16028 6180
rect 14869 6140 16028 6168
rect 14869 6137 14881 6140
rect 14823 6131 14881 6137
rect 16022 6128 16028 6140
rect 16080 6168 16086 6180
rect 16117 6171 16175 6177
rect 16117 6168 16129 6171
rect 16080 6140 16129 6168
rect 16080 6128 16086 6140
rect 16117 6137 16129 6140
rect 16163 6168 16175 6171
rect 16571 6171 16629 6177
rect 16571 6168 16583 6171
rect 16163 6140 16583 6168
rect 16163 6137 16175 6140
rect 16117 6131 16175 6137
rect 16571 6137 16583 6140
rect 16617 6168 16629 6171
rect 17034 6168 17040 6180
rect 16617 6140 17040 6168
rect 16617 6137 16629 6140
rect 16571 6131 16629 6137
rect 17034 6128 17040 6140
rect 17092 6128 17098 6180
rect 18230 6128 18236 6180
rect 18288 6168 18294 6180
rect 18785 6171 18843 6177
rect 18288 6140 18333 6168
rect 18288 6128 18294 6140
rect 18785 6137 18797 6171
rect 18831 6137 18843 6171
rect 18785 6131 18843 6137
rect 20901 6171 20959 6177
rect 20901 6137 20913 6171
rect 20947 6168 20959 6171
rect 21450 6168 21456 6180
rect 20947 6140 21456 6168
rect 20947 6137 20959 6140
rect 20901 6131 20959 6137
rect 13495 6072 13814 6100
rect 13495 6069 13507 6072
rect 13449 6063 13507 6069
rect 17310 6060 17316 6112
rect 17368 6100 17374 6112
rect 18800 6100 18828 6131
rect 21450 6128 21456 6140
rect 21508 6128 21514 6180
rect 21910 6128 21916 6180
rect 21968 6168 21974 6180
rect 22091 6171 22149 6177
rect 22091 6168 22103 6171
rect 21968 6140 22103 6168
rect 21968 6128 21974 6140
rect 22091 6137 22103 6140
rect 22137 6168 22149 6171
rect 22830 6168 22836 6180
rect 22137 6140 22836 6168
rect 22137 6137 22149 6140
rect 22091 6131 22149 6137
rect 22830 6128 22836 6140
rect 22888 6128 22894 6180
rect 21358 6100 21364 6112
rect 17368 6072 18828 6100
rect 21271 6072 21364 6100
rect 17368 6060 17374 6072
rect 21358 6060 21364 6072
rect 21416 6100 21422 6112
rect 21818 6100 21824 6112
rect 21416 6072 21824 6100
rect 21416 6060 21422 6072
rect 21818 6060 21824 6072
rect 21876 6060 21882 6112
rect 23032 6100 23060 6208
rect 23385 6205 23397 6208
rect 23431 6205 23443 6239
rect 23385 6199 23443 6205
rect 23106 6128 23112 6180
rect 23164 6168 23170 6180
rect 23584 6168 23612 6276
rect 23753 6273 23765 6276
rect 23799 6304 23811 6307
rect 23799 6276 24992 6304
rect 23799 6273 23811 6276
rect 23753 6267 23811 6273
rect 23164 6140 23612 6168
rect 23845 6171 23903 6177
rect 23164 6128 23170 6140
rect 23845 6137 23857 6171
rect 23891 6137 23903 6171
rect 24394 6168 24400 6180
rect 24355 6140 24400 6168
rect 23845 6131 23903 6137
rect 23860 6100 23888 6131
rect 24394 6128 24400 6140
rect 24452 6128 24458 6180
rect 23032 6072 23888 6100
rect 24964 6100 24992 6276
rect 25148 6168 25176 6412
rect 26602 6400 26608 6452
rect 26660 6440 26666 6452
rect 26881 6443 26939 6449
rect 26881 6440 26893 6443
rect 26660 6412 26893 6440
rect 26660 6400 26666 6412
rect 26881 6409 26893 6412
rect 26927 6409 26939 6443
rect 27338 6440 27344 6452
rect 27299 6412 27344 6440
rect 26881 6403 26939 6409
rect 27338 6400 27344 6412
rect 27396 6400 27402 6452
rect 28813 6443 28871 6449
rect 28813 6409 28825 6443
rect 28859 6440 28871 6443
rect 28902 6440 28908 6452
rect 28859 6412 28908 6440
rect 28859 6409 28871 6412
rect 28813 6403 28871 6409
rect 28902 6400 28908 6412
rect 28960 6400 28966 6452
rect 29454 6440 29460 6452
rect 29415 6412 29460 6440
rect 29454 6400 29460 6412
rect 29512 6400 29518 6452
rect 31938 6400 31944 6452
rect 31996 6440 32002 6452
rect 33321 6443 33379 6449
rect 33321 6440 33333 6443
rect 31996 6412 33333 6440
rect 31996 6400 32002 6412
rect 33321 6409 33333 6412
rect 33367 6409 33379 6443
rect 33321 6403 33379 6409
rect 34054 6400 34060 6452
rect 34112 6440 34118 6452
rect 34241 6443 34299 6449
rect 34241 6440 34253 6443
rect 34112 6412 34253 6440
rect 34112 6400 34118 6412
rect 34241 6409 34253 6412
rect 34287 6409 34299 6443
rect 34606 6440 34612 6452
rect 34567 6412 34612 6440
rect 34241 6403 34299 6409
rect 34606 6400 34612 6412
rect 34664 6400 34670 6452
rect 35894 6440 35900 6452
rect 35855 6412 35900 6440
rect 35894 6400 35900 6412
rect 35952 6400 35958 6452
rect 36354 6440 36360 6452
rect 36315 6412 36360 6440
rect 36354 6400 36360 6412
rect 36412 6400 36418 6452
rect 36998 6440 37004 6452
rect 36959 6412 37004 6440
rect 36998 6400 37004 6412
rect 37056 6400 37062 6452
rect 26513 6375 26571 6381
rect 26513 6341 26525 6375
rect 26559 6372 26571 6375
rect 26786 6372 26792 6384
rect 26559 6344 26792 6372
rect 26559 6341 26571 6344
rect 26513 6335 26571 6341
rect 26786 6332 26792 6344
rect 26844 6332 26850 6384
rect 30190 6332 30196 6384
rect 30248 6372 30254 6384
rect 36587 6375 36645 6381
rect 36587 6372 36599 6375
rect 30248 6344 36599 6372
rect 30248 6332 30254 6344
rect 25314 6304 25320 6316
rect 25275 6276 25320 6304
rect 25314 6264 25320 6276
rect 25372 6264 25378 6316
rect 25961 6307 26019 6313
rect 25961 6273 25973 6307
rect 26007 6304 26019 6307
rect 26694 6304 26700 6316
rect 26007 6276 26700 6304
rect 26007 6273 26019 6276
rect 25961 6267 26019 6273
rect 25409 6171 25467 6177
rect 25409 6168 25421 6171
rect 25148 6140 25421 6168
rect 25409 6137 25421 6140
rect 25455 6137 25467 6171
rect 25409 6131 25467 6137
rect 25976 6100 26004 6267
rect 26694 6264 26700 6276
rect 26752 6264 26758 6316
rect 28261 6307 28319 6313
rect 28261 6273 28273 6307
rect 28307 6304 28319 6307
rect 30466 6304 30472 6316
rect 28307 6276 30472 6304
rect 28307 6273 28319 6276
rect 28261 6267 28319 6273
rect 30466 6264 30472 6276
rect 30524 6264 30530 6316
rect 30668 6313 30696 6344
rect 36587 6341 36599 6344
rect 36633 6341 36645 6375
rect 36587 6335 36645 6341
rect 30653 6307 30711 6313
rect 30653 6273 30665 6307
rect 30699 6273 30711 6307
rect 30926 6304 30932 6316
rect 30887 6276 30932 6304
rect 30653 6267 30711 6273
rect 30926 6264 30932 6276
rect 30984 6264 30990 6316
rect 31846 6264 31852 6316
rect 31904 6304 31910 6316
rect 32125 6307 32183 6313
rect 32125 6304 32137 6307
rect 31904 6276 32137 6304
rect 31904 6264 31910 6276
rect 32125 6273 32137 6276
rect 32171 6304 32183 6307
rect 33689 6307 33747 6313
rect 33689 6304 33701 6307
rect 32171 6276 33701 6304
rect 32171 6273 32183 6276
rect 32125 6267 32183 6273
rect 33689 6273 33701 6276
rect 33735 6273 33747 6307
rect 33689 6267 33747 6273
rect 34977 6307 35035 6313
rect 34977 6273 34989 6307
rect 35023 6304 35035 6307
rect 35250 6304 35256 6316
rect 35023 6276 35256 6304
rect 35023 6273 35035 6276
rect 34977 6267 35035 6273
rect 35250 6264 35256 6276
rect 35308 6264 35314 6316
rect 35342 6264 35348 6316
rect 35400 6304 35406 6316
rect 35400 6276 35445 6304
rect 35400 6264 35406 6276
rect 27338 6196 27344 6248
rect 27396 6236 27402 6248
rect 27525 6239 27583 6245
rect 27525 6236 27537 6239
rect 27396 6208 27537 6236
rect 27396 6196 27402 6208
rect 27525 6205 27537 6208
rect 27571 6205 27583 6239
rect 27525 6199 27583 6205
rect 28077 6239 28135 6245
rect 28077 6205 28089 6239
rect 28123 6236 28135 6239
rect 28442 6236 28448 6248
rect 28123 6208 28448 6236
rect 28123 6205 28135 6208
rect 28077 6199 28135 6205
rect 28442 6196 28448 6208
rect 28500 6196 28506 6248
rect 29273 6239 29331 6245
rect 29273 6205 29285 6239
rect 29319 6236 29331 6239
rect 29733 6239 29791 6245
rect 29733 6236 29745 6239
rect 29319 6208 29745 6236
rect 29319 6205 29331 6208
rect 29273 6199 29331 6205
rect 29733 6205 29745 6208
rect 29779 6205 29791 6239
rect 29733 6199 29791 6205
rect 36516 6239 36574 6245
rect 36516 6205 36528 6239
rect 36562 6236 36574 6239
rect 36998 6236 37004 6248
rect 36562 6208 37004 6236
rect 36562 6205 36574 6208
rect 36516 6199 36574 6205
rect 27062 6128 27068 6180
rect 27120 6168 27126 6180
rect 28534 6168 28540 6180
rect 27120 6140 28540 6168
rect 27120 6128 27126 6140
rect 28534 6128 28540 6140
rect 28592 6168 28598 6180
rect 29288 6168 29316 6199
rect 36998 6196 37004 6208
rect 37056 6196 37062 6248
rect 30742 6168 30748 6180
rect 28592 6140 29316 6168
rect 30703 6140 30748 6168
rect 28592 6128 28598 6140
rect 30742 6128 30748 6140
rect 30800 6128 30806 6180
rect 32446 6171 32504 6177
rect 32446 6168 32458 6171
rect 31956 6140 32458 6168
rect 24964 6072 26004 6100
rect 29822 6060 29828 6112
rect 29880 6100 29886 6112
rect 30285 6103 30343 6109
rect 30285 6100 30297 6103
rect 29880 6072 30297 6100
rect 29880 6060 29886 6072
rect 30285 6069 30297 6072
rect 30331 6100 30343 6103
rect 30650 6100 30656 6112
rect 30331 6072 30656 6100
rect 30331 6069 30343 6072
rect 30285 6063 30343 6069
rect 30650 6060 30656 6072
rect 30708 6100 30714 6112
rect 31956 6109 31984 6140
rect 32446 6137 32458 6140
rect 32492 6137 32504 6171
rect 32446 6131 32504 6137
rect 35069 6171 35127 6177
rect 35069 6137 35081 6171
rect 35115 6137 35127 6171
rect 35069 6131 35127 6137
rect 31573 6103 31631 6109
rect 31573 6100 31585 6103
rect 30708 6072 31585 6100
rect 30708 6060 30714 6072
rect 31573 6069 31585 6072
rect 31619 6100 31631 6103
rect 31941 6103 31999 6109
rect 31941 6100 31953 6103
rect 31619 6072 31953 6100
rect 31619 6069 31631 6072
rect 31573 6063 31631 6069
rect 31941 6069 31953 6072
rect 31987 6069 31999 6103
rect 33042 6100 33048 6112
rect 33003 6072 33048 6100
rect 31941 6063 31999 6069
rect 33042 6060 33048 6072
rect 33100 6060 33106 6112
rect 34606 6060 34612 6112
rect 34664 6100 34670 6112
rect 35084 6100 35112 6131
rect 34664 6072 35112 6100
rect 34664 6060 34670 6072
rect 1104 6010 38824 6032
rect 1104 5958 14315 6010
rect 14367 5958 14379 6010
rect 14431 5958 14443 6010
rect 14495 5958 14507 6010
rect 14559 5958 27648 6010
rect 27700 5958 27712 6010
rect 27764 5958 27776 6010
rect 27828 5958 27840 6010
rect 27892 5958 38824 6010
rect 1104 5936 38824 5958
rect 3142 5896 3148 5908
rect 3103 5868 3148 5896
rect 3142 5856 3148 5868
rect 3200 5856 3206 5908
rect 3513 5899 3571 5905
rect 3513 5865 3525 5899
rect 3559 5896 3571 5899
rect 3786 5896 3792 5908
rect 3559 5868 3792 5896
rect 3559 5865 3571 5868
rect 3513 5859 3571 5865
rect 3786 5856 3792 5868
rect 3844 5896 3850 5908
rect 5626 5896 5632 5908
rect 3844 5868 4844 5896
rect 5587 5868 5632 5896
rect 3844 5856 3850 5868
rect 2406 5788 2412 5840
rect 2464 5828 2470 5840
rect 2546 5831 2604 5837
rect 2546 5828 2558 5831
rect 2464 5800 2558 5828
rect 2464 5788 2470 5800
rect 2546 5797 2558 5800
rect 2592 5797 2604 5831
rect 2546 5791 2604 5797
rect 3970 5788 3976 5840
rect 4028 5828 4034 5840
rect 4816 5837 4844 5868
rect 5626 5856 5632 5868
rect 5684 5856 5690 5908
rect 9953 5899 10011 5905
rect 9953 5865 9965 5899
rect 9999 5896 10011 5899
rect 10318 5896 10324 5908
rect 9999 5868 10324 5896
rect 9999 5865 10011 5868
rect 9953 5859 10011 5865
rect 10318 5856 10324 5868
rect 10376 5856 10382 5908
rect 11790 5896 11796 5908
rect 11751 5868 11796 5896
rect 11790 5856 11796 5868
rect 11848 5856 11854 5908
rect 15010 5896 15016 5908
rect 14971 5868 15016 5896
rect 15010 5856 15016 5868
rect 15068 5856 15074 5908
rect 15562 5856 15568 5908
rect 15620 5896 15626 5908
rect 15933 5899 15991 5905
rect 15933 5896 15945 5899
rect 15620 5868 15945 5896
rect 15620 5856 15626 5868
rect 15933 5865 15945 5868
rect 15979 5865 15991 5899
rect 17402 5896 17408 5908
rect 15933 5859 15991 5865
rect 16868 5868 17408 5896
rect 4249 5831 4307 5837
rect 4249 5828 4261 5831
rect 4028 5800 4261 5828
rect 4028 5788 4034 5800
rect 4249 5797 4261 5800
rect 4295 5797 4307 5831
rect 4249 5791 4307 5797
rect 4801 5831 4859 5837
rect 4801 5797 4813 5831
rect 4847 5828 4859 5831
rect 5994 5828 6000 5840
rect 4847 5800 6000 5828
rect 4847 5797 4859 5800
rect 4801 5791 4859 5797
rect 5994 5788 6000 5800
rect 6052 5788 6058 5840
rect 6638 5828 6644 5840
rect 6599 5800 6644 5828
rect 6638 5788 6644 5800
rect 6696 5788 6702 5840
rect 7193 5831 7251 5837
rect 7193 5797 7205 5831
rect 7239 5828 7251 5831
rect 8110 5828 8116 5840
rect 7239 5800 8116 5828
rect 7239 5797 7251 5800
rect 7193 5791 7251 5797
rect 8110 5788 8116 5800
rect 8168 5788 8174 5840
rect 8205 5831 8263 5837
rect 8205 5797 8217 5831
rect 8251 5828 8263 5831
rect 8386 5828 8392 5840
rect 8251 5800 8392 5828
rect 8251 5797 8263 5800
rect 8205 5791 8263 5797
rect 8386 5788 8392 5800
rect 8444 5788 8450 5840
rect 10134 5788 10140 5840
rect 10192 5828 10198 5840
rect 10597 5831 10655 5837
rect 10597 5828 10609 5831
rect 10192 5800 10609 5828
rect 10192 5788 10198 5800
rect 10597 5797 10609 5800
rect 10643 5828 10655 5831
rect 10686 5828 10692 5840
rect 10643 5800 10692 5828
rect 10643 5797 10655 5800
rect 10597 5791 10655 5797
rect 10686 5788 10692 5800
rect 10744 5788 10750 5840
rect 12158 5828 12164 5840
rect 12119 5800 12164 5828
rect 12158 5788 12164 5800
rect 12216 5788 12222 5840
rect 14369 5831 14427 5837
rect 14369 5797 14381 5831
rect 14415 5828 14427 5831
rect 16206 5828 16212 5840
rect 14415 5800 16212 5828
rect 14415 5797 14427 5800
rect 14369 5791 14427 5797
rect 16206 5788 16212 5800
rect 16264 5788 16270 5840
rect 16868 5837 16896 5868
rect 17402 5856 17408 5868
rect 17460 5856 17466 5908
rect 18046 5896 18052 5908
rect 18007 5868 18052 5896
rect 18046 5856 18052 5868
rect 18104 5896 18110 5908
rect 18506 5896 18512 5908
rect 18104 5868 18512 5896
rect 18104 5856 18110 5868
rect 18506 5856 18512 5868
rect 18564 5856 18570 5908
rect 18598 5856 18604 5908
rect 18656 5896 18662 5908
rect 18785 5899 18843 5905
rect 18785 5896 18797 5899
rect 18656 5868 18797 5896
rect 18656 5856 18662 5868
rect 18785 5865 18797 5868
rect 18831 5865 18843 5899
rect 22370 5896 22376 5908
rect 22331 5868 22376 5896
rect 18785 5859 18843 5865
rect 22370 5856 22376 5868
rect 22428 5856 22434 5908
rect 22462 5856 22468 5908
rect 22520 5896 22526 5908
rect 22649 5899 22707 5905
rect 22649 5896 22661 5899
rect 22520 5868 22661 5896
rect 22520 5856 22526 5868
rect 22649 5865 22661 5868
rect 22695 5865 22707 5899
rect 23106 5896 23112 5908
rect 23067 5868 23112 5896
rect 22649 5859 22707 5865
rect 23106 5856 23112 5868
rect 23164 5856 23170 5908
rect 24854 5896 24860 5908
rect 24815 5868 24860 5896
rect 24854 5856 24860 5868
rect 24912 5856 24918 5908
rect 29822 5856 29828 5908
rect 29880 5896 29886 5908
rect 29917 5899 29975 5905
rect 29917 5896 29929 5899
rect 29880 5868 29929 5896
rect 29880 5856 29886 5868
rect 29917 5865 29929 5868
rect 29963 5865 29975 5899
rect 31110 5896 31116 5908
rect 31071 5868 31116 5896
rect 29917 5859 29975 5865
rect 31110 5856 31116 5868
rect 31168 5856 31174 5908
rect 34882 5896 34888 5908
rect 34843 5868 34888 5896
rect 34882 5856 34888 5868
rect 34940 5856 34946 5908
rect 35250 5896 35256 5908
rect 35211 5868 35256 5896
rect 35250 5856 35256 5868
rect 35308 5856 35314 5908
rect 16853 5831 16911 5837
rect 16853 5797 16865 5831
rect 16899 5797 16911 5831
rect 16853 5791 16911 5797
rect 16945 5831 17003 5837
rect 16945 5797 16957 5831
rect 16991 5828 17003 5831
rect 17034 5828 17040 5840
rect 16991 5800 17040 5828
rect 16991 5797 17003 5800
rect 16945 5791 17003 5797
rect 17034 5788 17040 5800
rect 17092 5828 17098 5840
rect 18417 5831 18475 5837
rect 18417 5828 18429 5831
rect 17092 5800 18429 5828
rect 17092 5788 17098 5800
rect 18417 5797 18429 5800
rect 18463 5797 18475 5831
rect 18417 5791 18475 5797
rect 21815 5831 21873 5837
rect 21815 5797 21827 5831
rect 21861 5828 21873 5831
rect 21910 5828 21916 5840
rect 21861 5800 21916 5828
rect 21861 5797 21873 5800
rect 21815 5791 21873 5797
rect 21910 5788 21916 5800
rect 21968 5788 21974 5840
rect 23382 5828 23388 5840
rect 23343 5800 23388 5828
rect 23382 5788 23388 5800
rect 23440 5788 23446 5840
rect 25130 5828 25136 5840
rect 24780 5800 25136 5828
rect 24780 5772 24808 5800
rect 25130 5788 25136 5800
rect 25188 5788 25194 5840
rect 27246 5828 27252 5840
rect 27159 5800 27252 5828
rect 27246 5788 27252 5800
rect 27304 5828 27310 5840
rect 28902 5828 28908 5840
rect 27304 5800 28908 5828
rect 27304 5788 27310 5800
rect 28902 5788 28908 5800
rect 28960 5788 28966 5840
rect 30837 5831 30895 5837
rect 30837 5797 30849 5831
rect 30883 5828 30895 5831
rect 31938 5828 31944 5840
rect 30883 5800 31944 5828
rect 30883 5797 30895 5800
rect 30837 5791 30895 5797
rect 13906 5760 13912 5772
rect 13867 5732 13912 5760
rect 13906 5720 13912 5732
rect 13964 5720 13970 5772
rect 14090 5720 14096 5772
rect 14148 5760 14154 5772
rect 14185 5763 14243 5769
rect 14185 5760 14197 5763
rect 14148 5732 14197 5760
rect 14148 5720 14154 5732
rect 14185 5729 14197 5732
rect 14231 5760 14243 5763
rect 15470 5760 15476 5772
rect 14231 5732 15476 5760
rect 14231 5729 14243 5732
rect 14185 5723 14243 5729
rect 15470 5720 15476 5732
rect 15528 5720 15534 5772
rect 15562 5720 15568 5772
rect 15620 5760 15626 5772
rect 15749 5763 15807 5769
rect 15749 5760 15761 5763
rect 15620 5732 15761 5760
rect 15620 5720 15626 5732
rect 15749 5729 15761 5732
rect 15795 5729 15807 5763
rect 19242 5760 19248 5772
rect 19203 5732 19248 5760
rect 15749 5723 15807 5729
rect 19242 5720 19248 5732
rect 19300 5720 19306 5772
rect 19794 5760 19800 5772
rect 19755 5732 19800 5760
rect 19794 5720 19800 5732
rect 19852 5720 19858 5772
rect 24762 5760 24768 5772
rect 24723 5732 24768 5760
rect 24762 5720 24768 5732
rect 24820 5720 24826 5772
rect 25222 5760 25228 5772
rect 25183 5732 25228 5760
rect 25222 5720 25228 5732
rect 25280 5720 25286 5772
rect 30469 5763 30527 5769
rect 30469 5729 30481 5763
rect 30515 5760 30527 5763
rect 30742 5760 30748 5772
rect 30515 5732 30748 5760
rect 30515 5729 30527 5732
rect 30469 5723 30527 5729
rect 30742 5720 30748 5732
rect 30800 5760 30806 5772
rect 30852 5760 30880 5791
rect 31938 5788 31944 5800
rect 31996 5828 32002 5840
rect 32309 5831 32367 5837
rect 32309 5828 32321 5831
rect 31996 5800 32321 5828
rect 31996 5788 32002 5800
rect 32309 5797 32321 5800
rect 32355 5797 32367 5831
rect 32309 5791 32367 5797
rect 33042 5788 33048 5840
rect 33100 5828 33106 5840
rect 33962 5828 33968 5840
rect 33100 5800 33968 5828
rect 33100 5788 33106 5800
rect 33962 5788 33968 5800
rect 34020 5788 34026 5840
rect 34517 5831 34575 5837
rect 34517 5797 34529 5831
rect 34563 5828 34575 5831
rect 35342 5828 35348 5840
rect 34563 5800 35348 5828
rect 34563 5797 34575 5800
rect 34517 5791 34575 5797
rect 35342 5788 35348 5800
rect 35400 5788 35406 5840
rect 30800 5732 30880 5760
rect 30800 5720 30806 5732
rect 2222 5692 2228 5704
rect 2183 5664 2228 5692
rect 2222 5652 2228 5664
rect 2280 5652 2286 5704
rect 2498 5652 2504 5704
rect 2556 5692 2562 5704
rect 3786 5692 3792 5704
rect 2556 5664 3792 5692
rect 2556 5652 2562 5664
rect 3786 5652 3792 5664
rect 3844 5692 3850 5704
rect 4157 5695 4215 5701
rect 4157 5692 4169 5695
rect 3844 5664 4169 5692
rect 3844 5652 3850 5664
rect 4157 5661 4169 5664
rect 4203 5661 4215 5695
rect 4157 5655 4215 5661
rect 6549 5695 6607 5701
rect 6549 5661 6561 5695
rect 6595 5661 6607 5695
rect 8102 5695 8160 5701
rect 8102 5692 8114 5695
rect 6549 5655 6607 5661
rect 8036 5664 8114 5692
rect 1762 5556 1768 5568
rect 1723 5528 1768 5556
rect 1762 5516 1768 5528
rect 1820 5516 1826 5568
rect 2133 5559 2191 5565
rect 2133 5525 2145 5559
rect 2179 5556 2191 5559
rect 2590 5556 2596 5568
rect 2179 5528 2596 5556
rect 2179 5525 2191 5528
rect 2133 5519 2191 5525
rect 2590 5516 2596 5528
rect 2648 5556 2654 5568
rect 3326 5556 3332 5568
rect 2648 5528 3332 5556
rect 2648 5516 2654 5528
rect 3326 5516 3332 5528
rect 3384 5516 3390 5568
rect 3694 5516 3700 5568
rect 3752 5556 3758 5568
rect 3789 5559 3847 5565
rect 3789 5556 3801 5559
rect 3752 5528 3801 5556
rect 3752 5516 3758 5528
rect 3789 5525 3801 5528
rect 3835 5525 3847 5559
rect 3789 5519 3847 5525
rect 6178 5516 6184 5568
rect 6236 5556 6242 5568
rect 6273 5559 6331 5565
rect 6273 5556 6285 5559
rect 6236 5528 6285 5556
rect 6236 5516 6242 5528
rect 6273 5525 6285 5528
rect 6319 5556 6331 5559
rect 6564 5556 6592 5655
rect 8036 5568 8064 5664
rect 8102 5661 8114 5664
rect 8148 5661 8160 5695
rect 8102 5655 8160 5661
rect 8757 5695 8815 5701
rect 8757 5661 8769 5695
rect 8803 5692 8815 5695
rect 9306 5692 9312 5704
rect 8803 5664 9312 5692
rect 8803 5661 8815 5664
rect 8757 5655 8815 5661
rect 9306 5652 9312 5664
rect 9364 5652 9370 5704
rect 10321 5695 10379 5701
rect 10321 5661 10333 5695
rect 10367 5692 10379 5695
rect 10502 5692 10508 5704
rect 10367 5664 10508 5692
rect 10367 5661 10379 5664
rect 10321 5655 10379 5661
rect 10502 5652 10508 5664
rect 10560 5652 10566 5704
rect 10781 5695 10839 5701
rect 10781 5661 10793 5695
rect 10827 5661 10839 5695
rect 10781 5655 10839 5661
rect 9324 5624 9352 5652
rect 10796 5624 10824 5655
rect 11790 5652 11796 5704
rect 11848 5692 11854 5704
rect 12069 5695 12127 5701
rect 12069 5692 12081 5695
rect 11848 5664 12081 5692
rect 11848 5652 11854 5664
rect 12069 5661 12081 5664
rect 12115 5661 12127 5695
rect 12342 5692 12348 5704
rect 12303 5664 12348 5692
rect 12069 5655 12127 5661
rect 12342 5652 12348 5664
rect 12400 5652 12406 5704
rect 14642 5652 14648 5704
rect 14700 5692 14706 5704
rect 14737 5695 14795 5701
rect 14737 5692 14749 5695
rect 14700 5664 14749 5692
rect 14700 5652 14706 5664
rect 14737 5661 14749 5664
rect 14783 5692 14795 5695
rect 18138 5692 18144 5704
rect 14783 5664 18144 5692
rect 14783 5661 14795 5664
rect 14737 5655 14795 5661
rect 18138 5652 18144 5664
rect 18196 5652 18202 5704
rect 19981 5695 20039 5701
rect 19981 5661 19993 5695
rect 20027 5692 20039 5695
rect 21266 5692 21272 5704
rect 20027 5664 21272 5692
rect 20027 5661 20039 5664
rect 19981 5655 20039 5661
rect 21266 5652 21272 5664
rect 21324 5652 21330 5704
rect 21450 5692 21456 5704
rect 21411 5664 21456 5692
rect 21450 5652 21456 5664
rect 21508 5652 21514 5704
rect 23290 5692 23296 5704
rect 23251 5664 23296 5692
rect 23290 5652 23296 5664
rect 23348 5652 23354 5704
rect 23937 5695 23995 5701
rect 23937 5661 23949 5695
rect 23983 5692 23995 5695
rect 24394 5692 24400 5704
rect 23983 5664 24400 5692
rect 23983 5661 23995 5664
rect 23937 5655 23995 5661
rect 24394 5652 24400 5664
rect 24452 5652 24458 5704
rect 27154 5692 27160 5704
rect 27115 5664 27160 5692
rect 27154 5652 27160 5664
rect 27212 5652 27218 5704
rect 27801 5695 27859 5701
rect 27801 5661 27813 5695
rect 27847 5692 27859 5695
rect 28718 5692 28724 5704
rect 27847 5664 28724 5692
rect 27847 5661 27859 5664
rect 27801 5655 27859 5661
rect 28718 5652 28724 5664
rect 28776 5652 28782 5704
rect 28810 5652 28816 5704
rect 28868 5692 28874 5704
rect 29549 5695 29607 5701
rect 29549 5692 29561 5695
rect 28868 5664 29561 5692
rect 28868 5652 28874 5664
rect 29549 5661 29561 5664
rect 29595 5661 29607 5695
rect 29549 5655 29607 5661
rect 32217 5695 32275 5701
rect 32217 5661 32229 5695
rect 32263 5692 32275 5695
rect 33410 5692 33416 5704
rect 32263 5664 33416 5692
rect 32263 5661 32275 5664
rect 32217 5655 32275 5661
rect 33410 5652 33416 5664
rect 33468 5652 33474 5704
rect 33870 5692 33876 5704
rect 33783 5664 33876 5692
rect 33870 5652 33876 5664
rect 33928 5692 33934 5704
rect 35345 5695 35403 5701
rect 35345 5692 35357 5695
rect 33928 5664 35357 5692
rect 33928 5652 33934 5664
rect 35345 5661 35357 5664
rect 35391 5661 35403 5695
rect 35345 5655 35403 5661
rect 9324 5596 10824 5624
rect 15470 5584 15476 5636
rect 15528 5624 15534 5636
rect 15930 5624 15936 5636
rect 15528 5596 15936 5624
rect 15528 5584 15534 5596
rect 15930 5584 15936 5596
rect 15988 5624 15994 5636
rect 17218 5624 17224 5636
rect 15988 5596 17224 5624
rect 15988 5584 15994 5596
rect 17218 5584 17224 5596
rect 17276 5584 17282 5636
rect 17402 5624 17408 5636
rect 17363 5596 17408 5624
rect 17402 5584 17408 5596
rect 17460 5584 17466 5636
rect 28736 5624 28764 5652
rect 30926 5624 30932 5636
rect 28736 5596 30932 5624
rect 30926 5584 30932 5596
rect 30984 5584 30990 5636
rect 32766 5624 32772 5636
rect 32727 5596 32772 5624
rect 32766 5584 32772 5596
rect 32824 5584 32830 5636
rect 8018 5556 8024 5568
rect 6319 5528 6592 5556
rect 7931 5528 8024 5556
rect 6319 5525 6331 5528
rect 6273 5519 6331 5525
rect 8018 5516 8024 5528
rect 8076 5556 8082 5568
rect 9030 5556 9036 5568
rect 8076 5528 9036 5556
rect 8076 5516 8082 5528
rect 9030 5516 9036 5528
rect 9088 5516 9094 5568
rect 11882 5516 11888 5568
rect 11940 5556 11946 5568
rect 12986 5556 12992 5568
rect 11940 5528 12992 5556
rect 11940 5516 11946 5528
rect 12986 5516 12992 5528
rect 13044 5516 13050 5568
rect 13354 5556 13360 5568
rect 13315 5528 13360 5556
rect 13354 5516 13360 5528
rect 13412 5516 13418 5568
rect 15286 5516 15292 5568
rect 15344 5556 15350 5568
rect 15565 5559 15623 5565
rect 15565 5556 15577 5559
rect 15344 5528 15577 5556
rect 15344 5516 15350 5528
rect 15565 5525 15577 5528
rect 15611 5525 15623 5559
rect 15565 5519 15623 5525
rect 16298 5516 16304 5568
rect 16356 5556 16362 5568
rect 16485 5559 16543 5565
rect 16485 5556 16497 5559
rect 16356 5528 16497 5556
rect 16356 5516 16362 5528
rect 16485 5525 16497 5528
rect 16531 5556 16543 5559
rect 16758 5556 16764 5568
rect 16531 5528 16764 5556
rect 16531 5525 16543 5528
rect 16485 5519 16543 5525
rect 16758 5516 16764 5528
rect 16816 5516 16822 5568
rect 24210 5556 24216 5568
rect 24171 5528 24216 5556
rect 24210 5516 24216 5528
rect 24268 5516 24274 5568
rect 24302 5516 24308 5568
rect 24360 5556 24366 5568
rect 24673 5559 24731 5565
rect 24673 5556 24685 5559
rect 24360 5528 24685 5556
rect 24360 5516 24366 5528
rect 24673 5525 24685 5528
rect 24719 5556 24731 5559
rect 25038 5556 25044 5568
rect 24719 5528 25044 5556
rect 24719 5525 24731 5528
rect 24673 5519 24731 5525
rect 25038 5516 25044 5528
rect 25096 5516 25102 5568
rect 28626 5516 28632 5568
rect 28684 5556 28690 5568
rect 28721 5559 28779 5565
rect 28721 5556 28733 5559
rect 28684 5528 28733 5556
rect 28684 5516 28690 5528
rect 28721 5525 28733 5528
rect 28767 5525 28779 5559
rect 28721 5519 28779 5525
rect 1104 5466 38824 5488
rect 1104 5414 7648 5466
rect 7700 5414 7712 5466
rect 7764 5414 7776 5466
rect 7828 5414 7840 5466
rect 7892 5414 20982 5466
rect 21034 5414 21046 5466
rect 21098 5414 21110 5466
rect 21162 5414 21174 5466
rect 21226 5414 34315 5466
rect 34367 5414 34379 5466
rect 34431 5414 34443 5466
rect 34495 5414 34507 5466
rect 34559 5414 38824 5466
rect 1104 5392 38824 5414
rect 3326 5352 3332 5364
rect 3287 5324 3332 5352
rect 3326 5312 3332 5324
rect 3384 5312 3390 5364
rect 3970 5352 3976 5364
rect 3931 5324 3976 5352
rect 3970 5312 3976 5324
rect 4028 5312 4034 5364
rect 4706 5352 4712 5364
rect 4667 5324 4712 5352
rect 4706 5312 4712 5324
rect 4764 5312 4770 5364
rect 6549 5355 6607 5361
rect 6549 5321 6561 5355
rect 6595 5352 6607 5355
rect 6638 5352 6644 5364
rect 6595 5324 6644 5352
rect 6595 5321 6607 5324
rect 6549 5315 6607 5321
rect 6638 5312 6644 5324
rect 6696 5352 6702 5364
rect 8113 5355 8171 5361
rect 8113 5352 8125 5355
rect 6696 5324 8125 5352
rect 6696 5312 6702 5324
rect 8113 5321 8125 5324
rect 8159 5321 8171 5355
rect 8386 5352 8392 5364
rect 8347 5324 8392 5352
rect 8113 5315 8171 5321
rect 1535 5287 1593 5293
rect 1535 5253 1547 5287
rect 1581 5284 1593 5287
rect 3694 5284 3700 5296
rect 1581 5256 3700 5284
rect 1581 5253 1593 5256
rect 1535 5247 1593 5253
rect 3694 5244 3700 5256
rect 3752 5244 3758 5296
rect 1762 5176 1768 5228
rect 1820 5216 1826 5228
rect 2130 5216 2136 5228
rect 1820 5188 2136 5216
rect 1820 5176 1826 5188
rect 2130 5176 2136 5188
rect 2188 5216 2194 5228
rect 2409 5219 2467 5225
rect 2409 5216 2421 5219
rect 2188 5188 2421 5216
rect 2188 5176 2194 5188
rect 2409 5185 2421 5188
rect 2455 5185 2467 5219
rect 2409 5179 2467 5185
rect 2682 5176 2688 5228
rect 2740 5216 2746 5228
rect 4295 5219 4353 5225
rect 4295 5216 4307 5219
rect 2740 5188 4307 5216
rect 2740 5176 2746 5188
rect 4295 5185 4307 5188
rect 4341 5185 4353 5219
rect 4724 5216 4752 5312
rect 8128 5284 8156 5315
rect 8386 5312 8392 5324
rect 8444 5312 8450 5364
rect 10134 5352 10140 5364
rect 10095 5324 10140 5352
rect 10134 5312 10140 5324
rect 10192 5312 10198 5364
rect 11885 5355 11943 5361
rect 11885 5321 11897 5355
rect 11931 5352 11943 5355
rect 12526 5352 12532 5364
rect 11931 5324 12532 5352
rect 11931 5321 11943 5324
rect 11885 5315 11943 5321
rect 8757 5287 8815 5293
rect 8757 5284 8769 5287
rect 8128 5256 8769 5284
rect 8757 5253 8769 5256
rect 8803 5284 8815 5287
rect 9122 5284 9128 5296
rect 8803 5256 9128 5284
rect 8803 5253 8815 5256
rect 8757 5247 8815 5253
rect 9122 5244 9128 5256
rect 9180 5244 9186 5296
rect 4295 5179 4353 5185
rect 4448 5188 4752 5216
rect 7193 5219 7251 5225
rect 1486 5157 1492 5160
rect 1464 5151 1492 5157
rect 1464 5148 1476 5151
rect 1399 5120 1476 5148
rect 1464 5117 1476 5120
rect 1544 5148 1550 5160
rect 1857 5151 1915 5157
rect 1857 5148 1869 5151
rect 1544 5120 1869 5148
rect 1464 5111 1492 5117
rect 1486 5108 1492 5111
rect 1544 5108 1550 5120
rect 1857 5117 1869 5120
rect 1903 5148 1915 5151
rect 3970 5148 3976 5160
rect 1903 5120 3976 5148
rect 1903 5117 1915 5120
rect 1857 5111 1915 5117
rect 3970 5108 3976 5120
rect 4028 5108 4034 5160
rect 4208 5151 4266 5157
rect 4208 5117 4220 5151
rect 4254 5148 4266 5151
rect 4448 5148 4476 5188
rect 7193 5185 7205 5219
rect 7239 5216 7251 5219
rect 7466 5216 7472 5228
rect 7239 5188 7472 5216
rect 7239 5185 7251 5188
rect 7193 5179 7251 5185
rect 7466 5176 7472 5188
rect 7524 5176 7530 5228
rect 9306 5216 9312 5228
rect 9267 5188 9312 5216
rect 9306 5176 9312 5188
rect 9364 5176 9370 5228
rect 10597 5219 10655 5225
rect 10597 5185 10609 5219
rect 10643 5216 10655 5219
rect 11900 5216 11928 5315
rect 12526 5312 12532 5324
rect 12584 5312 12590 5364
rect 14090 5352 14096 5364
rect 14051 5324 14096 5352
rect 14090 5312 14096 5324
rect 14148 5352 14154 5364
rect 14369 5355 14427 5361
rect 14369 5352 14381 5355
rect 14148 5324 14381 5352
rect 14148 5312 14154 5324
rect 14369 5321 14381 5324
rect 14415 5321 14427 5355
rect 17034 5352 17040 5364
rect 16995 5324 17040 5352
rect 14369 5315 14427 5321
rect 12158 5244 12164 5296
rect 12216 5284 12222 5296
rect 12253 5287 12311 5293
rect 12253 5284 12265 5287
rect 12216 5256 12265 5284
rect 12216 5244 12222 5256
rect 12253 5253 12265 5256
rect 12299 5284 12311 5287
rect 13725 5287 13783 5293
rect 13725 5284 13737 5287
rect 12299 5256 13737 5284
rect 12299 5253 12311 5256
rect 12253 5247 12311 5253
rect 13725 5253 13737 5256
rect 13771 5253 13783 5287
rect 13725 5247 13783 5253
rect 10643 5188 11928 5216
rect 12805 5219 12863 5225
rect 10643 5185 10655 5188
rect 10597 5179 10655 5185
rect 12805 5185 12817 5219
rect 12851 5216 12863 5219
rect 13354 5216 13360 5228
rect 12851 5188 13360 5216
rect 12851 5185 12863 5188
rect 12805 5179 12863 5185
rect 13354 5176 13360 5188
rect 13412 5176 13418 5228
rect 14384 5216 14412 5315
rect 17034 5312 17040 5324
rect 17092 5312 17098 5364
rect 19242 5352 19248 5364
rect 19203 5324 19248 5352
rect 19242 5312 19248 5324
rect 19300 5312 19306 5364
rect 22189 5355 22247 5361
rect 22189 5321 22201 5355
rect 22235 5352 22247 5355
rect 23109 5355 23167 5361
rect 23109 5352 23121 5355
rect 22235 5324 23121 5352
rect 22235 5321 22247 5324
rect 22189 5315 22247 5321
rect 23109 5321 23121 5324
rect 23155 5352 23167 5355
rect 23382 5352 23388 5364
rect 23155 5324 23388 5352
rect 23155 5321 23167 5324
rect 23109 5315 23167 5321
rect 23382 5312 23388 5324
rect 23440 5312 23446 5364
rect 25222 5352 25228 5364
rect 25183 5324 25228 5352
rect 25222 5312 25228 5324
rect 25280 5352 25286 5364
rect 26510 5352 26516 5364
rect 25280 5324 26516 5352
rect 25280 5312 25286 5324
rect 26510 5312 26516 5324
rect 26568 5352 26574 5364
rect 26568 5324 27108 5352
rect 26568 5312 26574 5324
rect 21450 5244 21456 5296
rect 21508 5284 21514 5296
rect 22465 5287 22523 5293
rect 22465 5284 22477 5287
rect 21508 5256 22477 5284
rect 21508 5244 21514 5256
rect 22465 5253 22477 5256
rect 22511 5253 22523 5287
rect 26605 5287 26663 5293
rect 22465 5247 22523 5253
rect 22572 5256 26004 5284
rect 15286 5216 15292 5228
rect 14384 5188 15056 5216
rect 15247 5188 15292 5216
rect 4254 5120 4476 5148
rect 4254 5117 4266 5120
rect 4208 5111 4266 5117
rect 4522 5108 4528 5160
rect 4580 5148 4586 5160
rect 5077 5151 5135 5157
rect 5077 5148 5089 5151
rect 4580 5120 5089 5148
rect 4580 5108 4586 5120
rect 5077 5117 5089 5120
rect 5123 5148 5135 5151
rect 5442 5148 5448 5160
rect 5123 5120 5448 5148
rect 5123 5117 5135 5120
rect 5077 5111 5135 5117
rect 5442 5108 5448 5120
rect 5500 5108 5506 5160
rect 5721 5151 5779 5157
rect 5721 5117 5733 5151
rect 5767 5148 5779 5151
rect 5994 5148 6000 5160
rect 5767 5120 6000 5148
rect 5767 5117 5779 5120
rect 5721 5111 5779 5117
rect 5994 5108 6000 5120
rect 6052 5108 6058 5160
rect 15028 5157 15056 5188
rect 15286 5176 15292 5188
rect 15344 5216 15350 5228
rect 16117 5219 16175 5225
rect 16117 5216 16129 5219
rect 15344 5188 16129 5216
rect 15344 5176 15350 5188
rect 16117 5185 16129 5188
rect 16163 5185 16175 5219
rect 16117 5179 16175 5185
rect 17218 5176 17224 5228
rect 17276 5216 17282 5228
rect 20717 5219 20775 5225
rect 20717 5216 20729 5219
rect 17276 5188 20729 5216
rect 17276 5176 17282 5188
rect 14829 5151 14887 5157
rect 14829 5117 14841 5151
rect 14875 5117 14887 5151
rect 14829 5111 14887 5117
rect 15013 5151 15071 5157
rect 15013 5117 15025 5151
rect 15059 5148 15071 5151
rect 17773 5151 17831 5157
rect 17773 5148 17785 5151
rect 15059 5120 17785 5148
rect 15059 5117 15071 5120
rect 15013 5111 15071 5117
rect 17773 5117 17785 5120
rect 17819 5117 17831 5151
rect 18046 5148 18052 5160
rect 18007 5120 18052 5148
rect 17773 5111 17831 5117
rect 2317 5083 2375 5089
rect 2317 5049 2329 5083
rect 2363 5080 2375 5083
rect 2498 5080 2504 5092
rect 2363 5052 2504 5080
rect 2363 5049 2375 5052
rect 2317 5043 2375 5049
rect 2498 5040 2504 5052
rect 2556 5080 2562 5092
rect 2771 5083 2829 5089
rect 2771 5080 2783 5083
rect 2556 5052 2783 5080
rect 2556 5040 2562 5052
rect 2771 5049 2783 5052
rect 2817 5080 2829 5083
rect 7514 5083 7572 5089
rect 2817 5052 3740 5080
rect 2817 5049 2829 5052
rect 2771 5043 2829 5049
rect 3712 5021 3740 5052
rect 7514 5049 7526 5083
rect 7560 5049 7572 5083
rect 9030 5080 9036 5092
rect 8991 5052 9036 5080
rect 7514 5043 7572 5049
rect 3697 5015 3755 5021
rect 3697 4981 3709 5015
rect 3743 5012 3755 5015
rect 3878 5012 3884 5024
rect 3743 4984 3884 5012
rect 3743 4981 3755 4984
rect 3697 4975 3755 4981
rect 3878 4972 3884 4984
rect 3936 5012 3942 5024
rect 4430 5012 4436 5024
rect 3936 4984 4436 5012
rect 3936 4972 3942 4984
rect 4430 4972 4436 4984
rect 4488 4972 4494 5024
rect 5445 5015 5503 5021
rect 5445 4981 5457 5015
rect 5491 5012 5503 5015
rect 5626 5012 5632 5024
rect 5491 4984 5632 5012
rect 5491 4981 5503 4984
rect 5445 4975 5503 4981
rect 5626 4972 5632 4984
rect 5684 4972 5690 5024
rect 5718 4972 5724 5024
rect 5776 5012 5782 5024
rect 7009 5015 7067 5021
rect 7009 5012 7021 5015
rect 5776 4984 7021 5012
rect 5776 4972 5782 4984
rect 7009 4981 7021 4984
rect 7055 5012 7067 5015
rect 7098 5012 7104 5024
rect 7055 4984 7104 5012
rect 7055 4981 7067 4984
rect 7009 4975 7067 4981
rect 7098 4972 7104 4984
rect 7156 5012 7162 5024
rect 7529 5012 7557 5043
rect 9030 5040 9036 5052
rect 9088 5040 9094 5092
rect 9122 5040 9128 5092
rect 9180 5080 9186 5092
rect 9180 5052 9225 5080
rect 9180 5040 9186 5052
rect 10226 5040 10232 5092
rect 10284 5080 10290 5092
rect 10505 5083 10563 5089
rect 10505 5080 10517 5083
rect 10284 5052 10517 5080
rect 10284 5040 10290 5052
rect 10505 5049 10517 5052
rect 10551 5080 10563 5083
rect 10959 5083 11017 5089
rect 10959 5080 10971 5083
rect 10551 5052 10971 5080
rect 10551 5049 10563 5052
rect 10505 5043 10563 5049
rect 10959 5049 10971 5052
rect 11005 5080 11017 5083
rect 11005 5052 12756 5080
rect 11005 5049 11017 5052
rect 10959 5043 11017 5049
rect 11514 5012 11520 5024
rect 7156 4984 7557 5012
rect 11475 4984 11520 5012
rect 7156 4972 7162 4984
rect 11514 4972 11520 4984
rect 11572 4972 11578 5024
rect 12728 5021 12756 5052
rect 14642 5040 14648 5092
rect 14700 5080 14706 5092
rect 14844 5080 14872 5111
rect 15194 5080 15200 5092
rect 14700 5052 15200 5080
rect 14700 5040 14706 5052
rect 15194 5040 15200 5052
rect 15252 5040 15258 5092
rect 16022 5080 16028 5092
rect 15983 5052 16028 5080
rect 16022 5040 16028 5052
rect 16080 5080 16086 5092
rect 16438 5083 16496 5089
rect 16438 5080 16450 5083
rect 16080 5052 16450 5080
rect 16080 5040 16086 5052
rect 16438 5049 16450 5052
rect 16484 5049 16496 5083
rect 17788 5080 17816 5111
rect 18046 5108 18052 5120
rect 18104 5108 18110 5160
rect 19720 5157 19748 5188
rect 20717 5185 20729 5188
rect 20763 5185 20775 5219
rect 21266 5216 21272 5228
rect 21227 5188 21272 5216
rect 20717 5179 20775 5185
rect 18509 5151 18567 5157
rect 18509 5117 18521 5151
rect 18555 5117 18567 5151
rect 18509 5111 18567 5117
rect 19705 5151 19763 5157
rect 19705 5117 19717 5151
rect 19751 5117 19763 5151
rect 19705 5111 19763 5117
rect 18524 5080 18552 5111
rect 19794 5108 19800 5160
rect 19852 5148 19858 5160
rect 20165 5151 20223 5157
rect 20165 5148 20177 5151
rect 19852 5120 20177 5148
rect 19852 5108 19858 5120
rect 20165 5117 20177 5120
rect 20211 5117 20223 5151
rect 20732 5148 20760 5179
rect 21266 5176 21272 5188
rect 21324 5176 21330 5228
rect 22572 5148 22600 5256
rect 23014 5176 23020 5228
rect 23072 5216 23078 5228
rect 23385 5219 23443 5225
rect 23385 5216 23397 5219
rect 23072 5188 23397 5216
rect 23072 5176 23078 5188
rect 23385 5185 23397 5188
rect 23431 5216 23443 5219
rect 23753 5219 23811 5225
rect 23753 5216 23765 5219
rect 23431 5188 23765 5216
rect 23431 5185 23443 5188
rect 23385 5179 23443 5185
rect 23753 5185 23765 5188
rect 23799 5185 23811 5219
rect 23753 5179 23811 5185
rect 20732 5120 22600 5148
rect 25685 5151 25743 5157
rect 20165 5111 20223 5117
rect 25685 5117 25697 5151
rect 25731 5148 25743 5151
rect 25866 5148 25872 5160
rect 25731 5120 25872 5148
rect 25731 5117 25743 5120
rect 25685 5111 25743 5117
rect 25866 5108 25872 5120
rect 25924 5108 25930 5160
rect 25976 5148 26004 5256
rect 26605 5253 26617 5287
rect 26651 5253 26663 5287
rect 27080 5284 27108 5324
rect 27154 5312 27160 5364
rect 27212 5352 27218 5364
rect 28534 5352 28540 5364
rect 27212 5324 28540 5352
rect 27212 5312 27218 5324
rect 28534 5312 28540 5324
rect 28592 5352 28598 5364
rect 28629 5355 28687 5361
rect 28629 5352 28641 5355
rect 28592 5324 28641 5352
rect 28592 5312 28598 5324
rect 28629 5321 28641 5324
rect 28675 5321 28687 5355
rect 31938 5352 31944 5364
rect 31899 5324 31944 5352
rect 28629 5315 28687 5321
rect 31938 5312 31944 5324
rect 31996 5312 32002 5364
rect 33410 5352 33416 5364
rect 33371 5324 33416 5352
rect 33410 5312 33416 5324
rect 33468 5312 33474 5364
rect 33870 5352 33876 5364
rect 33831 5324 33876 5352
rect 33870 5312 33876 5324
rect 33928 5312 33934 5364
rect 33962 5312 33968 5364
rect 34020 5352 34026 5364
rect 34149 5355 34207 5361
rect 34149 5352 34161 5355
rect 34020 5324 34161 5352
rect 34020 5312 34026 5324
rect 34149 5321 34161 5324
rect 34195 5321 34207 5355
rect 34149 5315 34207 5321
rect 27433 5287 27491 5293
rect 27433 5284 27445 5287
rect 27080 5256 27445 5284
rect 26605 5247 26663 5253
rect 27433 5253 27445 5256
rect 27479 5253 27491 5287
rect 29457 5287 29515 5293
rect 29457 5284 29469 5287
rect 27433 5247 27491 5253
rect 28092 5256 29469 5284
rect 26620 5216 26648 5247
rect 27157 5219 27215 5225
rect 27157 5216 27169 5219
rect 26620 5188 27169 5216
rect 27157 5185 27169 5188
rect 27203 5216 27215 5219
rect 27246 5216 27252 5228
rect 27203 5188 27252 5216
rect 27203 5185 27215 5188
rect 27157 5179 27215 5185
rect 27246 5176 27252 5188
rect 27304 5176 27310 5228
rect 27448 5216 27476 5247
rect 28092 5216 28120 5256
rect 29457 5253 29469 5256
rect 29503 5253 29515 5287
rect 29457 5247 29515 5253
rect 27448 5188 28120 5216
rect 26878 5148 26884 5160
rect 25976 5120 26884 5148
rect 26878 5108 26884 5120
rect 26936 5108 26942 5160
rect 27522 5108 27528 5160
rect 27580 5148 27586 5160
rect 28092 5157 28120 5188
rect 28353 5219 28411 5225
rect 28353 5185 28365 5219
rect 28399 5216 28411 5219
rect 29914 5216 29920 5228
rect 28399 5188 29920 5216
rect 28399 5185 28411 5188
rect 28353 5179 28411 5185
rect 29914 5176 29920 5188
rect 29972 5176 29978 5228
rect 30926 5176 30932 5228
rect 30984 5216 30990 5228
rect 32769 5219 32827 5225
rect 32769 5216 32781 5219
rect 30984 5188 32781 5216
rect 30984 5176 30990 5188
rect 32769 5185 32781 5188
rect 32815 5185 32827 5219
rect 32769 5179 32827 5185
rect 27617 5151 27675 5157
rect 27617 5148 27629 5151
rect 27580 5120 27629 5148
rect 27580 5108 27586 5120
rect 27617 5117 27629 5120
rect 27663 5117 27675 5151
rect 27617 5111 27675 5117
rect 28077 5151 28135 5157
rect 28077 5117 28089 5151
rect 28123 5117 28135 5151
rect 28077 5111 28135 5117
rect 29178 5108 29184 5160
rect 29236 5148 29242 5160
rect 29273 5151 29331 5157
rect 29273 5148 29285 5151
rect 29236 5120 29285 5148
rect 29236 5108 29242 5120
rect 29273 5117 29285 5120
rect 29319 5148 29331 5151
rect 30101 5151 30159 5157
rect 30101 5148 30113 5151
rect 29319 5120 30113 5148
rect 29319 5117 29331 5120
rect 29273 5111 29331 5117
rect 30101 5117 30113 5120
rect 30147 5117 30159 5151
rect 30650 5148 30656 5160
rect 30611 5120 30656 5148
rect 30101 5111 30159 5117
rect 30650 5108 30656 5120
rect 30708 5108 30714 5160
rect 31573 5151 31631 5157
rect 31573 5117 31585 5151
rect 31619 5148 31631 5151
rect 32217 5151 32275 5157
rect 32217 5148 32229 5151
rect 31619 5120 32229 5148
rect 31619 5117 31631 5120
rect 31573 5111 31631 5117
rect 32217 5117 32229 5120
rect 32263 5148 32275 5151
rect 32306 5148 32312 5160
rect 32263 5120 32312 5148
rect 32263 5117 32275 5120
rect 32217 5111 32275 5117
rect 32306 5108 32312 5120
rect 32364 5108 32370 5160
rect 35342 5108 35348 5160
rect 35400 5148 35406 5160
rect 35472 5151 35530 5157
rect 35472 5148 35484 5151
rect 35400 5120 35484 5148
rect 35400 5108 35406 5120
rect 35472 5117 35484 5120
rect 35518 5148 35530 5151
rect 35897 5151 35955 5157
rect 35897 5148 35909 5151
rect 35518 5120 35909 5148
rect 35518 5117 35530 5120
rect 35472 5111 35530 5117
rect 35897 5117 35909 5120
rect 35943 5117 35955 5151
rect 35897 5111 35955 5117
rect 20438 5080 20444 5092
rect 17788 5052 18552 5080
rect 20399 5052 20444 5080
rect 16438 5043 16496 5049
rect 20438 5040 20444 5052
rect 20496 5040 20502 5092
rect 23845 5083 23903 5089
rect 23845 5049 23857 5083
rect 23891 5080 23903 5083
rect 24210 5080 24216 5092
rect 23891 5052 24216 5080
rect 23891 5049 23903 5052
rect 23845 5043 23903 5049
rect 24210 5040 24216 5052
rect 24268 5040 24274 5092
rect 24394 5080 24400 5092
rect 24307 5052 24400 5080
rect 24394 5040 24400 5052
rect 24452 5080 24458 5092
rect 24946 5080 24952 5092
rect 24452 5052 24952 5080
rect 24452 5040 24458 5052
rect 24946 5040 24952 5052
rect 25004 5040 25010 5092
rect 26006 5083 26064 5089
rect 26006 5080 26018 5083
rect 25700 5052 26018 5080
rect 25700 5024 25728 5052
rect 26006 5049 26018 5052
rect 26052 5049 26064 5083
rect 30974 5083 31032 5089
rect 30974 5080 30986 5083
rect 26006 5043 26064 5049
rect 30484 5052 30986 5080
rect 12713 5015 12771 5021
rect 12713 4981 12725 5015
rect 12759 5012 12771 5015
rect 13170 5012 13176 5024
rect 12759 4984 13176 5012
rect 12759 4981 12771 4984
rect 12713 4975 12771 4981
rect 13170 4972 13176 4984
rect 13228 4972 13234 5024
rect 15562 5012 15568 5024
rect 15523 4984 15568 5012
rect 15562 4972 15568 4984
rect 15620 4972 15626 5024
rect 16758 4972 16764 5024
rect 16816 5012 16822 5024
rect 17313 5015 17371 5021
rect 17313 5012 17325 5015
rect 16816 4984 17325 5012
rect 16816 4972 16822 4984
rect 17313 4981 17325 4984
rect 17359 4981 17371 5015
rect 18138 5012 18144 5024
rect 18099 4984 18144 5012
rect 17313 4975 17371 4981
rect 18138 4972 18144 4984
rect 18196 4972 18202 5024
rect 21177 5015 21235 5021
rect 21177 4981 21189 5015
rect 21223 5012 21235 5015
rect 21542 5012 21548 5024
rect 21223 4984 21548 5012
rect 21223 4981 21235 4984
rect 21177 4975 21235 4981
rect 21542 4972 21548 4984
rect 21600 5012 21606 5024
rect 21637 5015 21695 5021
rect 21637 5012 21649 5015
rect 21600 4984 21649 5012
rect 21600 4972 21606 4984
rect 21637 4981 21649 4984
rect 21683 5012 21695 5015
rect 21910 5012 21916 5024
rect 21683 4984 21916 5012
rect 21683 4981 21695 4984
rect 21637 4975 21695 4981
rect 21910 4972 21916 4984
rect 21968 4972 21974 5024
rect 24762 4972 24768 5024
rect 24820 5012 24826 5024
rect 24857 5015 24915 5021
rect 24857 5012 24869 5015
rect 24820 4984 24869 5012
rect 24820 4972 24826 4984
rect 24857 4981 24869 4984
rect 24903 5012 24915 5015
rect 25222 5012 25228 5024
rect 24903 4984 25228 5012
rect 24903 4981 24915 4984
rect 24857 4975 24915 4981
rect 25222 4972 25228 4984
rect 25280 4972 25286 5024
rect 25593 5015 25651 5021
rect 25593 4981 25605 5015
rect 25639 5012 25651 5015
rect 25682 5012 25688 5024
rect 25639 4984 25688 5012
rect 25639 4981 25651 4984
rect 25593 4975 25651 4981
rect 25682 4972 25688 4984
rect 25740 4972 25746 5024
rect 28810 4972 28816 5024
rect 28868 5012 28874 5024
rect 28997 5015 29055 5021
rect 28997 5012 29009 5015
rect 28868 4984 29009 5012
rect 28868 4972 28874 4984
rect 28997 4981 29009 4984
rect 29043 4981 29055 5015
rect 29822 5012 29828 5024
rect 29783 4984 29828 5012
rect 28997 4975 29055 4981
rect 29822 4972 29828 4984
rect 29880 5012 29886 5024
rect 30484 5021 30512 5052
rect 30974 5049 30986 5052
rect 31020 5049 31032 5083
rect 32490 5080 32496 5092
rect 32451 5052 32496 5080
rect 30974 5043 31032 5049
rect 32490 5040 32496 5052
rect 32548 5040 32554 5092
rect 32585 5083 32643 5089
rect 32585 5049 32597 5083
rect 32631 5049 32643 5083
rect 32585 5043 32643 5049
rect 35575 5083 35633 5089
rect 35575 5049 35587 5083
rect 35621 5080 35633 5083
rect 39574 5080 39580 5092
rect 35621 5052 39580 5080
rect 35621 5049 35633 5052
rect 35575 5043 35633 5049
rect 30469 5015 30527 5021
rect 30469 5012 30481 5015
rect 29880 4984 30481 5012
rect 29880 4972 29886 4984
rect 30469 4981 30481 4984
rect 30515 4981 30527 5015
rect 30469 4975 30527 4981
rect 32306 4972 32312 5024
rect 32364 5012 32370 5024
rect 32600 5012 32628 5043
rect 39574 5040 39580 5052
rect 39632 5040 39638 5092
rect 32364 4984 32628 5012
rect 32364 4972 32370 4984
rect 1104 4922 38824 4944
rect 1104 4870 14315 4922
rect 14367 4870 14379 4922
rect 14431 4870 14443 4922
rect 14495 4870 14507 4922
rect 14559 4870 27648 4922
rect 27700 4870 27712 4922
rect 27764 4870 27776 4922
rect 27828 4870 27840 4922
rect 27892 4870 38824 4922
rect 1104 4848 38824 4870
rect 2133 4811 2191 4817
rect 2133 4777 2145 4811
rect 2179 4808 2191 4811
rect 2222 4808 2228 4820
rect 2179 4780 2228 4808
rect 2179 4777 2191 4780
rect 2133 4771 2191 4777
rect 2222 4768 2228 4780
rect 2280 4768 2286 4820
rect 4157 4811 4215 4817
rect 4157 4808 4169 4811
rect 2424 4780 4169 4808
rect 2038 4632 2044 4684
rect 2096 4672 2102 4684
rect 2225 4675 2283 4681
rect 2225 4672 2237 4675
rect 2096 4644 2237 4672
rect 2096 4632 2102 4644
rect 2225 4641 2237 4644
rect 2271 4672 2283 4675
rect 2424 4672 2452 4780
rect 4157 4777 4169 4780
rect 4203 4777 4215 4811
rect 4157 4771 4215 4777
rect 7929 4811 7987 4817
rect 7929 4777 7941 4811
rect 7975 4808 7987 4811
rect 8018 4808 8024 4820
rect 7975 4780 8024 4808
rect 7975 4777 7987 4780
rect 7929 4771 7987 4777
rect 8018 4768 8024 4780
rect 8076 4768 8082 4820
rect 9306 4768 9312 4820
rect 9364 4808 9370 4820
rect 9861 4811 9919 4817
rect 9861 4808 9873 4811
rect 9364 4780 9873 4808
rect 9364 4768 9370 4780
rect 9861 4777 9873 4780
rect 9907 4777 9919 4811
rect 10226 4808 10232 4820
rect 10187 4780 10232 4808
rect 9861 4771 9919 4777
rect 2498 4700 2504 4752
rect 2556 4740 2562 4752
rect 3786 4740 3792 4752
rect 2556 4712 2601 4740
rect 3747 4712 3792 4740
rect 2556 4700 2562 4712
rect 3786 4700 3792 4712
rect 3844 4700 3850 4752
rect 5718 4700 5724 4752
rect 5776 4740 5782 4752
rect 5950 4743 6008 4749
rect 5950 4740 5962 4743
rect 5776 4712 5962 4740
rect 5776 4700 5782 4712
rect 5950 4709 5962 4712
rect 5996 4709 6008 4743
rect 5950 4703 6008 4709
rect 8757 4743 8815 4749
rect 8757 4709 8769 4743
rect 8803 4740 8815 4743
rect 9214 4740 9220 4752
rect 8803 4712 9220 4740
rect 8803 4709 8815 4712
rect 8757 4703 8815 4709
rect 9214 4700 9220 4712
rect 9272 4700 9278 4752
rect 2271 4644 2452 4672
rect 4065 4675 4123 4681
rect 2271 4641 2283 4644
rect 2225 4635 2283 4641
rect 4065 4641 4077 4675
rect 4111 4672 4123 4675
rect 4522 4672 4528 4684
rect 4111 4644 4528 4672
rect 4111 4641 4123 4644
rect 4065 4635 4123 4641
rect 1578 4564 1584 4616
rect 1636 4604 1642 4616
rect 4080 4604 4108 4635
rect 4522 4632 4528 4644
rect 4580 4632 4586 4684
rect 4617 4675 4675 4681
rect 4617 4641 4629 4675
rect 4663 4672 4675 4675
rect 4982 4672 4988 4684
rect 4663 4644 4988 4672
rect 4663 4641 4675 4644
rect 4617 4635 4675 4641
rect 4982 4632 4988 4644
rect 5040 4672 5046 4684
rect 5166 4672 5172 4684
rect 5040 4644 5172 4672
rect 5040 4632 5046 4644
rect 5166 4632 5172 4644
rect 5224 4632 5230 4684
rect 8297 4675 8355 4681
rect 8297 4641 8309 4675
rect 8343 4672 8355 4675
rect 8386 4672 8392 4684
rect 8343 4644 8392 4672
rect 8343 4641 8355 4644
rect 8297 4635 8355 4641
rect 8386 4632 8392 4644
rect 8444 4632 8450 4684
rect 8570 4672 8576 4684
rect 8531 4644 8576 4672
rect 8570 4632 8576 4644
rect 8628 4632 8634 4684
rect 5626 4604 5632 4616
rect 1636 4576 4108 4604
rect 5587 4576 5632 4604
rect 1636 4564 1642 4576
rect 5626 4564 5632 4576
rect 5684 4564 5690 4616
rect 9030 4604 9036 4616
rect 7621 4576 9036 4604
rect 4246 4496 4252 4548
rect 4304 4536 4310 4548
rect 7621 4536 7649 4576
rect 9030 4564 9036 4576
rect 9088 4564 9094 4616
rect 9876 4604 9904 4771
rect 10226 4768 10232 4780
rect 10284 4768 10290 4820
rect 13906 4808 13912 4820
rect 13867 4780 13912 4808
rect 13906 4768 13912 4780
rect 13964 4768 13970 4820
rect 14642 4808 14648 4820
rect 14603 4780 14648 4808
rect 14642 4768 14648 4780
rect 14700 4768 14706 4820
rect 15838 4768 15844 4820
rect 15896 4808 15902 4820
rect 17129 4811 17187 4817
rect 17129 4808 17141 4811
rect 15896 4780 17141 4808
rect 15896 4768 15902 4780
rect 17129 4777 17141 4780
rect 17175 4777 17187 4811
rect 19794 4808 19800 4820
rect 19755 4780 19800 4808
rect 17129 4771 17187 4777
rect 19794 4768 19800 4780
rect 19852 4808 19858 4820
rect 20165 4811 20223 4817
rect 20165 4808 20177 4811
rect 19852 4780 20177 4808
rect 19852 4768 19858 4780
rect 20165 4777 20177 4780
rect 20211 4777 20223 4811
rect 21542 4808 21548 4820
rect 21503 4780 21548 4808
rect 20165 4771 20223 4777
rect 21542 4768 21548 4780
rect 21600 4768 21606 4820
rect 22002 4808 22008 4820
rect 21963 4780 22008 4808
rect 22002 4768 22008 4780
rect 22060 4768 22066 4820
rect 22557 4811 22615 4817
rect 22557 4777 22569 4811
rect 22603 4808 22615 4811
rect 24210 4808 24216 4820
rect 22603 4780 24216 4808
rect 22603 4777 22615 4780
rect 22557 4771 22615 4777
rect 24210 4768 24216 4780
rect 24268 4768 24274 4820
rect 26697 4811 26755 4817
rect 26697 4777 26709 4811
rect 26743 4808 26755 4811
rect 27338 4808 27344 4820
rect 26743 4780 27344 4808
rect 26743 4777 26755 4780
rect 26697 4771 26755 4777
rect 27338 4768 27344 4780
rect 27396 4768 27402 4820
rect 28718 4768 28724 4820
rect 28776 4808 28782 4820
rect 29273 4811 29331 4817
rect 29273 4808 29285 4811
rect 28776 4780 29285 4808
rect 28776 4768 28782 4780
rect 29273 4777 29285 4780
rect 29319 4808 29331 4811
rect 29362 4808 29368 4820
rect 29319 4780 29368 4808
rect 29319 4777 29331 4780
rect 29273 4771 29331 4777
rect 29362 4768 29368 4780
rect 29420 4768 29426 4820
rect 29730 4768 29736 4820
rect 29788 4808 29794 4820
rect 29788 4780 30052 4808
rect 29788 4768 29794 4780
rect 10965 4743 11023 4749
rect 10965 4709 10977 4743
rect 11011 4740 11023 4743
rect 11241 4743 11299 4749
rect 11241 4740 11253 4743
rect 11011 4712 11253 4740
rect 11011 4709 11023 4712
rect 10965 4703 11023 4709
rect 11241 4709 11253 4712
rect 11287 4740 11299 4743
rect 11514 4740 11520 4752
rect 11287 4712 11520 4740
rect 11287 4709 11299 4712
rect 11241 4703 11299 4709
rect 11514 4700 11520 4712
rect 11572 4700 11578 4752
rect 15289 4743 15347 4749
rect 15289 4709 15301 4743
rect 15335 4740 15347 4743
rect 15930 4740 15936 4752
rect 15335 4712 15936 4740
rect 15335 4709 15347 4712
rect 15289 4703 15347 4709
rect 15930 4700 15936 4712
rect 15988 4700 15994 4752
rect 23290 4740 23296 4752
rect 23251 4712 23296 4740
rect 23290 4700 23296 4712
rect 23348 4700 23354 4752
rect 23474 4700 23480 4752
rect 23532 4740 23538 4752
rect 23569 4743 23627 4749
rect 23569 4740 23581 4743
rect 23532 4712 23581 4740
rect 23532 4700 23538 4712
rect 23569 4709 23581 4712
rect 23615 4709 23627 4743
rect 23569 4703 23627 4709
rect 24854 4700 24860 4752
rect 24912 4740 24918 4752
rect 25087 4743 25145 4749
rect 25087 4740 25099 4743
rect 24912 4712 25099 4740
rect 24912 4700 24918 4712
rect 25087 4709 25099 4712
rect 25133 4709 25145 4743
rect 25087 4703 25145 4709
rect 25222 4700 25228 4752
rect 25280 4740 25286 4752
rect 28163 4743 28221 4749
rect 25280 4712 27844 4740
rect 25280 4700 25286 4712
rect 10042 4672 10048 4684
rect 10003 4644 10048 4672
rect 10042 4632 10048 4644
rect 10100 4632 10106 4684
rect 13078 4672 13084 4684
rect 13039 4644 13084 4672
rect 13078 4632 13084 4644
rect 13136 4632 13142 4684
rect 13265 4675 13323 4681
rect 13265 4672 13277 4675
rect 13182 4644 13277 4672
rect 11149 4607 11207 4613
rect 11149 4604 11161 4607
rect 9876 4576 11161 4604
rect 11149 4573 11161 4576
rect 11195 4573 11207 4607
rect 11149 4567 11207 4573
rect 11425 4607 11483 4613
rect 11425 4573 11437 4607
rect 11471 4604 11483 4607
rect 12342 4604 12348 4616
rect 11471 4576 12348 4604
rect 11471 4573 11483 4576
rect 11425 4567 11483 4573
rect 4304 4508 7649 4536
rect 4304 4496 4310 4508
rect 8018 4496 8024 4548
rect 8076 4536 8082 4548
rect 11440 4536 11468 4567
rect 12342 4564 12348 4576
rect 12400 4564 12406 4616
rect 12986 4564 12992 4616
rect 13044 4604 13050 4616
rect 13182 4604 13210 4644
rect 13265 4641 13277 4644
rect 13311 4672 13323 4675
rect 13446 4672 13452 4684
rect 13311 4644 13452 4672
rect 13311 4641 13323 4644
rect 13265 4635 13323 4641
rect 13446 4632 13452 4644
rect 13504 4632 13510 4684
rect 15010 4632 15016 4684
rect 15068 4672 15074 4684
rect 15473 4675 15531 4681
rect 15473 4672 15485 4675
rect 15068 4644 15485 4672
rect 15068 4632 15074 4644
rect 15473 4641 15485 4644
rect 15519 4641 15531 4675
rect 16942 4672 16948 4684
rect 16855 4644 16948 4672
rect 15473 4635 15531 4641
rect 16942 4632 16948 4644
rect 17000 4672 17006 4684
rect 17681 4675 17739 4681
rect 17681 4672 17693 4675
rect 17000 4644 17693 4672
rect 17000 4632 17006 4644
rect 17681 4641 17693 4644
rect 17727 4641 17739 4675
rect 18785 4675 18843 4681
rect 18785 4672 18797 4675
rect 17681 4635 17739 4641
rect 18432 4644 18797 4672
rect 13354 4604 13360 4616
rect 13044 4576 13210 4604
rect 13315 4576 13360 4604
rect 13044 4564 13050 4576
rect 13354 4564 13360 4576
rect 13412 4564 13418 4616
rect 15286 4564 15292 4616
rect 15344 4604 15350 4616
rect 15841 4607 15899 4613
rect 15841 4604 15853 4607
rect 15344 4576 15853 4604
rect 15344 4564 15350 4576
rect 15841 4573 15853 4576
rect 15887 4604 15899 4607
rect 16298 4604 16304 4616
rect 15887 4576 16304 4604
rect 15887 4573 15899 4576
rect 15841 4567 15899 4573
rect 16298 4564 16304 4576
rect 16356 4604 16362 4616
rect 16393 4607 16451 4613
rect 16393 4604 16405 4607
rect 16356 4576 16405 4604
rect 16356 4564 16362 4576
rect 16393 4573 16405 4576
rect 16439 4573 16451 4607
rect 16393 4567 16451 4573
rect 16577 4607 16635 4613
rect 16577 4573 16589 4607
rect 16623 4604 16635 4607
rect 17402 4604 17408 4616
rect 16623 4576 17408 4604
rect 16623 4573 16635 4576
rect 16577 4567 16635 4573
rect 17402 4564 17408 4576
rect 17460 4604 17466 4616
rect 18432 4613 18460 4644
rect 18785 4641 18797 4644
rect 18831 4672 18843 4675
rect 18874 4672 18880 4684
rect 18831 4644 18880 4672
rect 18831 4641 18843 4644
rect 18785 4635 18843 4641
rect 18874 4632 18880 4644
rect 18932 4632 18938 4684
rect 19061 4675 19119 4681
rect 19061 4641 19073 4675
rect 19107 4672 19119 4675
rect 19150 4672 19156 4684
rect 19107 4644 19156 4672
rect 19107 4641 19119 4644
rect 19061 4635 19119 4641
rect 19150 4632 19156 4644
rect 19208 4632 19214 4684
rect 19521 4675 19579 4681
rect 19521 4641 19533 4675
rect 19567 4672 19579 4675
rect 24946 4672 24952 4684
rect 19567 4644 21772 4672
rect 24907 4644 24952 4672
rect 19567 4641 19579 4644
rect 19521 4635 19579 4641
rect 18417 4607 18475 4613
rect 18417 4604 18429 4607
rect 17460 4576 18429 4604
rect 17460 4564 17466 4576
rect 18417 4573 18429 4576
rect 18463 4573 18475 4607
rect 18417 4567 18475 4573
rect 20438 4564 20444 4616
rect 20496 4604 20502 4616
rect 21634 4604 21640 4616
rect 20496 4576 21640 4604
rect 20496 4564 20502 4576
rect 21634 4564 21640 4576
rect 21692 4564 21698 4616
rect 8076 4508 11468 4536
rect 12161 4539 12219 4545
rect 8076 4496 8082 4508
rect 12161 4505 12173 4539
rect 12207 4536 12219 4539
rect 13004 4536 13032 4564
rect 12207 4508 13032 4536
rect 12207 4505 12219 4508
rect 12161 4499 12219 4505
rect 16758 4496 16764 4548
rect 16816 4536 16822 4548
rect 18877 4539 18935 4545
rect 18877 4536 18889 4539
rect 16816 4508 18889 4536
rect 16816 4496 16822 4508
rect 18877 4505 18889 4508
rect 18923 4536 18935 4539
rect 19242 4536 19248 4548
rect 18923 4508 19248 4536
rect 18923 4505 18935 4508
rect 18877 4499 18935 4505
rect 19242 4496 19248 4508
rect 19300 4496 19306 4548
rect 21744 4536 21772 4644
rect 24946 4632 24952 4644
rect 25004 4632 25010 4684
rect 25958 4632 25964 4684
rect 26016 4672 26022 4684
rect 26513 4675 26571 4681
rect 26513 4672 26525 4675
rect 26016 4644 26525 4672
rect 26016 4632 26022 4644
rect 26513 4641 26525 4644
rect 26559 4672 26571 4675
rect 26786 4672 26792 4684
rect 26559 4644 26792 4672
rect 26559 4641 26571 4644
rect 26513 4635 26571 4641
rect 26786 4632 26792 4644
rect 26844 4632 26850 4684
rect 27816 4672 27844 4712
rect 28163 4709 28175 4743
rect 28209 4740 28221 4743
rect 28442 4740 28448 4752
rect 28209 4712 28448 4740
rect 28209 4709 28221 4712
rect 28163 4703 28221 4709
rect 28442 4700 28448 4712
rect 28500 4740 28506 4752
rect 29822 4740 29828 4752
rect 28500 4712 29828 4740
rect 28500 4700 28506 4712
rect 29822 4700 29828 4712
rect 29880 4749 29886 4752
rect 29880 4743 29928 4749
rect 29880 4709 29882 4743
rect 29916 4709 29928 4743
rect 30024 4740 30052 4780
rect 30650 4768 30656 4820
rect 30708 4808 30714 4820
rect 30745 4811 30803 4817
rect 30745 4808 30757 4811
rect 30708 4780 30757 4808
rect 30708 4768 30714 4780
rect 30745 4777 30757 4780
rect 30791 4777 30803 4811
rect 33873 4811 33931 4817
rect 33873 4808 33885 4811
rect 30745 4771 30803 4777
rect 30852 4780 33885 4808
rect 30852 4740 30880 4780
rect 33873 4777 33885 4780
rect 33919 4777 33931 4811
rect 33873 4771 33931 4777
rect 32306 4740 32312 4752
rect 30024 4712 30880 4740
rect 32267 4712 32312 4740
rect 29880 4703 29928 4709
rect 29880 4700 29886 4703
rect 32306 4700 32312 4712
rect 32364 4700 32370 4752
rect 30650 4672 30656 4684
rect 27816 4644 30656 4672
rect 30650 4632 30656 4644
rect 30708 4632 30714 4684
rect 33689 4675 33747 4681
rect 33689 4641 33701 4675
rect 33735 4672 33747 4675
rect 34146 4672 34152 4684
rect 33735 4644 34152 4672
rect 33735 4641 33747 4644
rect 33689 4635 33747 4641
rect 34146 4632 34152 4644
rect 34204 4632 34210 4684
rect 34768 4675 34826 4681
rect 34768 4641 34780 4675
rect 34814 4672 34826 4675
rect 35342 4672 35348 4684
rect 34814 4644 35348 4672
rect 34814 4641 34826 4644
rect 34768 4635 34826 4641
rect 35342 4632 35348 4644
rect 35400 4672 35406 4684
rect 35802 4672 35808 4684
rect 35400 4644 35808 4672
rect 35400 4632 35406 4644
rect 35802 4632 35808 4644
rect 35860 4632 35866 4684
rect 23474 4564 23480 4616
rect 23532 4604 23538 4616
rect 23934 4604 23940 4616
rect 23532 4576 23577 4604
rect 23895 4576 23940 4604
rect 23532 4564 23538 4576
rect 23934 4564 23940 4576
rect 23992 4564 23998 4616
rect 27614 4604 27620 4616
rect 27575 4576 27620 4604
rect 27614 4564 27620 4576
rect 27672 4564 27678 4616
rect 27801 4607 27859 4613
rect 27801 4573 27813 4607
rect 27847 4604 27859 4607
rect 27982 4604 27988 4616
rect 27847 4576 27988 4604
rect 27847 4573 27859 4576
rect 27801 4567 27859 4573
rect 27982 4564 27988 4576
rect 28040 4564 28046 4616
rect 29086 4564 29092 4616
rect 29144 4604 29150 4616
rect 29549 4607 29607 4613
rect 29549 4604 29561 4607
rect 29144 4576 29561 4604
rect 29144 4564 29150 4576
rect 29549 4573 29561 4576
rect 29595 4573 29607 4607
rect 29549 4567 29607 4573
rect 32217 4607 32275 4613
rect 32217 4573 32229 4607
rect 32263 4604 32275 4607
rect 32858 4604 32864 4616
rect 32263 4576 32864 4604
rect 32263 4573 32275 4576
rect 32217 4567 32275 4573
rect 32858 4564 32864 4576
rect 32916 4564 32922 4616
rect 29178 4536 29184 4548
rect 21744 4508 29184 4536
rect 29178 4496 29184 4508
rect 29236 4496 29242 4548
rect 29638 4496 29644 4548
rect 29696 4536 29702 4548
rect 32766 4536 32772 4548
rect 29696 4508 32772 4536
rect 29696 4496 29702 4508
rect 32766 4496 32772 4508
rect 32824 4496 32830 4548
rect 1673 4471 1731 4477
rect 1673 4437 1685 4471
rect 1719 4468 1731 4471
rect 1946 4468 1952 4480
rect 1719 4440 1952 4468
rect 1719 4437 1731 4440
rect 1673 4431 1731 4437
rect 1946 4428 1952 4440
rect 2004 4428 2010 4480
rect 3142 4468 3148 4480
rect 3103 4440 3148 4468
rect 3142 4428 3148 4440
rect 3200 4428 3206 4480
rect 5261 4471 5319 4477
rect 5261 4437 5273 4471
rect 5307 4468 5319 4471
rect 5994 4468 6000 4480
rect 5307 4440 6000 4468
rect 5307 4437 5319 4440
rect 5261 4431 5319 4437
rect 5994 4428 6000 4440
rect 6052 4428 6058 4480
rect 6549 4471 6607 4477
rect 6549 4437 6561 4471
rect 6595 4468 6607 4471
rect 6825 4471 6883 4477
rect 6825 4468 6837 4471
rect 6595 4440 6837 4468
rect 6595 4437 6607 4440
rect 6549 4431 6607 4437
rect 6825 4437 6837 4440
rect 6871 4468 6883 4471
rect 7006 4468 7012 4480
rect 6871 4440 7012 4468
rect 6871 4437 6883 4440
rect 6825 4431 6883 4437
rect 7006 4428 7012 4440
rect 7064 4428 7070 4480
rect 7285 4471 7343 4477
rect 7285 4437 7297 4471
rect 7331 4468 7343 4471
rect 7466 4468 7472 4480
rect 7331 4440 7472 4468
rect 7331 4437 7343 4440
rect 7285 4431 7343 4437
rect 7466 4428 7472 4440
rect 7524 4428 7530 4480
rect 10597 4471 10655 4477
rect 10597 4437 10609 4471
rect 10643 4468 10655 4471
rect 10778 4468 10784 4480
rect 10643 4440 10784 4468
rect 10643 4437 10655 4440
rect 10597 4431 10655 4437
rect 10778 4428 10784 4440
rect 10836 4428 10842 4480
rect 12529 4471 12587 4477
rect 12529 4437 12541 4471
rect 12575 4468 12587 4471
rect 12710 4468 12716 4480
rect 12575 4440 12716 4468
rect 12575 4437 12587 4440
rect 12529 4431 12587 4437
rect 12710 4428 12716 4440
rect 12768 4428 12774 4480
rect 15010 4468 15016 4480
rect 14971 4440 15016 4468
rect 15010 4428 15016 4440
rect 15068 4428 15074 4480
rect 18138 4468 18144 4480
rect 18099 4440 18144 4468
rect 18138 4428 18144 4440
rect 18196 4428 18202 4480
rect 25777 4471 25835 4477
rect 25777 4437 25789 4471
rect 25823 4468 25835 4471
rect 25866 4468 25872 4480
rect 25823 4440 25872 4468
rect 25823 4437 25835 4440
rect 25777 4431 25835 4437
rect 25866 4428 25872 4440
rect 25924 4428 25930 4480
rect 27246 4468 27252 4480
rect 27207 4440 27252 4468
rect 27246 4428 27252 4440
rect 27304 4428 27310 4480
rect 28718 4468 28724 4480
rect 28679 4440 28724 4468
rect 28718 4428 28724 4440
rect 28776 4428 28782 4480
rect 30466 4468 30472 4480
rect 30427 4440 30472 4468
rect 30466 4428 30472 4440
rect 30524 4428 30530 4480
rect 32490 4428 32496 4480
rect 32548 4468 32554 4480
rect 33137 4471 33195 4477
rect 33137 4468 33149 4471
rect 32548 4440 33149 4468
rect 32548 4428 32554 4440
rect 33137 4437 33149 4440
rect 33183 4437 33195 4471
rect 33137 4431 33195 4437
rect 33962 4428 33968 4480
rect 34020 4468 34026 4480
rect 34839 4471 34897 4477
rect 34839 4468 34851 4471
rect 34020 4440 34851 4468
rect 34020 4428 34026 4440
rect 34839 4437 34851 4440
rect 34885 4437 34897 4471
rect 34839 4431 34897 4437
rect 1104 4378 38824 4400
rect 1104 4326 7648 4378
rect 7700 4326 7712 4378
rect 7764 4326 7776 4378
rect 7828 4326 7840 4378
rect 7892 4326 20982 4378
rect 21034 4326 21046 4378
rect 21098 4326 21110 4378
rect 21162 4326 21174 4378
rect 21226 4326 34315 4378
rect 34367 4326 34379 4378
rect 34431 4326 34443 4378
rect 34495 4326 34507 4378
rect 34559 4326 38824 4378
rect 1104 4304 38824 4326
rect 2498 4264 2504 4276
rect 2459 4236 2504 4264
rect 2498 4224 2504 4236
rect 2556 4224 2562 4276
rect 3050 4224 3056 4276
rect 3108 4264 3114 4276
rect 3108 4236 3372 4264
rect 3108 4224 3114 4236
rect 2130 4128 2136 4140
rect 2091 4100 2136 4128
rect 2130 4088 2136 4100
rect 2188 4088 2194 4140
rect 2869 4131 2927 4137
rect 2869 4097 2881 4131
rect 2915 4128 2927 4131
rect 3050 4128 3056 4140
rect 2915 4100 3056 4128
rect 2915 4097 2927 4100
rect 2869 4091 2927 4097
rect 3050 4088 3056 4100
rect 3108 4088 3114 4140
rect 3344 4137 3372 4236
rect 5626 4224 5632 4276
rect 5684 4264 5690 4276
rect 6089 4267 6147 4273
rect 6089 4264 6101 4267
rect 5684 4236 6101 4264
rect 5684 4224 5690 4236
rect 6089 4233 6101 4236
rect 6135 4233 6147 4267
rect 8110 4264 8116 4276
rect 8023 4236 8116 4264
rect 6089 4227 6147 4233
rect 8110 4224 8116 4236
rect 8168 4264 8174 4276
rect 8570 4264 8576 4276
rect 8168 4236 8576 4264
rect 8168 4224 8174 4236
rect 8570 4224 8576 4236
rect 8628 4224 8634 4276
rect 14001 4267 14059 4273
rect 14001 4233 14013 4267
rect 14047 4264 14059 4267
rect 14826 4264 14832 4276
rect 14047 4236 14832 4264
rect 14047 4233 14059 4236
rect 14001 4227 14059 4233
rect 14826 4224 14832 4236
rect 14884 4264 14890 4276
rect 16574 4264 16580 4276
rect 14884 4236 16580 4264
rect 14884 4224 14890 4236
rect 16574 4224 16580 4236
rect 16632 4224 16638 4276
rect 16758 4224 16764 4276
rect 16816 4224 16822 4276
rect 21913 4267 21971 4273
rect 21913 4233 21925 4267
rect 21959 4264 21971 4267
rect 23017 4267 23075 4273
rect 23017 4264 23029 4267
rect 21959 4236 23029 4264
rect 21959 4233 21971 4236
rect 21913 4227 21971 4233
rect 23017 4233 23029 4236
rect 23063 4264 23075 4267
rect 23106 4264 23112 4276
rect 23063 4236 23112 4264
rect 23063 4233 23075 4236
rect 23017 4227 23075 4233
rect 23106 4224 23112 4236
rect 23164 4264 23170 4276
rect 23382 4264 23388 4276
rect 23164 4236 23388 4264
rect 23164 4224 23170 4236
rect 23382 4224 23388 4236
rect 23440 4224 23446 4276
rect 26513 4267 26571 4273
rect 26513 4233 26525 4267
rect 26559 4264 26571 4267
rect 27246 4264 27252 4276
rect 26559 4236 27252 4264
rect 26559 4233 26571 4236
rect 26513 4227 26571 4233
rect 27246 4224 27252 4236
rect 27304 4264 27310 4276
rect 27522 4264 27528 4276
rect 27304 4236 27528 4264
rect 27304 4224 27310 4236
rect 27522 4224 27528 4236
rect 27580 4224 27586 4276
rect 28442 4264 28448 4276
rect 27632 4236 28448 4264
rect 4617 4199 4675 4205
rect 4617 4165 4629 4199
rect 4663 4196 4675 4199
rect 5534 4196 5540 4208
rect 4663 4168 5540 4196
rect 4663 4165 4675 4168
rect 4617 4159 4675 4165
rect 3329 4131 3387 4137
rect 3329 4097 3341 4131
rect 3375 4097 3387 4131
rect 3329 4091 3387 4097
rect 1670 4060 1676 4072
rect 1631 4032 1676 4060
rect 1670 4020 1676 4032
rect 1728 4020 1734 4072
rect 1946 4060 1952 4072
rect 1907 4032 1952 4060
rect 1946 4020 1952 4032
rect 2004 4020 2010 4072
rect 5000 4069 5028 4168
rect 5534 4156 5540 4168
rect 5592 4156 5598 4208
rect 11790 4156 11796 4208
rect 11848 4196 11854 4208
rect 12529 4199 12587 4205
rect 12529 4196 12541 4199
rect 11848 4168 12541 4196
rect 11848 4156 11854 4168
rect 12529 4165 12541 4168
rect 12575 4165 12587 4199
rect 12529 4159 12587 4165
rect 13078 4156 13084 4208
rect 13136 4196 13142 4208
rect 13541 4199 13599 4205
rect 13541 4196 13553 4199
rect 13136 4168 13553 4196
rect 13136 4156 13142 4168
rect 13541 4165 13553 4168
rect 13587 4196 13599 4199
rect 15654 4196 15660 4208
rect 13587 4168 15660 4196
rect 13587 4165 13599 4168
rect 13541 4159 13599 4165
rect 15654 4156 15660 4168
rect 15712 4156 15718 4208
rect 16669 4199 16727 4205
rect 16669 4165 16681 4199
rect 16715 4196 16727 4199
rect 16776 4196 16804 4224
rect 16715 4168 16804 4196
rect 17037 4199 17095 4205
rect 16715 4165 16727 4168
rect 16669 4159 16727 4165
rect 17037 4165 17049 4199
rect 17083 4196 17095 4199
rect 18782 4196 18788 4208
rect 17083 4168 18788 4196
rect 17083 4165 17095 4168
rect 17037 4159 17095 4165
rect 18782 4156 18788 4168
rect 18840 4156 18846 4208
rect 21634 4156 21640 4208
rect 21692 4196 21698 4208
rect 22557 4199 22615 4205
rect 22557 4196 22569 4199
rect 21692 4168 22569 4196
rect 21692 4156 21698 4168
rect 22557 4165 22569 4168
rect 22603 4165 22615 4199
rect 24762 4196 24768 4208
rect 22557 4159 22615 4165
rect 23768 4168 24768 4196
rect 5258 4128 5264 4140
rect 5219 4100 5264 4128
rect 5258 4088 5264 4100
rect 5316 4088 5322 4140
rect 6086 4088 6092 4140
rect 6144 4128 6150 4140
rect 7561 4131 7619 4137
rect 7561 4128 7573 4131
rect 6144 4100 7573 4128
rect 6144 4088 6150 4100
rect 7561 4097 7573 4100
rect 7607 4128 7619 4131
rect 8018 4128 8024 4140
rect 7607 4100 8024 4128
rect 7607 4097 7619 4100
rect 7561 4091 7619 4097
rect 8018 4088 8024 4100
rect 8076 4088 8082 4140
rect 10226 4088 10232 4140
rect 10284 4128 10290 4140
rect 10597 4131 10655 4137
rect 10597 4128 10609 4131
rect 10284 4100 10609 4128
rect 10284 4088 10290 4100
rect 10597 4097 10609 4100
rect 10643 4097 10655 4131
rect 10597 4091 10655 4097
rect 12452 4100 13814 4128
rect 4985 4063 5043 4069
rect 4985 4029 4997 4063
rect 5031 4029 5043 4063
rect 5166 4060 5172 4072
rect 5127 4032 5172 4060
rect 4985 4023 5043 4029
rect 5166 4020 5172 4032
rect 5224 4020 5230 4072
rect 8478 4060 8484 4072
rect 8439 4032 8484 4060
rect 8478 4020 8484 4032
rect 8536 4020 8542 4072
rect 9033 4063 9091 4069
rect 9033 4060 9045 4063
rect 8772 4032 9045 4060
rect 3142 3952 3148 4004
rect 3200 3992 3206 4004
rect 6917 3995 6975 4001
rect 6917 3992 6929 3995
rect 3200 3964 3245 3992
rect 6564 3964 6929 3992
rect 3200 3952 3206 3964
rect 6564 3936 6592 3964
rect 6917 3961 6929 3964
rect 6963 3961 6975 3995
rect 6917 3955 6975 3961
rect 7006 3952 7012 4004
rect 7064 3992 7070 4004
rect 7064 3964 7109 3992
rect 7064 3952 7070 3964
rect 4154 3884 4160 3936
rect 4212 3924 4218 3936
rect 4212 3896 4257 3924
rect 4212 3884 4218 3896
rect 4430 3884 4436 3936
rect 4488 3924 4494 3936
rect 5718 3924 5724 3936
rect 4488 3896 5724 3924
rect 4488 3884 4494 3896
rect 5718 3884 5724 3896
rect 5776 3884 5782 3936
rect 6546 3924 6552 3936
rect 6507 3896 6552 3924
rect 6546 3884 6552 3896
rect 6604 3884 6610 3936
rect 8662 3884 8668 3936
rect 8720 3924 8726 3936
rect 8772 3933 8800 4032
rect 9033 4029 9045 4032
rect 9079 4060 9091 4063
rect 10134 4060 10140 4072
rect 9079 4032 10140 4060
rect 9079 4029 9091 4032
rect 9033 4023 9091 4029
rect 10134 4020 10140 4032
rect 10192 4020 10198 4072
rect 10502 4060 10508 4072
rect 10463 4032 10508 4060
rect 10502 4020 10508 4032
rect 10560 4020 10566 4072
rect 10778 4060 10784 4072
rect 10739 4032 10784 4060
rect 10778 4020 10784 4032
rect 10836 4020 10842 4072
rect 12452 4069 12480 4100
rect 12069 4063 12127 4069
rect 12069 4029 12081 4063
rect 12115 4060 12127 4063
rect 12437 4063 12495 4069
rect 12437 4060 12449 4063
rect 12115 4032 12449 4060
rect 12115 4029 12127 4032
rect 12069 4023 12127 4029
rect 12437 4029 12449 4032
rect 12483 4029 12495 4063
rect 12710 4060 12716 4072
rect 12671 4032 12716 4060
rect 12437 4023 12495 4029
rect 12710 4020 12716 4032
rect 12768 4020 12774 4072
rect 9677 3995 9735 4001
rect 9677 3961 9689 3995
rect 9723 3992 9735 3995
rect 9858 3992 9864 4004
rect 9723 3964 9864 3992
rect 9723 3961 9735 3964
rect 9677 3955 9735 3961
rect 9858 3952 9864 3964
rect 9916 3992 9922 4004
rect 10796 3992 10824 4020
rect 11238 3992 11244 4004
rect 9916 3964 10824 3992
rect 11199 3964 11244 3992
rect 9916 3952 9922 3964
rect 11238 3952 11244 3964
rect 11296 3952 11302 4004
rect 11790 3992 11796 4004
rect 11751 3964 11796 3992
rect 11790 3952 11796 3964
rect 11848 3952 11854 4004
rect 13786 3992 13814 4100
rect 14182 4088 14188 4140
rect 14240 4128 14246 4140
rect 14369 4131 14427 4137
rect 14369 4128 14381 4131
rect 14240 4100 14381 4128
rect 14240 4088 14246 4100
rect 14369 4097 14381 4100
rect 14415 4128 14427 4131
rect 15562 4128 15568 4140
rect 14415 4100 15148 4128
rect 15523 4100 15568 4128
rect 14415 4097 14427 4100
rect 14369 4091 14427 4097
rect 14826 4060 14832 4072
rect 14787 4032 14832 4060
rect 14826 4020 14832 4032
rect 14884 4020 14890 4072
rect 14918 4020 14924 4072
rect 14976 4060 14982 4072
rect 15120 4069 15148 4100
rect 15562 4088 15568 4100
rect 15620 4088 15626 4140
rect 16301 4131 16359 4137
rect 16301 4097 16313 4131
rect 16347 4128 16359 4131
rect 16761 4131 16819 4137
rect 16761 4128 16773 4131
rect 16347 4100 16773 4128
rect 16347 4097 16359 4100
rect 16301 4091 16359 4097
rect 16761 4097 16773 4100
rect 16807 4128 16819 4131
rect 16850 4128 16856 4140
rect 16807 4100 16856 4128
rect 16807 4097 16819 4100
rect 16761 4091 16819 4097
rect 16850 4088 16856 4100
rect 16908 4088 16914 4140
rect 19334 4088 19340 4140
rect 19392 4128 19398 4140
rect 20165 4131 20223 4137
rect 20165 4128 20177 4131
rect 19392 4100 20177 4128
rect 19392 4088 19398 4100
rect 20165 4097 20177 4100
rect 20211 4128 20223 4131
rect 20346 4128 20352 4140
rect 20211 4100 20352 4128
rect 20211 4097 20223 4100
rect 20165 4091 20223 4097
rect 20346 4088 20352 4100
rect 20404 4088 20410 4140
rect 22002 4088 22008 4140
rect 22060 4128 22066 4140
rect 23768 4137 23796 4168
rect 24762 4156 24768 4168
rect 24820 4156 24826 4208
rect 26786 4196 26792 4208
rect 26747 4168 26792 4196
rect 26786 4156 26792 4168
rect 26844 4156 26850 4208
rect 22189 4131 22247 4137
rect 22189 4128 22201 4131
rect 22060 4100 22201 4128
rect 22060 4088 22066 4100
rect 22189 4097 22201 4100
rect 22235 4097 22247 4131
rect 23753 4131 23811 4137
rect 23753 4128 23765 4131
rect 23731 4100 23765 4128
rect 22189 4091 22247 4097
rect 23753 4097 23765 4100
rect 23799 4097 23811 4131
rect 23753 4091 23811 4097
rect 23934 4088 23940 4140
rect 23992 4128 23998 4140
rect 24029 4131 24087 4137
rect 24029 4128 24041 4131
rect 23992 4100 24041 4128
rect 23992 4088 23998 4100
rect 24029 4097 24041 4100
rect 24075 4097 24087 4131
rect 27632 4128 27660 4236
rect 28442 4224 28448 4236
rect 28500 4224 28506 4276
rect 29086 4264 29092 4276
rect 29047 4236 29092 4264
rect 29086 4224 29092 4236
rect 29144 4224 29150 4276
rect 29822 4224 29828 4276
rect 29880 4264 29886 4276
rect 30285 4267 30343 4273
rect 30285 4264 30297 4267
rect 29880 4236 30297 4264
rect 29880 4224 29886 4236
rect 30285 4233 30297 4236
rect 30331 4233 30343 4267
rect 30285 4227 30343 4233
rect 32217 4267 32275 4273
rect 32217 4233 32229 4267
rect 32263 4264 32275 4267
rect 32306 4264 32312 4276
rect 32263 4236 32312 4264
rect 32263 4233 32275 4236
rect 32217 4227 32275 4233
rect 32306 4224 32312 4236
rect 32364 4224 32370 4276
rect 32858 4264 32864 4276
rect 32819 4236 32864 4264
rect 32858 4224 32864 4236
rect 32916 4264 32922 4276
rect 33962 4264 33968 4276
rect 32916 4236 33968 4264
rect 32916 4224 32922 4236
rect 33962 4224 33968 4236
rect 34020 4224 34026 4276
rect 30650 4196 30656 4208
rect 28966 4168 30052 4196
rect 30611 4168 30656 4196
rect 24029 4091 24087 4097
rect 25970 4100 27660 4128
rect 28077 4131 28135 4137
rect 15105 4063 15163 4069
rect 14976 4032 15021 4060
rect 14976 4020 14982 4032
rect 15105 4029 15117 4063
rect 15151 4060 15163 4063
rect 16025 4063 16083 4069
rect 16025 4060 16037 4063
rect 15151 4032 16037 4060
rect 15151 4029 15163 4032
rect 15105 4023 15163 4029
rect 16025 4029 16037 4032
rect 16071 4029 16083 4063
rect 16390 4060 16396 4072
rect 16351 4032 16396 4060
rect 16025 4023 16083 4029
rect 16390 4020 16396 4032
rect 16448 4020 16454 4072
rect 16574 4069 16580 4072
rect 16540 4063 16580 4069
rect 16540 4029 16552 4063
rect 16540 4023 16580 4029
rect 16574 4020 16580 4023
rect 16632 4020 16638 4072
rect 17954 4020 17960 4072
rect 18012 4060 18018 4072
rect 18049 4063 18107 4069
rect 18049 4060 18061 4063
rect 18012 4032 18061 4060
rect 18012 4020 18018 4032
rect 18049 4029 18061 4032
rect 18095 4029 18107 4063
rect 18049 4023 18107 4029
rect 18138 4020 18144 4072
rect 18196 4060 18202 4072
rect 18509 4063 18567 4069
rect 18509 4060 18521 4063
rect 18196 4032 18521 4060
rect 18196 4020 18202 4032
rect 18509 4029 18521 4032
rect 18555 4029 18567 4063
rect 18874 4060 18880 4072
rect 18835 4032 18880 4060
rect 18509 4023 18567 4029
rect 18874 4020 18880 4032
rect 18932 4020 18938 4072
rect 19245 4063 19303 4069
rect 19245 4029 19257 4063
rect 19291 4029 19303 4063
rect 19245 4023 19303 4029
rect 19521 4063 19579 4069
rect 19521 4029 19533 4063
rect 19567 4060 19579 4063
rect 20993 4063 21051 4069
rect 20993 4060 21005 4063
rect 19567 4032 21005 4060
rect 19567 4029 19579 4032
rect 19521 4023 19579 4029
rect 20993 4029 21005 4032
rect 21039 4060 21051 4063
rect 21082 4060 21088 4072
rect 21039 4032 21088 4060
rect 21039 4029 21051 4032
rect 20993 4023 21051 4029
rect 17773 3995 17831 4001
rect 17773 3992 17785 3995
rect 13786 3964 17785 3992
rect 17773 3961 17785 3964
rect 17819 3992 17831 3995
rect 19260 3992 19288 4023
rect 21082 4020 21088 4032
rect 21140 4020 21146 4072
rect 17819 3964 19288 3992
rect 20901 3995 20959 4001
rect 17819 3961 17831 3964
rect 17773 3955 17831 3961
rect 20901 3961 20913 3995
rect 20947 3992 20959 3995
rect 21355 3995 21413 4001
rect 21355 3992 21367 3995
rect 20947 3964 21367 3992
rect 20947 3961 20959 3964
rect 20901 3955 20959 3961
rect 21355 3961 21367 3964
rect 21401 3992 21413 3995
rect 22020 3992 22048 4088
rect 25133 4063 25191 4069
rect 23400 4032 23520 4060
rect 23400 4004 23428 4032
rect 23382 3992 23388 4004
rect 21401 3964 22048 3992
rect 23343 3964 23388 3992
rect 21401 3961 21413 3964
rect 21355 3955 21413 3961
rect 23382 3952 23388 3964
rect 23440 3952 23446 4004
rect 23492 3992 23520 4032
rect 25133 4029 25145 4063
rect 25179 4060 25191 4063
rect 25593 4063 25651 4069
rect 25593 4060 25605 4063
rect 25179 4032 25605 4060
rect 25179 4029 25191 4032
rect 25133 4023 25191 4029
rect 25593 4029 25605 4032
rect 25639 4060 25651 4063
rect 25774 4060 25780 4072
rect 25639 4032 25780 4060
rect 25639 4029 25651 4032
rect 25593 4023 25651 4029
rect 25774 4020 25780 4032
rect 25832 4020 25838 4072
rect 23845 3995 23903 4001
rect 23845 3992 23857 3995
rect 23492 3964 23857 3992
rect 23845 3961 23857 3964
rect 23891 3961 23903 3995
rect 23845 3955 23903 3961
rect 25501 3995 25559 4001
rect 25501 3961 25513 3995
rect 25547 3992 25559 3995
rect 25682 3992 25688 4004
rect 25547 3964 25688 3992
rect 25547 3961 25559 3964
rect 25501 3955 25559 3961
rect 25682 3952 25688 3964
rect 25740 3992 25746 4004
rect 25970 4001 25998 4100
rect 28077 4097 28089 4131
rect 28123 4128 28135 4131
rect 28966 4128 28994 4168
rect 28123 4100 28994 4128
rect 28123 4097 28135 4100
rect 28077 4091 28135 4097
rect 29362 4088 29368 4140
rect 29420 4128 29426 4140
rect 29420 4100 29465 4128
rect 29420 4088 29426 4100
rect 30024 4069 30052 4168
rect 30650 4156 30656 4168
rect 30708 4156 30714 4208
rect 33410 4156 33416 4208
rect 33468 4196 33474 4208
rect 33551 4199 33609 4205
rect 33551 4196 33563 4199
rect 33468 4168 33563 4196
rect 33468 4156 33474 4168
rect 33551 4165 33563 4168
rect 33597 4165 33609 4199
rect 33551 4159 33609 4165
rect 30009 4063 30067 4069
rect 30009 4029 30021 4063
rect 30055 4060 30067 4063
rect 30282 4060 30288 4072
rect 30055 4032 30288 4060
rect 30055 4029 30067 4032
rect 30009 4023 30067 4029
rect 30282 4020 30288 4032
rect 30340 4020 30346 4072
rect 30650 4020 30656 4072
rect 30708 4060 30714 4072
rect 30837 4063 30895 4069
rect 30837 4060 30849 4063
rect 30708 4032 30849 4060
rect 30708 4020 30714 4032
rect 30837 4029 30849 4032
rect 30883 4029 30895 4063
rect 31294 4060 31300 4072
rect 31255 4032 31300 4060
rect 30837 4023 30895 4029
rect 31294 4020 31300 4032
rect 31352 4020 31358 4072
rect 31478 4020 31484 4072
rect 31536 4060 31542 4072
rect 33480 4063 33538 4069
rect 33480 4060 33492 4063
rect 31536 4032 33492 4060
rect 31536 4020 31542 4032
rect 33480 4029 33492 4032
rect 33526 4060 33538 4063
rect 33873 4063 33931 4069
rect 33873 4060 33885 4063
rect 33526 4032 33885 4060
rect 33526 4029 33538 4032
rect 33480 4023 33538 4029
rect 33873 4029 33885 4032
rect 33919 4029 33931 4063
rect 33873 4023 33931 4029
rect 25955 3995 26013 4001
rect 25955 3992 25967 3995
rect 25740 3964 25967 3992
rect 25740 3952 25746 3964
rect 25955 3961 25967 3964
rect 26001 3961 26013 3995
rect 25955 3955 26013 3961
rect 27433 3995 27491 4001
rect 27433 3961 27445 3995
rect 27479 3961 27491 3995
rect 27433 3955 27491 3961
rect 8757 3927 8815 3933
rect 8757 3924 8769 3927
rect 8720 3896 8769 3924
rect 8720 3884 8726 3896
rect 8757 3893 8769 3896
rect 8803 3893 8815 3927
rect 10042 3924 10048 3936
rect 10003 3896 10048 3924
rect 8757 3887 8815 3893
rect 10042 3884 10048 3896
rect 10100 3884 10106 3936
rect 10226 3884 10232 3936
rect 10284 3924 10290 3936
rect 10321 3927 10379 3933
rect 10321 3924 10333 3927
rect 10284 3896 10333 3924
rect 10284 3884 10290 3896
rect 10321 3893 10333 3896
rect 10367 3893 10379 3927
rect 10321 3887 10379 3893
rect 10870 3884 10876 3936
rect 10928 3924 10934 3936
rect 12069 3927 12127 3933
rect 12069 3924 12081 3927
rect 10928 3896 12081 3924
rect 10928 3884 10934 3896
rect 12069 3893 12081 3896
rect 12115 3924 12127 3927
rect 12161 3927 12219 3933
rect 12161 3924 12173 3927
rect 12115 3896 12173 3924
rect 12115 3893 12127 3896
rect 12069 3887 12127 3893
rect 12161 3893 12173 3896
rect 12207 3893 12219 3927
rect 12161 3887 12219 3893
rect 12618 3884 12624 3936
rect 12676 3924 12682 3936
rect 12897 3927 12955 3933
rect 12897 3924 12909 3927
rect 12676 3896 12909 3924
rect 12676 3884 12682 3896
rect 12897 3893 12909 3896
rect 12943 3893 12955 3927
rect 12897 3887 12955 3893
rect 14737 3927 14795 3933
rect 14737 3893 14749 3927
rect 14783 3924 14795 3927
rect 14918 3924 14924 3936
rect 14783 3896 14924 3924
rect 14783 3893 14795 3896
rect 14737 3887 14795 3893
rect 14918 3884 14924 3896
rect 14976 3884 14982 3936
rect 15930 3924 15936 3936
rect 15891 3896 15936 3924
rect 15930 3884 15936 3896
rect 15988 3884 15994 3936
rect 16025 3927 16083 3933
rect 16025 3893 16037 3927
rect 16071 3924 16083 3927
rect 16942 3924 16948 3936
rect 16071 3896 16948 3924
rect 16071 3893 16083 3896
rect 16025 3887 16083 3893
rect 16942 3884 16948 3896
rect 17000 3884 17006 3936
rect 17402 3924 17408 3936
rect 17363 3896 17408 3924
rect 17402 3884 17408 3896
rect 17460 3884 17466 3936
rect 19150 3884 19156 3936
rect 19208 3924 19214 3936
rect 19797 3927 19855 3933
rect 19797 3924 19809 3927
rect 19208 3896 19809 3924
rect 19208 3884 19214 3896
rect 19797 3893 19809 3896
rect 19843 3893 19855 3927
rect 24762 3924 24768 3936
rect 24723 3896 24768 3924
rect 19797 3887 19855 3893
rect 24762 3884 24768 3896
rect 24820 3884 24826 3936
rect 27249 3927 27307 3933
rect 27249 3893 27261 3927
rect 27295 3924 27307 3927
rect 27448 3924 27476 3955
rect 27522 3952 27528 4004
rect 27580 3992 27586 4004
rect 27580 3964 27625 3992
rect 27580 3952 27586 3964
rect 28718 3952 28724 4004
rect 28776 3992 28782 4004
rect 29362 3992 29368 4004
rect 28776 3964 29368 3992
rect 28776 3952 28782 3964
rect 29362 3952 29368 3964
rect 29420 3992 29426 4004
rect 29457 3995 29515 4001
rect 29457 3992 29469 3995
rect 29420 3964 29469 3992
rect 29420 3952 29426 3964
rect 29457 3961 29469 3964
rect 29503 3961 29515 3995
rect 32401 3995 32459 4001
rect 32401 3992 32413 3995
rect 29457 3955 29515 3961
rect 30795 3964 32413 3992
rect 30795 3924 30823 3964
rect 32401 3961 32413 3964
rect 32447 3961 32459 3995
rect 32401 3955 32459 3961
rect 30926 3924 30932 3936
rect 27295 3896 30823 3924
rect 30887 3896 30932 3924
rect 27295 3893 27307 3896
rect 27249 3887 27307 3893
rect 30926 3884 30932 3896
rect 30984 3884 30990 3936
rect 34146 3884 34152 3936
rect 34204 3924 34210 3936
rect 34241 3927 34299 3933
rect 34241 3924 34253 3927
rect 34204 3896 34253 3924
rect 34204 3884 34210 3896
rect 34241 3893 34253 3896
rect 34287 3893 34299 3927
rect 34241 3887 34299 3893
rect 35161 3927 35219 3933
rect 35161 3893 35173 3927
rect 35207 3924 35219 3927
rect 35342 3924 35348 3936
rect 35207 3896 35348 3924
rect 35207 3893 35219 3896
rect 35161 3887 35219 3893
rect 35342 3884 35348 3896
rect 35400 3884 35406 3936
rect 1104 3834 38824 3856
rect 1104 3782 14315 3834
rect 14367 3782 14379 3834
rect 14431 3782 14443 3834
rect 14495 3782 14507 3834
rect 14559 3782 27648 3834
rect 27700 3782 27712 3834
rect 27764 3782 27776 3834
rect 27828 3782 27840 3834
rect 27892 3782 38824 3834
rect 1104 3760 38824 3782
rect 1670 3720 1676 3732
rect 1631 3692 1676 3720
rect 1670 3680 1676 3692
rect 1728 3680 1734 3732
rect 2038 3720 2044 3732
rect 1999 3692 2044 3720
rect 2038 3680 2044 3692
rect 2096 3680 2102 3732
rect 2222 3720 2228 3732
rect 2183 3692 2228 3720
rect 2222 3680 2228 3692
rect 2280 3680 2286 3732
rect 3142 3720 3148 3732
rect 3103 3692 3148 3720
rect 3142 3680 3148 3692
rect 3200 3680 3206 3732
rect 4341 3723 4399 3729
rect 4341 3689 4353 3723
rect 4387 3720 4399 3723
rect 4522 3720 4528 3732
rect 4387 3692 4528 3720
rect 4387 3689 4399 3692
rect 4341 3683 4399 3689
rect 4522 3680 4528 3692
rect 4580 3680 4586 3732
rect 4801 3723 4859 3729
rect 4801 3689 4813 3723
rect 4847 3720 4859 3723
rect 5166 3720 5172 3732
rect 4847 3692 5172 3720
rect 4847 3689 4859 3692
rect 4801 3683 4859 3689
rect 1946 3612 1952 3664
rect 2004 3652 2010 3664
rect 2866 3652 2872 3664
rect 2004 3624 2872 3652
rect 2004 3612 2010 3624
rect 2409 3587 2467 3593
rect 2409 3553 2421 3587
rect 2455 3584 2467 3587
rect 2498 3584 2504 3596
rect 2455 3556 2504 3584
rect 2455 3553 2467 3556
rect 2409 3547 2467 3553
rect 2498 3544 2504 3556
rect 2556 3544 2562 3596
rect 2700 3593 2728 3624
rect 2866 3612 2872 3624
rect 2924 3652 2930 3664
rect 4154 3652 4160 3664
rect 2924 3624 4160 3652
rect 2924 3612 2930 3624
rect 4154 3612 4160 3624
rect 4212 3652 4218 3664
rect 4816 3652 4844 3683
rect 5166 3680 5172 3692
rect 5224 3680 5230 3732
rect 5905 3723 5963 3729
rect 5905 3689 5917 3723
rect 5951 3720 5963 3723
rect 6546 3720 6552 3732
rect 5951 3692 6552 3720
rect 5951 3689 5963 3692
rect 5905 3683 5963 3689
rect 6546 3680 6552 3692
rect 6604 3680 6610 3732
rect 7190 3720 7196 3732
rect 7151 3692 7196 3720
rect 7190 3680 7196 3692
rect 7248 3680 7254 3732
rect 8110 3680 8116 3732
rect 8168 3720 8174 3732
rect 8665 3723 8723 3729
rect 8665 3720 8677 3723
rect 8168 3692 8677 3720
rect 8168 3680 8174 3692
rect 8665 3689 8677 3692
rect 8711 3689 8723 3723
rect 9950 3720 9956 3732
rect 9911 3692 9956 3720
rect 8665 3683 8723 3689
rect 9950 3680 9956 3692
rect 10008 3680 10014 3732
rect 11238 3680 11244 3732
rect 11296 3720 11302 3732
rect 11793 3723 11851 3729
rect 11793 3720 11805 3723
rect 11296 3692 11805 3720
rect 11296 3680 11302 3692
rect 11793 3689 11805 3692
rect 11839 3689 11851 3723
rect 11793 3683 11851 3689
rect 14093 3723 14151 3729
rect 14093 3689 14105 3723
rect 14139 3720 14151 3723
rect 15470 3720 15476 3732
rect 14139 3692 15476 3720
rect 14139 3689 14151 3692
rect 14093 3683 14151 3689
rect 15470 3680 15476 3692
rect 15528 3680 15534 3732
rect 15654 3680 15660 3732
rect 15712 3720 15718 3732
rect 18966 3720 18972 3732
rect 15712 3692 18972 3720
rect 15712 3680 15718 3692
rect 18966 3680 18972 3692
rect 19024 3680 19030 3732
rect 20346 3720 20352 3732
rect 20307 3692 20352 3720
rect 20346 3680 20352 3692
rect 20404 3680 20410 3732
rect 21082 3720 21088 3732
rect 21043 3692 21088 3720
rect 21082 3680 21088 3692
rect 21140 3680 21146 3732
rect 23474 3680 23480 3732
rect 23532 3720 23538 3732
rect 24946 3720 24952 3732
rect 23532 3692 23577 3720
rect 24907 3692 24952 3720
rect 23532 3680 23538 3692
rect 24946 3680 24952 3692
rect 25004 3680 25010 3732
rect 25038 3680 25044 3732
rect 25096 3720 25102 3732
rect 25547 3723 25605 3729
rect 25547 3720 25559 3723
rect 25096 3692 25559 3720
rect 25096 3680 25102 3692
rect 25547 3689 25559 3692
rect 25593 3689 25605 3723
rect 25547 3683 25605 3689
rect 25958 3680 25964 3732
rect 26016 3720 26022 3732
rect 26329 3723 26387 3729
rect 26329 3720 26341 3723
rect 26016 3692 26341 3720
rect 26016 3680 26022 3692
rect 26329 3689 26341 3692
rect 26375 3720 26387 3723
rect 26878 3720 26884 3732
rect 26375 3692 26884 3720
rect 26375 3689 26387 3692
rect 26329 3683 26387 3689
rect 26878 3680 26884 3692
rect 26936 3680 26942 3732
rect 27893 3723 27951 3729
rect 27893 3689 27905 3723
rect 27939 3720 27951 3723
rect 27982 3720 27988 3732
rect 27939 3692 27988 3720
rect 27939 3689 27951 3692
rect 27893 3683 27951 3689
rect 27982 3680 27988 3692
rect 28040 3680 28046 3732
rect 28626 3680 28632 3732
rect 28684 3720 28690 3732
rect 29362 3720 29368 3732
rect 28684 3692 29040 3720
rect 29323 3692 29368 3720
rect 28684 3680 28690 3692
rect 4212 3624 4844 3652
rect 4212 3612 4218 3624
rect 5994 3612 6000 3664
rect 6052 3652 6058 3664
rect 8386 3652 8392 3664
rect 6052 3624 8392 3652
rect 6052 3612 6058 3624
rect 7208 3596 7236 3624
rect 8386 3612 8392 3624
rect 8444 3612 8450 3664
rect 2685 3587 2743 3593
rect 2685 3553 2697 3587
rect 2731 3553 2743 3587
rect 2685 3547 2743 3553
rect 4062 3544 4068 3596
rect 4120 3584 4126 3596
rect 4960 3587 5018 3593
rect 4960 3584 4972 3587
rect 4120 3556 4972 3584
rect 4120 3544 4126 3556
rect 4960 3553 4972 3556
rect 5006 3584 5018 3587
rect 5074 3584 5080 3596
rect 5006 3556 5080 3584
rect 5006 3553 5018 3556
rect 4960 3547 5018 3553
rect 5074 3544 5080 3556
rect 5132 3544 5138 3596
rect 7190 3584 7196 3596
rect 7103 3556 7196 3584
rect 7190 3544 7196 3556
rect 7248 3544 7254 3596
rect 7377 3587 7435 3593
rect 7377 3553 7389 3587
rect 7423 3553 7435 3587
rect 7377 3547 7435 3553
rect 6825 3519 6883 3525
rect 6825 3485 6837 3519
rect 6871 3516 6883 3519
rect 7392 3516 7420 3547
rect 8110 3544 8116 3596
rect 8168 3584 8174 3596
rect 8481 3587 8539 3593
rect 8481 3584 8493 3587
rect 8168 3556 8493 3584
rect 8168 3544 8174 3556
rect 8481 3553 8493 3556
rect 8527 3553 8539 3587
rect 8481 3547 8539 3553
rect 9493 3587 9551 3593
rect 9493 3553 9505 3587
rect 9539 3584 9551 3587
rect 9766 3584 9772 3596
rect 9539 3556 9772 3584
rect 9539 3553 9551 3556
rect 9493 3547 9551 3553
rect 9766 3544 9772 3556
rect 9824 3544 9830 3596
rect 9968 3584 9996 3680
rect 10502 3612 10508 3664
rect 10560 3652 10566 3664
rect 10597 3655 10655 3661
rect 10597 3652 10609 3655
rect 10560 3624 10609 3652
rect 10560 3612 10566 3624
rect 10597 3621 10609 3624
rect 10643 3652 10655 3655
rect 15286 3652 15292 3664
rect 10643 3624 11560 3652
rect 15247 3624 15292 3652
rect 10643 3621 10655 3624
rect 10597 3615 10655 3621
rect 10870 3584 10876 3596
rect 9876 3556 9996 3584
rect 10831 3556 10876 3584
rect 9876 3516 9904 3556
rect 10870 3544 10876 3556
rect 10928 3544 10934 3596
rect 11532 3593 11560 3624
rect 15286 3612 15292 3624
rect 15344 3612 15350 3664
rect 16393 3655 16451 3661
rect 16393 3652 16405 3655
rect 15396 3624 16405 3652
rect 11517 3587 11575 3593
rect 11517 3553 11529 3587
rect 11563 3584 11575 3587
rect 12250 3584 12256 3596
rect 11563 3556 12256 3584
rect 11563 3553 11575 3556
rect 11517 3547 11575 3553
rect 12250 3544 12256 3556
rect 12308 3584 12314 3596
rect 12345 3587 12403 3593
rect 12345 3584 12357 3587
rect 12308 3556 12357 3584
rect 12308 3544 12314 3556
rect 12345 3553 12357 3556
rect 12391 3553 12403 3587
rect 12345 3547 12403 3553
rect 12621 3587 12679 3593
rect 12621 3553 12633 3587
rect 12667 3584 12679 3587
rect 12710 3584 12716 3596
rect 12667 3556 12716 3584
rect 12667 3553 12679 3556
rect 12621 3547 12679 3553
rect 12710 3544 12716 3556
rect 12768 3544 12774 3596
rect 13906 3584 13912 3596
rect 13819 3556 13912 3584
rect 13906 3544 13912 3556
rect 13964 3584 13970 3596
rect 14369 3587 14427 3593
rect 14369 3584 14381 3587
rect 13964 3556 14381 3584
rect 13964 3544 13970 3556
rect 14369 3553 14381 3556
rect 14415 3553 14427 3587
rect 14369 3547 14427 3553
rect 15194 3544 15200 3596
rect 15252 3584 15258 3596
rect 15396 3584 15424 3624
rect 16393 3621 16405 3624
rect 16439 3652 16451 3655
rect 16574 3652 16580 3664
rect 16439 3624 16580 3652
rect 16439 3621 16451 3624
rect 16393 3615 16451 3621
rect 16574 3612 16580 3624
rect 16632 3612 16638 3664
rect 17402 3612 17408 3664
rect 17460 3652 17466 3664
rect 17460 3624 18552 3652
rect 17460 3612 17466 3624
rect 16758 3584 16764 3596
rect 15252 3556 15424 3584
rect 15488 3556 16764 3584
rect 15252 3544 15258 3556
rect 6871 3488 9904 3516
rect 6871 3485 6883 3488
rect 6825 3479 6883 3485
rect 10042 3476 10048 3528
rect 10100 3516 10106 3528
rect 12805 3519 12863 3525
rect 12805 3516 12817 3519
rect 10100 3488 12817 3516
rect 10100 3476 10106 3488
rect 12805 3485 12817 3488
rect 12851 3485 12863 3519
rect 15488 3516 15516 3556
rect 16758 3544 16764 3556
rect 16816 3544 16822 3596
rect 16853 3587 16911 3593
rect 16853 3553 16865 3587
rect 16899 3584 16911 3587
rect 16942 3584 16948 3596
rect 16899 3556 16948 3584
rect 16899 3553 16911 3556
rect 16853 3547 16911 3553
rect 16942 3544 16948 3556
rect 17000 3584 17006 3596
rect 17954 3584 17960 3596
rect 17000 3556 17960 3584
rect 17000 3544 17006 3556
rect 17954 3544 17960 3556
rect 18012 3544 18018 3596
rect 18138 3584 18144 3596
rect 18099 3556 18144 3584
rect 18138 3544 18144 3556
rect 18196 3544 18202 3596
rect 18524 3593 18552 3624
rect 22002 3612 22008 3664
rect 22060 3652 22066 3664
rect 22142 3655 22200 3661
rect 22142 3652 22154 3655
rect 22060 3624 22154 3652
rect 22060 3612 22066 3624
rect 22142 3621 22154 3624
rect 22188 3621 22200 3655
rect 22142 3615 22200 3621
rect 23109 3655 23167 3661
rect 23109 3621 23121 3655
rect 23155 3652 23167 3655
rect 23934 3652 23940 3664
rect 23155 3624 23940 3652
rect 23155 3621 23167 3624
rect 23109 3615 23167 3621
rect 23934 3612 23940 3624
rect 23992 3612 23998 3664
rect 24029 3655 24087 3661
rect 24029 3621 24041 3655
rect 24075 3652 24087 3655
rect 24210 3652 24216 3664
rect 24075 3624 24216 3652
rect 24075 3621 24087 3624
rect 24029 3615 24087 3621
rect 24210 3612 24216 3624
rect 24268 3612 24274 3664
rect 27249 3655 27307 3661
rect 27249 3621 27261 3655
rect 27295 3652 27307 3655
rect 28902 3652 28908 3664
rect 27295 3624 28908 3652
rect 27295 3621 27307 3624
rect 27249 3615 27307 3621
rect 28902 3612 28908 3624
rect 28960 3612 28966 3664
rect 29012 3652 29040 3692
rect 29362 3680 29368 3692
rect 29420 3680 29426 3732
rect 33275 3723 33333 3729
rect 33275 3720 33287 3723
rect 29472 3692 33287 3720
rect 29472 3652 29500 3692
rect 33275 3689 33287 3692
rect 33321 3689 33333 3723
rect 33275 3683 33333 3689
rect 29012 3624 29500 3652
rect 29733 3655 29791 3661
rect 29733 3621 29745 3655
rect 29779 3652 29791 3655
rect 30466 3652 30472 3664
rect 29779 3624 30472 3652
rect 29779 3621 29791 3624
rect 29733 3615 29791 3621
rect 30466 3612 30472 3624
rect 30524 3612 30530 3664
rect 30929 3655 30987 3661
rect 30929 3621 30941 3655
rect 30975 3652 30987 3655
rect 31294 3652 31300 3664
rect 30975 3624 31300 3652
rect 30975 3621 30987 3624
rect 30929 3615 30987 3621
rect 31294 3612 31300 3624
rect 31352 3612 31358 3664
rect 18509 3587 18567 3593
rect 18509 3553 18521 3587
rect 18555 3553 18567 3587
rect 18877 3587 18935 3593
rect 18877 3584 18889 3587
rect 18509 3547 18567 3553
rect 18800 3556 18889 3584
rect 15654 3516 15660 3528
rect 12805 3479 12863 3485
rect 14108 3488 15516 3516
rect 15615 3488 15660 3516
rect 14108 3460 14136 3488
rect 15654 3476 15660 3488
rect 15712 3476 15718 3528
rect 17218 3516 17224 3528
rect 17131 3488 17224 3516
rect 17218 3476 17224 3488
rect 17276 3516 17282 3528
rect 18800 3516 18828 3556
rect 18877 3553 18889 3556
rect 18923 3553 18935 3587
rect 25406 3584 25412 3596
rect 25367 3556 25412 3584
rect 18877 3547 18935 3553
rect 25406 3544 25412 3556
rect 25464 3544 25470 3596
rect 26786 3584 26792 3596
rect 26747 3556 26792 3584
rect 26786 3544 26792 3556
rect 26844 3544 26850 3596
rect 27062 3584 27068 3596
rect 27023 3556 27068 3584
rect 27062 3544 27068 3556
rect 27120 3544 27126 3596
rect 28128 3587 28186 3593
rect 28128 3553 28140 3587
rect 28174 3584 28186 3587
rect 28350 3584 28356 3596
rect 28174 3556 28356 3584
rect 28174 3553 28186 3556
rect 28128 3547 28186 3553
rect 28350 3544 28356 3556
rect 28408 3544 28414 3596
rect 30282 3544 30288 3596
rect 30340 3584 30346 3596
rect 32192 3587 32250 3593
rect 32192 3584 32204 3587
rect 30340 3556 32204 3584
rect 30340 3544 30346 3556
rect 32192 3553 32204 3556
rect 32238 3584 32250 3587
rect 32674 3584 32680 3596
rect 32238 3556 32680 3584
rect 32238 3553 32250 3556
rect 32192 3547 32250 3553
rect 32674 3544 32680 3556
rect 32732 3544 32738 3596
rect 33226 3593 33232 3596
rect 33204 3587 33232 3593
rect 33204 3553 33216 3587
rect 33284 3584 33290 3596
rect 38102 3584 38108 3596
rect 33284 3556 38108 3584
rect 33204 3547 33232 3553
rect 33226 3544 33232 3547
rect 33284 3544 33290 3556
rect 38102 3544 38108 3556
rect 38160 3544 38166 3596
rect 17276 3488 18828 3516
rect 19153 3519 19211 3525
rect 17276 3476 17282 3488
rect 19153 3485 19165 3519
rect 19199 3516 19211 3519
rect 21637 3519 21695 3525
rect 21637 3516 21649 3519
rect 19199 3488 21649 3516
rect 19199 3485 19211 3488
rect 19153 3479 19211 3485
rect 21637 3485 21649 3488
rect 21683 3516 21695 3519
rect 21821 3519 21879 3525
rect 21821 3516 21833 3519
rect 21683 3488 21833 3516
rect 21683 3485 21695 3488
rect 21637 3479 21695 3485
rect 21821 3485 21833 3488
rect 21867 3485 21879 3519
rect 24578 3516 24584 3528
rect 24539 3488 24584 3516
rect 21821 3479 21879 3485
rect 24578 3476 24584 3488
rect 24636 3476 24642 3528
rect 24762 3476 24768 3528
rect 24820 3516 24826 3528
rect 28215 3519 28273 3525
rect 28215 3516 28227 3519
rect 24820 3488 28227 3516
rect 24820 3476 24826 3488
rect 28215 3485 28227 3488
rect 28261 3485 28273 3519
rect 28215 3479 28273 3485
rect 28718 3476 28724 3528
rect 28776 3516 28782 3528
rect 29638 3516 29644 3528
rect 28776 3488 29644 3516
rect 28776 3476 28782 3488
rect 29638 3476 29644 3488
rect 29696 3476 29702 3528
rect 6457 3451 6515 3457
rect 6457 3417 6469 3451
rect 6503 3448 6515 3451
rect 7374 3448 7380 3460
rect 6503 3420 7380 3448
rect 6503 3417 6515 3420
rect 6457 3411 6515 3417
rect 7374 3408 7380 3420
rect 7432 3408 7438 3460
rect 12434 3448 12440 3460
rect 12395 3420 12440 3448
rect 12434 3408 12440 3420
rect 12492 3408 12498 3460
rect 13817 3451 13875 3457
rect 13817 3417 13829 3451
rect 13863 3448 13875 3451
rect 14090 3448 14096 3460
rect 13863 3420 14096 3448
rect 13863 3417 13875 3420
rect 13817 3411 13875 3417
rect 14090 3408 14096 3420
rect 14148 3408 14154 3460
rect 15562 3448 15568 3460
rect 15523 3420 15568 3448
rect 15562 3408 15568 3420
rect 15620 3408 15626 3460
rect 16666 3408 16672 3460
rect 16724 3448 16730 3460
rect 18782 3448 18788 3460
rect 16724 3420 18788 3448
rect 16724 3408 16730 3420
rect 18782 3408 18788 3420
rect 18840 3448 18846 3460
rect 19794 3448 19800 3460
rect 18840 3420 19800 3448
rect 18840 3408 18846 3420
rect 19794 3408 19800 3420
rect 19852 3408 19858 3460
rect 22741 3451 22799 3457
rect 22741 3417 22753 3451
rect 22787 3448 22799 3451
rect 24210 3448 24216 3460
rect 22787 3420 24216 3448
rect 22787 3417 22799 3420
rect 22741 3411 22799 3417
rect 24210 3408 24216 3420
rect 24268 3408 24274 3460
rect 32263 3451 32321 3457
rect 32263 3417 32275 3451
rect 32309 3448 32321 3451
rect 39574 3448 39580 3460
rect 32309 3420 39580 3448
rect 32309 3417 32321 3420
rect 32263 3411 32321 3417
rect 39574 3408 39580 3420
rect 39632 3408 39638 3460
rect 5031 3383 5089 3389
rect 5031 3349 5043 3383
rect 5077 3380 5089 3383
rect 10318 3380 10324 3392
rect 5077 3352 10324 3380
rect 5077 3349 5089 3352
rect 5031 3343 5089 3349
rect 10318 3340 10324 3352
rect 10376 3340 10382 3392
rect 12250 3380 12256 3392
rect 12211 3352 12256 3380
rect 12250 3340 12256 3352
rect 12308 3340 12314 3392
rect 12618 3340 12624 3392
rect 12676 3380 12682 3392
rect 13357 3383 13415 3389
rect 13357 3380 13369 3383
rect 12676 3352 13369 3380
rect 12676 3340 12682 3352
rect 13357 3349 13369 3352
rect 13403 3349 13415 3383
rect 13357 3343 13415 3349
rect 13630 3340 13636 3392
rect 13688 3380 13694 3392
rect 15013 3383 15071 3389
rect 15013 3380 15025 3383
rect 13688 3352 15025 3380
rect 13688 3340 13694 3352
rect 15013 3349 15025 3352
rect 15059 3380 15071 3383
rect 15194 3380 15200 3392
rect 15059 3352 15200 3380
rect 15059 3349 15071 3352
rect 15013 3343 15071 3349
rect 15194 3340 15200 3352
rect 15252 3380 15258 3392
rect 15427 3383 15485 3389
rect 15427 3380 15439 3383
rect 15252 3352 15439 3380
rect 15252 3340 15258 3352
rect 15427 3349 15439 3352
rect 15473 3349 15485 3383
rect 15746 3380 15752 3392
rect 15707 3352 15752 3380
rect 15427 3343 15485 3349
rect 15746 3340 15752 3352
rect 15804 3340 15810 3392
rect 15838 3340 15844 3392
rect 15896 3380 15902 3392
rect 17402 3380 17408 3392
rect 15896 3352 17408 3380
rect 15896 3340 15902 3352
rect 17402 3340 17408 3352
rect 17460 3380 17466 3392
rect 17497 3383 17555 3389
rect 17497 3380 17509 3383
rect 17460 3352 17509 3380
rect 17460 3340 17466 3352
rect 17497 3349 17509 3352
rect 17543 3349 17555 3383
rect 17497 3343 17555 3349
rect 18874 3340 18880 3392
rect 18932 3380 18938 3392
rect 19521 3383 19579 3389
rect 19521 3380 19533 3383
rect 18932 3352 19533 3380
rect 18932 3340 18938 3352
rect 19521 3349 19533 3352
rect 19567 3380 19579 3383
rect 20622 3380 20628 3392
rect 19567 3352 20628 3380
rect 19567 3349 19579 3352
rect 19521 3343 19579 3349
rect 20622 3340 20628 3352
rect 20680 3340 20686 3392
rect 25961 3383 26019 3389
rect 25961 3349 25973 3383
rect 26007 3380 26019 3383
rect 26050 3380 26056 3392
rect 26007 3352 26056 3380
rect 26007 3349 26019 3352
rect 25961 3343 26019 3349
rect 26050 3340 26056 3352
rect 26108 3340 26114 3392
rect 1104 3290 38824 3312
rect 1104 3238 7648 3290
rect 7700 3238 7712 3290
rect 7764 3238 7776 3290
rect 7828 3238 7840 3290
rect 7892 3238 20982 3290
rect 21034 3238 21046 3290
rect 21098 3238 21110 3290
rect 21162 3238 21174 3290
rect 21226 3238 34315 3290
rect 34367 3238 34379 3290
rect 34431 3238 34443 3290
rect 34495 3238 34507 3290
rect 34559 3238 38824 3290
rect 1104 3216 38824 3238
rect 2498 3176 2504 3188
rect 2459 3148 2504 3176
rect 2498 3136 2504 3148
rect 2556 3136 2562 3188
rect 2866 3176 2872 3188
rect 2827 3148 2872 3176
rect 2866 3136 2872 3148
rect 2924 3136 2930 3188
rect 4062 3176 4068 3188
rect 4023 3148 4068 3176
rect 4062 3136 4068 3148
rect 4120 3136 4126 3188
rect 4709 3179 4767 3185
rect 4709 3145 4721 3179
rect 4755 3176 4767 3179
rect 6086 3176 6092 3188
rect 4755 3148 6092 3176
rect 4755 3145 4767 3148
rect 4709 3139 4767 3145
rect 106 3068 112 3120
rect 164 3108 170 3120
rect 2179 3111 2237 3117
rect 2179 3108 2191 3111
rect 164 3080 2191 3108
rect 164 3068 170 3080
rect 2179 3077 2191 3080
rect 2225 3077 2237 3111
rect 2179 3071 2237 3077
rect 3050 3040 3056 3052
rect 3011 3012 3056 3040
rect 3050 3000 3056 3012
rect 3108 3000 3114 3052
rect 1949 2975 2007 2981
rect 1949 2941 1961 2975
rect 1995 2972 2007 2975
rect 2108 2975 2166 2981
rect 2108 2972 2120 2975
rect 1995 2944 2120 2972
rect 1995 2941 2007 2944
rect 1949 2935 2007 2941
rect 2108 2941 2120 2944
rect 2154 2972 2166 2975
rect 2958 2972 2964 2984
rect 2154 2944 2964 2972
rect 2154 2941 2166 2944
rect 2108 2935 2166 2941
rect 2958 2932 2964 2944
rect 3016 2932 3022 2984
rect 4208 2975 4266 2981
rect 4208 2941 4220 2975
rect 4254 2972 4266 2975
rect 4724 2972 4752 3139
rect 6086 3136 6092 3148
rect 6144 3136 6150 3188
rect 8110 3176 8116 3188
rect 8071 3148 8116 3176
rect 8110 3136 8116 3148
rect 8168 3136 8174 3188
rect 8297 3179 8355 3185
rect 8297 3145 8309 3179
rect 8343 3176 8355 3179
rect 9401 3179 9459 3185
rect 9401 3176 9413 3179
rect 8343 3148 9413 3176
rect 8343 3145 8355 3148
rect 8297 3139 8355 3145
rect 9401 3145 9413 3148
rect 9447 3176 9459 3179
rect 10781 3179 10839 3185
rect 10781 3176 10793 3179
rect 9447 3148 10793 3176
rect 9447 3145 9459 3148
rect 9401 3139 9459 3145
rect 10781 3145 10793 3148
rect 10827 3176 10839 3179
rect 10870 3176 10876 3188
rect 10827 3148 10876 3176
rect 10827 3145 10839 3148
rect 10781 3139 10839 3145
rect 10870 3136 10876 3148
rect 10928 3136 10934 3188
rect 11333 3179 11391 3185
rect 11333 3145 11345 3179
rect 11379 3176 11391 3179
rect 11882 3176 11888 3188
rect 11379 3148 11888 3176
rect 11379 3145 11391 3148
rect 11333 3139 11391 3145
rect 11882 3136 11888 3148
rect 11940 3136 11946 3188
rect 13909 3179 13967 3185
rect 13909 3145 13921 3179
rect 13955 3176 13967 3179
rect 14001 3179 14059 3185
rect 14001 3176 14013 3179
rect 13955 3148 14013 3176
rect 13955 3145 13967 3148
rect 13909 3139 13967 3145
rect 14001 3145 14013 3148
rect 14047 3176 14059 3179
rect 17218 3176 17224 3188
rect 14047 3148 17224 3176
rect 14047 3145 14059 3148
rect 14001 3139 14059 3145
rect 17218 3136 17224 3148
rect 17276 3136 17282 3188
rect 17954 3136 17960 3188
rect 18012 3176 18018 3188
rect 19797 3179 19855 3185
rect 19797 3176 19809 3179
rect 18012 3148 19809 3176
rect 18012 3136 18018 3148
rect 19797 3145 19809 3148
rect 19843 3145 19855 3179
rect 19797 3139 19855 3145
rect 21913 3179 21971 3185
rect 21913 3145 21925 3179
rect 21959 3176 21971 3179
rect 22002 3176 22008 3188
rect 21959 3148 22008 3176
rect 21959 3145 21971 3148
rect 21913 3139 21971 3145
rect 22002 3136 22008 3148
rect 22060 3136 22066 3188
rect 23106 3176 23112 3188
rect 23067 3148 23112 3176
rect 23106 3136 23112 3148
rect 23164 3136 23170 3188
rect 28718 3176 28724 3188
rect 28679 3148 28724 3176
rect 28718 3136 28724 3148
rect 28776 3136 28782 3188
rect 30377 3179 30435 3185
rect 30377 3145 30389 3179
rect 30423 3176 30435 3179
rect 30466 3176 30472 3188
rect 30423 3148 30472 3176
rect 30423 3145 30435 3148
rect 30377 3139 30435 3145
rect 30466 3136 30472 3148
rect 30524 3136 30530 3188
rect 31987 3179 32045 3185
rect 31987 3145 31999 3179
rect 32033 3176 32045 3179
rect 32490 3176 32496 3188
rect 32033 3148 32496 3176
rect 32033 3145 32045 3148
rect 31987 3139 32045 3145
rect 32490 3136 32496 3148
rect 32548 3136 32554 3188
rect 32674 3176 32680 3188
rect 32635 3148 32680 3176
rect 32674 3136 32680 3148
rect 32732 3136 32738 3188
rect 33226 3176 33232 3188
rect 33187 3148 33232 3176
rect 33226 3136 33232 3148
rect 33284 3136 33290 3188
rect 9306 3108 9312 3120
rect 6196 3080 9312 3108
rect 5902 3040 5908 3052
rect 5863 3012 5908 3040
rect 5902 3000 5908 3012
rect 5960 3000 5966 3052
rect 4254 2944 4752 2972
rect 5077 2975 5135 2981
rect 4254 2941 4266 2944
rect 4208 2935 4266 2941
rect 5077 2941 5089 2975
rect 5123 2972 5135 2975
rect 5813 2975 5871 2981
rect 5813 2972 5825 2975
rect 5123 2944 5825 2972
rect 5123 2941 5135 2944
rect 5077 2935 5135 2941
rect 5813 2941 5825 2944
rect 5859 2972 5871 2975
rect 6196 2972 6224 3080
rect 9306 3068 9312 3080
rect 9364 3068 9370 3120
rect 10226 3108 10232 3120
rect 9692 3080 10232 3108
rect 7466 3040 7472 3052
rect 7427 3012 7472 3040
rect 7466 3000 7472 3012
rect 7524 3000 7530 3052
rect 9122 3040 9128 3052
rect 8496 3012 9128 3040
rect 5859 2944 6224 2972
rect 6273 2975 6331 2981
rect 5859 2941 5871 2944
rect 5813 2935 5871 2941
rect 6273 2941 6285 2975
rect 6319 2972 6331 2975
rect 6641 2975 6699 2981
rect 6641 2972 6653 2975
rect 6319 2944 6653 2972
rect 6319 2941 6331 2944
rect 6273 2935 6331 2941
rect 6641 2941 6653 2944
rect 6687 2972 6699 2975
rect 7190 2972 7196 2984
rect 6687 2944 7196 2972
rect 6687 2941 6699 2944
rect 6641 2935 6699 2941
rect 7190 2932 7196 2944
rect 7248 2932 7254 2984
rect 7374 2972 7380 2984
rect 7287 2944 7380 2972
rect 7374 2932 7380 2944
rect 7432 2972 7438 2984
rect 8496 2972 8524 3012
rect 9122 3000 9128 3012
rect 9180 3000 9186 3052
rect 9692 3049 9720 3080
rect 10226 3068 10232 3080
rect 10284 3068 10290 3120
rect 12710 3068 12716 3120
rect 12768 3068 12774 3120
rect 14829 3111 14887 3117
rect 14829 3077 14841 3111
rect 14875 3108 14887 3111
rect 14918 3108 14924 3120
rect 14875 3080 14924 3108
rect 14875 3077 14887 3080
rect 14829 3071 14887 3077
rect 14918 3068 14924 3080
rect 14976 3108 14982 3120
rect 15562 3108 15568 3120
rect 14976 3080 15568 3108
rect 14976 3068 14982 3080
rect 15562 3068 15568 3080
rect 15620 3108 15626 3120
rect 15749 3111 15807 3117
rect 15749 3108 15761 3111
rect 15620 3080 15761 3108
rect 15620 3068 15626 3080
rect 15749 3077 15761 3080
rect 15795 3077 15807 3111
rect 16850 3108 16856 3120
rect 16811 3080 16856 3108
rect 15749 3071 15807 3077
rect 9217 3043 9275 3049
rect 9217 3009 9229 3043
rect 9263 3040 9275 3043
rect 9677 3043 9735 3049
rect 9677 3040 9689 3043
rect 9263 3012 9689 3040
rect 9263 3009 9275 3012
rect 9217 3003 9275 3009
rect 9677 3009 9689 3012
rect 9723 3009 9735 3043
rect 9677 3003 9735 3009
rect 9766 3000 9772 3052
rect 9824 3040 9830 3052
rect 10045 3043 10103 3049
rect 10045 3040 10057 3043
rect 9824 3012 10057 3040
rect 9824 3000 9830 3012
rect 10045 3009 10057 3012
rect 10091 3009 10103 3043
rect 10045 3003 10103 3009
rect 10134 3000 10140 3052
rect 10192 3040 10198 3052
rect 11793 3043 11851 3049
rect 11793 3040 11805 3043
rect 10192 3012 11805 3040
rect 10192 3000 10198 3012
rect 11793 3009 11805 3012
rect 11839 3040 11851 3043
rect 12161 3043 12219 3049
rect 12161 3040 12173 3043
rect 11839 3012 12173 3040
rect 11839 3009 11851 3012
rect 11793 3003 11851 3009
rect 12161 3009 12173 3012
rect 12207 3040 12219 3043
rect 12728 3040 12756 3068
rect 12207 3012 12756 3040
rect 12207 3009 12219 3012
rect 12161 3003 12219 3009
rect 7432 2944 8524 2972
rect 7432 2932 7438 2944
rect 8570 2932 8576 2984
rect 8628 2972 8634 2984
rect 9309 2975 9367 2981
rect 8628 2944 8673 2972
rect 8628 2932 8634 2944
rect 9309 2941 9321 2975
rect 9355 2972 9367 2975
rect 9585 2975 9643 2981
rect 9585 2972 9597 2975
rect 9355 2944 9597 2972
rect 9355 2941 9367 2944
rect 9309 2935 9367 2941
rect 9585 2941 9597 2944
rect 9631 2941 9643 2975
rect 9858 2972 9864 2984
rect 9819 2944 9864 2972
rect 9585 2935 9643 2941
rect 9858 2932 9864 2944
rect 9916 2932 9922 2984
rect 11149 2975 11207 2981
rect 11149 2941 11161 2975
rect 11195 2972 11207 2975
rect 11238 2972 11244 2984
rect 11195 2944 11244 2972
rect 11195 2941 11207 2944
rect 11149 2935 11207 2941
rect 11238 2932 11244 2944
rect 11296 2932 11302 2984
rect 12250 2932 12256 2984
rect 12308 2972 12314 2984
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 12308 2944 12449 2972
rect 12308 2932 12314 2944
rect 12437 2941 12449 2944
rect 12483 2941 12495 2975
rect 12437 2935 12495 2941
rect 4295 2907 4353 2913
rect 4295 2873 4307 2907
rect 4341 2904 4353 2907
rect 9766 2904 9772 2916
rect 4341 2876 9772 2904
rect 4341 2873 4353 2876
rect 4295 2867 4353 2873
rect 9766 2864 9772 2876
rect 9824 2864 9830 2916
rect 7098 2796 7104 2848
rect 7156 2836 7162 2848
rect 8297 2839 8355 2845
rect 8297 2836 8309 2839
rect 7156 2808 8309 2836
rect 7156 2796 7162 2808
rect 8297 2805 8309 2808
rect 8343 2805 8355 2839
rect 8478 2836 8484 2848
rect 8439 2808 8484 2836
rect 8297 2799 8355 2805
rect 8478 2796 8484 2808
rect 8536 2796 8542 2848
rect 8754 2836 8760 2848
rect 8715 2808 8760 2836
rect 8754 2796 8760 2808
rect 8812 2796 8818 2848
rect 9030 2836 9036 2848
rect 8991 2808 9036 2836
rect 9030 2796 9036 2808
rect 9088 2836 9094 2848
rect 9217 2839 9275 2845
rect 9217 2836 9229 2839
rect 9088 2808 9229 2836
rect 9088 2796 9094 2808
rect 9217 2805 9229 2808
rect 9263 2805 9275 2839
rect 12452 2836 12480 2935
rect 12526 2932 12532 2984
rect 12584 2972 12590 2984
rect 12728 2981 12756 3012
rect 13173 3043 13231 3049
rect 13173 3009 13185 3043
rect 13219 3040 13231 3043
rect 13906 3040 13912 3052
rect 13219 3012 13912 3040
rect 13219 3009 13231 3012
rect 13173 3003 13231 3009
rect 13906 3000 13912 3012
rect 13964 3000 13970 3052
rect 15764 3040 15792 3071
rect 16850 3068 16856 3080
rect 16908 3108 16914 3120
rect 18233 3111 18291 3117
rect 18233 3108 18245 3111
rect 16908 3080 18245 3108
rect 16908 3068 16914 3080
rect 18233 3077 18245 3080
rect 18279 3108 18291 3111
rect 19150 3108 19156 3120
rect 18279 3080 19156 3108
rect 18279 3077 18291 3080
rect 18233 3071 18291 3077
rect 17681 3043 17739 3049
rect 17681 3040 17693 3043
rect 15764 3012 17693 3040
rect 17681 3009 17693 3012
rect 17727 3040 17739 3043
rect 18138 3040 18144 3052
rect 17727 3012 18144 3040
rect 17727 3009 17739 3012
rect 17681 3003 17739 3009
rect 18138 3000 18144 3012
rect 18196 3040 18202 3052
rect 18601 3043 18659 3049
rect 18601 3040 18613 3043
rect 18196 3012 18613 3040
rect 18196 3000 18202 3012
rect 18601 3009 18613 3012
rect 18647 3009 18659 3043
rect 18601 3003 18659 3009
rect 12713 2975 12771 2981
rect 12584 2944 12629 2972
rect 12584 2932 12590 2944
rect 12713 2941 12725 2975
rect 12759 2941 12771 2975
rect 12713 2935 12771 2941
rect 12802 2932 12808 2984
rect 12860 2972 12866 2984
rect 14277 2975 14335 2981
rect 14277 2972 14289 2975
rect 12860 2944 14289 2972
rect 12860 2932 12866 2944
rect 14277 2941 14289 2944
rect 14323 2972 14335 2975
rect 14461 2975 14519 2981
rect 14461 2972 14473 2975
rect 14323 2944 14473 2972
rect 14323 2941 14335 2944
rect 14277 2935 14335 2941
rect 14461 2941 14473 2944
rect 14507 2941 14519 2975
rect 14461 2935 14519 2941
rect 16485 2975 16543 2981
rect 16485 2941 16497 2975
rect 16531 2941 16543 2975
rect 16485 2935 16543 2941
rect 12544 2904 12572 2932
rect 13449 2907 13507 2913
rect 13449 2904 13461 2907
rect 12544 2876 13461 2904
rect 13449 2873 13461 2876
rect 13495 2873 13507 2907
rect 15654 2904 15660 2916
rect 13449 2867 13507 2873
rect 15396 2876 15660 2904
rect 14001 2839 14059 2845
rect 14001 2836 14013 2839
rect 12452 2808 14013 2836
rect 9217 2799 9275 2805
rect 14001 2805 14013 2808
rect 14047 2805 14059 2839
rect 14001 2799 14059 2805
rect 15102 2796 15108 2848
rect 15160 2836 15166 2848
rect 15396 2845 15424 2876
rect 15654 2864 15660 2876
rect 15712 2904 15718 2916
rect 16209 2907 16267 2913
rect 16209 2904 16221 2907
rect 15712 2876 16221 2904
rect 15712 2864 15718 2876
rect 16209 2873 16221 2876
rect 16255 2904 16267 2907
rect 16500 2904 16528 2935
rect 16255 2876 16528 2904
rect 16255 2873 16267 2876
rect 16209 2867 16267 2873
rect 16666 2864 16672 2916
rect 16724 2904 16730 2916
rect 17218 2904 17224 2916
rect 16724 2876 17224 2904
rect 16724 2864 16730 2876
rect 17218 2864 17224 2876
rect 17276 2864 17282 2916
rect 18616 2904 18644 3003
rect 18782 2972 18788 2984
rect 18743 2944 18788 2972
rect 18782 2932 18788 2944
rect 18840 2932 18846 2984
rect 19076 2981 19104 3080
rect 19150 3068 19156 3080
rect 19208 3108 19214 3120
rect 20073 3111 20131 3117
rect 20073 3108 20085 3111
rect 19208 3080 20085 3108
rect 19208 3068 19214 3080
rect 20073 3077 20085 3080
rect 20119 3108 20131 3111
rect 20165 3111 20223 3117
rect 20165 3108 20177 3111
rect 20119 3080 20177 3108
rect 20119 3077 20131 3080
rect 20073 3071 20131 3077
rect 20165 3077 20177 3080
rect 20211 3077 20223 3111
rect 20165 3071 20223 3077
rect 20346 3068 20352 3120
rect 20404 3108 20410 3120
rect 20441 3111 20499 3117
rect 20441 3108 20453 3111
rect 20404 3080 20453 3108
rect 20404 3068 20410 3080
rect 20441 3077 20453 3080
rect 20487 3077 20499 3111
rect 20441 3071 20499 3077
rect 24578 3068 24584 3120
rect 24636 3108 24642 3120
rect 24765 3111 24823 3117
rect 24765 3108 24777 3111
rect 24636 3080 24777 3108
rect 24636 3068 24642 3080
rect 24765 3077 24777 3080
rect 24811 3077 24823 3111
rect 24765 3071 24823 3077
rect 25498 3068 25504 3120
rect 25556 3108 25562 3120
rect 32398 3108 32404 3120
rect 25556 3080 26740 3108
rect 25556 3068 25562 3080
rect 19518 3040 19524 3052
rect 19479 3012 19524 3040
rect 19518 3000 19524 3012
rect 19576 3000 19582 3052
rect 19702 3000 19708 3052
rect 19760 3040 19766 3052
rect 20809 3043 20867 3049
rect 20809 3040 20821 3043
rect 19760 3012 20821 3040
rect 19760 3000 19766 3012
rect 20809 3009 20821 3012
rect 20855 3009 20867 3043
rect 20809 3003 20867 3009
rect 22741 3043 22799 3049
rect 22741 3009 22753 3043
rect 22787 3040 22799 3043
rect 23382 3040 23388 3052
rect 22787 3012 23388 3040
rect 22787 3009 22799 3012
rect 22741 3003 22799 3009
rect 23382 3000 23388 3012
rect 23440 3000 23446 3052
rect 23477 3043 23535 3049
rect 23477 3009 23489 3043
rect 23523 3040 23535 3043
rect 24213 3043 24271 3049
rect 24213 3040 24225 3043
rect 23523 3012 24225 3040
rect 23523 3009 23535 3012
rect 23477 3003 23535 3009
rect 24213 3009 24225 3012
rect 24259 3040 24271 3043
rect 24259 3012 26280 3040
rect 24259 3009 24271 3012
rect 24213 3003 24271 3009
rect 18877 2975 18935 2981
rect 18877 2941 18889 2975
rect 18923 2941 18935 2975
rect 18877 2935 18935 2941
rect 19061 2975 19119 2981
rect 19061 2941 19073 2975
rect 19107 2941 19119 2975
rect 19061 2935 19119 2941
rect 18892 2904 18920 2935
rect 19794 2932 19800 2984
rect 19852 2972 19858 2984
rect 20346 2972 20352 2984
rect 19852 2944 20352 2972
rect 19852 2932 19858 2944
rect 20346 2932 20352 2944
rect 20404 2932 20410 2984
rect 20625 2975 20683 2981
rect 20625 2941 20637 2975
rect 20671 2941 20683 2975
rect 20625 2935 20683 2941
rect 22649 2975 22707 2981
rect 22649 2941 22661 2975
rect 22695 2972 22707 2975
rect 23106 2972 23112 2984
rect 22695 2944 23112 2972
rect 22695 2941 22707 2944
rect 22649 2935 22707 2941
rect 19978 2904 19984 2916
rect 18616 2876 19984 2904
rect 19978 2864 19984 2876
rect 20036 2864 20042 2916
rect 20073 2907 20131 2913
rect 20073 2873 20085 2907
rect 20119 2904 20131 2907
rect 20530 2904 20536 2916
rect 20119 2876 20536 2904
rect 20119 2873 20131 2876
rect 20073 2867 20131 2873
rect 20530 2864 20536 2876
rect 20588 2904 20594 2916
rect 20640 2904 20668 2935
rect 23106 2932 23112 2944
rect 23164 2932 23170 2984
rect 25958 2972 25964 2984
rect 25919 2944 25964 2972
rect 25958 2932 25964 2944
rect 26016 2932 26022 2984
rect 26050 2932 26056 2984
rect 26108 2972 26114 2984
rect 26145 2975 26203 2981
rect 26145 2972 26157 2975
rect 26108 2944 26157 2972
rect 26108 2932 26114 2944
rect 26145 2941 26157 2944
rect 26191 2941 26203 2975
rect 26145 2935 26203 2941
rect 20588 2876 20668 2904
rect 24305 2907 24363 2913
rect 20588 2864 20594 2876
rect 24305 2873 24317 2907
rect 24351 2873 24363 2907
rect 24305 2867 24363 2873
rect 15381 2839 15439 2845
rect 15381 2836 15393 2839
rect 15160 2808 15393 2836
rect 15160 2796 15166 2808
rect 15381 2805 15393 2808
rect 15427 2805 15439 2839
rect 15381 2799 15439 2805
rect 16574 2796 16580 2848
rect 16632 2836 16638 2848
rect 18598 2836 18604 2848
rect 16632 2808 18604 2836
rect 16632 2796 16638 2808
rect 18598 2796 18604 2808
rect 18656 2796 18662 2848
rect 20346 2796 20352 2848
rect 20404 2836 20410 2848
rect 21361 2839 21419 2845
rect 21361 2836 21373 2839
rect 20404 2808 21373 2836
rect 20404 2796 20410 2808
rect 21361 2805 21373 2808
rect 21407 2805 21419 2839
rect 24026 2836 24032 2848
rect 23987 2808 24032 2836
rect 21361 2799 21419 2805
rect 24026 2796 24032 2808
rect 24084 2836 24090 2848
rect 24320 2836 24348 2867
rect 25406 2836 25412 2848
rect 24084 2808 24348 2836
rect 25367 2808 25412 2836
rect 24084 2796 24090 2808
rect 25406 2796 25412 2808
rect 25464 2796 25470 2848
rect 25774 2836 25780 2848
rect 25735 2808 25780 2836
rect 25774 2796 25780 2808
rect 25832 2796 25838 2848
rect 26160 2836 26188 2935
rect 26252 2904 26280 3012
rect 26712 2972 26740 3080
rect 27816 3080 29132 3108
rect 32359 3080 32404 3108
rect 26789 3043 26847 3049
rect 26789 3009 26801 3043
rect 26835 3040 26847 3043
rect 26881 3043 26939 3049
rect 26881 3040 26893 3043
rect 26835 3012 26893 3040
rect 26835 3009 26847 3012
rect 26789 3003 26847 3009
rect 26881 3009 26893 3012
rect 26927 3040 26939 3043
rect 27062 3040 27068 3052
rect 26927 3012 27068 3040
rect 26927 3009 26939 3012
rect 26881 3003 26939 3009
rect 27062 3000 27068 3012
rect 27120 3040 27126 3052
rect 27157 3043 27215 3049
rect 27157 3040 27169 3043
rect 27120 3012 27169 3040
rect 27120 3000 27126 3012
rect 27157 3009 27169 3012
rect 27203 3040 27215 3043
rect 27816 3040 27844 3080
rect 27982 3040 27988 3052
rect 27203 3012 27844 3040
rect 27943 3012 27988 3040
rect 27203 3009 27215 3012
rect 27157 3003 27215 3009
rect 27249 2975 27307 2981
rect 27249 2972 27261 2975
rect 26712 2944 27261 2972
rect 27249 2941 27261 2944
rect 27295 2972 27307 2975
rect 27338 2972 27344 2984
rect 27295 2944 27344 2972
rect 27295 2941 27307 2944
rect 27249 2935 27307 2941
rect 27338 2932 27344 2944
rect 27396 2932 27402 2984
rect 27816 2981 27844 3012
rect 27982 3000 27988 3012
rect 28040 3000 28046 3052
rect 29104 3049 29132 3080
rect 32398 3068 32404 3080
rect 32456 3068 32462 3120
rect 29089 3043 29147 3049
rect 29089 3009 29101 3043
rect 29135 3040 29147 3043
rect 30009 3043 30067 3049
rect 29135 3012 29868 3040
rect 29135 3009 29147 3012
rect 29089 3003 29147 3009
rect 27801 2975 27859 2981
rect 27801 2941 27813 2975
rect 27847 2941 27859 2975
rect 27801 2935 27859 2941
rect 28074 2932 28080 2984
rect 28132 2972 28138 2984
rect 29270 2972 29276 2984
rect 28132 2944 29276 2972
rect 28132 2932 28138 2944
rect 29270 2932 29276 2944
rect 29328 2932 29334 2984
rect 29840 2981 29868 3012
rect 30009 3009 30021 3043
rect 30055 3040 30067 3043
rect 30742 3040 30748 3052
rect 30055 3012 30748 3040
rect 30055 3009 30067 3012
rect 30009 3003 30067 3009
rect 30742 3000 30748 3012
rect 30800 3000 30806 3052
rect 29825 2975 29883 2981
rect 29825 2941 29837 2975
rect 29871 2972 29883 2975
rect 29914 2972 29920 2984
rect 29871 2944 29920 2972
rect 29871 2941 29883 2944
rect 29825 2935 29883 2941
rect 29914 2932 29920 2944
rect 29972 2972 29978 2984
rect 31294 2972 31300 2984
rect 29972 2944 31300 2972
rect 29972 2932 29978 2944
rect 31294 2932 31300 2944
rect 31352 2932 31358 2984
rect 31916 2975 31974 2981
rect 31916 2941 31928 2975
rect 31962 2972 31974 2975
rect 32416 2972 32444 3068
rect 31962 2944 32444 2972
rect 31962 2941 31974 2944
rect 31916 2935 31974 2941
rect 30837 2907 30895 2913
rect 30837 2904 30849 2907
rect 26252 2876 30849 2904
rect 30837 2873 30849 2876
rect 30883 2873 30895 2907
rect 30837 2867 30895 2873
rect 26881 2839 26939 2845
rect 26881 2836 26893 2839
rect 26160 2808 26893 2836
rect 26881 2805 26893 2808
rect 26927 2805 26939 2839
rect 28350 2836 28356 2848
rect 28263 2808 28356 2836
rect 26881 2799 26939 2805
rect 28350 2796 28356 2808
rect 28408 2836 28414 2848
rect 30190 2836 30196 2848
rect 28408 2808 30196 2836
rect 28408 2796 28414 2808
rect 30190 2796 30196 2808
rect 30248 2796 30254 2848
rect 1104 2746 38824 2768
rect 1104 2694 14315 2746
rect 14367 2694 14379 2746
rect 14431 2694 14443 2746
rect 14495 2694 14507 2746
rect 14559 2694 27648 2746
rect 27700 2694 27712 2746
rect 27764 2694 27776 2746
rect 27828 2694 27840 2746
rect 27892 2694 38824 2746
rect 1104 2672 38824 2694
rect 2133 2635 2191 2641
rect 2133 2601 2145 2635
rect 2179 2632 2191 2635
rect 2866 2632 2872 2644
rect 2179 2604 2872 2632
rect 2179 2601 2191 2604
rect 2133 2595 2191 2601
rect 2866 2592 2872 2604
rect 2924 2592 2930 2644
rect 3099 2635 3157 2641
rect 3099 2601 3111 2635
rect 3145 2632 3157 2635
rect 4246 2632 4252 2644
rect 3145 2604 4252 2632
rect 3145 2601 3157 2604
rect 3099 2595 3157 2601
rect 4246 2592 4252 2604
rect 4304 2592 4310 2644
rect 4387 2635 4445 2641
rect 4387 2601 4399 2635
rect 4433 2632 4445 2635
rect 6178 2632 6184 2644
rect 4433 2604 6184 2632
rect 4433 2601 4445 2604
rect 4387 2595 4445 2601
rect 6178 2592 6184 2604
rect 6236 2592 6242 2644
rect 7009 2635 7067 2641
rect 7009 2601 7021 2635
rect 7055 2632 7067 2635
rect 9585 2635 9643 2641
rect 7055 2604 9536 2632
rect 7055 2601 7067 2604
rect 7009 2595 7067 2601
rect 3513 2567 3571 2573
rect 3513 2533 3525 2567
rect 3559 2564 3571 2567
rect 4798 2564 4804 2576
rect 3559 2536 4804 2564
rect 3559 2533 3571 2536
rect 3513 2527 3571 2533
rect 1949 2499 2007 2505
rect 1949 2465 1961 2499
rect 1995 2496 2007 2499
rect 2498 2496 2504 2508
rect 1995 2468 2504 2496
rect 1995 2465 2007 2468
rect 1949 2459 2007 2465
rect 2498 2456 2504 2468
rect 2556 2456 2562 2508
rect 3028 2499 3086 2505
rect 3028 2465 3040 2499
rect 3074 2496 3086 2499
rect 3528 2496 3556 2527
rect 4798 2524 4804 2536
rect 4856 2524 4862 2576
rect 7837 2567 7895 2573
rect 7300 2536 7788 2564
rect 7300 2508 7328 2536
rect 3074 2468 3556 2496
rect 3074 2465 3086 2468
rect 3028 2459 3086 2465
rect 3970 2456 3976 2508
rect 4028 2496 4034 2508
rect 4284 2499 4342 2505
rect 4284 2496 4296 2499
rect 4028 2468 4296 2496
rect 4028 2456 4034 2468
rect 4284 2465 4296 2468
rect 4330 2496 4342 2499
rect 4709 2499 4767 2505
rect 4709 2496 4721 2499
rect 4330 2468 4721 2496
rect 4330 2465 4342 2468
rect 4284 2459 4342 2465
rect 4709 2465 4721 2468
rect 4755 2465 4767 2499
rect 4709 2459 4767 2465
rect 5905 2499 5963 2505
rect 5905 2465 5917 2499
rect 5951 2465 5963 2499
rect 5905 2459 5963 2465
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 5169 2431 5227 2437
rect 5169 2428 5181 2431
rect 1360 2400 5181 2428
rect 1360 2388 1366 2400
rect 5169 2397 5181 2400
rect 5215 2428 5227 2431
rect 5920 2428 5948 2459
rect 5994 2456 6000 2508
rect 6052 2496 6058 2508
rect 6052 2468 6097 2496
rect 6052 2456 6058 2468
rect 6638 2456 6644 2508
rect 6696 2496 6702 2508
rect 7098 2496 7104 2508
rect 6696 2468 7104 2496
rect 6696 2456 6702 2468
rect 7098 2456 7104 2468
rect 7156 2456 7162 2508
rect 7193 2499 7251 2505
rect 7193 2465 7205 2499
rect 7239 2496 7251 2499
rect 7282 2496 7288 2508
rect 7239 2468 7288 2496
rect 7239 2465 7251 2468
rect 7193 2459 7251 2465
rect 7282 2456 7288 2468
rect 7340 2456 7346 2508
rect 7374 2456 7380 2508
rect 7432 2496 7438 2508
rect 7760 2496 7788 2536
rect 7837 2533 7849 2567
rect 7883 2564 7895 2567
rect 8110 2564 8116 2576
rect 7883 2536 8116 2564
rect 7883 2533 7895 2536
rect 7837 2527 7895 2533
rect 8110 2524 8116 2536
rect 8168 2524 8174 2576
rect 9030 2564 9036 2576
rect 8220 2536 9036 2564
rect 8220 2505 8248 2536
rect 9030 2524 9036 2536
rect 9088 2524 9094 2576
rect 8205 2499 8263 2505
rect 8205 2496 8217 2499
rect 7432 2468 7477 2496
rect 7760 2468 8217 2496
rect 7432 2456 7438 2468
rect 8205 2465 8217 2468
rect 8251 2465 8263 2499
rect 8205 2459 8263 2465
rect 8665 2499 8723 2505
rect 8665 2465 8677 2499
rect 8711 2496 8723 2499
rect 9214 2496 9220 2508
rect 8711 2468 9220 2496
rect 8711 2465 8723 2468
rect 8665 2459 8723 2465
rect 9214 2456 9220 2468
rect 9272 2456 9278 2508
rect 9508 2496 9536 2604
rect 9585 2601 9597 2635
rect 9631 2632 9643 2635
rect 9858 2632 9864 2644
rect 9631 2604 9864 2632
rect 9631 2601 9643 2604
rect 9585 2595 9643 2601
rect 9858 2592 9864 2604
rect 9916 2592 9922 2644
rect 12710 2632 12716 2644
rect 10428 2604 12716 2632
rect 10428 2505 10456 2604
rect 12710 2592 12716 2604
rect 12768 2592 12774 2644
rect 12805 2635 12863 2641
rect 12805 2601 12817 2635
rect 12851 2632 12863 2635
rect 12986 2632 12992 2644
rect 12851 2604 12992 2632
rect 12851 2601 12863 2604
rect 12805 2595 12863 2601
rect 12986 2592 12992 2604
rect 13044 2592 13050 2644
rect 14461 2635 14519 2641
rect 14461 2632 14473 2635
rect 13096 2604 14473 2632
rect 11701 2567 11759 2573
rect 11701 2533 11713 2567
rect 11747 2564 11759 2567
rect 11790 2564 11796 2576
rect 11747 2536 11796 2564
rect 11747 2533 11759 2536
rect 11701 2527 11759 2533
rect 11790 2524 11796 2536
rect 11848 2564 11854 2576
rect 12526 2564 12532 2576
rect 11848 2536 12532 2564
rect 11848 2524 11854 2536
rect 12526 2524 12532 2536
rect 12584 2524 12590 2576
rect 12894 2524 12900 2576
rect 12952 2564 12958 2576
rect 13096 2564 13124 2604
rect 14461 2601 14473 2604
rect 14507 2601 14519 2635
rect 14461 2595 14519 2601
rect 14921 2635 14979 2641
rect 14921 2601 14933 2635
rect 14967 2632 14979 2635
rect 15286 2632 15292 2644
rect 14967 2604 15292 2632
rect 14967 2601 14979 2604
rect 14921 2595 14979 2601
rect 12952 2536 13124 2564
rect 13357 2567 13415 2573
rect 12952 2524 12958 2536
rect 13357 2533 13369 2567
rect 13403 2564 13415 2567
rect 13817 2567 13875 2573
rect 13817 2564 13829 2567
rect 13403 2536 13829 2564
rect 13403 2533 13415 2536
rect 13357 2527 13415 2533
rect 13817 2533 13829 2536
rect 13863 2564 13875 2567
rect 14936 2564 14964 2595
rect 15286 2592 15292 2604
rect 15344 2592 15350 2644
rect 16868 2604 18828 2632
rect 13863 2536 14964 2564
rect 13863 2533 13875 2536
rect 13817 2527 13875 2533
rect 16482 2524 16488 2576
rect 16540 2564 16546 2576
rect 16868 2564 16896 2604
rect 17218 2564 17224 2576
rect 16540 2536 16896 2564
rect 17179 2536 17224 2564
rect 16540 2524 16546 2536
rect 9953 2499 10011 2505
rect 9953 2496 9965 2499
rect 9508 2468 9965 2496
rect 9953 2465 9965 2468
rect 9999 2496 10011 2499
rect 10413 2499 10471 2505
rect 10413 2496 10425 2499
rect 9999 2468 10425 2496
rect 9999 2465 10011 2468
rect 9953 2459 10011 2465
rect 10413 2465 10425 2468
rect 10459 2465 10471 2499
rect 10413 2459 10471 2465
rect 10689 2499 10747 2505
rect 10689 2465 10701 2499
rect 10735 2496 10747 2499
rect 11057 2499 11115 2505
rect 11057 2496 11069 2499
rect 10735 2468 11069 2496
rect 10735 2465 10747 2468
rect 10689 2459 10747 2465
rect 11057 2465 11069 2468
rect 11103 2496 11115 2499
rect 12345 2499 12403 2505
rect 12345 2496 12357 2499
rect 11103 2468 12357 2496
rect 11103 2465 11115 2468
rect 11057 2459 11115 2465
rect 12345 2465 12357 2468
rect 12391 2496 12403 2499
rect 12434 2496 12440 2508
rect 12391 2468 12440 2496
rect 12391 2465 12403 2468
rect 12345 2459 12403 2465
rect 12434 2456 12440 2468
rect 12492 2456 12498 2508
rect 12618 2496 12624 2508
rect 12579 2468 12624 2496
rect 12618 2456 12624 2468
rect 12676 2456 12682 2508
rect 15838 2496 15844 2508
rect 12728 2468 13814 2496
rect 5215 2400 8524 2428
rect 5215 2397 5227 2400
rect 5169 2391 5227 2397
rect 106 2320 112 2372
rect 164 2360 170 2372
rect 7009 2363 7067 2369
rect 7009 2360 7021 2363
rect 164 2332 7021 2360
rect 164 2320 170 2332
rect 7009 2329 7021 2332
rect 7055 2329 7067 2363
rect 7009 2323 7067 2329
rect 2498 2292 2504 2304
rect 2459 2264 2504 2292
rect 2498 2252 2504 2264
rect 2556 2252 2562 2304
rect 6270 2292 6276 2304
rect 6231 2264 6276 2292
rect 6270 2252 6276 2264
rect 6328 2252 6334 2304
rect 6638 2292 6644 2304
rect 6599 2264 6644 2292
rect 6638 2252 6644 2264
rect 6696 2252 6702 2304
rect 8496 2292 8524 2400
rect 8754 2388 8760 2440
rect 8812 2428 8818 2440
rect 11977 2431 12035 2437
rect 11977 2428 11989 2431
rect 8812 2400 11989 2428
rect 8812 2388 8818 2400
rect 11977 2397 11989 2400
rect 12023 2428 12035 2431
rect 12728 2428 12756 2468
rect 12023 2400 12756 2428
rect 13786 2428 13814 2468
rect 15120 2468 15844 2496
rect 14182 2428 14188 2440
rect 13786 2400 14188 2428
rect 12023 2397 12035 2400
rect 11977 2391 12035 2397
rect 14182 2388 14188 2400
rect 14240 2388 14246 2440
rect 8849 2363 8907 2369
rect 8849 2329 8861 2363
rect 8895 2360 8907 2363
rect 15120 2360 15148 2468
rect 15838 2456 15844 2468
rect 15896 2456 15902 2508
rect 15930 2456 15936 2508
rect 15988 2496 15994 2508
rect 16025 2499 16083 2505
rect 16025 2496 16037 2499
rect 15988 2468 16037 2496
rect 15988 2456 15994 2468
rect 16025 2465 16037 2468
rect 16071 2496 16083 2499
rect 16390 2496 16396 2508
rect 16071 2468 16396 2496
rect 16071 2465 16083 2468
rect 16025 2459 16083 2465
rect 16390 2456 16396 2468
rect 16448 2456 16454 2508
rect 16776 2505 16804 2536
rect 17218 2524 17224 2536
rect 17276 2524 17282 2576
rect 17770 2564 17776 2576
rect 17683 2536 17776 2564
rect 17770 2524 17776 2536
rect 17828 2564 17834 2576
rect 17828 2536 18460 2564
rect 17828 2524 17834 2536
rect 18432 2508 18460 2536
rect 16761 2499 16819 2505
rect 16761 2465 16773 2499
rect 16807 2465 16819 2499
rect 16761 2459 16819 2465
rect 16853 2499 16911 2505
rect 16853 2465 16865 2499
rect 16899 2465 16911 2499
rect 16853 2459 16911 2465
rect 18141 2499 18199 2505
rect 18141 2465 18153 2499
rect 18187 2496 18199 2499
rect 18322 2496 18328 2508
rect 18187 2468 18328 2496
rect 18187 2465 18199 2468
rect 18141 2459 18199 2465
rect 16868 2428 16896 2459
rect 18322 2456 18328 2468
rect 18380 2456 18386 2508
rect 18414 2456 18420 2508
rect 18472 2496 18478 2508
rect 18598 2496 18604 2508
rect 18472 2468 18517 2496
rect 18559 2468 18604 2496
rect 18472 2456 18478 2468
rect 18598 2456 18604 2468
rect 18656 2456 18662 2508
rect 18800 2496 18828 2604
rect 18966 2592 18972 2644
rect 19024 2632 19030 2644
rect 20073 2635 20131 2641
rect 20073 2632 20085 2635
rect 19024 2604 20085 2632
rect 19024 2592 19030 2604
rect 20073 2601 20085 2604
rect 20119 2601 20131 2635
rect 20530 2632 20536 2644
rect 20491 2604 20536 2632
rect 20073 2595 20131 2601
rect 20530 2592 20536 2604
rect 20588 2592 20594 2644
rect 20622 2592 20628 2644
rect 20680 2632 20686 2644
rect 21082 2632 21088 2644
rect 20680 2604 21088 2632
rect 20680 2592 20686 2604
rect 21082 2592 21088 2604
rect 21140 2632 21146 2644
rect 22189 2635 22247 2641
rect 22189 2632 22201 2635
rect 21140 2604 22201 2632
rect 21140 2592 21146 2604
rect 22189 2601 22201 2604
rect 22235 2601 22247 2635
rect 22189 2595 22247 2601
rect 22879 2635 22937 2641
rect 22879 2601 22891 2635
rect 22925 2632 22937 2635
rect 23474 2632 23480 2644
rect 22925 2604 23480 2632
rect 22925 2601 22937 2604
rect 22879 2595 22937 2601
rect 23474 2592 23480 2604
rect 23532 2592 23538 2644
rect 24578 2592 24584 2644
rect 24636 2632 24642 2644
rect 25409 2635 25467 2641
rect 25409 2632 25421 2635
rect 24636 2604 25421 2632
rect 24636 2592 24642 2604
rect 25409 2601 25421 2604
rect 25455 2601 25467 2635
rect 25409 2595 25467 2601
rect 26605 2635 26663 2641
rect 26605 2601 26617 2635
rect 26651 2632 26663 2635
rect 26786 2632 26792 2644
rect 26651 2604 26792 2632
rect 26651 2601 26663 2604
rect 26605 2595 26663 2601
rect 19978 2524 19984 2576
rect 20036 2564 20042 2576
rect 20901 2567 20959 2573
rect 20901 2564 20913 2567
rect 20036 2536 20913 2564
rect 20036 2524 20042 2536
rect 20901 2533 20913 2536
rect 20947 2564 20959 2567
rect 24026 2564 24032 2576
rect 20947 2536 21312 2564
rect 23987 2536 24032 2564
rect 20947 2533 20959 2536
rect 20901 2527 20959 2533
rect 19705 2499 19763 2505
rect 19705 2496 19717 2499
rect 18800 2468 19717 2496
rect 19705 2465 19717 2468
rect 19751 2465 19763 2499
rect 19705 2459 19763 2465
rect 19889 2499 19947 2505
rect 19889 2465 19901 2499
rect 19935 2465 19947 2499
rect 21082 2496 21088 2508
rect 21043 2468 21088 2496
rect 19889 2459 19947 2465
rect 8895 2332 15148 2360
rect 15212 2400 16896 2428
rect 8895 2329 8907 2332
rect 8849 2323 8907 2329
rect 15212 2304 15240 2400
rect 16942 2388 16948 2440
rect 17000 2428 17006 2440
rect 18785 2431 18843 2437
rect 18785 2428 18797 2431
rect 17000 2400 18797 2428
rect 17000 2388 17006 2400
rect 18785 2397 18797 2400
rect 18831 2397 18843 2431
rect 18785 2391 18843 2397
rect 16114 2320 16120 2372
rect 16172 2360 16178 2372
rect 19904 2360 19932 2459
rect 21082 2456 21088 2468
rect 21140 2456 21146 2508
rect 21284 2505 21312 2536
rect 24026 2524 24032 2536
rect 24084 2524 24090 2576
rect 25424 2564 25452 2595
rect 26786 2592 26792 2604
rect 26844 2592 26850 2644
rect 27338 2632 27344 2644
rect 27299 2604 27344 2632
rect 27338 2592 27344 2604
rect 27396 2592 27402 2644
rect 28905 2635 28963 2641
rect 28905 2632 28917 2635
rect 27908 2604 28917 2632
rect 25424 2536 26959 2564
rect 21269 2499 21327 2505
rect 21269 2465 21281 2499
rect 21315 2465 21327 2499
rect 21269 2459 21327 2465
rect 21453 2499 21511 2505
rect 21453 2465 21465 2499
rect 21499 2465 21511 2499
rect 21453 2459 21511 2465
rect 20530 2388 20536 2440
rect 20588 2428 20594 2440
rect 21468 2428 21496 2459
rect 22646 2456 22652 2508
rect 22704 2496 22710 2508
rect 22776 2499 22834 2505
rect 22776 2496 22788 2499
rect 22704 2468 22788 2496
rect 22704 2456 22710 2468
rect 22776 2465 22788 2468
rect 22822 2496 22834 2499
rect 23201 2499 23259 2505
rect 23201 2496 23213 2499
rect 22822 2468 23213 2496
rect 22822 2465 22834 2468
rect 22776 2459 22834 2465
rect 23201 2465 23213 2468
rect 23247 2465 23259 2499
rect 23201 2459 23259 2465
rect 23845 2499 23903 2505
rect 23845 2465 23857 2499
rect 23891 2496 23903 2499
rect 24210 2496 24216 2508
rect 23891 2468 24216 2496
rect 23891 2465 23903 2468
rect 23845 2459 23903 2465
rect 24210 2456 24216 2468
rect 24268 2496 24274 2508
rect 24673 2499 24731 2505
rect 24673 2496 24685 2499
rect 24268 2468 24685 2496
rect 24268 2456 24274 2468
rect 24673 2465 24685 2468
rect 24719 2496 24731 2499
rect 25041 2499 25099 2505
rect 25041 2496 25053 2499
rect 24719 2468 25053 2496
rect 24719 2465 24731 2468
rect 24673 2459 24731 2465
rect 25041 2465 25053 2468
rect 25087 2465 25099 2499
rect 25590 2496 25596 2508
rect 25551 2468 25596 2496
rect 25041 2459 25099 2465
rect 25590 2456 25596 2468
rect 25648 2496 25654 2508
rect 26931 2505 26959 2536
rect 26145 2499 26203 2505
rect 26145 2496 26157 2499
rect 25648 2468 26157 2496
rect 25648 2456 25654 2468
rect 26145 2465 26157 2468
rect 26191 2496 26203 2499
rect 26697 2499 26755 2505
rect 26697 2496 26709 2499
rect 26191 2468 26709 2496
rect 26191 2465 26203 2468
rect 26145 2459 26203 2465
rect 26697 2465 26709 2468
rect 26743 2465 26755 2499
rect 26697 2459 26755 2465
rect 26916 2499 26974 2505
rect 26916 2465 26928 2499
rect 26962 2465 26974 2499
rect 26916 2459 26974 2465
rect 27246 2456 27252 2508
rect 27304 2496 27310 2508
rect 27908 2505 27936 2604
rect 28905 2601 28917 2604
rect 28951 2601 28963 2635
rect 29270 2632 29276 2644
rect 29231 2604 29276 2632
rect 28905 2595 28963 2601
rect 29270 2592 29276 2604
rect 29328 2592 29334 2644
rect 29914 2632 29920 2644
rect 29875 2604 29920 2632
rect 29914 2592 29920 2604
rect 29972 2592 29978 2644
rect 30190 2592 30196 2644
rect 30248 2632 30254 2644
rect 32398 2632 32404 2644
rect 30248 2604 32404 2632
rect 30248 2592 30254 2604
rect 32398 2592 32404 2604
rect 32456 2592 32462 2644
rect 28629 2567 28687 2573
rect 28629 2533 28641 2567
rect 28675 2564 28687 2567
rect 28810 2564 28816 2576
rect 28675 2536 28816 2564
rect 28675 2533 28687 2536
rect 28629 2527 28687 2533
rect 28810 2524 28816 2536
rect 28868 2524 28874 2576
rect 29932 2564 29960 2592
rect 28920 2536 29960 2564
rect 27893 2499 27951 2505
rect 27893 2496 27905 2499
rect 27304 2468 27905 2496
rect 27304 2456 27310 2468
rect 27893 2465 27905 2468
rect 27939 2465 27951 2499
rect 28442 2496 28448 2508
rect 28355 2468 28448 2496
rect 27893 2459 27951 2465
rect 28442 2456 28448 2468
rect 28500 2496 28506 2508
rect 28920 2496 28948 2536
rect 28500 2468 28948 2496
rect 29733 2499 29791 2505
rect 28500 2456 28506 2468
rect 29733 2465 29745 2499
rect 29779 2465 29791 2499
rect 29733 2459 29791 2465
rect 30812 2499 30870 2505
rect 30812 2465 30824 2499
rect 30858 2496 30870 2499
rect 30858 2468 31064 2496
rect 30858 2465 30870 2468
rect 30812 2459 30870 2465
rect 20588 2400 21496 2428
rect 21913 2431 21971 2437
rect 20588 2388 20594 2400
rect 21913 2397 21925 2431
rect 21959 2428 21971 2431
rect 29748 2428 29776 2459
rect 30193 2431 30251 2437
rect 30193 2428 30205 2431
rect 21959 2400 30205 2428
rect 21959 2397 21971 2400
rect 21913 2391 21971 2397
rect 30193 2397 30205 2400
rect 30239 2397 30251 2431
rect 30193 2391 30251 2397
rect 25777 2363 25835 2369
rect 16172 2332 21036 2360
rect 16172 2320 16178 2332
rect 9030 2292 9036 2304
rect 8496 2264 9036 2292
rect 9030 2252 9036 2264
rect 9088 2252 9094 2304
rect 9214 2292 9220 2304
rect 9175 2264 9220 2292
rect 9214 2252 9220 2264
rect 9272 2252 9278 2304
rect 10134 2292 10140 2304
rect 10095 2264 10140 2292
rect 10134 2252 10140 2264
rect 10192 2252 10198 2304
rect 10226 2252 10232 2304
rect 10284 2292 10290 2304
rect 10689 2295 10747 2301
rect 10689 2292 10701 2295
rect 10284 2264 10701 2292
rect 10284 2252 10290 2264
rect 10689 2261 10701 2264
rect 10735 2292 10747 2295
rect 10781 2295 10839 2301
rect 10781 2292 10793 2295
rect 10735 2264 10793 2292
rect 10735 2261 10747 2264
rect 10689 2255 10747 2261
rect 10781 2261 10793 2264
rect 10827 2261 10839 2295
rect 13630 2292 13636 2304
rect 13591 2264 13636 2292
rect 10781 2255 10839 2261
rect 13630 2252 13636 2264
rect 13688 2292 13694 2304
rect 13955 2295 14013 2301
rect 13955 2292 13967 2295
rect 13688 2264 13967 2292
rect 13688 2252 13694 2264
rect 13955 2261 13967 2264
rect 14001 2261 14013 2295
rect 13955 2255 14013 2261
rect 14090 2252 14096 2304
rect 14148 2292 14154 2304
rect 15194 2292 15200 2304
rect 14148 2264 14193 2292
rect 15155 2264 15200 2292
rect 14148 2252 14154 2264
rect 15194 2252 15200 2264
rect 15252 2252 15258 2304
rect 16390 2252 16396 2304
rect 16448 2292 16454 2304
rect 18322 2292 18328 2304
rect 16448 2264 18328 2292
rect 16448 2252 16454 2264
rect 18322 2252 18328 2264
rect 18380 2252 18386 2304
rect 18598 2252 18604 2304
rect 18656 2292 18662 2304
rect 19337 2295 19395 2301
rect 19337 2292 19349 2295
rect 18656 2264 19349 2292
rect 18656 2252 18662 2264
rect 19337 2261 19349 2264
rect 19383 2261 19395 2295
rect 21008 2292 21036 2332
rect 25777 2329 25789 2363
rect 25823 2360 25835 2363
rect 26786 2360 26792 2372
rect 25823 2332 26792 2360
rect 25823 2329 25835 2332
rect 25777 2323 25835 2329
rect 26786 2320 26792 2332
rect 26844 2320 26850 2372
rect 27801 2363 27859 2369
rect 26931 2332 27752 2360
rect 22557 2295 22615 2301
rect 22557 2292 22569 2295
rect 21008 2264 22569 2292
rect 19337 2255 19395 2261
rect 22557 2261 22569 2264
rect 22603 2261 22615 2295
rect 22557 2255 22615 2261
rect 26697 2295 26755 2301
rect 26697 2261 26709 2295
rect 26743 2292 26755 2295
rect 26931 2292 26959 2332
rect 26743 2264 26959 2292
rect 27019 2295 27077 2301
rect 26743 2261 26755 2264
rect 26697 2255 26755 2261
rect 27019 2261 27031 2295
rect 27065 2292 27077 2295
rect 27246 2292 27252 2304
rect 27065 2264 27252 2292
rect 27065 2261 27077 2264
rect 27019 2255 27077 2261
rect 27246 2252 27252 2264
rect 27304 2252 27310 2304
rect 27724 2292 27752 2332
rect 27801 2329 27813 2363
rect 27847 2360 27859 2363
rect 28442 2360 28448 2372
rect 27847 2332 28448 2360
rect 27847 2329 27859 2332
rect 27801 2323 27859 2329
rect 28442 2320 28448 2332
rect 28500 2320 28506 2372
rect 28534 2320 28540 2372
rect 28592 2360 28598 2372
rect 30883 2363 30941 2369
rect 30883 2360 30895 2363
rect 28592 2332 30895 2360
rect 28592 2320 28598 2332
rect 30883 2329 30895 2332
rect 30929 2329 30941 2363
rect 30883 2323 30941 2329
rect 31036 2292 31064 2468
rect 31205 2295 31263 2301
rect 31205 2292 31217 2295
rect 27724 2264 31217 2292
rect 31205 2261 31217 2264
rect 31251 2261 31263 2295
rect 31205 2255 31263 2261
rect 1104 2202 38824 2224
rect 1104 2150 7648 2202
rect 7700 2150 7712 2202
rect 7764 2150 7776 2202
rect 7828 2150 7840 2202
rect 7892 2150 20982 2202
rect 21034 2150 21046 2202
rect 21098 2150 21110 2202
rect 21162 2150 21174 2202
rect 21226 2150 34315 2202
rect 34367 2150 34379 2202
rect 34431 2150 34443 2202
rect 34495 2150 34507 2202
rect 34559 2150 38824 2202
rect 1104 2128 38824 2150
rect 5994 2048 6000 2100
rect 6052 2088 6058 2100
rect 13630 2088 13636 2100
rect 6052 2060 13636 2088
rect 6052 2048 6058 2060
rect 13630 2048 13636 2060
rect 13688 2048 13694 2100
rect 6270 1980 6276 2032
rect 6328 2020 6334 2032
rect 7374 2020 7380 2032
rect 6328 1992 7380 2020
rect 6328 1980 6334 1992
rect 7374 1980 7380 1992
rect 7432 2020 7438 2032
rect 8662 2020 8668 2032
rect 7432 1992 8668 2020
rect 7432 1980 7438 1992
rect 8662 1980 8668 1992
rect 8720 1980 8726 2032
rect 10134 1980 10140 2032
rect 10192 2020 10198 2032
rect 14090 2020 14096 2032
rect 10192 1992 14096 2020
rect 10192 1980 10198 1992
rect 14090 1980 14096 1992
rect 14148 1980 14154 2032
rect 7098 76 7104 128
rect 7156 116 7162 128
rect 8478 116 8484 128
rect 7156 88 8484 116
rect 7156 76 7162 88
rect 8478 76 8484 88
rect 8536 76 8542 128
rect 10318 76 10324 128
rect 10376 116 10382 128
rect 12802 116 12808 128
rect 10376 88 12808 116
rect 10376 76 10382 88
rect 12802 76 12808 88
rect 12860 76 12866 128
rect 21358 76 21364 128
rect 21416 116 21422 128
rect 24486 116 24492 128
rect 21416 88 24492 116
rect 21416 76 21422 88
rect 24486 76 24492 88
rect 24544 76 24550 128
<< via1 >>
rect 14315 13574 14367 13626
rect 14379 13574 14431 13626
rect 14443 13574 14495 13626
rect 14507 13574 14559 13626
rect 27648 13574 27700 13626
rect 27712 13574 27764 13626
rect 27776 13574 27828 13626
rect 27840 13574 27892 13626
rect 112 13132 164 13184
rect 28264 13132 28316 13184
rect 7648 13030 7700 13082
rect 7712 13030 7764 13082
rect 7776 13030 7828 13082
rect 7840 13030 7892 13082
rect 20982 13030 21034 13082
rect 21046 13030 21098 13082
rect 21110 13030 21162 13082
rect 21174 13030 21226 13082
rect 34315 13030 34367 13082
rect 34379 13030 34431 13082
rect 34443 13030 34495 13082
rect 34507 13030 34559 13082
rect 19616 12928 19668 12980
rect 28264 12971 28316 12980
rect 28264 12937 28273 12971
rect 28273 12937 28307 12971
rect 28307 12937 28316 12971
rect 28264 12928 28316 12937
rect 34060 12928 34112 12980
rect 35624 12971 35676 12980
rect 35624 12937 35633 12971
rect 35633 12937 35667 12971
rect 35667 12937 35676 12971
rect 35624 12928 35676 12937
rect 8208 12724 8260 12776
rect 8392 12724 8444 12776
rect 28724 12724 28776 12776
rect 31392 12724 31444 12776
rect 34796 12724 34848 12776
rect 12900 12656 12952 12708
rect 16856 12656 16908 12708
rect 39580 12656 39632 12708
rect 112 12588 164 12640
rect 1768 12588 1820 12640
rect 7472 12631 7524 12640
rect 7472 12597 7481 12631
rect 7481 12597 7515 12631
rect 7515 12597 7524 12631
rect 7472 12588 7524 12597
rect 8024 12588 8076 12640
rect 19248 12588 19300 12640
rect 28724 12631 28776 12640
rect 28724 12597 28733 12631
rect 28733 12597 28767 12631
rect 28767 12597 28776 12631
rect 28724 12588 28776 12597
rect 14315 12486 14367 12538
rect 14379 12486 14431 12538
rect 14443 12486 14495 12538
rect 14507 12486 14559 12538
rect 27648 12486 27700 12538
rect 27712 12486 27764 12538
rect 27776 12486 27828 12538
rect 27840 12486 27892 12538
rect 2044 12248 2096 12300
rect 6552 12248 6604 12300
rect 8116 12248 8168 12300
rect 9588 12291 9640 12300
rect 9588 12257 9597 12291
rect 9597 12257 9631 12291
rect 9631 12257 9640 12291
rect 9588 12248 9640 12257
rect 10784 12248 10836 12300
rect 15660 12291 15712 12300
rect 15660 12257 15669 12291
rect 15669 12257 15703 12291
rect 15703 12257 15712 12291
rect 15660 12248 15712 12257
rect 17040 12248 17092 12300
rect 19248 12248 19300 12300
rect 19708 12248 19760 12300
rect 23480 12291 23532 12300
rect 23480 12257 23489 12291
rect 23489 12257 23523 12291
rect 23523 12257 23532 12291
rect 23480 12248 23532 12257
rect 25136 12248 25188 12300
rect 28080 12248 28132 12300
rect 2688 12223 2740 12232
rect 2688 12189 2697 12223
rect 2697 12189 2731 12223
rect 2731 12189 2740 12223
rect 2688 12180 2740 12189
rect 18144 12180 18196 12232
rect 1584 12155 1636 12164
rect 1584 12121 1593 12155
rect 1593 12121 1627 12155
rect 1627 12121 1636 12155
rect 1584 12112 1636 12121
rect 18604 12112 18656 12164
rect 6920 12044 6972 12096
rect 8852 12044 8904 12096
rect 9036 12044 9088 12096
rect 10508 12044 10560 12096
rect 16764 12044 16816 12096
rect 18420 12044 18472 12096
rect 19800 12044 19852 12096
rect 24124 12044 24176 12096
rect 24676 12087 24728 12096
rect 24676 12053 24685 12087
rect 24685 12053 24719 12087
rect 24719 12053 24728 12087
rect 24676 12044 24728 12053
rect 27528 12087 27580 12096
rect 27528 12053 27537 12087
rect 27537 12053 27571 12087
rect 27571 12053 27580 12087
rect 27528 12044 27580 12053
rect 7648 11942 7700 11994
rect 7712 11942 7764 11994
rect 7776 11942 7828 11994
rect 7840 11942 7892 11994
rect 20982 11942 21034 11994
rect 21046 11942 21098 11994
rect 21110 11942 21162 11994
rect 21174 11942 21226 11994
rect 34315 11942 34367 11994
rect 34379 11942 34431 11994
rect 34443 11942 34495 11994
rect 34507 11942 34559 11994
rect 1124 11840 1176 11892
rect 1952 11840 2004 11892
rect 4804 11840 4856 11892
rect 17040 11883 17092 11892
rect 17040 11849 17049 11883
rect 17049 11849 17083 11883
rect 17083 11849 17092 11883
rect 23020 11883 23072 11892
rect 17040 11840 17092 11849
rect 1676 11772 1728 11824
rect 6552 11815 6604 11824
rect 6552 11781 6561 11815
rect 6561 11781 6595 11815
rect 6595 11781 6604 11815
rect 6552 11772 6604 11781
rect 19708 11772 19760 11824
rect 2044 11747 2096 11756
rect 2044 11713 2053 11747
rect 2053 11713 2087 11747
rect 2087 11713 2096 11747
rect 2044 11704 2096 11713
rect 4528 11704 4580 11756
rect 9588 11704 9640 11756
rect 9864 11747 9916 11756
rect 9864 11713 9873 11747
rect 9873 11713 9907 11747
rect 9907 11713 9916 11747
rect 9864 11704 9916 11713
rect 15660 11704 15712 11756
rect 20352 11704 20404 11756
rect 7012 11679 7064 11688
rect 7012 11645 7021 11679
rect 7021 11645 7055 11679
rect 7055 11645 7064 11679
rect 7012 11636 7064 11645
rect 6276 11611 6328 11620
rect 6276 11577 6285 11611
rect 6285 11577 6319 11611
rect 6319 11577 6328 11611
rect 7472 11636 7524 11688
rect 9128 11636 9180 11688
rect 9312 11636 9364 11688
rect 11796 11636 11848 11688
rect 18236 11679 18288 11688
rect 18236 11645 18245 11679
rect 18245 11645 18279 11679
rect 18279 11645 18288 11679
rect 18236 11636 18288 11645
rect 18696 11679 18748 11688
rect 18696 11645 18705 11679
rect 18705 11645 18739 11679
rect 18739 11645 18748 11679
rect 18696 11636 18748 11645
rect 6276 11568 6328 11577
rect 17224 11568 17276 11620
rect 22376 11636 22428 11688
rect 23020 11849 23029 11883
rect 23029 11849 23063 11883
rect 23063 11849 23072 11883
rect 23020 11840 23072 11849
rect 35624 11883 35676 11892
rect 35624 11849 35633 11883
rect 35633 11849 35667 11883
rect 35667 11849 35676 11883
rect 35624 11840 35676 11849
rect 24400 11772 24452 11824
rect 26332 11704 26384 11756
rect 35440 11679 35492 11688
rect 21640 11568 21692 11620
rect 35440 11645 35449 11679
rect 35449 11645 35483 11679
rect 35483 11645 35492 11679
rect 35440 11636 35492 11645
rect 30932 11568 30984 11620
rect 2964 11500 3016 11552
rect 7104 11543 7156 11552
rect 7104 11509 7113 11543
rect 7113 11509 7147 11543
rect 7147 11509 7156 11543
rect 7104 11500 7156 11509
rect 8116 11500 8168 11552
rect 8668 11500 8720 11552
rect 8944 11500 8996 11552
rect 10324 11500 10376 11552
rect 10784 11500 10836 11552
rect 11796 11500 11848 11552
rect 14188 11500 14240 11552
rect 14832 11543 14884 11552
rect 14832 11509 14841 11543
rect 14841 11509 14875 11543
rect 14875 11509 14884 11543
rect 14832 11500 14884 11509
rect 17408 11500 17460 11552
rect 17960 11500 18012 11552
rect 19064 11500 19116 11552
rect 19248 11543 19300 11552
rect 19248 11509 19257 11543
rect 19257 11509 19291 11543
rect 19291 11509 19300 11543
rect 19248 11500 19300 11509
rect 19984 11500 20036 11552
rect 22928 11500 22980 11552
rect 23480 11500 23532 11552
rect 24308 11500 24360 11552
rect 25136 11500 25188 11552
rect 27344 11543 27396 11552
rect 27344 11509 27353 11543
rect 27353 11509 27387 11543
rect 27387 11509 27396 11543
rect 27344 11500 27396 11509
rect 28080 11500 28132 11552
rect 14315 11398 14367 11450
rect 14379 11398 14431 11450
rect 14443 11398 14495 11450
rect 14507 11398 14559 11450
rect 27648 11398 27700 11450
rect 27712 11398 27764 11450
rect 27776 11398 27828 11450
rect 27840 11398 27892 11450
rect 1676 11339 1728 11348
rect 1676 11305 1685 11339
rect 1685 11305 1719 11339
rect 1719 11305 1728 11339
rect 1676 11296 1728 11305
rect 5448 11296 5500 11348
rect 8576 11296 8628 11348
rect 8852 11339 8904 11348
rect 8852 11305 8861 11339
rect 8861 11305 8895 11339
rect 8895 11305 8904 11339
rect 8852 11296 8904 11305
rect 7196 11228 7248 11280
rect 14648 11228 14700 11280
rect 16856 11296 16908 11348
rect 19064 11296 19116 11348
rect 22928 11296 22980 11348
rect 23848 11296 23900 11348
rect 24492 11339 24544 11348
rect 24492 11305 24501 11339
rect 24501 11305 24535 11339
rect 24535 11305 24544 11339
rect 24492 11296 24544 11305
rect 37740 11296 37792 11348
rect 17500 11228 17552 11280
rect 17592 11228 17644 11280
rect 23020 11228 23072 11280
rect 2412 11203 2464 11212
rect 2412 11169 2421 11203
rect 2421 11169 2455 11203
rect 2455 11169 2464 11203
rect 2412 11160 2464 11169
rect 2872 11160 2924 11212
rect 4712 11160 4764 11212
rect 6184 11203 6236 11212
rect 2780 11135 2832 11144
rect 2780 11101 2789 11135
rect 2789 11101 2823 11135
rect 2823 11101 2832 11135
rect 2780 11092 2832 11101
rect 6184 11169 6193 11203
rect 6193 11169 6227 11203
rect 6227 11169 6236 11203
rect 6184 11160 6236 11169
rect 9588 11160 9640 11212
rect 9864 11160 9916 11212
rect 10968 11160 11020 11212
rect 13912 11160 13964 11212
rect 15844 11160 15896 11212
rect 16488 11160 16540 11212
rect 19340 11203 19392 11212
rect 19340 11169 19349 11203
rect 19349 11169 19383 11203
rect 19383 11169 19392 11203
rect 19340 11160 19392 11169
rect 8668 11092 8720 11144
rect 12256 11092 12308 11144
rect 18696 11092 18748 11144
rect 19800 11160 19852 11212
rect 19984 11160 20036 11212
rect 23480 11160 23532 11212
rect 24860 11160 24912 11212
rect 25228 11160 25280 11212
rect 26424 11203 26476 11212
rect 26424 11169 26433 11203
rect 26433 11169 26467 11203
rect 26467 11169 26476 11203
rect 26424 11160 26476 11169
rect 28632 11203 28684 11212
rect 23020 11092 23072 11144
rect 6368 11024 6420 11076
rect 7012 11024 7064 11076
rect 8484 11067 8536 11076
rect 3148 10999 3200 11008
rect 3148 10965 3157 10999
rect 3157 10965 3191 10999
rect 3191 10965 3200 10999
rect 3148 10956 3200 10965
rect 7196 10999 7248 11008
rect 7196 10965 7205 10999
rect 7205 10965 7239 10999
rect 7239 10965 7248 10999
rect 7196 10956 7248 10965
rect 8484 11033 8493 11067
rect 8493 11033 8527 11067
rect 8527 11033 8536 11067
rect 8484 11024 8536 11033
rect 10232 11024 10284 11076
rect 16396 11024 16448 11076
rect 21272 11024 21324 11076
rect 26976 11092 27028 11144
rect 28632 11169 28641 11203
rect 28641 11169 28675 11203
rect 28675 11169 28684 11203
rect 28632 11160 28684 11169
rect 30932 11203 30984 11212
rect 30932 11169 30941 11203
rect 30941 11169 30975 11203
rect 30975 11169 30984 11203
rect 30932 11160 30984 11169
rect 32588 11160 32640 11212
rect 32680 11160 32732 11212
rect 28540 11092 28592 11144
rect 28908 11135 28960 11144
rect 28908 11101 28917 11135
rect 28917 11101 28951 11135
rect 28951 11101 28960 11135
rect 28908 11092 28960 11101
rect 24216 11024 24268 11076
rect 9680 10956 9732 11008
rect 11888 10956 11940 11008
rect 12440 10956 12492 11008
rect 12624 10999 12676 11008
rect 12624 10965 12633 10999
rect 12633 10965 12667 10999
rect 12667 10965 12676 10999
rect 12624 10956 12676 10965
rect 13544 10956 13596 11008
rect 16028 10999 16080 11008
rect 16028 10965 16037 10999
rect 16037 10965 16071 10999
rect 16071 10965 16080 10999
rect 16028 10956 16080 10965
rect 17776 10956 17828 11008
rect 18236 10999 18288 11008
rect 18236 10965 18245 10999
rect 18245 10965 18279 10999
rect 18279 10965 18288 10999
rect 18236 10956 18288 10965
rect 20168 10956 20220 11008
rect 23296 10956 23348 11008
rect 25872 10999 25924 11008
rect 25872 10965 25881 10999
rect 25881 10965 25915 10999
rect 25915 10965 25924 10999
rect 25872 10956 25924 10965
rect 27068 10956 27120 11008
rect 27712 10999 27764 11008
rect 27712 10965 27721 10999
rect 27721 10965 27755 10999
rect 27755 10965 27764 10999
rect 27712 10956 27764 10965
rect 29276 10999 29328 11008
rect 29276 10965 29285 10999
rect 29285 10965 29319 10999
rect 29319 10965 29328 10999
rect 29276 10956 29328 10965
rect 31576 10956 31628 11008
rect 31668 10956 31720 11008
rect 7648 10854 7700 10906
rect 7712 10854 7764 10906
rect 7776 10854 7828 10906
rect 7840 10854 7892 10906
rect 20982 10854 21034 10906
rect 21046 10854 21098 10906
rect 21110 10854 21162 10906
rect 21174 10854 21226 10906
rect 34315 10854 34367 10906
rect 34379 10854 34431 10906
rect 34443 10854 34495 10906
rect 34507 10854 34559 10906
rect 6368 10752 6420 10804
rect 6552 10752 6604 10804
rect 9588 10752 9640 10804
rect 10968 10795 11020 10804
rect 10968 10761 10977 10795
rect 10977 10761 11011 10795
rect 11011 10761 11020 10795
rect 10968 10752 11020 10761
rect 21272 10752 21324 10804
rect 2872 10727 2924 10736
rect 2872 10693 2881 10727
rect 2881 10693 2915 10727
rect 2915 10693 2924 10727
rect 2872 10684 2924 10693
rect 2688 10616 2740 10668
rect 3056 10659 3108 10668
rect 3056 10625 3065 10659
rect 3065 10625 3099 10659
rect 3099 10625 3108 10659
rect 3056 10616 3108 10625
rect 4160 10684 4212 10736
rect 6276 10616 6328 10668
rect 6920 10616 6972 10668
rect 7932 10616 7984 10668
rect 8852 10616 8904 10668
rect 11888 10684 11940 10736
rect 13912 10727 13964 10736
rect 13912 10693 13921 10727
rect 13921 10693 13955 10727
rect 13955 10693 13964 10727
rect 13912 10684 13964 10693
rect 16028 10684 16080 10736
rect 16304 10684 16356 10736
rect 19800 10684 19852 10736
rect 22836 10684 22888 10736
rect 13636 10616 13688 10668
rect 1584 10591 1636 10600
rect 1584 10557 1593 10591
rect 1593 10557 1627 10591
rect 1627 10557 1636 10591
rect 1584 10548 1636 10557
rect 2872 10548 2924 10600
rect 5632 10591 5684 10600
rect 2136 10523 2188 10532
rect 2136 10489 2145 10523
rect 2145 10489 2179 10523
rect 2179 10489 2188 10523
rect 2136 10480 2188 10489
rect 3148 10523 3200 10532
rect 3148 10489 3157 10523
rect 3157 10489 3191 10523
rect 3191 10489 3200 10523
rect 3148 10480 3200 10489
rect 5632 10557 5641 10591
rect 5641 10557 5675 10591
rect 5675 10557 5684 10591
rect 5632 10548 5684 10557
rect 6184 10548 6236 10600
rect 1676 10412 1728 10464
rect 2412 10455 2464 10464
rect 2412 10421 2421 10455
rect 2421 10421 2455 10455
rect 2455 10421 2464 10455
rect 2412 10412 2464 10421
rect 4712 10455 4764 10464
rect 4712 10421 4721 10455
rect 4721 10421 4755 10455
rect 4755 10421 4764 10455
rect 4712 10412 4764 10421
rect 5080 10412 5132 10464
rect 6092 10480 6144 10532
rect 7196 10523 7248 10532
rect 7196 10489 7205 10523
rect 7205 10489 7239 10523
rect 7239 10489 7248 10523
rect 7196 10480 7248 10489
rect 7012 10412 7064 10464
rect 8392 10455 8444 10464
rect 8392 10421 8401 10455
rect 8401 10421 8435 10455
rect 8435 10421 8444 10455
rect 8392 10412 8444 10421
rect 9772 10412 9824 10464
rect 10968 10548 11020 10600
rect 11888 10591 11940 10600
rect 11888 10557 11897 10591
rect 11897 10557 11931 10591
rect 11931 10557 11940 10591
rect 11888 10548 11940 10557
rect 12256 10548 12308 10600
rect 12624 10548 12676 10600
rect 14096 10591 14148 10600
rect 14096 10557 14105 10591
rect 14105 10557 14139 10591
rect 14139 10557 14148 10591
rect 14648 10591 14700 10600
rect 14096 10548 14148 10557
rect 14648 10557 14657 10591
rect 14657 10557 14691 10591
rect 14691 10557 14700 10591
rect 14648 10548 14700 10557
rect 16672 10616 16724 10668
rect 13268 10523 13320 10532
rect 13268 10489 13277 10523
rect 13277 10489 13311 10523
rect 13311 10489 13320 10523
rect 13268 10480 13320 10489
rect 18880 10548 18932 10600
rect 19432 10548 19484 10600
rect 20168 10659 20220 10668
rect 20168 10625 20177 10659
rect 20177 10625 20211 10659
rect 20211 10625 20220 10659
rect 20168 10616 20220 10625
rect 22376 10548 22428 10600
rect 22560 10591 22612 10600
rect 26424 10752 26476 10804
rect 32588 10795 32640 10804
rect 32588 10761 32597 10795
rect 32597 10761 32631 10795
rect 32631 10761 32640 10795
rect 32588 10752 32640 10761
rect 35440 10752 35492 10804
rect 28816 10684 28868 10736
rect 29276 10684 29328 10736
rect 23848 10659 23900 10668
rect 23848 10625 23857 10659
rect 23857 10625 23891 10659
rect 23891 10625 23900 10659
rect 23848 10616 23900 10625
rect 24676 10616 24728 10668
rect 22560 10557 22604 10591
rect 22604 10557 22612 10591
rect 22560 10548 22612 10557
rect 24860 10591 24912 10600
rect 24860 10557 24869 10591
rect 24869 10557 24903 10591
rect 24903 10557 24912 10591
rect 24860 10548 24912 10557
rect 25412 10548 25464 10600
rect 25504 10548 25556 10600
rect 25872 10548 25924 10600
rect 26056 10591 26108 10600
rect 26056 10557 26065 10591
rect 26065 10557 26099 10591
rect 26099 10557 26108 10591
rect 26056 10548 26108 10557
rect 10784 10412 10836 10464
rect 11060 10412 11112 10464
rect 13820 10412 13872 10464
rect 14924 10412 14976 10464
rect 16028 10480 16080 10532
rect 16488 10480 16540 10532
rect 19248 10523 19300 10532
rect 19248 10489 19257 10523
rect 19257 10489 19291 10523
rect 19291 10489 19300 10523
rect 19248 10480 19300 10489
rect 20168 10480 20220 10532
rect 20812 10523 20864 10532
rect 20812 10489 20821 10523
rect 20821 10489 20855 10523
rect 20855 10489 20864 10523
rect 20812 10480 20864 10489
rect 22468 10480 22520 10532
rect 23940 10523 23992 10532
rect 15844 10412 15896 10464
rect 16120 10455 16172 10464
rect 16120 10421 16129 10455
rect 16129 10421 16163 10455
rect 16163 10421 16172 10455
rect 16120 10412 16172 10421
rect 16672 10455 16724 10464
rect 16672 10421 16681 10455
rect 16681 10421 16715 10455
rect 16715 10421 16724 10455
rect 16672 10412 16724 10421
rect 17776 10455 17828 10464
rect 17776 10421 17785 10455
rect 17785 10421 17819 10455
rect 17819 10421 17828 10455
rect 17776 10412 17828 10421
rect 19340 10412 19392 10464
rect 22928 10412 22980 10464
rect 23480 10455 23532 10464
rect 23480 10421 23489 10455
rect 23489 10421 23523 10455
rect 23523 10421 23532 10455
rect 23940 10489 23949 10523
rect 23949 10489 23983 10523
rect 23983 10489 23992 10523
rect 23940 10480 23992 10489
rect 24584 10480 24636 10532
rect 27528 10548 27580 10600
rect 27712 10548 27764 10600
rect 28816 10548 28868 10600
rect 30932 10684 30984 10736
rect 35256 10684 35308 10736
rect 31668 10659 31720 10668
rect 31668 10625 31677 10659
rect 31677 10625 31711 10659
rect 31711 10625 31720 10659
rect 31668 10616 31720 10625
rect 32680 10616 32732 10668
rect 35900 10548 35952 10600
rect 26332 10523 26384 10532
rect 26332 10489 26341 10523
rect 26341 10489 26375 10523
rect 26375 10489 26384 10523
rect 26332 10480 26384 10489
rect 29828 10480 29880 10532
rect 30012 10523 30064 10532
rect 30012 10489 30021 10523
rect 30021 10489 30055 10523
rect 30055 10489 30064 10523
rect 30012 10480 30064 10489
rect 31484 10523 31536 10532
rect 31484 10489 31493 10523
rect 31493 10489 31527 10523
rect 31527 10489 31536 10523
rect 31484 10480 31536 10489
rect 32496 10480 32548 10532
rect 23480 10412 23532 10421
rect 24768 10412 24820 10464
rect 25228 10412 25280 10464
rect 28632 10412 28684 10464
rect 29644 10412 29696 10464
rect 33508 10412 33560 10464
rect 14315 10310 14367 10362
rect 14379 10310 14431 10362
rect 14443 10310 14495 10362
rect 14507 10310 14559 10362
rect 27648 10310 27700 10362
rect 27712 10310 27764 10362
rect 27776 10310 27828 10362
rect 27840 10310 27892 10362
rect 1584 10208 1636 10260
rect 2228 10251 2280 10260
rect 2228 10217 2237 10251
rect 2237 10217 2271 10251
rect 2271 10217 2280 10251
rect 2228 10208 2280 10217
rect 3056 10208 3108 10260
rect 5724 10251 5776 10260
rect 5724 10217 5733 10251
rect 5733 10217 5767 10251
rect 5767 10217 5776 10251
rect 5724 10208 5776 10217
rect 7104 10251 7156 10260
rect 7104 10217 7113 10251
rect 7113 10217 7147 10251
rect 7147 10217 7156 10251
rect 7104 10208 7156 10217
rect 8668 10251 8720 10260
rect 8668 10217 8677 10251
rect 8677 10217 8711 10251
rect 8711 10217 8720 10251
rect 8668 10208 8720 10217
rect 10968 10208 11020 10260
rect 12440 10208 12492 10260
rect 13728 10251 13780 10260
rect 13728 10217 13737 10251
rect 13737 10217 13771 10251
rect 13771 10217 13780 10251
rect 13728 10208 13780 10217
rect 16580 10208 16632 10260
rect 17960 10251 18012 10260
rect 17960 10217 17969 10251
rect 17969 10217 18003 10251
rect 18003 10217 18012 10251
rect 17960 10208 18012 10217
rect 22744 10251 22796 10260
rect 22744 10217 22753 10251
rect 22753 10217 22787 10251
rect 22787 10217 22796 10251
rect 22744 10208 22796 10217
rect 27068 10251 27120 10260
rect 27068 10217 27077 10251
rect 27077 10217 27111 10251
rect 27111 10217 27120 10251
rect 27068 10208 27120 10217
rect 31668 10251 31720 10260
rect 31668 10217 31677 10251
rect 31677 10217 31711 10251
rect 31711 10217 31720 10251
rect 31668 10208 31720 10217
rect 2044 10140 2096 10192
rect 3976 10140 4028 10192
rect 6920 10140 6972 10192
rect 8208 10140 8260 10192
rect 9772 10183 9824 10192
rect 9772 10149 9781 10183
rect 9781 10149 9815 10183
rect 9815 10149 9824 10183
rect 9772 10140 9824 10149
rect 9864 10183 9916 10192
rect 9864 10149 9873 10183
rect 9873 10149 9907 10183
rect 9907 10149 9916 10183
rect 9864 10140 9916 10149
rect 15384 10140 15436 10192
rect 18236 10183 18288 10192
rect 18236 10149 18245 10183
rect 18245 10149 18279 10183
rect 18279 10149 18288 10183
rect 18236 10140 18288 10149
rect 21272 10140 21324 10192
rect 23940 10140 23992 10192
rect 27344 10140 27396 10192
rect 27712 10183 27764 10192
rect 27712 10149 27721 10183
rect 27721 10149 27755 10183
rect 27755 10149 27764 10183
rect 27712 10140 27764 10149
rect 28172 10140 28224 10192
rect 31576 10140 31628 10192
rect 32312 10183 32364 10192
rect 32312 10149 32321 10183
rect 32321 10149 32355 10183
rect 32355 10149 32364 10183
rect 33876 10183 33928 10192
rect 32312 10140 32364 10149
rect 33876 10149 33885 10183
rect 33885 10149 33919 10183
rect 33919 10149 33928 10183
rect 33876 10140 33928 10149
rect 2872 10072 2924 10124
rect 5540 10072 5592 10124
rect 3608 10004 3660 10056
rect 4160 10047 4212 10056
rect 4160 10013 4169 10047
rect 4169 10013 4203 10047
rect 4203 10013 4212 10047
rect 4160 10004 4212 10013
rect 4712 9979 4764 9988
rect 4712 9945 4721 9979
rect 4721 9945 4755 9979
rect 4755 9945 4764 9979
rect 4712 9936 4764 9945
rect 6276 10072 6328 10124
rect 12348 10115 12400 10124
rect 12348 10081 12357 10115
rect 12357 10081 12391 10115
rect 12391 10081 12400 10115
rect 12348 10072 12400 10081
rect 12532 10115 12584 10124
rect 12532 10081 12541 10115
rect 12541 10081 12575 10115
rect 12575 10081 12584 10115
rect 12532 10072 12584 10081
rect 6828 10004 6880 10056
rect 7932 10004 7984 10056
rect 10048 10047 10100 10056
rect 10048 10013 10057 10047
rect 10057 10013 10091 10047
rect 10091 10013 10100 10047
rect 10048 10004 10100 10013
rect 13360 10004 13412 10056
rect 13452 10004 13504 10056
rect 13820 10072 13872 10124
rect 14096 10072 14148 10124
rect 14648 10072 14700 10124
rect 17224 10072 17276 10124
rect 19524 10072 19576 10124
rect 22468 10115 22520 10124
rect 22468 10081 22477 10115
rect 22477 10081 22511 10115
rect 22511 10081 22520 10115
rect 22468 10072 22520 10081
rect 22836 10072 22888 10124
rect 24216 10115 24268 10124
rect 24216 10081 24225 10115
rect 24225 10081 24259 10115
rect 24259 10081 24268 10115
rect 24216 10072 24268 10081
rect 26240 10072 26292 10124
rect 28632 10072 28684 10124
rect 29644 10115 29696 10124
rect 29644 10081 29653 10115
rect 29653 10081 29687 10115
rect 29687 10081 29696 10115
rect 29644 10072 29696 10081
rect 12256 9936 12308 9988
rect 4988 9868 5040 9920
rect 5632 9868 5684 9920
rect 13084 9868 13136 9920
rect 14740 10004 14792 10056
rect 14832 10004 14884 10056
rect 16028 10047 16080 10056
rect 16028 10013 16037 10047
rect 16037 10013 16071 10047
rect 16071 10013 16080 10047
rect 16028 10004 16080 10013
rect 18144 10047 18196 10056
rect 18144 10013 18153 10047
rect 18153 10013 18187 10047
rect 18187 10013 18196 10047
rect 18144 10004 18196 10013
rect 20812 10004 20864 10056
rect 23204 10004 23256 10056
rect 24400 10047 24452 10056
rect 24400 10013 24409 10047
rect 24409 10013 24443 10047
rect 24443 10013 24452 10047
rect 24400 10004 24452 10013
rect 24492 10004 24544 10056
rect 29000 10004 29052 10056
rect 17776 9936 17828 9988
rect 21548 9979 21600 9988
rect 21548 9945 21557 9979
rect 21557 9945 21591 9979
rect 21591 9945 21600 9979
rect 21548 9936 21600 9945
rect 23480 9936 23532 9988
rect 31760 10072 31812 10124
rect 35256 10115 35308 10124
rect 35256 10081 35265 10115
rect 35265 10081 35299 10115
rect 35299 10081 35308 10115
rect 35256 10072 35308 10081
rect 32036 10004 32088 10056
rect 32496 10047 32548 10056
rect 32496 10013 32505 10047
rect 32505 10013 32539 10047
rect 32539 10013 32548 10047
rect 32496 10004 32548 10013
rect 14004 9868 14056 9920
rect 19892 9911 19944 9920
rect 19892 9877 19901 9911
rect 19901 9877 19935 9911
rect 19935 9877 19944 9911
rect 19892 9868 19944 9877
rect 20168 9911 20220 9920
rect 20168 9877 20177 9911
rect 20177 9877 20211 9911
rect 20211 9877 20220 9911
rect 20168 9868 20220 9877
rect 23388 9868 23440 9920
rect 23940 9868 23992 9920
rect 30564 9936 30616 9988
rect 33508 10004 33560 10056
rect 26056 9868 26108 9920
rect 26608 9868 26660 9920
rect 26792 9911 26844 9920
rect 26792 9877 26801 9911
rect 26801 9877 26835 9911
rect 26835 9877 26844 9911
rect 26792 9868 26844 9877
rect 28540 9868 28592 9920
rect 30656 9911 30708 9920
rect 30656 9877 30665 9911
rect 30665 9877 30699 9911
rect 30699 9877 30708 9911
rect 30656 9868 30708 9877
rect 34980 9868 35032 9920
rect 7648 9766 7700 9818
rect 7712 9766 7764 9818
rect 7776 9766 7828 9818
rect 7840 9766 7892 9818
rect 20982 9766 21034 9818
rect 21046 9766 21098 9818
rect 21110 9766 21162 9818
rect 21174 9766 21226 9818
rect 34315 9766 34367 9818
rect 34379 9766 34431 9818
rect 34443 9766 34495 9818
rect 34507 9766 34559 9818
rect 112 9664 164 9716
rect 6000 9664 6052 9716
rect 6276 9664 6328 9716
rect 8208 9707 8260 9716
rect 8208 9673 8217 9707
rect 8217 9673 8251 9707
rect 8251 9673 8260 9707
rect 8208 9664 8260 9673
rect 9772 9664 9824 9716
rect 10232 9664 10284 9716
rect 12348 9664 12400 9716
rect 15384 9707 15436 9716
rect 15384 9673 15393 9707
rect 15393 9673 15427 9707
rect 15427 9673 15436 9707
rect 15384 9664 15436 9673
rect 17224 9707 17276 9716
rect 17224 9673 17233 9707
rect 17233 9673 17267 9707
rect 17267 9673 17276 9707
rect 17224 9664 17276 9673
rect 21272 9664 21324 9716
rect 27712 9664 27764 9716
rect 30748 9664 30800 9716
rect 32312 9664 32364 9716
rect 8392 9596 8444 9648
rect 9864 9639 9916 9648
rect 9864 9605 9873 9639
rect 9873 9605 9907 9639
rect 9907 9605 9916 9639
rect 9864 9596 9916 9605
rect 12440 9596 12492 9648
rect 2780 9528 2832 9580
rect 4712 9571 4764 9580
rect 4712 9537 4721 9571
rect 4721 9537 4755 9571
rect 4755 9537 4764 9571
rect 4712 9528 4764 9537
rect 7104 9528 7156 9580
rect 8852 9571 8904 9580
rect 8852 9537 8861 9571
rect 8861 9537 8895 9571
rect 8895 9537 8904 9571
rect 12716 9596 12768 9648
rect 14096 9596 14148 9648
rect 14740 9596 14792 9648
rect 15016 9596 15068 9648
rect 17868 9596 17920 9648
rect 20168 9596 20220 9648
rect 21732 9596 21784 9648
rect 23388 9596 23440 9648
rect 27160 9596 27212 9648
rect 33876 9664 33928 9716
rect 35256 9707 35308 9716
rect 35256 9673 35265 9707
rect 35265 9673 35299 9707
rect 35299 9673 35308 9707
rect 35256 9664 35308 9673
rect 33508 9596 33560 9648
rect 35624 9639 35676 9648
rect 35624 9605 35633 9639
rect 35633 9605 35667 9639
rect 35667 9605 35676 9639
rect 35624 9596 35676 9605
rect 8852 9528 8904 9537
rect 12808 9571 12860 9580
rect 12808 9537 12817 9571
rect 12817 9537 12851 9571
rect 12851 9537 12860 9571
rect 12808 9528 12860 9537
rect 15384 9528 15436 9580
rect 17960 9528 18012 9580
rect 19248 9528 19300 9580
rect 20260 9528 20312 9580
rect 21640 9571 21692 9580
rect 21640 9537 21649 9571
rect 21649 9537 21683 9571
rect 21683 9537 21692 9571
rect 21640 9528 21692 9537
rect 21916 9571 21968 9580
rect 21916 9537 21925 9571
rect 21925 9537 21959 9571
rect 21959 9537 21968 9571
rect 21916 9528 21968 9537
rect 24216 9528 24268 9580
rect 24492 9528 24544 9580
rect 24584 9528 24636 9580
rect 27068 9528 27120 9580
rect 30656 9571 30708 9580
rect 30656 9537 30665 9571
rect 30665 9537 30699 9571
rect 30699 9537 30708 9571
rect 30656 9528 30708 9537
rect 30932 9571 30984 9580
rect 30932 9537 30941 9571
rect 30941 9537 30975 9571
rect 30975 9537 30984 9571
rect 30932 9528 30984 9537
rect 32496 9528 32548 9580
rect 32680 9571 32732 9580
rect 32680 9537 32689 9571
rect 32689 9537 32723 9571
rect 32723 9537 32732 9571
rect 32680 9528 32732 9537
rect 1400 9503 1452 9512
rect 1400 9469 1409 9503
rect 1409 9469 1443 9503
rect 1443 9469 1452 9503
rect 1952 9503 2004 9512
rect 1400 9460 1452 9469
rect 1952 9469 1961 9503
rect 1961 9469 1995 9503
rect 1995 9469 2004 9503
rect 1952 9460 2004 9469
rect 3976 9460 4028 9512
rect 3240 9392 3292 9444
rect 4436 9435 4488 9444
rect 112 9324 164 9376
rect 2504 9367 2556 9376
rect 2504 9333 2513 9367
rect 2513 9333 2547 9367
rect 2547 9333 2556 9367
rect 2504 9324 2556 9333
rect 3608 9324 3660 9376
rect 4436 9401 4445 9435
rect 4445 9401 4479 9435
rect 4479 9401 4488 9435
rect 4436 9392 4488 9401
rect 5540 9324 5592 9376
rect 5816 9324 5868 9376
rect 7288 9392 7340 9444
rect 8208 9392 8260 9444
rect 7104 9324 7156 9376
rect 8484 9324 8536 9376
rect 10048 9392 10100 9444
rect 11796 9503 11848 9512
rect 11796 9469 11805 9503
rect 11805 9469 11839 9503
rect 11839 9469 11848 9503
rect 11796 9460 11848 9469
rect 14648 9460 14700 9512
rect 16488 9503 16540 9512
rect 16488 9469 16497 9503
rect 16497 9469 16531 9503
rect 16531 9469 16540 9503
rect 16488 9460 16540 9469
rect 12992 9392 13044 9444
rect 10876 9367 10928 9376
rect 10876 9333 10885 9367
rect 10885 9333 10919 9367
rect 10919 9333 10928 9367
rect 10876 9324 10928 9333
rect 11704 9324 11756 9376
rect 12532 9324 12584 9376
rect 15016 9392 15068 9444
rect 18236 9460 18288 9512
rect 28632 9503 28684 9512
rect 28632 9469 28641 9503
rect 28641 9469 28675 9503
rect 28675 9469 28684 9503
rect 28632 9460 28684 9469
rect 28724 9460 28776 9512
rect 16948 9435 17000 9444
rect 16948 9401 16957 9435
rect 16957 9401 16991 9435
rect 16991 9401 17000 9435
rect 16948 9392 17000 9401
rect 17868 9435 17920 9444
rect 17868 9401 17877 9435
rect 17877 9401 17911 9435
rect 17911 9401 17920 9435
rect 17868 9392 17920 9401
rect 20076 9392 20128 9444
rect 21732 9435 21784 9444
rect 21732 9401 21741 9435
rect 21741 9401 21775 9435
rect 21775 9401 21784 9435
rect 21732 9392 21784 9401
rect 15568 9324 15620 9376
rect 18788 9324 18840 9376
rect 19524 9324 19576 9376
rect 19984 9324 20036 9376
rect 22468 9324 22520 9376
rect 22836 9324 22888 9376
rect 23204 9324 23256 9376
rect 23664 9324 23716 9376
rect 24124 9392 24176 9444
rect 25320 9435 25372 9444
rect 25320 9401 25329 9435
rect 25329 9401 25363 9435
rect 25363 9401 25372 9435
rect 25320 9392 25372 9401
rect 25688 9392 25740 9444
rect 27160 9392 27212 9444
rect 28356 9392 28408 9444
rect 35256 9460 35308 9512
rect 30748 9435 30800 9444
rect 30748 9401 30757 9435
rect 30757 9401 30791 9435
rect 30791 9401 30800 9435
rect 30748 9392 30800 9401
rect 26240 9324 26292 9376
rect 28264 9367 28316 9376
rect 28264 9333 28273 9367
rect 28273 9333 28307 9367
rect 28307 9333 28316 9367
rect 28264 9324 28316 9333
rect 28724 9324 28776 9376
rect 29644 9324 29696 9376
rect 30104 9367 30156 9376
rect 30104 9333 30113 9367
rect 30113 9333 30147 9367
rect 30147 9333 30156 9367
rect 30104 9324 30156 9333
rect 31760 9324 31812 9376
rect 33140 9324 33192 9376
rect 14315 9222 14367 9274
rect 14379 9222 14431 9274
rect 14443 9222 14495 9274
rect 14507 9222 14559 9274
rect 27648 9222 27700 9274
rect 27712 9222 27764 9274
rect 27776 9222 27828 9274
rect 27840 9222 27892 9274
rect 2044 9163 2096 9172
rect 2044 9129 2053 9163
rect 2053 9129 2087 9163
rect 2087 9129 2096 9163
rect 2044 9120 2096 9129
rect 2504 9120 2556 9172
rect 3240 9120 3292 9172
rect 4160 9120 4212 9172
rect 4436 9120 4488 9172
rect 6092 9163 6144 9172
rect 2780 9052 2832 9104
rect 3976 9052 4028 9104
rect 5816 9052 5868 9104
rect 6092 9129 6101 9163
rect 6101 9129 6135 9163
rect 6135 9129 6144 9163
rect 6092 9120 6144 9129
rect 6828 9163 6880 9172
rect 6828 9129 6837 9163
rect 6837 9129 6871 9163
rect 6871 9129 6880 9163
rect 6828 9120 6880 9129
rect 7288 9163 7340 9172
rect 7288 9129 7297 9163
rect 7297 9129 7331 9163
rect 7331 9129 7340 9163
rect 7288 9120 7340 9129
rect 8208 9120 8260 9172
rect 8852 9163 8904 9172
rect 8852 9129 8861 9163
rect 8861 9129 8895 9163
rect 8895 9129 8904 9163
rect 8852 9120 8904 9129
rect 13820 9163 13872 9172
rect 13820 9129 13829 9163
rect 13829 9129 13863 9163
rect 13863 9129 13872 9163
rect 13820 9120 13872 9129
rect 14832 9120 14884 9172
rect 7104 9052 7156 9104
rect 9864 9095 9916 9104
rect 9864 9061 9873 9095
rect 9873 9061 9907 9095
rect 9907 9061 9916 9095
rect 9864 9052 9916 9061
rect 11704 9052 11756 9104
rect 12992 9052 13044 9104
rect 14648 9052 14700 9104
rect 18144 9163 18196 9172
rect 18144 9129 18153 9163
rect 18153 9129 18187 9163
rect 18187 9129 18196 9163
rect 18144 9120 18196 9129
rect 18236 9120 18288 9172
rect 15476 9095 15528 9104
rect 15476 9061 15485 9095
rect 15485 9061 15519 9095
rect 15519 9061 15528 9095
rect 15476 9052 15528 9061
rect 16396 9095 16448 9104
rect 16396 9061 16405 9095
rect 16405 9061 16439 9095
rect 16439 9061 16448 9095
rect 16396 9052 16448 9061
rect 20076 9120 20128 9172
rect 20260 9163 20312 9172
rect 20260 9129 20269 9163
rect 20269 9129 20303 9163
rect 20303 9129 20312 9163
rect 20260 9120 20312 9129
rect 20812 9120 20864 9172
rect 21640 9120 21692 9172
rect 23480 9163 23532 9172
rect 23480 9129 23489 9163
rect 23489 9129 23523 9163
rect 23523 9129 23532 9163
rect 23480 9120 23532 9129
rect 24400 9163 24452 9172
rect 24400 9129 24409 9163
rect 24409 9129 24443 9163
rect 24443 9129 24452 9163
rect 24400 9120 24452 9129
rect 2228 9027 2280 9036
rect 2228 8993 2237 9027
rect 2237 8993 2271 9027
rect 2271 8993 2280 9027
rect 2228 8984 2280 8993
rect 4068 9027 4120 9036
rect 4068 8993 4077 9027
rect 4077 8993 4111 9027
rect 4111 8993 4120 9027
rect 5172 9027 5224 9036
rect 4068 8984 4120 8993
rect 5172 8993 5181 9027
rect 5181 8993 5215 9027
rect 5215 8993 5224 9027
rect 5172 8984 5224 8993
rect 5724 8984 5776 9036
rect 8116 8984 8168 9036
rect 13728 8984 13780 9036
rect 16856 9027 16908 9036
rect 16856 8993 16865 9027
rect 16865 8993 16899 9027
rect 16899 8993 16908 9027
rect 16856 8984 16908 8993
rect 17500 8984 17552 9036
rect 19064 9027 19116 9036
rect 19064 8993 19073 9027
rect 19073 8993 19107 9027
rect 19107 8993 19116 9027
rect 19064 8984 19116 8993
rect 22100 9052 22152 9104
rect 25320 9120 25372 9172
rect 28264 9120 28316 9172
rect 28908 9120 28960 9172
rect 29552 9163 29604 9172
rect 29552 9129 29561 9163
rect 29561 9129 29595 9163
rect 29595 9129 29604 9163
rect 29552 9120 29604 9129
rect 31576 9120 31628 9172
rect 32496 9163 32548 9172
rect 32496 9129 32505 9163
rect 32505 9129 32539 9163
rect 32539 9129 32548 9163
rect 32496 9120 32548 9129
rect 33140 9120 33192 9172
rect 25504 9052 25556 9104
rect 26976 9052 27028 9104
rect 28448 9095 28500 9104
rect 28448 9061 28457 9095
rect 28457 9061 28491 9095
rect 28491 9061 28500 9095
rect 28448 9052 28500 9061
rect 29000 9095 29052 9104
rect 29000 9061 29009 9095
rect 29009 9061 29043 9095
rect 29043 9061 29052 9095
rect 29000 9052 29052 9061
rect 30564 9095 30616 9104
rect 30564 9061 30573 9095
rect 30573 9061 30607 9095
rect 30607 9061 30616 9095
rect 30564 9052 30616 9061
rect 30840 9052 30892 9104
rect 31484 9052 31536 9104
rect 34612 9052 34664 9104
rect 6920 8959 6972 8968
rect 6920 8925 6929 8959
rect 6929 8925 6963 8959
rect 6963 8925 6972 8959
rect 6920 8916 6972 8925
rect 11060 8916 11112 8968
rect 11152 8916 11204 8968
rect 15108 8916 15160 8968
rect 16028 8959 16080 8968
rect 16028 8925 16037 8959
rect 16037 8925 16071 8959
rect 16071 8925 16080 8959
rect 16028 8916 16080 8925
rect 20720 8916 20772 8968
rect 21916 8916 21968 8968
rect 23112 8959 23164 8968
rect 23112 8925 23121 8959
rect 23121 8925 23155 8959
rect 23155 8925 23164 8959
rect 23112 8916 23164 8925
rect 23204 8916 23256 8968
rect 32036 8984 32088 9036
rect 33232 8984 33284 9036
rect 35900 9027 35952 9036
rect 35900 8993 35909 9027
rect 35909 8993 35943 9027
rect 35943 8993 35952 9027
rect 35900 8984 35952 8993
rect 26516 8959 26568 8968
rect 26516 8925 26525 8959
rect 26525 8925 26559 8959
rect 26559 8925 26568 8959
rect 26516 8916 26568 8925
rect 28356 8959 28408 8968
rect 28356 8925 28365 8959
rect 28365 8925 28399 8959
rect 28399 8925 28408 8959
rect 28356 8916 28408 8925
rect 30932 8916 30984 8968
rect 34704 8916 34756 8968
rect 36268 8916 36320 8968
rect 20 8848 72 8900
rect 8760 8848 8812 8900
rect 12808 8848 12860 8900
rect 15016 8848 15068 8900
rect 21548 8891 21600 8900
rect 21548 8857 21557 8891
rect 21557 8857 21591 8891
rect 21591 8857 21600 8891
rect 21548 8848 21600 8857
rect 23388 8848 23440 8900
rect 30104 8848 30156 8900
rect 36636 8848 36688 8900
rect 8300 8823 8352 8832
rect 8300 8789 8309 8823
rect 8309 8789 8343 8823
rect 8343 8789 8352 8823
rect 8300 8780 8352 8789
rect 12992 8823 13044 8832
rect 12992 8789 13001 8823
rect 13001 8789 13035 8823
rect 13035 8789 13044 8823
rect 12992 8780 13044 8789
rect 18972 8823 19024 8832
rect 18972 8789 18981 8823
rect 18981 8789 19015 8823
rect 19015 8789 19024 8823
rect 18972 8780 19024 8789
rect 21272 8780 21324 8832
rect 24676 8780 24728 8832
rect 39580 8780 39632 8832
rect 7648 8678 7700 8730
rect 7712 8678 7764 8730
rect 7776 8678 7828 8730
rect 7840 8678 7892 8730
rect 20982 8678 21034 8730
rect 21046 8678 21098 8730
rect 21110 8678 21162 8730
rect 21174 8678 21226 8730
rect 34315 8678 34367 8730
rect 34379 8678 34431 8730
rect 34443 8678 34495 8730
rect 34507 8678 34559 8730
rect 2228 8576 2280 8628
rect 3148 8619 3200 8628
rect 1860 8508 1912 8560
rect 3148 8585 3157 8619
rect 3157 8585 3191 8619
rect 3191 8585 3200 8619
rect 3148 8576 3200 8585
rect 4068 8576 4120 8628
rect 6828 8576 6880 8628
rect 2136 8440 2188 8492
rect 7196 8508 7248 8560
rect 3792 8440 3844 8492
rect 6000 8415 6052 8424
rect 6000 8381 6009 8415
rect 6009 8381 6043 8415
rect 6043 8381 6052 8415
rect 6000 8372 6052 8381
rect 6368 8372 6420 8424
rect 8208 8576 8260 8628
rect 9864 8619 9916 8628
rect 9864 8585 9873 8619
rect 9873 8585 9907 8619
rect 9907 8585 9916 8619
rect 9864 8576 9916 8585
rect 11060 8619 11112 8628
rect 11060 8585 11069 8619
rect 11069 8585 11103 8619
rect 11103 8585 11112 8619
rect 11060 8576 11112 8585
rect 11704 8576 11756 8628
rect 12992 8576 13044 8628
rect 15476 8576 15528 8628
rect 17500 8619 17552 8628
rect 17500 8585 17509 8619
rect 17509 8585 17543 8619
rect 17543 8585 17552 8619
rect 17500 8576 17552 8585
rect 19156 8576 19208 8628
rect 20168 8576 20220 8628
rect 22100 8619 22152 8628
rect 22100 8585 22109 8619
rect 22109 8585 22143 8619
rect 22143 8585 22152 8619
rect 22100 8576 22152 8585
rect 23112 8576 23164 8628
rect 25688 8619 25740 8628
rect 25688 8585 25697 8619
rect 25697 8585 25731 8619
rect 25731 8585 25740 8619
rect 25688 8576 25740 8585
rect 28448 8576 28500 8628
rect 30564 8576 30616 8628
rect 33232 8619 33284 8628
rect 33232 8585 33241 8619
rect 33241 8585 33275 8619
rect 33275 8585 33284 8619
rect 33232 8576 33284 8585
rect 34704 8576 34756 8628
rect 10416 8508 10468 8560
rect 11152 8508 11204 8560
rect 16396 8508 16448 8560
rect 8300 8440 8352 8492
rect 10692 8440 10744 8492
rect 13636 8440 13688 8492
rect 14648 8440 14700 8492
rect 19892 8508 19944 8560
rect 30840 8551 30892 8560
rect 17132 8483 17184 8492
rect 17132 8449 17141 8483
rect 17141 8449 17175 8483
rect 17175 8449 17184 8483
rect 17132 8440 17184 8449
rect 18880 8440 18932 8492
rect 18972 8440 19024 8492
rect 30840 8517 30849 8551
rect 30849 8517 30883 8551
rect 30883 8517 30892 8551
rect 30840 8508 30892 8517
rect 35900 8551 35952 8560
rect 35900 8517 35909 8551
rect 35909 8517 35943 8551
rect 35943 8517 35952 8551
rect 35900 8508 35952 8517
rect 21364 8440 21416 8492
rect 12624 8372 12676 8424
rect 18696 8372 18748 8424
rect 21272 8372 21324 8424
rect 26332 8440 26384 8492
rect 28356 8440 28408 8492
rect 29552 8483 29604 8492
rect 29552 8449 29561 8483
rect 29561 8449 29595 8483
rect 29595 8449 29604 8483
rect 29552 8440 29604 8449
rect 30012 8440 30064 8492
rect 31668 8483 31720 8492
rect 31668 8449 31677 8483
rect 31677 8449 31711 8483
rect 31711 8449 31720 8483
rect 31668 8440 31720 8449
rect 34612 8483 34664 8492
rect 23756 8372 23808 8424
rect 24584 8372 24636 8424
rect 24860 8372 24912 8424
rect 30748 8372 30800 8424
rect 34612 8449 34621 8483
rect 34621 8449 34655 8483
rect 34655 8449 34664 8483
rect 34612 8440 34664 8449
rect 34980 8483 35032 8492
rect 34980 8449 34989 8483
rect 34989 8449 35023 8483
rect 35023 8449 35032 8483
rect 34980 8440 35032 8449
rect 35256 8483 35308 8492
rect 35256 8449 35265 8483
rect 35265 8449 35299 8483
rect 35299 8449 35308 8483
rect 35256 8440 35308 8449
rect 35440 8440 35492 8492
rect 34152 8372 34204 8424
rect 3884 8304 3936 8356
rect 4528 8304 4580 8356
rect 5816 8304 5868 8356
rect 8668 8304 8720 8356
rect 10048 8347 10100 8356
rect 10048 8313 10057 8347
rect 10057 8313 10091 8347
rect 10091 8313 10100 8347
rect 10048 8304 10100 8313
rect 2504 8236 2556 8288
rect 3332 8236 3384 8288
rect 5264 8236 5316 8288
rect 6920 8236 6972 8288
rect 9864 8236 9916 8288
rect 16580 8347 16632 8356
rect 16580 8313 16589 8347
rect 16589 8313 16623 8347
rect 16623 8313 16632 8347
rect 16580 8304 16632 8313
rect 19524 8304 19576 8356
rect 13912 8236 13964 8288
rect 14740 8279 14792 8288
rect 14740 8245 14749 8279
rect 14749 8245 14783 8279
rect 14783 8245 14792 8279
rect 14740 8236 14792 8245
rect 15936 8236 15988 8288
rect 16856 8236 16908 8288
rect 20076 8304 20128 8356
rect 21824 8347 21876 8356
rect 21824 8313 21833 8347
rect 21833 8313 21867 8347
rect 21867 8313 21876 8347
rect 21824 8304 21876 8313
rect 24952 8304 25004 8356
rect 23480 8236 23532 8288
rect 26976 8304 27028 8356
rect 36636 8372 36688 8424
rect 29920 8279 29972 8288
rect 29920 8245 29929 8279
rect 29929 8245 29963 8279
rect 29963 8245 29972 8279
rect 29920 8236 29972 8245
rect 32496 8236 32548 8288
rect 34152 8236 34204 8288
rect 35992 8236 36044 8288
rect 38108 8236 38160 8288
rect 14315 8134 14367 8186
rect 14379 8134 14431 8186
rect 14443 8134 14495 8186
rect 14507 8134 14559 8186
rect 27648 8134 27700 8186
rect 27712 8134 27764 8186
rect 27776 8134 27828 8186
rect 27840 8134 27892 8186
rect 2136 8075 2188 8084
rect 2136 8041 2145 8075
rect 2145 8041 2179 8075
rect 2179 8041 2188 8075
rect 2136 8032 2188 8041
rect 3884 8075 3936 8084
rect 3884 8041 3893 8075
rect 3893 8041 3927 8075
rect 3927 8041 3936 8075
rect 3884 8032 3936 8041
rect 3976 8032 4028 8084
rect 4528 8032 4580 8084
rect 5172 8075 5224 8084
rect 5172 8041 5181 8075
rect 5181 8041 5215 8075
rect 5215 8041 5224 8075
rect 5172 8032 5224 8041
rect 5816 8075 5868 8084
rect 5816 8041 5825 8075
rect 5825 8041 5859 8075
rect 5859 8041 5868 8075
rect 5816 8032 5868 8041
rect 9680 8032 9732 8084
rect 11336 8075 11388 8084
rect 2412 8007 2464 8016
rect 2412 7973 2421 8007
rect 2421 7973 2455 8007
rect 2455 7973 2464 8007
rect 2412 7964 2464 7973
rect 3700 7896 3752 7948
rect 5448 7939 5500 7948
rect 5448 7905 5457 7939
rect 5457 7905 5491 7939
rect 5491 7905 5500 7939
rect 5448 7896 5500 7905
rect 8116 7964 8168 8016
rect 11336 8041 11345 8075
rect 11345 8041 11379 8075
rect 11379 8041 11388 8075
rect 11336 8032 11388 8041
rect 13728 8032 13780 8084
rect 14648 8075 14700 8084
rect 14648 8041 14657 8075
rect 14657 8041 14691 8075
rect 14691 8041 14700 8075
rect 14648 8032 14700 8041
rect 15108 8075 15160 8084
rect 15108 8041 15117 8075
rect 15117 8041 15151 8075
rect 15151 8041 15160 8075
rect 15108 8032 15160 8041
rect 16580 8032 16632 8084
rect 17776 8075 17828 8084
rect 17776 8041 17785 8075
rect 17785 8041 17819 8075
rect 17819 8041 17828 8075
rect 17776 8032 17828 8041
rect 18420 8032 18472 8084
rect 18972 8032 19024 8084
rect 19524 8032 19576 8084
rect 22652 8032 22704 8084
rect 23296 8032 23348 8084
rect 5908 7896 5960 7948
rect 8760 7939 8812 7948
rect 8760 7905 8769 7939
rect 8769 7905 8803 7939
rect 8803 7905 8812 7939
rect 8760 7896 8812 7905
rect 1952 7760 2004 7812
rect 3424 7828 3476 7880
rect 8208 7828 8260 7880
rect 8944 7828 8996 7880
rect 9864 8007 9916 8016
rect 9864 7973 9873 8007
rect 9873 7973 9907 8007
rect 9907 7973 9916 8007
rect 10416 8007 10468 8016
rect 9864 7964 9916 7973
rect 10416 7973 10425 8007
rect 10425 7973 10459 8007
rect 10459 7973 10468 8007
rect 10416 7964 10468 7973
rect 13820 8007 13872 8016
rect 13820 7973 13829 8007
rect 13829 7973 13863 8007
rect 13863 7973 13872 8007
rect 13820 7964 13872 7973
rect 15016 7964 15068 8016
rect 16028 8007 16080 8016
rect 16028 7973 16037 8007
rect 16037 7973 16071 8007
rect 16071 7973 16080 8007
rect 16028 7964 16080 7973
rect 17040 7964 17092 8016
rect 17868 7964 17920 8016
rect 20720 8007 20772 8016
rect 20720 7973 20729 8007
rect 20729 7973 20763 8007
rect 20763 7973 20772 8007
rect 20720 7964 20772 7973
rect 22836 7964 22888 8016
rect 23480 7964 23532 8016
rect 26516 8032 26568 8084
rect 26976 8032 27028 8084
rect 29920 8032 29972 8084
rect 24768 7964 24820 8016
rect 9864 7828 9916 7880
rect 11704 7896 11756 7948
rect 12716 7896 12768 7948
rect 16948 7896 17000 7948
rect 18696 7896 18748 7948
rect 18972 7939 19024 7948
rect 18972 7905 18981 7939
rect 18981 7905 19015 7939
rect 19015 7905 19024 7939
rect 18972 7896 19024 7905
rect 19432 7939 19484 7948
rect 19432 7905 19441 7939
rect 19441 7905 19475 7939
rect 19475 7905 19484 7939
rect 19432 7896 19484 7905
rect 21364 7939 21416 7948
rect 12072 7828 12124 7880
rect 13544 7828 13596 7880
rect 14648 7828 14700 7880
rect 15384 7871 15436 7880
rect 15384 7837 15393 7871
rect 15393 7837 15427 7871
rect 15427 7837 15436 7871
rect 15384 7828 15436 7837
rect 19064 7828 19116 7880
rect 21364 7905 21373 7939
rect 21373 7905 21407 7939
rect 21407 7905 21416 7939
rect 21364 7896 21416 7905
rect 22744 7939 22796 7948
rect 22744 7905 22753 7939
rect 22753 7905 22787 7939
rect 22787 7905 22796 7939
rect 22744 7896 22796 7905
rect 23664 7939 23716 7948
rect 23664 7905 23673 7939
rect 23673 7905 23707 7939
rect 23707 7905 23716 7939
rect 23664 7896 23716 7905
rect 26424 7896 26476 7948
rect 26608 7896 26660 7948
rect 28724 7964 28776 8016
rect 30656 8032 30708 8084
rect 30840 8075 30892 8084
rect 30840 8041 30849 8075
rect 30849 8041 30883 8075
rect 30883 8041 30892 8075
rect 30840 8032 30892 8041
rect 31668 8075 31720 8084
rect 31668 8041 31677 8075
rect 31677 8041 31711 8075
rect 31711 8041 31720 8075
rect 31668 8032 31720 8041
rect 32496 8075 32548 8084
rect 32496 8041 32505 8075
rect 32505 8041 32539 8075
rect 32539 8041 32548 8075
rect 32496 8032 32548 8041
rect 34704 8032 34756 8084
rect 34980 8032 35032 8084
rect 34152 7964 34204 8016
rect 34520 8007 34572 8016
rect 34520 7973 34529 8007
rect 34529 7973 34563 8007
rect 34563 7973 34572 8007
rect 34520 7964 34572 7973
rect 35256 7964 35308 8016
rect 35992 8007 36044 8016
rect 35992 7973 36001 8007
rect 36001 7973 36035 8007
rect 36035 7973 36044 8007
rect 35992 7964 36044 7973
rect 36084 8007 36136 8016
rect 36084 7973 36093 8007
rect 36093 7973 36127 8007
rect 36127 7973 36136 8007
rect 36084 7964 36136 7973
rect 5264 7760 5316 7812
rect 16488 7760 16540 7812
rect 21272 7828 21324 7880
rect 21640 7871 21692 7880
rect 21640 7837 21649 7871
rect 21649 7837 21683 7871
rect 21683 7837 21692 7871
rect 21640 7828 21692 7837
rect 24676 7828 24728 7880
rect 24308 7760 24360 7812
rect 28816 7939 28868 7948
rect 28816 7905 28825 7939
rect 28825 7905 28859 7939
rect 28859 7905 28868 7939
rect 28816 7896 28868 7905
rect 31852 7896 31904 7948
rect 29920 7871 29972 7880
rect 29920 7837 29929 7871
rect 29929 7837 29963 7871
rect 29963 7837 29972 7871
rect 29920 7828 29972 7837
rect 32128 7871 32180 7880
rect 32128 7837 32137 7871
rect 32137 7837 32171 7871
rect 32171 7837 32180 7871
rect 32128 7828 32180 7837
rect 33692 7828 33744 7880
rect 34520 7828 34572 7880
rect 36084 7828 36136 7880
rect 36268 7871 36320 7880
rect 36268 7837 36277 7871
rect 36277 7837 36311 7871
rect 36311 7837 36320 7871
rect 36268 7828 36320 7837
rect 30380 7760 30432 7812
rect 31760 7760 31812 7812
rect 36452 7760 36504 7812
rect 2688 7692 2740 7744
rect 10048 7692 10100 7744
rect 12624 7692 12676 7744
rect 20076 7735 20128 7744
rect 20076 7701 20085 7735
rect 20085 7701 20119 7735
rect 20119 7701 20128 7735
rect 20076 7692 20128 7701
rect 21548 7692 21600 7744
rect 24860 7692 24912 7744
rect 25504 7735 25556 7744
rect 25504 7701 25513 7735
rect 25513 7701 25547 7735
rect 25547 7701 25556 7735
rect 25504 7692 25556 7701
rect 27528 7692 27580 7744
rect 27712 7735 27764 7744
rect 27712 7701 27721 7735
rect 27721 7701 27755 7735
rect 27755 7701 27764 7735
rect 27712 7692 27764 7701
rect 33692 7692 33744 7744
rect 7648 7590 7700 7642
rect 7712 7590 7764 7642
rect 7776 7590 7828 7642
rect 7840 7590 7892 7642
rect 20982 7590 21034 7642
rect 21046 7590 21098 7642
rect 21110 7590 21162 7642
rect 21174 7590 21226 7642
rect 34315 7590 34367 7642
rect 34379 7590 34431 7642
rect 34443 7590 34495 7642
rect 34507 7590 34559 7642
rect 2412 7488 2464 7540
rect 2596 7488 2648 7540
rect 3700 7531 3752 7540
rect 3700 7497 3709 7531
rect 3709 7497 3743 7531
rect 3743 7497 3752 7531
rect 3700 7488 3752 7497
rect 4528 7488 4580 7540
rect 5448 7488 5500 7540
rect 8116 7531 8168 7540
rect 8116 7497 8125 7531
rect 8125 7497 8159 7531
rect 8159 7497 8168 7531
rect 8116 7488 8168 7497
rect 8668 7531 8720 7540
rect 8668 7497 8677 7531
rect 8677 7497 8711 7531
rect 8711 7497 8720 7531
rect 8668 7488 8720 7497
rect 11704 7531 11756 7540
rect 11704 7497 11713 7531
rect 11713 7497 11747 7531
rect 11747 7497 11756 7531
rect 11704 7488 11756 7497
rect 15016 7488 15068 7540
rect 16948 7488 17000 7540
rect 17776 7531 17828 7540
rect 17776 7497 17785 7531
rect 17785 7497 17819 7531
rect 17819 7497 17828 7531
rect 17776 7488 17828 7497
rect 18972 7488 19024 7540
rect 19432 7531 19484 7540
rect 19432 7497 19441 7531
rect 19441 7497 19475 7531
rect 19475 7497 19484 7531
rect 19432 7488 19484 7497
rect 19892 7531 19944 7540
rect 19892 7497 19901 7531
rect 19901 7497 19935 7531
rect 19935 7497 19944 7531
rect 19892 7488 19944 7497
rect 22744 7488 22796 7540
rect 24768 7531 24820 7540
rect 24768 7497 24777 7531
rect 24777 7497 24811 7531
rect 24811 7497 24820 7531
rect 24768 7488 24820 7497
rect 26792 7488 26844 7540
rect 26884 7488 26936 7540
rect 3884 7420 3936 7472
rect 13912 7420 13964 7472
rect 17040 7463 17092 7472
rect 17040 7429 17049 7463
rect 17049 7429 17083 7463
rect 17083 7429 17092 7463
rect 17040 7420 17092 7429
rect 17960 7420 18012 7472
rect 22836 7463 22888 7472
rect 22836 7429 22845 7463
rect 22845 7429 22879 7463
rect 22879 7429 22888 7463
rect 22836 7420 22888 7429
rect 22928 7420 22980 7472
rect 2688 7352 2740 7404
rect 5080 7352 5132 7404
rect 6276 7352 6328 7404
rect 6736 7352 6788 7404
rect 3424 7284 3476 7336
rect 3884 7327 3936 7336
rect 3884 7293 3893 7327
rect 3893 7293 3927 7327
rect 3927 7293 3936 7327
rect 3884 7284 3936 7293
rect 4528 7284 4580 7336
rect 4620 7284 4672 7336
rect 7104 7327 7156 7336
rect 7104 7293 7113 7327
rect 7113 7293 7147 7327
rect 7147 7293 7156 7327
rect 7104 7284 7156 7293
rect 9128 7352 9180 7404
rect 11336 7352 11388 7404
rect 13820 7352 13872 7404
rect 15384 7352 15436 7404
rect 16028 7395 16080 7404
rect 16028 7361 16037 7395
rect 16037 7361 16071 7395
rect 16071 7361 16080 7395
rect 16028 7352 16080 7361
rect 17132 7352 17184 7404
rect 18420 7352 18472 7404
rect 21180 7395 21232 7404
rect 21180 7361 21189 7395
rect 21189 7361 21223 7395
rect 21223 7361 21232 7395
rect 21180 7352 21232 7361
rect 21640 7395 21692 7404
rect 21640 7361 21649 7395
rect 21649 7361 21683 7395
rect 21683 7361 21692 7395
rect 21640 7352 21692 7361
rect 22652 7352 22704 7404
rect 25596 7352 25648 7404
rect 3332 7191 3384 7200
rect 3332 7157 3341 7191
rect 3341 7157 3375 7191
rect 3375 7157 3384 7191
rect 8668 7216 8720 7268
rect 9312 7216 9364 7268
rect 3332 7148 3384 7157
rect 5816 7148 5868 7200
rect 6920 7191 6972 7200
rect 6920 7157 6929 7191
rect 6929 7157 6963 7191
rect 6963 7157 6972 7191
rect 6920 7148 6972 7157
rect 9864 7148 9916 7200
rect 9956 7148 10008 7200
rect 11704 7284 11756 7336
rect 13360 7327 13412 7336
rect 13360 7293 13369 7327
rect 13369 7293 13403 7327
rect 13403 7293 13412 7327
rect 13360 7284 13412 7293
rect 15660 7284 15712 7336
rect 19892 7284 19944 7336
rect 20168 7284 20220 7336
rect 21364 7284 21416 7336
rect 10692 7191 10744 7200
rect 10692 7157 10701 7191
rect 10701 7157 10735 7191
rect 10735 7157 10744 7191
rect 10692 7148 10744 7157
rect 12072 7191 12124 7200
rect 12072 7157 12081 7191
rect 12081 7157 12115 7191
rect 12115 7157 12124 7191
rect 12072 7148 12124 7157
rect 13774 7216 13826 7268
rect 15752 7191 15804 7200
rect 15752 7157 15761 7191
rect 15761 7157 15795 7191
rect 15795 7157 15804 7191
rect 17316 7216 17368 7268
rect 20812 7259 20864 7268
rect 15752 7148 15804 7157
rect 17776 7148 17828 7200
rect 20812 7225 20821 7259
rect 20821 7225 20855 7259
rect 20855 7225 20864 7259
rect 20812 7216 20864 7225
rect 21548 7259 21600 7268
rect 21548 7225 21557 7259
rect 21557 7225 21591 7259
rect 21591 7225 21600 7259
rect 21548 7216 21600 7225
rect 22836 7216 22888 7268
rect 24676 7284 24728 7336
rect 26424 7284 26476 7336
rect 27528 7488 27580 7540
rect 33692 7531 33744 7540
rect 23756 7148 23808 7200
rect 26700 7216 26752 7268
rect 27712 7284 27764 7336
rect 33692 7497 33701 7531
rect 33701 7497 33735 7531
rect 33735 7497 33744 7531
rect 33692 7488 33744 7497
rect 32128 7352 32180 7404
rect 25504 7148 25556 7200
rect 26240 7148 26292 7200
rect 26516 7191 26568 7200
rect 26516 7157 26525 7191
rect 26525 7157 26559 7191
rect 26559 7157 26568 7191
rect 26516 7148 26568 7157
rect 26884 7191 26936 7200
rect 26884 7157 26893 7191
rect 26893 7157 26927 7191
rect 26927 7157 26936 7191
rect 26884 7148 26936 7157
rect 29460 7284 29512 7336
rect 29736 7327 29788 7336
rect 29736 7293 29745 7327
rect 29745 7293 29779 7327
rect 29779 7293 29788 7327
rect 29736 7284 29788 7293
rect 29920 7284 29972 7336
rect 31760 7327 31812 7336
rect 31760 7293 31769 7327
rect 31769 7293 31803 7327
rect 31803 7293 31812 7327
rect 31760 7284 31812 7293
rect 32404 7284 32456 7336
rect 34796 7488 34848 7540
rect 35992 7488 36044 7540
rect 36636 7531 36688 7540
rect 36636 7497 36645 7531
rect 36645 7497 36679 7531
rect 36679 7497 36688 7531
rect 36636 7488 36688 7497
rect 35900 7420 35952 7472
rect 33968 7352 34020 7404
rect 35072 7352 35124 7404
rect 35256 7395 35308 7404
rect 35256 7361 35265 7395
rect 35265 7361 35299 7395
rect 35299 7361 35308 7395
rect 35256 7352 35308 7361
rect 36084 7352 36136 7404
rect 36452 7327 36504 7336
rect 36452 7293 36461 7327
rect 36461 7293 36495 7327
rect 36495 7293 36504 7327
rect 36452 7284 36504 7293
rect 31944 7216 31996 7268
rect 28448 7148 28500 7200
rect 28816 7148 28868 7200
rect 29736 7148 29788 7200
rect 30656 7148 30708 7200
rect 32496 7216 32548 7268
rect 34980 7259 35032 7268
rect 34980 7225 34989 7259
rect 34989 7225 35023 7259
rect 35023 7225 35032 7259
rect 34980 7216 35032 7225
rect 35072 7259 35124 7268
rect 35072 7225 35081 7259
rect 35081 7225 35115 7259
rect 35115 7225 35124 7259
rect 35072 7216 35124 7225
rect 32680 7191 32732 7200
rect 32680 7157 32689 7191
rect 32689 7157 32723 7191
rect 32723 7157 32732 7191
rect 32680 7148 32732 7157
rect 37096 7148 37148 7200
rect 14315 7046 14367 7098
rect 14379 7046 14431 7098
rect 14443 7046 14495 7098
rect 14507 7046 14559 7098
rect 27648 7046 27700 7098
rect 27712 7046 27764 7098
rect 27776 7046 27828 7098
rect 27840 7046 27892 7098
rect 1952 6987 2004 6996
rect 1952 6953 1961 6987
rect 1961 6953 1995 6987
rect 1995 6953 2004 6987
rect 1952 6944 2004 6953
rect 3884 6987 3936 6996
rect 3884 6953 3893 6987
rect 3893 6953 3927 6987
rect 3927 6953 3936 6987
rect 3884 6944 3936 6953
rect 4068 6944 4120 6996
rect 3148 6876 3200 6928
rect 3976 6876 4028 6928
rect 6736 6944 6788 6996
rect 8024 6944 8076 6996
rect 9128 6987 9180 6996
rect 5908 6876 5960 6928
rect 9128 6953 9137 6987
rect 9137 6953 9171 6987
rect 9171 6953 9180 6987
rect 9128 6944 9180 6953
rect 9680 6944 9732 6996
rect 9864 6987 9916 6996
rect 9864 6953 9873 6987
rect 9873 6953 9907 6987
rect 9907 6953 9916 6987
rect 9864 6944 9916 6953
rect 10324 6944 10376 6996
rect 8392 6876 8444 6928
rect 13544 6944 13596 6996
rect 14648 6944 14700 6996
rect 16028 6944 16080 6996
rect 16764 6987 16816 6996
rect 16764 6953 16773 6987
rect 16773 6953 16807 6987
rect 16807 6953 16816 6987
rect 16764 6944 16816 6953
rect 20168 6987 20220 6996
rect 20168 6953 20177 6987
rect 20177 6953 20211 6987
rect 20211 6953 20220 6987
rect 20168 6944 20220 6953
rect 20812 6944 20864 6996
rect 21732 6944 21784 6996
rect 23756 6987 23808 6996
rect 23756 6953 23765 6987
rect 23765 6953 23799 6987
rect 23799 6953 23808 6987
rect 23756 6944 23808 6953
rect 10692 6876 10744 6928
rect 12624 6919 12676 6928
rect 12624 6885 12633 6919
rect 12633 6885 12667 6919
rect 12667 6885 12676 6919
rect 12624 6876 12676 6885
rect 13912 6876 13964 6928
rect 14188 6876 14240 6928
rect 15016 6876 15068 6928
rect 15660 6876 15712 6928
rect 17132 6919 17184 6928
rect 17132 6885 17141 6919
rect 17141 6885 17175 6919
rect 17175 6885 17184 6919
rect 17132 6876 17184 6885
rect 1860 6808 1912 6860
rect 3700 6808 3752 6860
rect 11980 6851 12032 6860
rect 2504 6783 2556 6792
rect 2504 6749 2513 6783
rect 2513 6749 2547 6783
rect 2547 6749 2556 6783
rect 2504 6740 2556 6749
rect 3056 6715 3108 6724
rect 3056 6681 3065 6715
rect 3065 6681 3099 6715
rect 3099 6681 3108 6715
rect 3056 6672 3108 6681
rect 3424 6647 3476 6656
rect 3424 6613 3433 6647
rect 3433 6613 3467 6647
rect 3467 6613 3476 6647
rect 3424 6604 3476 6613
rect 11980 6817 11989 6851
rect 11989 6817 12023 6851
rect 12023 6817 12032 6851
rect 11980 6808 12032 6817
rect 12716 6808 12768 6860
rect 13268 6808 13320 6860
rect 20352 6808 20404 6860
rect 21364 6808 21416 6860
rect 22836 6876 22888 6928
rect 21824 6808 21876 6860
rect 22468 6808 22520 6860
rect 24768 6944 24820 6996
rect 24216 6919 24268 6928
rect 24216 6885 24225 6919
rect 24225 6885 24259 6919
rect 24259 6885 24268 6919
rect 24216 6876 24268 6885
rect 24400 6876 24452 6928
rect 25320 6944 25372 6996
rect 25596 6987 25648 6996
rect 25596 6953 25605 6987
rect 25605 6953 25639 6987
rect 25639 6953 25648 6987
rect 25596 6944 25648 6953
rect 28448 6987 28500 6996
rect 28448 6953 28457 6987
rect 28457 6953 28491 6987
rect 28491 6953 28500 6987
rect 28448 6944 28500 6953
rect 30656 6987 30708 6996
rect 30656 6953 30665 6987
rect 30665 6953 30699 6987
rect 30699 6953 30708 6987
rect 30656 6944 30708 6953
rect 33968 6944 34020 6996
rect 34152 6987 34204 6996
rect 34152 6953 34161 6987
rect 34161 6953 34195 6987
rect 34195 6953 34204 6987
rect 34152 6944 34204 6953
rect 34980 6944 35032 6996
rect 24952 6876 25004 6928
rect 26608 6919 26660 6928
rect 26608 6885 26617 6919
rect 26617 6885 26651 6919
rect 26651 6885 26660 6919
rect 26608 6876 26660 6885
rect 26792 6876 26844 6928
rect 28908 6919 28960 6928
rect 28908 6885 28917 6919
rect 28917 6885 28951 6919
rect 28951 6885 28960 6919
rect 28908 6876 28960 6885
rect 32496 6919 32548 6928
rect 32496 6885 32499 6919
rect 32499 6885 32533 6919
rect 32533 6885 32548 6919
rect 32496 6876 32548 6885
rect 32680 6876 32732 6928
rect 34060 6876 34112 6928
rect 35072 6876 35124 6928
rect 35900 6876 35952 6928
rect 36268 6876 36320 6928
rect 29828 6808 29880 6860
rect 31116 6808 31168 6860
rect 31944 6808 31996 6860
rect 6000 6783 6052 6792
rect 5632 6604 5684 6656
rect 6000 6749 6009 6783
rect 6009 6749 6043 6783
rect 6043 6749 6052 6783
rect 6000 6740 6052 6749
rect 8116 6740 8168 6792
rect 11796 6740 11848 6792
rect 14188 6740 14240 6792
rect 14924 6740 14976 6792
rect 8208 6672 8260 6724
rect 17132 6740 17184 6792
rect 18604 6783 18656 6792
rect 18604 6749 18613 6783
rect 18613 6749 18647 6783
rect 18647 6749 18656 6783
rect 18604 6740 18656 6749
rect 18880 6783 18932 6792
rect 18880 6749 18889 6783
rect 18889 6749 18923 6783
rect 18923 6749 18932 6783
rect 18880 6740 18932 6749
rect 24308 6740 24360 6792
rect 24768 6783 24820 6792
rect 24768 6749 24777 6783
rect 24777 6749 24811 6783
rect 24811 6749 24820 6783
rect 24768 6740 24820 6749
rect 26700 6740 26752 6792
rect 28632 6740 28684 6792
rect 29644 6740 29696 6792
rect 17960 6672 18012 6724
rect 7196 6604 7248 6656
rect 12808 6604 12860 6656
rect 16212 6604 16264 6656
rect 18236 6604 18288 6656
rect 24400 6672 24452 6724
rect 35348 6740 35400 6792
rect 36360 6740 36412 6792
rect 37096 6740 37148 6792
rect 34888 6672 34940 6724
rect 36268 6672 36320 6724
rect 30196 6647 30248 6656
rect 30196 6613 30205 6647
rect 30205 6613 30239 6647
rect 30239 6613 30248 6647
rect 30196 6604 30248 6613
rect 30472 6604 30524 6656
rect 31760 6647 31812 6656
rect 31760 6613 31769 6647
rect 31769 6613 31803 6647
rect 31803 6613 31812 6647
rect 31760 6604 31812 6613
rect 34612 6604 34664 6656
rect 7648 6502 7700 6554
rect 7712 6502 7764 6554
rect 7776 6502 7828 6554
rect 7840 6502 7892 6554
rect 20982 6502 21034 6554
rect 21046 6502 21098 6554
rect 21110 6502 21162 6554
rect 21174 6502 21226 6554
rect 34315 6502 34367 6554
rect 34379 6502 34431 6554
rect 34443 6502 34495 6554
rect 34507 6502 34559 6554
rect 1860 6443 1912 6452
rect 1860 6409 1869 6443
rect 1869 6409 1903 6443
rect 1903 6409 1912 6443
rect 1860 6400 1912 6409
rect 2504 6400 2556 6452
rect 3792 6400 3844 6452
rect 5908 6400 5960 6452
rect 2596 6332 2648 6384
rect 3056 6375 3108 6384
rect 3056 6341 3065 6375
rect 3065 6341 3099 6375
rect 3099 6341 3108 6375
rect 3056 6332 3108 6341
rect 6368 6400 6420 6452
rect 8024 6400 8076 6452
rect 11704 6400 11756 6452
rect 13268 6400 13320 6452
rect 15752 6400 15804 6452
rect 17224 6400 17276 6452
rect 19800 6400 19852 6452
rect 20168 6400 20220 6452
rect 24216 6400 24268 6452
rect 15660 6375 15712 6384
rect 3424 6264 3476 6316
rect 4068 6264 4120 6316
rect 5264 6264 5316 6316
rect 4712 6196 4764 6248
rect 15660 6341 15669 6375
rect 15669 6341 15703 6375
rect 15703 6341 15712 6375
rect 15660 6332 15712 6341
rect 18236 6332 18288 6384
rect 10048 6264 10100 6316
rect 17408 6307 17460 6316
rect 17408 6273 17417 6307
rect 17417 6273 17451 6307
rect 17451 6273 17460 6307
rect 17408 6264 17460 6273
rect 17960 6264 18012 6316
rect 18512 6264 18564 6316
rect 19340 6264 19392 6316
rect 22836 6332 22888 6384
rect 23296 6332 23348 6384
rect 24768 6332 24820 6384
rect 21732 6307 21784 6316
rect 7196 6196 7248 6248
rect 2504 6128 2556 6180
rect 2596 6171 2648 6180
rect 2596 6137 2605 6171
rect 2605 6137 2639 6171
rect 2639 6137 2648 6171
rect 2596 6128 2648 6137
rect 4436 6128 4488 6180
rect 9312 6128 9364 6180
rect 10232 6128 10284 6180
rect 3332 6060 3384 6112
rect 3884 6103 3936 6112
rect 3884 6069 3893 6103
rect 3893 6069 3927 6103
rect 3927 6069 3936 6103
rect 3884 6060 3936 6069
rect 3976 6060 4028 6112
rect 5264 6103 5316 6112
rect 5264 6069 5273 6103
rect 5273 6069 5307 6103
rect 5307 6069 5316 6103
rect 5264 6060 5316 6069
rect 7104 6103 7156 6112
rect 7104 6069 7113 6103
rect 7113 6069 7147 6103
rect 7147 6069 7156 6103
rect 7104 6060 7156 6069
rect 8392 6060 8444 6112
rect 9220 6103 9272 6112
rect 9220 6069 9229 6103
rect 9229 6069 9263 6103
rect 9263 6069 9272 6103
rect 9220 6060 9272 6069
rect 10692 6103 10744 6112
rect 10692 6069 10701 6103
rect 10701 6069 10735 6103
rect 10735 6069 10744 6103
rect 10692 6060 10744 6069
rect 11980 6103 12032 6112
rect 11980 6069 11989 6103
rect 11989 6069 12023 6103
rect 12023 6069 12032 6103
rect 11980 6060 12032 6069
rect 12532 6103 12584 6112
rect 12532 6069 12541 6103
rect 12541 6069 12575 6103
rect 12575 6069 12584 6103
rect 12532 6060 12584 6069
rect 12808 6196 12860 6248
rect 12992 6239 13044 6248
rect 12992 6205 13001 6239
rect 13001 6205 13035 6239
rect 13035 6205 13044 6239
rect 12992 6196 13044 6205
rect 14648 6196 14700 6248
rect 16212 6239 16264 6248
rect 16212 6205 16221 6239
rect 16221 6205 16255 6239
rect 16255 6205 16264 6239
rect 16212 6196 16264 6205
rect 20168 6239 20220 6248
rect 20168 6205 20177 6239
rect 20177 6205 20211 6239
rect 20211 6205 20220 6239
rect 20168 6196 20220 6205
rect 21732 6273 21741 6307
rect 21741 6273 21775 6307
rect 21775 6273 21784 6307
rect 21732 6264 21784 6273
rect 22376 6196 22428 6248
rect 13084 6060 13136 6112
rect 13176 6060 13228 6112
rect 16028 6128 16080 6180
rect 17040 6128 17092 6180
rect 18236 6171 18288 6180
rect 18236 6137 18245 6171
rect 18245 6137 18279 6171
rect 18279 6137 18288 6171
rect 18236 6128 18288 6137
rect 17316 6060 17368 6112
rect 21456 6128 21508 6180
rect 21916 6128 21968 6180
rect 22836 6128 22888 6180
rect 21364 6103 21416 6112
rect 21364 6069 21373 6103
rect 21373 6069 21407 6103
rect 21407 6069 21416 6103
rect 21364 6060 21416 6069
rect 21824 6060 21876 6112
rect 23112 6128 23164 6180
rect 24400 6171 24452 6180
rect 24400 6137 24409 6171
rect 24409 6137 24443 6171
rect 24443 6137 24452 6171
rect 24400 6128 24452 6137
rect 26608 6400 26660 6452
rect 27344 6443 27396 6452
rect 27344 6409 27353 6443
rect 27353 6409 27387 6443
rect 27387 6409 27396 6443
rect 27344 6400 27396 6409
rect 28908 6400 28960 6452
rect 29460 6443 29512 6452
rect 29460 6409 29469 6443
rect 29469 6409 29503 6443
rect 29503 6409 29512 6443
rect 29460 6400 29512 6409
rect 31944 6400 31996 6452
rect 34060 6400 34112 6452
rect 34612 6443 34664 6452
rect 34612 6409 34621 6443
rect 34621 6409 34655 6443
rect 34655 6409 34664 6443
rect 34612 6400 34664 6409
rect 35900 6443 35952 6452
rect 35900 6409 35909 6443
rect 35909 6409 35943 6443
rect 35943 6409 35952 6443
rect 35900 6400 35952 6409
rect 36360 6443 36412 6452
rect 36360 6409 36369 6443
rect 36369 6409 36403 6443
rect 36403 6409 36412 6443
rect 36360 6400 36412 6409
rect 37004 6443 37056 6452
rect 37004 6409 37013 6443
rect 37013 6409 37047 6443
rect 37047 6409 37056 6443
rect 37004 6400 37056 6409
rect 26792 6332 26844 6384
rect 30196 6332 30248 6384
rect 25320 6307 25372 6316
rect 25320 6273 25329 6307
rect 25329 6273 25363 6307
rect 25363 6273 25372 6307
rect 25320 6264 25372 6273
rect 26700 6264 26752 6316
rect 30472 6264 30524 6316
rect 30932 6307 30984 6316
rect 30932 6273 30941 6307
rect 30941 6273 30975 6307
rect 30975 6273 30984 6307
rect 30932 6264 30984 6273
rect 31852 6264 31904 6316
rect 35256 6264 35308 6316
rect 35348 6307 35400 6316
rect 35348 6273 35357 6307
rect 35357 6273 35391 6307
rect 35391 6273 35400 6307
rect 35348 6264 35400 6273
rect 27344 6196 27396 6248
rect 28448 6196 28500 6248
rect 27068 6128 27120 6180
rect 28540 6128 28592 6180
rect 37004 6196 37056 6248
rect 30748 6171 30800 6180
rect 30748 6137 30757 6171
rect 30757 6137 30791 6171
rect 30791 6137 30800 6171
rect 30748 6128 30800 6137
rect 29828 6060 29880 6112
rect 30656 6060 30708 6112
rect 33048 6103 33100 6112
rect 33048 6069 33057 6103
rect 33057 6069 33091 6103
rect 33091 6069 33100 6103
rect 33048 6060 33100 6069
rect 34612 6060 34664 6112
rect 14315 5958 14367 6010
rect 14379 5958 14431 6010
rect 14443 5958 14495 6010
rect 14507 5958 14559 6010
rect 27648 5958 27700 6010
rect 27712 5958 27764 6010
rect 27776 5958 27828 6010
rect 27840 5958 27892 6010
rect 3148 5899 3200 5908
rect 3148 5865 3157 5899
rect 3157 5865 3191 5899
rect 3191 5865 3200 5899
rect 3148 5856 3200 5865
rect 3792 5856 3844 5908
rect 5632 5899 5684 5908
rect 2412 5788 2464 5840
rect 3976 5788 4028 5840
rect 5632 5865 5641 5899
rect 5641 5865 5675 5899
rect 5675 5865 5684 5899
rect 5632 5856 5684 5865
rect 10324 5856 10376 5908
rect 11796 5899 11848 5908
rect 11796 5865 11805 5899
rect 11805 5865 11839 5899
rect 11839 5865 11848 5899
rect 11796 5856 11848 5865
rect 15016 5899 15068 5908
rect 15016 5865 15025 5899
rect 15025 5865 15059 5899
rect 15059 5865 15068 5899
rect 15016 5856 15068 5865
rect 15568 5856 15620 5908
rect 6000 5788 6052 5840
rect 6644 5831 6696 5840
rect 6644 5797 6653 5831
rect 6653 5797 6687 5831
rect 6687 5797 6696 5831
rect 6644 5788 6696 5797
rect 8116 5788 8168 5840
rect 8392 5788 8444 5840
rect 10140 5788 10192 5840
rect 10692 5788 10744 5840
rect 12164 5831 12216 5840
rect 12164 5797 12173 5831
rect 12173 5797 12207 5831
rect 12207 5797 12216 5831
rect 12164 5788 12216 5797
rect 16212 5788 16264 5840
rect 17408 5856 17460 5908
rect 18052 5899 18104 5908
rect 18052 5865 18061 5899
rect 18061 5865 18095 5899
rect 18095 5865 18104 5899
rect 18052 5856 18104 5865
rect 18512 5856 18564 5908
rect 18604 5856 18656 5908
rect 22376 5899 22428 5908
rect 22376 5865 22385 5899
rect 22385 5865 22419 5899
rect 22419 5865 22428 5899
rect 22376 5856 22428 5865
rect 22468 5856 22520 5908
rect 23112 5899 23164 5908
rect 23112 5865 23121 5899
rect 23121 5865 23155 5899
rect 23155 5865 23164 5899
rect 23112 5856 23164 5865
rect 24860 5899 24912 5908
rect 24860 5865 24869 5899
rect 24869 5865 24903 5899
rect 24903 5865 24912 5899
rect 24860 5856 24912 5865
rect 29828 5856 29880 5908
rect 31116 5899 31168 5908
rect 31116 5865 31125 5899
rect 31125 5865 31159 5899
rect 31159 5865 31168 5899
rect 31116 5856 31168 5865
rect 34888 5899 34940 5908
rect 34888 5865 34897 5899
rect 34897 5865 34931 5899
rect 34931 5865 34940 5899
rect 34888 5856 34940 5865
rect 35256 5899 35308 5908
rect 35256 5865 35265 5899
rect 35265 5865 35299 5899
rect 35299 5865 35308 5899
rect 35256 5856 35308 5865
rect 17040 5788 17092 5840
rect 21916 5788 21968 5840
rect 23388 5831 23440 5840
rect 23388 5797 23397 5831
rect 23397 5797 23431 5831
rect 23431 5797 23440 5831
rect 23388 5788 23440 5797
rect 25136 5788 25188 5840
rect 27252 5831 27304 5840
rect 27252 5797 27261 5831
rect 27261 5797 27295 5831
rect 27295 5797 27304 5831
rect 27252 5788 27304 5797
rect 28908 5788 28960 5840
rect 13912 5763 13964 5772
rect 13912 5729 13921 5763
rect 13921 5729 13955 5763
rect 13955 5729 13964 5763
rect 13912 5720 13964 5729
rect 14096 5720 14148 5772
rect 15476 5720 15528 5772
rect 15568 5720 15620 5772
rect 19248 5763 19300 5772
rect 19248 5729 19257 5763
rect 19257 5729 19291 5763
rect 19291 5729 19300 5763
rect 19248 5720 19300 5729
rect 19800 5763 19852 5772
rect 19800 5729 19809 5763
rect 19809 5729 19843 5763
rect 19843 5729 19852 5763
rect 19800 5720 19852 5729
rect 24768 5763 24820 5772
rect 24768 5729 24777 5763
rect 24777 5729 24811 5763
rect 24811 5729 24820 5763
rect 24768 5720 24820 5729
rect 25228 5763 25280 5772
rect 25228 5729 25237 5763
rect 25237 5729 25271 5763
rect 25271 5729 25280 5763
rect 25228 5720 25280 5729
rect 30748 5720 30800 5772
rect 31944 5788 31996 5840
rect 33048 5788 33100 5840
rect 33968 5831 34020 5840
rect 33968 5797 33977 5831
rect 33977 5797 34011 5831
rect 34011 5797 34020 5831
rect 33968 5788 34020 5797
rect 35348 5788 35400 5840
rect 2228 5695 2280 5704
rect 2228 5661 2237 5695
rect 2237 5661 2271 5695
rect 2271 5661 2280 5695
rect 2228 5652 2280 5661
rect 2504 5652 2556 5704
rect 3792 5652 3844 5704
rect 1768 5559 1820 5568
rect 1768 5525 1777 5559
rect 1777 5525 1811 5559
rect 1811 5525 1820 5559
rect 1768 5516 1820 5525
rect 2596 5516 2648 5568
rect 3332 5516 3384 5568
rect 3700 5516 3752 5568
rect 6184 5516 6236 5568
rect 9312 5652 9364 5704
rect 10508 5695 10560 5704
rect 10508 5661 10517 5695
rect 10517 5661 10551 5695
rect 10551 5661 10560 5695
rect 10508 5652 10560 5661
rect 11796 5652 11848 5704
rect 12348 5695 12400 5704
rect 12348 5661 12357 5695
rect 12357 5661 12391 5695
rect 12391 5661 12400 5695
rect 12348 5652 12400 5661
rect 14648 5652 14700 5704
rect 18144 5652 18196 5704
rect 21272 5695 21324 5704
rect 21272 5661 21281 5695
rect 21281 5661 21315 5695
rect 21315 5661 21324 5695
rect 21272 5652 21324 5661
rect 21456 5695 21508 5704
rect 21456 5661 21465 5695
rect 21465 5661 21499 5695
rect 21499 5661 21508 5695
rect 21456 5652 21508 5661
rect 23296 5695 23348 5704
rect 23296 5661 23305 5695
rect 23305 5661 23339 5695
rect 23339 5661 23348 5695
rect 23296 5652 23348 5661
rect 24400 5652 24452 5704
rect 27160 5695 27212 5704
rect 27160 5661 27169 5695
rect 27169 5661 27203 5695
rect 27203 5661 27212 5695
rect 27160 5652 27212 5661
rect 28724 5652 28776 5704
rect 28816 5652 28868 5704
rect 33416 5652 33468 5704
rect 33876 5695 33928 5704
rect 33876 5661 33885 5695
rect 33885 5661 33919 5695
rect 33919 5661 33928 5695
rect 33876 5652 33928 5661
rect 15476 5584 15528 5636
rect 15936 5584 15988 5636
rect 17224 5584 17276 5636
rect 17408 5627 17460 5636
rect 17408 5593 17417 5627
rect 17417 5593 17451 5627
rect 17451 5593 17460 5627
rect 17408 5584 17460 5593
rect 30932 5584 30984 5636
rect 32772 5627 32824 5636
rect 32772 5593 32781 5627
rect 32781 5593 32815 5627
rect 32815 5593 32824 5627
rect 32772 5584 32824 5593
rect 8024 5516 8076 5568
rect 9036 5516 9088 5568
rect 11888 5516 11940 5568
rect 12992 5559 13044 5568
rect 12992 5525 13001 5559
rect 13001 5525 13035 5559
rect 13035 5525 13044 5559
rect 12992 5516 13044 5525
rect 13360 5559 13412 5568
rect 13360 5525 13369 5559
rect 13369 5525 13403 5559
rect 13403 5525 13412 5559
rect 13360 5516 13412 5525
rect 15292 5516 15344 5568
rect 16304 5516 16356 5568
rect 16764 5516 16816 5568
rect 24216 5559 24268 5568
rect 24216 5525 24225 5559
rect 24225 5525 24259 5559
rect 24259 5525 24268 5559
rect 24216 5516 24268 5525
rect 24308 5516 24360 5568
rect 25044 5516 25096 5568
rect 28632 5516 28684 5568
rect 7648 5414 7700 5466
rect 7712 5414 7764 5466
rect 7776 5414 7828 5466
rect 7840 5414 7892 5466
rect 20982 5414 21034 5466
rect 21046 5414 21098 5466
rect 21110 5414 21162 5466
rect 21174 5414 21226 5466
rect 34315 5414 34367 5466
rect 34379 5414 34431 5466
rect 34443 5414 34495 5466
rect 34507 5414 34559 5466
rect 3332 5355 3384 5364
rect 3332 5321 3341 5355
rect 3341 5321 3375 5355
rect 3375 5321 3384 5355
rect 3332 5312 3384 5321
rect 3976 5355 4028 5364
rect 3976 5321 3985 5355
rect 3985 5321 4019 5355
rect 4019 5321 4028 5355
rect 3976 5312 4028 5321
rect 4712 5355 4764 5364
rect 4712 5321 4721 5355
rect 4721 5321 4755 5355
rect 4755 5321 4764 5355
rect 4712 5312 4764 5321
rect 6644 5312 6696 5364
rect 8392 5355 8444 5364
rect 3700 5244 3752 5296
rect 1768 5176 1820 5228
rect 2136 5176 2188 5228
rect 2688 5176 2740 5228
rect 8392 5321 8401 5355
rect 8401 5321 8435 5355
rect 8435 5321 8444 5355
rect 8392 5312 8444 5321
rect 10140 5355 10192 5364
rect 10140 5321 10149 5355
rect 10149 5321 10183 5355
rect 10183 5321 10192 5355
rect 10140 5312 10192 5321
rect 9128 5244 9180 5296
rect 1492 5151 1544 5160
rect 1492 5117 1510 5151
rect 1510 5117 1544 5151
rect 1492 5108 1544 5117
rect 3976 5108 4028 5160
rect 7472 5176 7524 5228
rect 9312 5219 9364 5228
rect 9312 5185 9321 5219
rect 9321 5185 9355 5219
rect 9355 5185 9364 5219
rect 9312 5176 9364 5185
rect 12532 5312 12584 5364
rect 14096 5355 14148 5364
rect 14096 5321 14105 5355
rect 14105 5321 14139 5355
rect 14139 5321 14148 5355
rect 14096 5312 14148 5321
rect 17040 5355 17092 5364
rect 12164 5244 12216 5296
rect 13360 5176 13412 5228
rect 17040 5321 17049 5355
rect 17049 5321 17083 5355
rect 17083 5321 17092 5355
rect 17040 5312 17092 5321
rect 19248 5355 19300 5364
rect 19248 5321 19257 5355
rect 19257 5321 19291 5355
rect 19291 5321 19300 5355
rect 19248 5312 19300 5321
rect 23388 5312 23440 5364
rect 25228 5355 25280 5364
rect 25228 5321 25237 5355
rect 25237 5321 25271 5355
rect 25271 5321 25280 5355
rect 25228 5312 25280 5321
rect 26516 5312 26568 5364
rect 21456 5244 21508 5296
rect 15292 5219 15344 5228
rect 4528 5108 4580 5160
rect 5448 5151 5500 5160
rect 5448 5117 5457 5151
rect 5457 5117 5491 5151
rect 5491 5117 5500 5151
rect 5448 5108 5500 5117
rect 6000 5108 6052 5160
rect 15292 5185 15301 5219
rect 15301 5185 15335 5219
rect 15335 5185 15344 5219
rect 15292 5176 15344 5185
rect 17224 5176 17276 5228
rect 18052 5151 18104 5160
rect 2504 5040 2556 5092
rect 9036 5083 9088 5092
rect 3884 4972 3936 5024
rect 4436 4972 4488 5024
rect 5632 4972 5684 5024
rect 5724 4972 5776 5024
rect 7104 4972 7156 5024
rect 9036 5049 9045 5083
rect 9045 5049 9079 5083
rect 9079 5049 9088 5083
rect 9036 5040 9088 5049
rect 9128 5083 9180 5092
rect 9128 5049 9137 5083
rect 9137 5049 9171 5083
rect 9171 5049 9180 5083
rect 9128 5040 9180 5049
rect 10232 5040 10284 5092
rect 11520 5015 11572 5024
rect 11520 4981 11529 5015
rect 11529 4981 11563 5015
rect 11563 4981 11572 5015
rect 11520 4972 11572 4981
rect 14648 5040 14700 5092
rect 15200 5040 15252 5092
rect 16028 5083 16080 5092
rect 16028 5049 16037 5083
rect 16037 5049 16071 5083
rect 16071 5049 16080 5083
rect 16028 5040 16080 5049
rect 18052 5117 18061 5151
rect 18061 5117 18095 5151
rect 18095 5117 18104 5151
rect 18052 5108 18104 5117
rect 21272 5219 21324 5228
rect 19800 5108 19852 5160
rect 21272 5185 21281 5219
rect 21281 5185 21315 5219
rect 21315 5185 21324 5219
rect 21272 5176 21324 5185
rect 23020 5176 23072 5228
rect 25872 5108 25924 5160
rect 27160 5312 27212 5364
rect 28540 5312 28592 5364
rect 31944 5355 31996 5364
rect 31944 5321 31953 5355
rect 31953 5321 31987 5355
rect 31987 5321 31996 5355
rect 31944 5312 31996 5321
rect 33416 5355 33468 5364
rect 33416 5321 33425 5355
rect 33425 5321 33459 5355
rect 33459 5321 33468 5355
rect 33416 5312 33468 5321
rect 33876 5355 33928 5364
rect 33876 5321 33885 5355
rect 33885 5321 33919 5355
rect 33919 5321 33928 5355
rect 33876 5312 33928 5321
rect 33968 5312 34020 5364
rect 27252 5176 27304 5228
rect 26884 5108 26936 5160
rect 27528 5108 27580 5160
rect 29920 5176 29972 5228
rect 30932 5176 30984 5228
rect 29184 5108 29236 5160
rect 30656 5151 30708 5160
rect 30656 5117 30665 5151
rect 30665 5117 30699 5151
rect 30699 5117 30708 5151
rect 30656 5108 30708 5117
rect 32312 5108 32364 5160
rect 35348 5108 35400 5160
rect 20444 5083 20496 5092
rect 20444 5049 20453 5083
rect 20453 5049 20487 5083
rect 20487 5049 20496 5083
rect 20444 5040 20496 5049
rect 24216 5040 24268 5092
rect 24400 5083 24452 5092
rect 24400 5049 24409 5083
rect 24409 5049 24443 5083
rect 24443 5049 24452 5083
rect 24400 5040 24452 5049
rect 24952 5040 25004 5092
rect 13176 5015 13228 5024
rect 13176 4981 13185 5015
rect 13185 4981 13219 5015
rect 13219 4981 13228 5015
rect 13176 4972 13228 4981
rect 15568 5015 15620 5024
rect 15568 4981 15577 5015
rect 15577 4981 15611 5015
rect 15611 4981 15620 5015
rect 15568 4972 15620 4981
rect 16764 4972 16816 5024
rect 18144 5015 18196 5024
rect 18144 4981 18153 5015
rect 18153 4981 18187 5015
rect 18187 4981 18196 5015
rect 18144 4972 18196 4981
rect 21548 4972 21600 5024
rect 21916 4972 21968 5024
rect 24768 4972 24820 5024
rect 25228 4972 25280 5024
rect 25688 4972 25740 5024
rect 28816 4972 28868 5024
rect 29828 5015 29880 5024
rect 29828 4981 29837 5015
rect 29837 4981 29871 5015
rect 29871 4981 29880 5015
rect 32496 5083 32548 5092
rect 32496 5049 32505 5083
rect 32505 5049 32539 5083
rect 32539 5049 32548 5083
rect 32496 5040 32548 5049
rect 29828 4972 29880 4981
rect 32312 4972 32364 5024
rect 39580 5040 39632 5092
rect 14315 4870 14367 4922
rect 14379 4870 14431 4922
rect 14443 4870 14495 4922
rect 14507 4870 14559 4922
rect 27648 4870 27700 4922
rect 27712 4870 27764 4922
rect 27776 4870 27828 4922
rect 27840 4870 27892 4922
rect 2228 4768 2280 4820
rect 2044 4632 2096 4684
rect 8024 4768 8076 4820
rect 9312 4768 9364 4820
rect 10232 4811 10284 4820
rect 2504 4743 2556 4752
rect 2504 4709 2513 4743
rect 2513 4709 2547 4743
rect 2547 4709 2556 4743
rect 3792 4743 3844 4752
rect 2504 4700 2556 4709
rect 3792 4709 3801 4743
rect 3801 4709 3835 4743
rect 3835 4709 3844 4743
rect 3792 4700 3844 4709
rect 5724 4700 5776 4752
rect 9220 4700 9272 4752
rect 1584 4564 1636 4616
rect 4528 4632 4580 4684
rect 4988 4632 5040 4684
rect 5172 4632 5224 4684
rect 8392 4632 8444 4684
rect 8576 4675 8628 4684
rect 8576 4641 8585 4675
rect 8585 4641 8619 4675
rect 8619 4641 8628 4675
rect 8576 4632 8628 4641
rect 5632 4607 5684 4616
rect 5632 4573 5641 4607
rect 5641 4573 5675 4607
rect 5675 4573 5684 4607
rect 5632 4564 5684 4573
rect 9036 4607 9088 4616
rect 4252 4496 4304 4548
rect 9036 4573 9045 4607
rect 9045 4573 9079 4607
rect 9079 4573 9088 4607
rect 9036 4564 9088 4573
rect 10232 4777 10241 4811
rect 10241 4777 10275 4811
rect 10275 4777 10284 4811
rect 10232 4768 10284 4777
rect 13912 4811 13964 4820
rect 13912 4777 13921 4811
rect 13921 4777 13955 4811
rect 13955 4777 13964 4811
rect 13912 4768 13964 4777
rect 14648 4811 14700 4820
rect 14648 4777 14657 4811
rect 14657 4777 14691 4811
rect 14691 4777 14700 4811
rect 14648 4768 14700 4777
rect 15844 4768 15896 4820
rect 19800 4811 19852 4820
rect 19800 4777 19809 4811
rect 19809 4777 19843 4811
rect 19843 4777 19852 4811
rect 19800 4768 19852 4777
rect 21548 4811 21600 4820
rect 21548 4777 21557 4811
rect 21557 4777 21591 4811
rect 21591 4777 21600 4811
rect 21548 4768 21600 4777
rect 22008 4811 22060 4820
rect 22008 4777 22017 4811
rect 22017 4777 22051 4811
rect 22051 4777 22060 4811
rect 22008 4768 22060 4777
rect 24216 4768 24268 4820
rect 27344 4768 27396 4820
rect 28724 4768 28776 4820
rect 29368 4768 29420 4820
rect 29736 4768 29788 4820
rect 11520 4700 11572 4752
rect 15936 4700 15988 4752
rect 23296 4743 23348 4752
rect 23296 4709 23305 4743
rect 23305 4709 23339 4743
rect 23339 4709 23348 4743
rect 23296 4700 23348 4709
rect 23480 4700 23532 4752
rect 24860 4700 24912 4752
rect 25228 4700 25280 4752
rect 10048 4675 10100 4684
rect 10048 4641 10057 4675
rect 10057 4641 10091 4675
rect 10091 4641 10100 4675
rect 10048 4632 10100 4641
rect 13084 4675 13136 4684
rect 13084 4641 13093 4675
rect 13093 4641 13127 4675
rect 13127 4641 13136 4675
rect 13084 4632 13136 4641
rect 8024 4496 8076 4548
rect 12348 4564 12400 4616
rect 12992 4564 13044 4616
rect 13452 4632 13504 4684
rect 15016 4632 15068 4684
rect 16948 4675 17000 4684
rect 16948 4641 16957 4675
rect 16957 4641 16991 4675
rect 16991 4641 17000 4675
rect 16948 4632 17000 4641
rect 13360 4607 13412 4616
rect 13360 4573 13369 4607
rect 13369 4573 13403 4607
rect 13403 4573 13412 4607
rect 13360 4564 13412 4573
rect 15292 4564 15344 4616
rect 16304 4564 16356 4616
rect 17408 4564 17460 4616
rect 18880 4632 18932 4684
rect 19156 4632 19208 4684
rect 24952 4675 25004 4684
rect 20444 4564 20496 4616
rect 21640 4607 21692 4616
rect 21640 4573 21649 4607
rect 21649 4573 21683 4607
rect 21683 4573 21692 4607
rect 21640 4564 21692 4573
rect 16764 4539 16816 4548
rect 16764 4505 16773 4539
rect 16773 4505 16807 4539
rect 16807 4505 16816 4539
rect 16764 4496 16816 4505
rect 19248 4496 19300 4548
rect 24952 4641 24961 4675
rect 24961 4641 24995 4675
rect 24995 4641 25004 4675
rect 24952 4632 25004 4641
rect 25964 4632 26016 4684
rect 26792 4632 26844 4684
rect 28448 4700 28500 4752
rect 29828 4700 29880 4752
rect 30656 4768 30708 4820
rect 32312 4743 32364 4752
rect 32312 4709 32321 4743
rect 32321 4709 32355 4743
rect 32355 4709 32364 4743
rect 32312 4700 32364 4709
rect 30656 4632 30708 4684
rect 34152 4632 34204 4684
rect 35348 4632 35400 4684
rect 35808 4632 35860 4684
rect 23480 4607 23532 4616
rect 23480 4573 23489 4607
rect 23489 4573 23523 4607
rect 23523 4573 23532 4607
rect 23940 4607 23992 4616
rect 23480 4564 23532 4573
rect 23940 4573 23949 4607
rect 23949 4573 23983 4607
rect 23983 4573 23992 4607
rect 23940 4564 23992 4573
rect 27620 4607 27672 4616
rect 27620 4573 27629 4607
rect 27629 4573 27663 4607
rect 27663 4573 27672 4607
rect 27620 4564 27672 4573
rect 27988 4564 28040 4616
rect 29092 4564 29144 4616
rect 32864 4564 32916 4616
rect 29184 4496 29236 4548
rect 29644 4496 29696 4548
rect 32772 4539 32824 4548
rect 32772 4505 32781 4539
rect 32781 4505 32815 4539
rect 32815 4505 32824 4539
rect 32772 4496 32824 4505
rect 1952 4428 2004 4480
rect 3148 4471 3200 4480
rect 3148 4437 3157 4471
rect 3157 4437 3191 4471
rect 3191 4437 3200 4471
rect 3148 4428 3200 4437
rect 6000 4428 6052 4480
rect 7012 4428 7064 4480
rect 7472 4428 7524 4480
rect 10784 4428 10836 4480
rect 12716 4428 12768 4480
rect 15016 4471 15068 4480
rect 15016 4437 15025 4471
rect 15025 4437 15059 4471
rect 15059 4437 15068 4471
rect 15016 4428 15068 4437
rect 18144 4471 18196 4480
rect 18144 4437 18153 4471
rect 18153 4437 18187 4471
rect 18187 4437 18196 4471
rect 18144 4428 18196 4437
rect 25872 4428 25924 4480
rect 27252 4471 27304 4480
rect 27252 4437 27261 4471
rect 27261 4437 27295 4471
rect 27295 4437 27304 4471
rect 27252 4428 27304 4437
rect 28724 4471 28776 4480
rect 28724 4437 28733 4471
rect 28733 4437 28767 4471
rect 28767 4437 28776 4471
rect 28724 4428 28776 4437
rect 30472 4471 30524 4480
rect 30472 4437 30481 4471
rect 30481 4437 30515 4471
rect 30515 4437 30524 4471
rect 30472 4428 30524 4437
rect 32496 4428 32548 4480
rect 33968 4428 34020 4480
rect 7648 4326 7700 4378
rect 7712 4326 7764 4378
rect 7776 4326 7828 4378
rect 7840 4326 7892 4378
rect 20982 4326 21034 4378
rect 21046 4326 21098 4378
rect 21110 4326 21162 4378
rect 21174 4326 21226 4378
rect 34315 4326 34367 4378
rect 34379 4326 34431 4378
rect 34443 4326 34495 4378
rect 34507 4326 34559 4378
rect 2504 4267 2556 4276
rect 2504 4233 2513 4267
rect 2513 4233 2547 4267
rect 2547 4233 2556 4267
rect 2504 4224 2556 4233
rect 3056 4224 3108 4276
rect 2136 4131 2188 4140
rect 2136 4097 2145 4131
rect 2145 4097 2179 4131
rect 2179 4097 2188 4131
rect 2136 4088 2188 4097
rect 3056 4131 3108 4140
rect 3056 4097 3065 4131
rect 3065 4097 3099 4131
rect 3099 4097 3108 4131
rect 3056 4088 3108 4097
rect 5632 4224 5684 4276
rect 8116 4267 8168 4276
rect 8116 4233 8125 4267
rect 8125 4233 8159 4267
rect 8159 4233 8168 4267
rect 8116 4224 8168 4233
rect 8576 4224 8628 4276
rect 14832 4224 14884 4276
rect 16580 4224 16632 4276
rect 16764 4224 16816 4276
rect 23112 4224 23164 4276
rect 23388 4224 23440 4276
rect 27252 4224 27304 4276
rect 27528 4224 27580 4276
rect 28448 4267 28500 4276
rect 1676 4063 1728 4072
rect 1676 4029 1685 4063
rect 1685 4029 1719 4063
rect 1719 4029 1728 4063
rect 1676 4020 1728 4029
rect 1952 4063 2004 4072
rect 1952 4029 1961 4063
rect 1961 4029 1995 4063
rect 1995 4029 2004 4063
rect 1952 4020 2004 4029
rect 5540 4156 5592 4208
rect 11796 4156 11848 4208
rect 13084 4156 13136 4208
rect 15660 4156 15712 4208
rect 18788 4156 18840 4208
rect 21640 4156 21692 4208
rect 5264 4131 5316 4140
rect 5264 4097 5273 4131
rect 5273 4097 5307 4131
rect 5307 4097 5316 4131
rect 5264 4088 5316 4097
rect 6092 4088 6144 4140
rect 8024 4088 8076 4140
rect 10232 4088 10284 4140
rect 5172 4063 5224 4072
rect 5172 4029 5181 4063
rect 5181 4029 5215 4063
rect 5215 4029 5224 4063
rect 5172 4020 5224 4029
rect 8484 4063 8536 4072
rect 8484 4029 8493 4063
rect 8493 4029 8527 4063
rect 8527 4029 8536 4063
rect 8484 4020 8536 4029
rect 3148 3995 3200 4004
rect 3148 3961 3157 3995
rect 3157 3961 3191 3995
rect 3191 3961 3200 3995
rect 3148 3952 3200 3961
rect 7012 3995 7064 4004
rect 7012 3961 7021 3995
rect 7021 3961 7055 3995
rect 7055 3961 7064 3995
rect 7012 3952 7064 3961
rect 4160 3927 4212 3936
rect 4160 3893 4169 3927
rect 4169 3893 4203 3927
rect 4203 3893 4212 3927
rect 4160 3884 4212 3893
rect 4436 3884 4488 3936
rect 5724 3927 5776 3936
rect 5724 3893 5733 3927
rect 5733 3893 5767 3927
rect 5767 3893 5776 3927
rect 5724 3884 5776 3893
rect 6552 3927 6604 3936
rect 6552 3893 6561 3927
rect 6561 3893 6595 3927
rect 6595 3893 6604 3927
rect 6552 3884 6604 3893
rect 8668 3884 8720 3936
rect 10140 4020 10192 4072
rect 10508 4063 10560 4072
rect 10508 4029 10517 4063
rect 10517 4029 10551 4063
rect 10551 4029 10560 4063
rect 10508 4020 10560 4029
rect 10784 4063 10836 4072
rect 10784 4029 10793 4063
rect 10793 4029 10827 4063
rect 10827 4029 10836 4063
rect 10784 4020 10836 4029
rect 12716 4063 12768 4072
rect 12716 4029 12725 4063
rect 12725 4029 12759 4063
rect 12759 4029 12768 4063
rect 12716 4020 12768 4029
rect 9864 3952 9916 4004
rect 11244 3995 11296 4004
rect 11244 3961 11253 3995
rect 11253 3961 11287 3995
rect 11287 3961 11296 3995
rect 11244 3952 11296 3961
rect 11796 3995 11848 4004
rect 11796 3961 11805 3995
rect 11805 3961 11839 3995
rect 11839 3961 11848 3995
rect 11796 3952 11848 3961
rect 14188 4088 14240 4140
rect 15568 4131 15620 4140
rect 14832 4063 14884 4072
rect 14832 4029 14841 4063
rect 14841 4029 14875 4063
rect 14875 4029 14884 4063
rect 14832 4020 14884 4029
rect 14924 4063 14976 4072
rect 14924 4029 14933 4063
rect 14933 4029 14967 4063
rect 14967 4029 14976 4063
rect 15568 4097 15577 4131
rect 15577 4097 15611 4131
rect 15611 4097 15620 4131
rect 15568 4088 15620 4097
rect 16856 4088 16908 4140
rect 19340 4088 19392 4140
rect 20352 4088 20404 4140
rect 22008 4088 22060 4140
rect 24768 4156 24820 4208
rect 26792 4199 26844 4208
rect 26792 4165 26801 4199
rect 26801 4165 26835 4199
rect 26835 4165 26844 4199
rect 26792 4156 26844 4165
rect 23940 4088 23992 4140
rect 28448 4233 28457 4267
rect 28457 4233 28491 4267
rect 28491 4233 28500 4267
rect 28448 4224 28500 4233
rect 29092 4267 29144 4276
rect 29092 4233 29101 4267
rect 29101 4233 29135 4267
rect 29135 4233 29144 4267
rect 29092 4224 29144 4233
rect 29828 4224 29880 4276
rect 32312 4224 32364 4276
rect 32864 4267 32916 4276
rect 32864 4233 32873 4267
rect 32873 4233 32907 4267
rect 32907 4233 32916 4267
rect 32864 4224 32916 4233
rect 33968 4224 34020 4276
rect 30656 4199 30708 4208
rect 14924 4020 14976 4029
rect 16396 4063 16448 4072
rect 16396 4029 16405 4063
rect 16405 4029 16439 4063
rect 16439 4029 16448 4063
rect 16396 4020 16448 4029
rect 16580 4063 16632 4072
rect 16580 4029 16586 4063
rect 16586 4029 16632 4063
rect 16580 4020 16632 4029
rect 17960 4020 18012 4072
rect 18144 4020 18196 4072
rect 18880 4063 18932 4072
rect 18880 4029 18889 4063
rect 18889 4029 18923 4063
rect 18923 4029 18932 4063
rect 18880 4020 18932 4029
rect 21088 4020 21140 4072
rect 23388 3995 23440 4004
rect 23388 3961 23397 3995
rect 23397 3961 23431 3995
rect 23431 3961 23440 3995
rect 23388 3952 23440 3961
rect 25780 4020 25832 4072
rect 25688 3952 25740 4004
rect 29368 4131 29420 4140
rect 29368 4097 29377 4131
rect 29377 4097 29411 4131
rect 29411 4097 29420 4131
rect 29368 4088 29420 4097
rect 30656 4165 30665 4199
rect 30665 4165 30699 4199
rect 30699 4165 30708 4199
rect 30656 4156 30708 4165
rect 33416 4156 33468 4208
rect 30288 4020 30340 4072
rect 30656 4020 30708 4072
rect 31300 4063 31352 4072
rect 31300 4029 31309 4063
rect 31309 4029 31343 4063
rect 31343 4029 31352 4063
rect 31300 4020 31352 4029
rect 31484 4020 31536 4072
rect 10048 3927 10100 3936
rect 10048 3893 10057 3927
rect 10057 3893 10091 3927
rect 10091 3893 10100 3927
rect 10048 3884 10100 3893
rect 10232 3884 10284 3936
rect 10876 3884 10928 3936
rect 12624 3884 12676 3936
rect 14924 3884 14976 3936
rect 15936 3927 15988 3936
rect 15936 3893 15945 3927
rect 15945 3893 15979 3927
rect 15979 3893 15988 3927
rect 15936 3884 15988 3893
rect 16948 3884 17000 3936
rect 17408 3927 17460 3936
rect 17408 3893 17417 3927
rect 17417 3893 17451 3927
rect 17451 3893 17460 3927
rect 17408 3884 17460 3893
rect 19156 3884 19208 3936
rect 24768 3927 24820 3936
rect 24768 3893 24777 3927
rect 24777 3893 24811 3927
rect 24811 3893 24820 3927
rect 24768 3884 24820 3893
rect 27528 3995 27580 4004
rect 27528 3961 27537 3995
rect 27537 3961 27571 3995
rect 27571 3961 27580 3995
rect 27528 3952 27580 3961
rect 28724 3952 28776 4004
rect 29368 3952 29420 4004
rect 30932 3927 30984 3936
rect 30932 3893 30941 3927
rect 30941 3893 30975 3927
rect 30975 3893 30984 3927
rect 30932 3884 30984 3893
rect 34152 3884 34204 3936
rect 35348 3884 35400 3936
rect 14315 3782 14367 3834
rect 14379 3782 14431 3834
rect 14443 3782 14495 3834
rect 14507 3782 14559 3834
rect 27648 3782 27700 3834
rect 27712 3782 27764 3834
rect 27776 3782 27828 3834
rect 27840 3782 27892 3834
rect 1676 3723 1728 3732
rect 1676 3689 1685 3723
rect 1685 3689 1719 3723
rect 1719 3689 1728 3723
rect 1676 3680 1728 3689
rect 2044 3723 2096 3732
rect 2044 3689 2053 3723
rect 2053 3689 2087 3723
rect 2087 3689 2096 3723
rect 2044 3680 2096 3689
rect 2228 3723 2280 3732
rect 2228 3689 2237 3723
rect 2237 3689 2271 3723
rect 2271 3689 2280 3723
rect 2228 3680 2280 3689
rect 3148 3723 3200 3732
rect 3148 3689 3157 3723
rect 3157 3689 3191 3723
rect 3191 3689 3200 3723
rect 3148 3680 3200 3689
rect 4528 3680 4580 3732
rect 1952 3612 2004 3664
rect 2504 3544 2556 3596
rect 2872 3612 2924 3664
rect 4160 3612 4212 3664
rect 5172 3680 5224 3732
rect 6552 3680 6604 3732
rect 7196 3723 7248 3732
rect 7196 3689 7205 3723
rect 7205 3689 7239 3723
rect 7239 3689 7248 3723
rect 7196 3680 7248 3689
rect 8116 3680 8168 3732
rect 9956 3723 10008 3732
rect 9956 3689 9965 3723
rect 9965 3689 9999 3723
rect 9999 3689 10008 3723
rect 9956 3680 10008 3689
rect 11244 3680 11296 3732
rect 15476 3680 15528 3732
rect 15660 3680 15712 3732
rect 18972 3680 19024 3732
rect 20352 3723 20404 3732
rect 20352 3689 20361 3723
rect 20361 3689 20395 3723
rect 20395 3689 20404 3723
rect 20352 3680 20404 3689
rect 21088 3723 21140 3732
rect 21088 3689 21097 3723
rect 21097 3689 21131 3723
rect 21131 3689 21140 3723
rect 21088 3680 21140 3689
rect 23480 3723 23532 3732
rect 23480 3689 23489 3723
rect 23489 3689 23523 3723
rect 23523 3689 23532 3723
rect 24952 3723 25004 3732
rect 23480 3680 23532 3689
rect 24952 3689 24961 3723
rect 24961 3689 24995 3723
rect 24995 3689 25004 3723
rect 24952 3680 25004 3689
rect 25044 3680 25096 3732
rect 25964 3680 26016 3732
rect 26884 3680 26936 3732
rect 27988 3680 28040 3732
rect 28632 3680 28684 3732
rect 29368 3723 29420 3732
rect 6000 3612 6052 3664
rect 8392 3612 8444 3664
rect 4068 3544 4120 3596
rect 5080 3544 5132 3596
rect 7196 3587 7248 3596
rect 7196 3553 7205 3587
rect 7205 3553 7239 3587
rect 7239 3553 7248 3587
rect 7196 3544 7248 3553
rect 8116 3544 8168 3596
rect 9772 3587 9824 3596
rect 9772 3553 9781 3587
rect 9781 3553 9815 3587
rect 9815 3553 9824 3587
rect 9772 3544 9824 3553
rect 10508 3612 10560 3664
rect 15292 3655 15344 3664
rect 10876 3587 10928 3596
rect 10876 3553 10885 3587
rect 10885 3553 10919 3587
rect 10919 3553 10928 3587
rect 10876 3544 10928 3553
rect 15292 3621 15301 3655
rect 15301 3621 15335 3655
rect 15335 3621 15344 3655
rect 15292 3612 15344 3621
rect 12256 3544 12308 3596
rect 12716 3544 12768 3596
rect 13912 3587 13964 3596
rect 13912 3553 13921 3587
rect 13921 3553 13955 3587
rect 13955 3553 13964 3587
rect 13912 3544 13964 3553
rect 15200 3544 15252 3596
rect 16580 3612 16632 3664
rect 17408 3612 17460 3664
rect 10048 3476 10100 3528
rect 16764 3544 16816 3596
rect 16948 3544 17000 3596
rect 17960 3587 18012 3596
rect 17960 3553 17969 3587
rect 17969 3553 18003 3587
rect 18003 3553 18012 3587
rect 17960 3544 18012 3553
rect 18144 3587 18196 3596
rect 18144 3553 18153 3587
rect 18153 3553 18187 3587
rect 18187 3553 18196 3587
rect 18144 3544 18196 3553
rect 22008 3612 22060 3664
rect 23940 3655 23992 3664
rect 23940 3621 23949 3655
rect 23949 3621 23983 3655
rect 23983 3621 23992 3655
rect 23940 3612 23992 3621
rect 24216 3612 24268 3664
rect 28908 3612 28960 3664
rect 29368 3689 29377 3723
rect 29377 3689 29411 3723
rect 29411 3689 29420 3723
rect 29368 3680 29420 3689
rect 30472 3612 30524 3664
rect 31300 3612 31352 3664
rect 15660 3519 15712 3528
rect 15660 3485 15669 3519
rect 15669 3485 15703 3519
rect 15703 3485 15712 3519
rect 15660 3476 15712 3485
rect 17224 3519 17276 3528
rect 17224 3485 17233 3519
rect 17233 3485 17267 3519
rect 17267 3485 17276 3519
rect 25412 3587 25464 3596
rect 25412 3553 25421 3587
rect 25421 3553 25455 3587
rect 25455 3553 25464 3587
rect 25412 3544 25464 3553
rect 26792 3587 26844 3596
rect 26792 3553 26801 3587
rect 26801 3553 26835 3587
rect 26835 3553 26844 3587
rect 26792 3544 26844 3553
rect 27068 3587 27120 3596
rect 27068 3553 27077 3587
rect 27077 3553 27111 3587
rect 27111 3553 27120 3587
rect 27068 3544 27120 3553
rect 28356 3544 28408 3596
rect 30288 3587 30340 3596
rect 30288 3553 30297 3587
rect 30297 3553 30331 3587
rect 30331 3553 30340 3587
rect 30288 3544 30340 3553
rect 32680 3544 32732 3596
rect 33232 3587 33284 3596
rect 33232 3553 33250 3587
rect 33250 3553 33284 3587
rect 33232 3544 33284 3553
rect 38108 3544 38160 3596
rect 17224 3476 17276 3485
rect 24584 3519 24636 3528
rect 24584 3485 24593 3519
rect 24593 3485 24627 3519
rect 24627 3485 24636 3519
rect 24584 3476 24636 3485
rect 24768 3476 24820 3528
rect 28724 3476 28776 3528
rect 29644 3519 29696 3528
rect 29644 3485 29653 3519
rect 29653 3485 29687 3519
rect 29687 3485 29696 3519
rect 29644 3476 29696 3485
rect 7380 3408 7432 3460
rect 12440 3451 12492 3460
rect 12440 3417 12449 3451
rect 12449 3417 12483 3451
rect 12483 3417 12492 3451
rect 12440 3408 12492 3417
rect 14096 3408 14148 3460
rect 15568 3451 15620 3460
rect 15568 3417 15577 3451
rect 15577 3417 15611 3451
rect 15611 3417 15620 3451
rect 15568 3408 15620 3417
rect 16672 3408 16724 3460
rect 18788 3408 18840 3460
rect 19800 3451 19852 3460
rect 19800 3417 19809 3451
rect 19809 3417 19843 3451
rect 19843 3417 19852 3451
rect 19800 3408 19852 3417
rect 24216 3408 24268 3460
rect 39580 3408 39632 3460
rect 10324 3340 10376 3392
rect 12256 3383 12308 3392
rect 12256 3349 12265 3383
rect 12265 3349 12299 3383
rect 12299 3349 12308 3383
rect 12256 3340 12308 3349
rect 12624 3340 12676 3392
rect 13636 3340 13688 3392
rect 15200 3340 15252 3392
rect 15752 3383 15804 3392
rect 15752 3349 15761 3383
rect 15761 3349 15795 3383
rect 15795 3349 15804 3383
rect 15752 3340 15804 3349
rect 15844 3340 15896 3392
rect 17408 3340 17460 3392
rect 18880 3340 18932 3392
rect 20628 3340 20680 3392
rect 26056 3340 26108 3392
rect 7648 3238 7700 3290
rect 7712 3238 7764 3290
rect 7776 3238 7828 3290
rect 7840 3238 7892 3290
rect 20982 3238 21034 3290
rect 21046 3238 21098 3290
rect 21110 3238 21162 3290
rect 21174 3238 21226 3290
rect 34315 3238 34367 3290
rect 34379 3238 34431 3290
rect 34443 3238 34495 3290
rect 34507 3238 34559 3290
rect 2504 3179 2556 3188
rect 2504 3145 2513 3179
rect 2513 3145 2547 3179
rect 2547 3145 2556 3179
rect 2504 3136 2556 3145
rect 2872 3179 2924 3188
rect 2872 3145 2881 3179
rect 2881 3145 2915 3179
rect 2915 3145 2924 3179
rect 2872 3136 2924 3145
rect 4068 3179 4120 3188
rect 4068 3145 4077 3179
rect 4077 3145 4111 3179
rect 4111 3145 4120 3179
rect 4068 3136 4120 3145
rect 112 3068 164 3120
rect 3056 3043 3108 3052
rect 3056 3009 3065 3043
rect 3065 3009 3099 3043
rect 3099 3009 3108 3043
rect 3056 3000 3108 3009
rect 2964 2932 3016 2984
rect 6092 3136 6144 3188
rect 8116 3179 8168 3188
rect 8116 3145 8125 3179
rect 8125 3145 8159 3179
rect 8159 3145 8168 3179
rect 8116 3136 8168 3145
rect 10876 3136 10928 3188
rect 11888 3136 11940 3188
rect 17224 3136 17276 3188
rect 17960 3136 18012 3188
rect 22008 3136 22060 3188
rect 23112 3179 23164 3188
rect 23112 3145 23121 3179
rect 23121 3145 23155 3179
rect 23155 3145 23164 3179
rect 23112 3136 23164 3145
rect 28724 3179 28776 3188
rect 28724 3145 28733 3179
rect 28733 3145 28767 3179
rect 28767 3145 28776 3179
rect 28724 3136 28776 3145
rect 30472 3136 30524 3188
rect 32496 3136 32548 3188
rect 32680 3179 32732 3188
rect 32680 3145 32689 3179
rect 32689 3145 32723 3179
rect 32723 3145 32732 3179
rect 32680 3136 32732 3145
rect 33232 3179 33284 3188
rect 33232 3145 33241 3179
rect 33241 3145 33275 3179
rect 33275 3145 33284 3179
rect 33232 3136 33284 3145
rect 5908 3043 5960 3052
rect 5908 3009 5917 3043
rect 5917 3009 5951 3043
rect 5951 3009 5960 3043
rect 5908 3000 5960 3009
rect 9312 3068 9364 3120
rect 7472 3043 7524 3052
rect 7472 3009 7481 3043
rect 7481 3009 7515 3043
rect 7515 3009 7524 3043
rect 7472 3000 7524 3009
rect 7196 2975 7248 2984
rect 7196 2941 7205 2975
rect 7205 2941 7239 2975
rect 7239 2941 7248 2975
rect 7196 2932 7248 2941
rect 7380 2975 7432 2984
rect 7380 2941 7389 2975
rect 7389 2941 7423 2975
rect 7423 2941 7432 2975
rect 9128 3000 9180 3052
rect 10232 3068 10284 3120
rect 12716 3068 12768 3120
rect 14924 3068 14976 3120
rect 15568 3068 15620 3120
rect 16856 3111 16908 3120
rect 9772 3000 9824 3052
rect 10140 3000 10192 3052
rect 7380 2932 7432 2941
rect 8576 2975 8628 2984
rect 8576 2941 8585 2975
rect 8585 2941 8619 2975
rect 8619 2941 8628 2975
rect 8576 2932 8628 2941
rect 9864 2975 9916 2984
rect 9864 2941 9873 2975
rect 9873 2941 9907 2975
rect 9907 2941 9916 2975
rect 9864 2932 9916 2941
rect 11244 2932 11296 2984
rect 12256 2932 12308 2984
rect 9772 2864 9824 2916
rect 7104 2796 7156 2848
rect 8484 2839 8536 2848
rect 8484 2805 8493 2839
rect 8493 2805 8527 2839
rect 8527 2805 8536 2839
rect 8484 2796 8536 2805
rect 8760 2839 8812 2848
rect 8760 2805 8769 2839
rect 8769 2805 8803 2839
rect 8803 2805 8812 2839
rect 8760 2796 8812 2805
rect 9036 2839 9088 2848
rect 9036 2805 9045 2839
rect 9045 2805 9079 2839
rect 9079 2805 9088 2839
rect 9036 2796 9088 2805
rect 12532 2975 12584 2984
rect 12532 2941 12541 2975
rect 12541 2941 12575 2975
rect 12575 2941 12584 2975
rect 13912 3000 13964 3052
rect 16856 3077 16865 3111
rect 16865 3077 16899 3111
rect 16899 3077 16908 3111
rect 16856 3068 16908 3077
rect 18144 3000 18196 3052
rect 12532 2932 12584 2941
rect 12808 2932 12860 2984
rect 15108 2796 15160 2848
rect 15660 2864 15712 2916
rect 16672 2864 16724 2916
rect 17224 2864 17276 2916
rect 18788 2975 18840 2984
rect 18788 2941 18797 2975
rect 18797 2941 18831 2975
rect 18831 2941 18840 2975
rect 18788 2932 18840 2941
rect 19156 3068 19208 3120
rect 20352 3068 20404 3120
rect 24584 3068 24636 3120
rect 25504 3068 25556 3120
rect 32404 3111 32456 3120
rect 19524 3043 19576 3052
rect 19524 3009 19533 3043
rect 19533 3009 19567 3043
rect 19567 3009 19576 3043
rect 19524 3000 19576 3009
rect 19708 3000 19760 3052
rect 23388 3000 23440 3052
rect 19800 2932 19852 2984
rect 20352 2975 20404 2984
rect 20352 2941 20361 2975
rect 20361 2941 20395 2975
rect 20395 2941 20404 2975
rect 20352 2932 20404 2941
rect 19984 2864 20036 2916
rect 20536 2864 20588 2916
rect 23112 2932 23164 2984
rect 25964 2975 26016 2984
rect 25964 2941 25973 2975
rect 25973 2941 26007 2975
rect 26007 2941 26016 2975
rect 25964 2932 26016 2941
rect 26056 2932 26108 2984
rect 16580 2796 16632 2848
rect 18604 2796 18656 2848
rect 20352 2796 20404 2848
rect 24032 2839 24084 2848
rect 24032 2805 24041 2839
rect 24041 2805 24075 2839
rect 24075 2805 24084 2839
rect 25412 2839 25464 2848
rect 24032 2796 24084 2805
rect 25412 2805 25421 2839
rect 25421 2805 25455 2839
rect 25455 2805 25464 2839
rect 25412 2796 25464 2805
rect 25780 2839 25832 2848
rect 25780 2805 25789 2839
rect 25789 2805 25823 2839
rect 25823 2805 25832 2839
rect 25780 2796 25832 2805
rect 27068 3000 27120 3052
rect 27988 3043 28040 3052
rect 27344 2932 27396 2984
rect 27988 3009 27997 3043
rect 27997 3009 28031 3043
rect 28031 3009 28040 3043
rect 27988 3000 28040 3009
rect 32404 3077 32413 3111
rect 32413 3077 32447 3111
rect 32447 3077 32456 3111
rect 32404 3068 32456 3077
rect 28080 2932 28132 2984
rect 29276 2975 29328 2984
rect 29276 2941 29285 2975
rect 29285 2941 29319 2975
rect 29319 2941 29328 2975
rect 29276 2932 29328 2941
rect 30748 3000 30800 3052
rect 29920 2932 29972 2984
rect 31300 2932 31352 2984
rect 28356 2839 28408 2848
rect 28356 2805 28365 2839
rect 28365 2805 28399 2839
rect 28399 2805 28408 2839
rect 28356 2796 28408 2805
rect 30196 2796 30248 2848
rect 14315 2694 14367 2746
rect 14379 2694 14431 2746
rect 14443 2694 14495 2746
rect 14507 2694 14559 2746
rect 27648 2694 27700 2746
rect 27712 2694 27764 2746
rect 27776 2694 27828 2746
rect 27840 2694 27892 2746
rect 2872 2592 2924 2644
rect 4252 2592 4304 2644
rect 6184 2592 6236 2644
rect 2504 2456 2556 2508
rect 4804 2524 4856 2576
rect 3976 2456 4028 2508
rect 1308 2388 1360 2440
rect 6000 2499 6052 2508
rect 6000 2465 6009 2499
rect 6009 2465 6043 2499
rect 6043 2465 6052 2499
rect 6000 2456 6052 2465
rect 6644 2456 6696 2508
rect 7104 2499 7156 2508
rect 7104 2465 7113 2499
rect 7113 2465 7147 2499
rect 7147 2465 7156 2499
rect 7104 2456 7156 2465
rect 7288 2456 7340 2508
rect 7380 2499 7432 2508
rect 7380 2465 7389 2499
rect 7389 2465 7423 2499
rect 7423 2465 7432 2499
rect 8116 2524 8168 2576
rect 9036 2524 9088 2576
rect 7380 2456 7432 2465
rect 9220 2456 9272 2508
rect 9864 2592 9916 2644
rect 12716 2592 12768 2644
rect 12992 2592 13044 2644
rect 11796 2524 11848 2576
rect 12532 2524 12584 2576
rect 12900 2524 12952 2576
rect 15292 2592 15344 2644
rect 16488 2524 16540 2576
rect 17224 2567 17276 2576
rect 12440 2456 12492 2508
rect 12624 2499 12676 2508
rect 12624 2465 12633 2499
rect 12633 2465 12667 2499
rect 12667 2465 12676 2499
rect 12624 2456 12676 2465
rect 112 2320 164 2372
rect 2504 2295 2556 2304
rect 2504 2261 2513 2295
rect 2513 2261 2547 2295
rect 2547 2261 2556 2295
rect 2504 2252 2556 2261
rect 6276 2295 6328 2304
rect 6276 2261 6285 2295
rect 6285 2261 6319 2295
rect 6319 2261 6328 2295
rect 6276 2252 6328 2261
rect 6644 2295 6696 2304
rect 6644 2261 6653 2295
rect 6653 2261 6687 2295
rect 6687 2261 6696 2295
rect 6644 2252 6696 2261
rect 8760 2388 8812 2440
rect 14188 2431 14240 2440
rect 14188 2397 14197 2431
rect 14197 2397 14231 2431
rect 14231 2397 14240 2431
rect 14188 2388 14240 2397
rect 15844 2456 15896 2508
rect 15936 2456 15988 2508
rect 16396 2499 16448 2508
rect 16396 2465 16405 2499
rect 16405 2465 16439 2499
rect 16439 2465 16448 2499
rect 16396 2456 16448 2465
rect 17224 2533 17233 2567
rect 17233 2533 17267 2567
rect 17267 2533 17276 2567
rect 17224 2524 17276 2533
rect 17776 2567 17828 2576
rect 17776 2533 17785 2567
rect 17785 2533 17819 2567
rect 17819 2533 17828 2567
rect 17776 2524 17828 2533
rect 18328 2499 18380 2508
rect 18328 2465 18337 2499
rect 18337 2465 18371 2499
rect 18371 2465 18380 2499
rect 18328 2456 18380 2465
rect 18420 2499 18472 2508
rect 18420 2465 18429 2499
rect 18429 2465 18463 2499
rect 18463 2465 18472 2499
rect 18604 2499 18656 2508
rect 18420 2456 18472 2465
rect 18604 2465 18613 2499
rect 18613 2465 18647 2499
rect 18647 2465 18656 2499
rect 18604 2456 18656 2465
rect 18972 2592 19024 2644
rect 20536 2635 20588 2644
rect 20536 2601 20545 2635
rect 20545 2601 20579 2635
rect 20579 2601 20588 2635
rect 20536 2592 20588 2601
rect 20628 2592 20680 2644
rect 21088 2592 21140 2644
rect 23480 2592 23532 2644
rect 24584 2592 24636 2644
rect 19984 2524 20036 2576
rect 24032 2567 24084 2576
rect 21088 2499 21140 2508
rect 16948 2388 17000 2440
rect 16120 2320 16172 2372
rect 21088 2465 21097 2499
rect 21097 2465 21131 2499
rect 21131 2465 21140 2499
rect 21088 2456 21140 2465
rect 24032 2533 24041 2567
rect 24041 2533 24075 2567
rect 24075 2533 24084 2567
rect 24032 2524 24084 2533
rect 26792 2592 26844 2644
rect 27344 2635 27396 2644
rect 27344 2601 27353 2635
rect 27353 2601 27387 2635
rect 27387 2601 27396 2635
rect 27344 2592 27396 2601
rect 20536 2388 20588 2440
rect 22652 2456 22704 2508
rect 24216 2456 24268 2508
rect 25596 2499 25648 2508
rect 25596 2465 25605 2499
rect 25605 2465 25639 2499
rect 25639 2465 25648 2499
rect 25596 2456 25648 2465
rect 27252 2456 27304 2508
rect 29276 2635 29328 2644
rect 29276 2601 29285 2635
rect 29285 2601 29319 2635
rect 29319 2601 29328 2635
rect 29276 2592 29328 2601
rect 29920 2635 29972 2644
rect 29920 2601 29929 2635
rect 29929 2601 29963 2635
rect 29963 2601 29972 2635
rect 29920 2592 29972 2601
rect 30196 2592 30248 2644
rect 32404 2592 32456 2644
rect 28816 2524 28868 2576
rect 28448 2499 28500 2508
rect 28448 2465 28457 2499
rect 28457 2465 28491 2499
rect 28491 2465 28500 2499
rect 28448 2456 28500 2465
rect 9036 2252 9088 2304
rect 9220 2295 9272 2304
rect 9220 2261 9229 2295
rect 9229 2261 9263 2295
rect 9263 2261 9272 2295
rect 9220 2252 9272 2261
rect 10140 2295 10192 2304
rect 10140 2261 10149 2295
rect 10149 2261 10183 2295
rect 10183 2261 10192 2295
rect 10140 2252 10192 2261
rect 10232 2252 10284 2304
rect 13636 2295 13688 2304
rect 13636 2261 13645 2295
rect 13645 2261 13679 2295
rect 13679 2261 13688 2295
rect 13636 2252 13688 2261
rect 14096 2295 14148 2304
rect 14096 2261 14105 2295
rect 14105 2261 14139 2295
rect 14139 2261 14148 2295
rect 15200 2295 15252 2304
rect 14096 2252 14148 2261
rect 15200 2261 15209 2295
rect 15209 2261 15243 2295
rect 15243 2261 15252 2295
rect 15200 2252 15252 2261
rect 16396 2252 16448 2304
rect 18328 2252 18380 2304
rect 18604 2252 18656 2304
rect 26792 2320 26844 2372
rect 27252 2252 27304 2304
rect 28448 2320 28500 2372
rect 28540 2320 28592 2372
rect 7648 2150 7700 2202
rect 7712 2150 7764 2202
rect 7776 2150 7828 2202
rect 7840 2150 7892 2202
rect 20982 2150 21034 2202
rect 21046 2150 21098 2202
rect 21110 2150 21162 2202
rect 21174 2150 21226 2202
rect 34315 2150 34367 2202
rect 34379 2150 34431 2202
rect 34443 2150 34495 2202
rect 34507 2150 34559 2202
rect 6000 2048 6052 2100
rect 13636 2048 13688 2100
rect 6276 1980 6328 2032
rect 7380 1980 7432 2032
rect 8668 1980 8720 2032
rect 10140 1980 10192 2032
rect 14096 1980 14148 2032
rect 7104 76 7156 128
rect 8484 76 8536 128
rect 10324 76 10376 128
rect 12808 76 12860 128
rect 21364 76 21416 128
rect 24492 76 24544 128
<< metal2 >>
rect 1766 15586 1822 16000
rect 5354 15586 5410 16000
rect 9034 15586 9090 16000
rect 12622 15586 12678 16000
rect 1766 15558 1900 15586
rect 1766 15520 1822 15558
rect 1122 15056 1178 15065
rect 1122 14991 1178 15000
rect 110 13696 166 13705
rect 110 13631 166 13640
rect 124 13190 152 13631
rect 112 13184 164 13190
rect 112 13126 164 13132
rect 112 12640 164 12646
rect 112 12582 164 12588
rect 124 11801 152 12582
rect 1136 11898 1164 14991
rect 1768 12640 1820 12646
rect 1768 12582 1820 12588
rect 1582 12472 1638 12481
rect 1582 12407 1638 12416
rect 1596 12170 1624 12407
rect 1584 12164 1636 12170
rect 1584 12106 1636 12112
rect 1124 11892 1176 11898
rect 1124 11834 1176 11840
rect 1676 11824 1728 11830
rect 110 11792 166 11801
rect 1676 11766 1728 11772
rect 110 11727 166 11736
rect 1688 11354 1716 11766
rect 1676 11348 1728 11354
rect 1504 11308 1676 11336
rect 1398 10296 1454 10305
rect 1398 10231 1454 10240
rect 110 9888 166 9897
rect 110 9823 166 9832
rect 124 9722 152 9823
rect 112 9716 164 9722
rect 112 9658 164 9664
rect 1412 9518 1440 10231
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 112 9376 164 9382
rect 112 9318 164 9324
rect 124 8945 152 9318
rect 110 8936 166 8945
rect 20 8900 72 8906
rect 110 8871 166 8880
rect 20 8842 72 8848
rect 32 7993 60 8842
rect 18 7984 74 7993
rect 18 7919 74 7928
rect 1504 5817 1532 11308
rect 1676 11290 1728 11296
rect 1780 10713 1808 12582
rect 1766 10704 1822 10713
rect 1766 10639 1822 10648
rect 1584 10600 1636 10606
rect 1584 10542 1636 10548
rect 1596 10266 1624 10542
rect 1676 10464 1728 10470
rect 1676 10406 1728 10412
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 1490 5808 1546 5817
rect 1490 5743 1546 5752
rect 1504 5166 1532 5743
rect 1492 5160 1544 5166
rect 1492 5102 1544 5108
rect 1596 4622 1624 10202
rect 1688 5001 1716 10406
rect 1780 6848 1808 10639
rect 1872 8566 1900 15558
rect 5354 15558 5672 15586
rect 5354 15520 5410 15558
rect 1950 14240 2006 14249
rect 1950 14175 2006 14184
rect 1964 11898 1992 14175
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 1952 11892 2004 11898
rect 1952 11834 2004 11840
rect 2056 11762 2084 12242
rect 2688 12232 2740 12238
rect 2688 12174 2740 12180
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 2056 11665 2084 11698
rect 2042 11656 2098 11665
rect 2042 11591 2098 11600
rect 2412 11212 2464 11218
rect 2412 11154 2464 11160
rect 2136 10532 2188 10538
rect 2136 10474 2188 10480
rect 2044 10192 2096 10198
rect 2044 10134 2096 10140
rect 1950 9616 2006 9625
rect 1950 9551 2006 9560
rect 1964 9518 1992 9551
rect 1952 9512 2004 9518
rect 1952 9454 2004 9460
rect 2056 9178 2084 10134
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 1860 8560 1912 8566
rect 1860 8502 1912 8508
rect 2148 8498 2176 10474
rect 2424 10470 2452 11154
rect 2700 10674 2728 12174
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2872 11212 2924 11218
rect 2872 11154 2924 11160
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 2688 10668 2740 10674
rect 2688 10610 2740 10616
rect 2412 10464 2464 10470
rect 2412 10406 2464 10412
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 2240 9042 2268 10202
rect 2792 9586 2820 11086
rect 2884 10742 2912 11154
rect 2872 10736 2924 10742
rect 2872 10678 2924 10684
rect 2884 10606 2912 10678
rect 2872 10600 2924 10606
rect 2872 10542 2924 10548
rect 2884 10130 2912 10542
rect 2976 10305 3004 11494
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 3056 10668 3108 10674
rect 3056 10610 3108 10616
rect 2962 10296 3018 10305
rect 3068 10266 3096 10610
rect 3160 10538 3188 10950
rect 4160 10736 4212 10742
rect 4160 10678 4212 10684
rect 3148 10532 3200 10538
rect 3148 10474 3200 10480
rect 2962 10231 3018 10240
rect 3056 10260 3108 10266
rect 2872 10124 2924 10130
rect 2872 10066 2924 10072
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 2504 9376 2556 9382
rect 2504 9318 2556 9324
rect 2516 9178 2544 9318
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2228 9036 2280 9042
rect 2228 8978 2280 8984
rect 2240 8634 2268 8978
rect 2228 8628 2280 8634
rect 2228 8570 2280 8576
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 2148 8090 2176 8434
rect 2516 8294 2544 9114
rect 2792 9110 2820 9522
rect 2780 9104 2832 9110
rect 2780 9046 2832 9052
rect 2504 8288 2556 8294
rect 2504 8230 2556 8236
rect 2136 8084 2188 8090
rect 2136 8026 2188 8032
rect 2412 8016 2464 8022
rect 2412 7958 2464 7964
rect 1952 7812 2004 7818
rect 1952 7754 2004 7760
rect 1964 7002 1992 7754
rect 2424 7546 2452 7958
rect 2688 7744 2740 7750
rect 2688 7686 2740 7692
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 1860 6860 1912 6866
rect 1780 6820 1860 6848
rect 1860 6802 1912 6808
rect 1872 6458 1900 6802
rect 2504 6792 2556 6798
rect 2504 6734 2556 6740
rect 2516 6458 2544 6734
rect 1860 6452 1912 6458
rect 1860 6394 1912 6400
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2608 6390 2636 7482
rect 2700 7410 2728 7686
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 2596 6384 2648 6390
rect 2596 6326 2648 6332
rect 2504 6180 2556 6186
rect 2504 6122 2556 6128
rect 2596 6180 2648 6186
rect 2596 6122 2648 6128
rect 2412 5840 2464 5846
rect 2412 5782 2464 5788
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 1768 5568 1820 5574
rect 1768 5510 1820 5516
rect 1780 5234 1808 5510
rect 1768 5228 1820 5234
rect 1768 5170 1820 5176
rect 2136 5228 2188 5234
rect 2136 5170 2188 5176
rect 1674 4992 1730 5001
rect 1674 4927 1730 4936
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 1688 4078 1716 4927
rect 2044 4684 2096 4690
rect 2044 4626 2096 4632
rect 1952 4480 2004 4486
rect 1952 4422 2004 4428
rect 1964 4078 1992 4422
rect 1676 4072 1728 4078
rect 1676 4014 1728 4020
rect 1952 4072 2004 4078
rect 1952 4014 2004 4020
rect 1688 3738 1716 4014
rect 1676 3732 1728 3738
rect 1676 3674 1728 3680
rect 1964 3670 1992 4014
rect 2056 3738 2084 4626
rect 2148 4146 2176 5170
rect 2240 4826 2268 5646
rect 2424 5080 2452 5782
rect 2516 5710 2544 6122
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 2608 5574 2636 6122
rect 2596 5568 2648 5574
rect 2596 5510 2648 5516
rect 2700 5234 2728 7346
rect 2778 6760 2834 6769
rect 2778 6695 2834 6704
rect 2688 5228 2740 5234
rect 2688 5170 2740 5176
rect 2504 5092 2556 5098
rect 2424 5052 2504 5080
rect 2504 5034 2556 5040
rect 2228 4820 2280 4826
rect 2228 4762 2280 4768
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 2240 3738 2268 4762
rect 2516 4758 2544 5034
rect 2504 4752 2556 4758
rect 2504 4694 2556 4700
rect 2516 4282 2544 4694
rect 2504 4276 2556 4282
rect 2504 4218 2556 4224
rect 2792 4154 2820 6695
rect 2976 5681 3004 10231
rect 3056 10202 3108 10208
rect 3160 8634 3188 10474
rect 3976 10192 4028 10198
rect 3976 10134 4028 10140
rect 3608 10056 3660 10062
rect 3608 9998 3660 10004
rect 3240 9444 3292 9450
rect 3240 9386 3292 9392
rect 3252 9178 3280 9386
rect 3620 9382 3648 9998
rect 3988 9518 4016 10134
rect 4172 10062 4200 10678
rect 4540 10305 4568 11698
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4724 10470 4752 11154
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4526 10296 4582 10305
rect 4526 10231 4582 10240
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 3332 8288 3384 8294
rect 3332 8230 3384 8236
rect 3344 7206 3372 8230
rect 3424 7880 3476 7886
rect 3424 7822 3476 7828
rect 3436 7342 3464 7822
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3148 6928 3200 6934
rect 3148 6870 3200 6876
rect 3056 6724 3108 6730
rect 3056 6666 3108 6672
rect 3068 6390 3096 6666
rect 3056 6384 3108 6390
rect 3056 6326 3108 6332
rect 2962 5672 3018 5681
rect 2962 5607 3018 5616
rect 3068 4282 3096 6326
rect 3160 5914 3188 6870
rect 3344 6118 3372 7142
rect 3436 6662 3464 7278
rect 3620 6769 3648 9318
rect 3698 9208 3754 9217
rect 3698 9143 3754 9152
rect 3712 7954 3740 9143
rect 3988 9110 4016 9454
rect 4172 9178 4200 9998
rect 4540 9568 4568 10231
rect 4724 9994 4752 10406
rect 4712 9988 4764 9994
rect 4712 9930 4764 9936
rect 4724 9586 4752 9930
rect 4712 9580 4764 9586
rect 4540 9540 4660 9568
rect 4436 9444 4488 9450
rect 4436 9386 4488 9392
rect 4448 9178 4476 9386
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 4436 9172 4488 9178
rect 4436 9114 4488 9120
rect 3976 9104 4028 9110
rect 3976 9046 4028 9052
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 4080 8634 4108 8978
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 3700 7948 3752 7954
rect 3700 7890 3752 7896
rect 3712 7546 3740 7890
rect 3700 7540 3752 7546
rect 3700 7482 3752 7488
rect 3700 6860 3752 6866
rect 3700 6802 3752 6808
rect 3606 6760 3662 6769
rect 3606 6695 3662 6704
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3436 6322 3464 6598
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 3712 5574 3740 6802
rect 3804 6458 3832 8434
rect 3884 8356 3936 8362
rect 3884 8298 3936 8304
rect 4528 8356 4580 8362
rect 4528 8298 4580 8304
rect 3896 8090 3924 8298
rect 4540 8090 4568 8298
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3976 8084 4028 8090
rect 3976 8026 4028 8032
rect 4528 8084 4580 8090
rect 4528 8026 4580 8032
rect 3896 7478 3924 8026
rect 3884 7472 3936 7478
rect 3988 7449 4016 8026
rect 4540 7546 4568 8026
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 3884 7414 3936 7420
rect 3974 7440 4030 7449
rect 3974 7375 4030 7384
rect 4540 7342 4568 7482
rect 4632 7342 4660 9540
rect 4712 9522 4764 9528
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 4528 7336 4580 7342
rect 4528 7278 4580 7284
rect 4620 7336 4672 7342
rect 4620 7278 4672 7284
rect 3896 7002 3924 7278
rect 3884 6996 3936 7002
rect 3884 6938 3936 6944
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 3976 6928 4028 6934
rect 3976 6870 4028 6876
rect 3792 6452 3844 6458
rect 3792 6394 3844 6400
rect 3804 5914 3832 6394
rect 3988 6118 4016 6870
rect 4080 6322 4108 6938
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 4712 6248 4764 6254
rect 4712 6190 4764 6196
rect 4436 6180 4488 6186
rect 4436 6122 4488 6128
rect 3884 6112 3936 6118
rect 3884 6054 3936 6060
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3332 5568 3384 5574
rect 3332 5510 3384 5516
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 3344 5370 3372 5510
rect 3332 5364 3384 5370
rect 3332 5306 3384 5312
rect 3712 5302 3740 5510
rect 3700 5296 3752 5302
rect 3700 5238 3752 5244
rect 3804 4758 3832 5646
rect 3896 5030 3924 6054
rect 3988 5846 4016 6054
rect 3976 5840 4028 5846
rect 3976 5782 4028 5788
rect 3988 5370 4016 5782
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 3976 5160 4028 5166
rect 3976 5102 4028 5108
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 3792 4752 3844 4758
rect 3792 4694 3844 4700
rect 3148 4480 3200 4486
rect 3148 4422 3200 4428
rect 3056 4276 3108 4282
rect 2516 4126 2820 4154
rect 2976 4236 3056 4264
rect 2044 3732 2096 3738
rect 2044 3674 2096 3680
rect 2228 3732 2280 3738
rect 2228 3674 2280 3680
rect 1952 3664 2004 3670
rect 1952 3606 2004 3612
rect 2516 3602 2544 4126
rect 2872 3664 2924 3670
rect 2872 3606 2924 3612
rect 2504 3596 2556 3602
rect 2504 3538 2556 3544
rect 110 3224 166 3233
rect 2516 3194 2544 3538
rect 2884 3194 2912 3606
rect 110 3159 166 3168
rect 2504 3188 2556 3194
rect 124 3126 152 3159
rect 2504 3130 2556 3136
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 112 3120 164 3126
rect 112 3062 164 3068
rect 2884 2650 2912 3130
rect 2976 2990 3004 4236
rect 3056 4218 3108 4224
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 3068 3058 3096 4082
rect 3160 4010 3188 4422
rect 3148 4004 3200 4010
rect 3148 3946 3200 3952
rect 3160 3738 3188 3946
rect 3148 3732 3200 3738
rect 3148 3674 3200 3680
rect 3056 3052 3108 3058
rect 3056 2994 3108 3000
rect 2964 2984 3016 2990
rect 2964 2926 3016 2932
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 3988 2514 4016 5102
rect 4448 5030 4476 6122
rect 4724 5370 4752 6190
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4528 5160 4580 5166
rect 4528 5102 4580 5108
rect 4436 5024 4488 5030
rect 4436 4966 4488 4972
rect 4252 4548 4304 4554
rect 4252 4490 4304 4496
rect 4160 3936 4212 3942
rect 4160 3878 4212 3884
rect 4172 3670 4200 3878
rect 4160 3664 4212 3670
rect 4160 3606 4212 3612
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 4080 3194 4108 3538
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 4264 2650 4292 4490
rect 4448 3942 4476 4966
rect 4540 4690 4568 5102
rect 4528 4684 4580 4690
rect 4528 4626 4580 4632
rect 4436 3936 4488 3942
rect 4436 3878 4488 3884
rect 4252 2644 4304 2650
rect 4252 2586 4304 2592
rect 2504 2508 2556 2514
rect 2504 2450 2556 2456
rect 3976 2508 4028 2514
rect 3976 2450 4028 2456
rect 1308 2440 1360 2446
rect 1308 2382 1360 2388
rect 112 2372 164 2378
rect 112 2314 164 2320
rect 124 2281 152 2314
rect 110 2272 166 2281
rect 110 2207 166 2216
rect 1320 82 1348 2382
rect 2516 2310 2544 2450
rect 2504 2304 2556 2310
rect 2504 2246 2556 2252
rect 2516 1737 2544 2246
rect 2502 1728 2558 1737
rect 2502 1663 2558 1672
rect 1398 82 1454 480
rect 1320 54 1454 82
rect 1398 0 1454 54
rect 4250 82 4306 480
rect 4448 82 4476 3878
rect 4540 3738 4568 4626
rect 4528 3732 4580 3738
rect 4528 3674 4580 3680
rect 4816 2582 4844 11834
rect 5644 11801 5672 15558
rect 8588 15558 9090 15586
rect 7622 13084 7918 13104
rect 7678 13082 7702 13084
rect 7758 13082 7782 13084
rect 7838 13082 7862 13084
rect 7700 13030 7702 13082
rect 7764 13030 7776 13082
rect 7838 13030 7840 13082
rect 7678 13028 7702 13030
rect 7758 13028 7782 13030
rect 7838 13028 7862 13030
rect 7622 13008 7918 13028
rect 8208 12776 8260 12782
rect 8392 12776 8444 12782
rect 8260 12736 8392 12764
rect 8208 12718 8260 12724
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 6552 12300 6604 12306
rect 6552 12242 6604 12248
rect 6564 11830 6592 12242
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6552 11824 6604 11830
rect 5630 11792 5686 11801
rect 6552 11766 6604 11772
rect 5630 11727 5686 11736
rect 6276 11620 6328 11626
rect 6276 11562 6328 11568
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5080 10464 5132 10470
rect 5080 10406 5132 10412
rect 4988 9920 5040 9926
rect 4988 9862 5040 9868
rect 5000 4690 5028 9862
rect 5092 7410 5120 10406
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 5184 8090 5212 8978
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 5276 7818 5304 8230
rect 5460 7954 5488 11290
rect 6184 11212 6236 11218
rect 6184 11154 6236 11160
rect 6196 10606 6224 11154
rect 6288 10674 6316 11562
rect 6368 11076 6420 11082
rect 6368 11018 6420 11024
rect 6380 10810 6408 11018
rect 6564 10810 6592 11766
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 6932 10674 6960 12038
rect 7484 11694 7512 12582
rect 7622 11996 7918 12016
rect 7678 11994 7702 11996
rect 7758 11994 7782 11996
rect 7838 11994 7862 11996
rect 7700 11942 7702 11994
rect 7764 11942 7776 11994
rect 7838 11942 7840 11994
rect 7678 11940 7702 11942
rect 7758 11940 7782 11942
rect 7838 11940 7862 11942
rect 7622 11920 7918 11940
rect 7012 11688 7064 11694
rect 7012 11630 7064 11636
rect 7472 11688 7524 11694
rect 7472 11630 7524 11636
rect 7024 11082 7052 11630
rect 7104 11552 7156 11558
rect 7104 11494 7156 11500
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 6276 10668 6328 10674
rect 6276 10610 6328 10616
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 5632 10600 5684 10606
rect 5632 10542 5684 10548
rect 6184 10600 6236 10606
rect 6184 10542 6236 10548
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5552 9382 5580 10066
rect 5644 9926 5672 10542
rect 6092 10532 6144 10538
rect 6092 10474 6144 10480
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5264 7812 5316 7818
rect 5264 7754 5316 7760
rect 5460 7546 5488 7890
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 5276 6118 5304 6258
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 5078 5264 5134 5273
rect 5078 5199 5134 5208
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 5092 3602 5120 5199
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5184 4078 5212 4626
rect 5276 4146 5304 6054
rect 5446 5672 5502 5681
rect 5446 5607 5502 5616
rect 5460 5166 5488 5607
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5552 4214 5580 9318
rect 5736 9042 5764 10202
rect 5998 9752 6054 9761
rect 5998 9687 6000 9696
rect 6052 9687 6054 9696
rect 6000 9658 6052 9664
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5828 9110 5856 9318
rect 5816 9104 5868 9110
rect 5816 9046 5868 9052
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5828 8362 5856 9046
rect 6012 8430 6040 9658
rect 6104 9178 6132 10474
rect 6288 10130 6316 10610
rect 6932 10198 6960 10610
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 6920 10192 6972 10198
rect 6920 10134 6972 10140
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 6288 9722 6316 10066
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 6000 8424 6052 8430
rect 6000 8366 6052 8372
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 5828 8090 5856 8298
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 5828 7206 5856 8026
rect 5908 7948 5960 7954
rect 5908 7890 5960 7896
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5920 6934 5948 7890
rect 6288 7410 6316 9658
rect 6366 9480 6422 9489
rect 6366 9415 6422 9424
rect 6380 8430 6408 9415
rect 6840 9178 6868 9998
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6840 8634 6868 9114
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 5908 6928 5960 6934
rect 5908 6870 5960 6876
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5644 5914 5672 6598
rect 5920 6458 5948 6870
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 6012 5846 6040 6734
rect 6380 6458 6408 8366
rect 6932 8294 6960 8910
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6748 7002 6776 7346
rect 6932 7206 6960 8230
rect 7024 7970 7052 10406
rect 7116 10266 7144 11494
rect 7196 11280 7248 11286
rect 7196 11222 7248 11228
rect 7208 11014 7236 11222
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 7208 10538 7236 10950
rect 7622 10908 7918 10928
rect 7678 10906 7702 10908
rect 7758 10906 7782 10908
rect 7838 10906 7862 10908
rect 7700 10854 7702 10906
rect 7764 10854 7776 10906
rect 7838 10854 7840 10906
rect 7678 10852 7702 10854
rect 7758 10852 7782 10854
rect 7838 10852 7862 10854
rect 7622 10832 7918 10852
rect 7932 10668 7984 10674
rect 7932 10610 7984 10616
rect 7196 10532 7248 10538
rect 7196 10474 7248 10480
rect 7104 10260 7156 10266
rect 7104 10202 7156 10208
rect 7116 9586 7144 10202
rect 7944 10062 7972 10610
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 7622 9820 7918 9840
rect 7678 9818 7702 9820
rect 7758 9818 7782 9820
rect 7838 9818 7862 9820
rect 7700 9766 7702 9818
rect 7764 9766 7776 9818
rect 7838 9766 7840 9818
rect 7678 9764 7702 9766
rect 7758 9764 7782 9766
rect 7838 9764 7862 9766
rect 7622 9744 7918 9764
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 7288 9444 7340 9450
rect 7288 9386 7340 9392
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7116 9110 7144 9318
rect 7300 9178 7328 9386
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7104 9104 7156 9110
rect 7104 9046 7156 9052
rect 7622 8732 7918 8752
rect 7678 8730 7702 8732
rect 7758 8730 7782 8732
rect 7838 8730 7862 8732
rect 7700 8678 7702 8730
rect 7764 8678 7776 8730
rect 7838 8678 7840 8730
rect 7678 8676 7702 8678
rect 7758 8676 7782 8678
rect 7838 8676 7862 8678
rect 7622 8656 7918 8676
rect 7196 8560 7248 8566
rect 7248 8520 7328 8548
rect 7196 8502 7248 8508
rect 7102 7984 7158 7993
rect 7024 7942 7102 7970
rect 7102 7919 7158 7928
rect 7116 7342 7144 7919
rect 7104 7336 7156 7342
rect 7104 7278 7156 7284
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6736 6996 6788 7002
rect 6736 6938 6788 6944
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 6368 6452 6420 6458
rect 6368 6394 6420 6400
rect 7208 6254 7236 6598
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 6000 5840 6052 5846
rect 6000 5782 6052 5788
rect 6644 5840 6696 5846
rect 6644 5782 6696 5788
rect 6184 5568 6236 5574
rect 6184 5510 6236 5516
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5644 4622 5672 4966
rect 5736 4758 5764 4966
rect 5724 4752 5776 4758
rect 5724 4694 5776 4700
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5644 4282 5672 4558
rect 5632 4276 5684 4282
rect 5632 4218 5684 4224
rect 5540 4208 5592 4214
rect 5540 4150 5592 4156
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 5172 4072 5224 4078
rect 5172 4014 5224 4020
rect 5184 3738 5212 4014
rect 5736 3942 5764 4694
rect 6012 4486 6040 5102
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 5906 4176 5962 4185
rect 5906 4111 5962 4120
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5080 3596 5132 3602
rect 5080 3538 5132 3544
rect 5920 3058 5948 4111
rect 6012 3670 6040 4422
rect 6092 4140 6144 4146
rect 6092 4082 6144 4088
rect 6000 3664 6052 3670
rect 6000 3606 6052 3612
rect 6104 3194 6132 4082
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 6196 2650 6224 5510
rect 6656 5370 6684 5782
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 7116 5030 7144 6054
rect 7104 5024 7156 5030
rect 7104 4966 7156 4972
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 7024 4010 7052 4422
rect 7012 4004 7064 4010
rect 7012 3946 7064 3952
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 6564 3738 6592 3878
rect 7208 3738 7236 6190
rect 6552 3732 6604 3738
rect 6552 3674 6604 3680
rect 7196 3732 7248 3738
rect 7196 3674 7248 3680
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 7208 2990 7236 3538
rect 7196 2984 7248 2990
rect 7196 2926 7248 2932
rect 7104 2848 7156 2854
rect 7104 2790 7156 2796
rect 6184 2644 6236 2650
rect 6184 2586 6236 2592
rect 4804 2576 4856 2582
rect 4804 2518 4856 2524
rect 7116 2514 7144 2790
rect 7300 2514 7328 8520
rect 7622 7644 7918 7664
rect 7678 7642 7702 7644
rect 7758 7642 7782 7644
rect 7838 7642 7862 7644
rect 7700 7590 7702 7642
rect 7764 7590 7776 7642
rect 7838 7590 7840 7642
rect 7678 7588 7702 7590
rect 7758 7588 7782 7590
rect 7838 7588 7862 7590
rect 7622 7568 7918 7588
rect 8036 7002 8064 12582
rect 8116 12300 8168 12306
rect 8116 12242 8168 12248
rect 8128 11558 8156 12242
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 8128 9081 8156 11494
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 8220 9722 8248 10134
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 8220 9450 8248 9658
rect 8208 9444 8260 9450
rect 8208 9386 8260 9392
rect 8220 9178 8248 9386
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 8114 9072 8170 9081
rect 8114 9007 8116 9016
rect 8168 9007 8170 9016
rect 8116 8978 8168 8984
rect 8128 8947 8156 8978
rect 8312 8922 8340 12736
rect 8392 12718 8444 12724
rect 8588 11354 8616 15558
rect 9034 15520 9090 15558
rect 12544 15558 12678 15586
rect 9588 12300 9640 12306
rect 9588 12242 9640 12248
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 8852 12096 8904 12102
rect 8852 12038 8904 12044
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8680 11150 8708 11494
rect 8864 11354 8892 12038
rect 8944 11552 8996 11558
rect 8944 11494 8996 11500
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8404 9654 8432 10406
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 8496 9382 8524 11018
rect 8680 10266 8708 11086
rect 8864 10674 8892 11290
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8852 9580 8904 9586
rect 8852 9522 8904 9528
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8864 9178 8892 9522
rect 8852 9172 8904 9178
rect 8852 9114 8904 9120
rect 8220 8894 8340 8922
rect 8760 8900 8812 8906
rect 8220 8634 8248 8894
rect 8760 8842 8812 8848
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 8312 8498 8340 8774
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 8668 8356 8720 8362
rect 8668 8298 8720 8304
rect 8116 8016 8168 8022
rect 8116 7958 8168 7964
rect 8128 7546 8156 7958
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8024 6996 8076 7002
rect 8024 6938 8076 6944
rect 7622 6556 7918 6576
rect 7678 6554 7702 6556
rect 7758 6554 7782 6556
rect 7838 6554 7862 6556
rect 7700 6502 7702 6554
rect 7764 6502 7776 6554
rect 7838 6502 7840 6554
rect 7678 6500 7702 6502
rect 7758 6500 7782 6502
rect 7838 6500 7862 6502
rect 7622 6480 7918 6500
rect 8036 6458 8064 6938
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 8128 5846 8156 6734
rect 8220 6730 8248 7822
rect 8680 7546 8708 8298
rect 8772 7954 8800 8842
rect 8760 7948 8812 7954
rect 8760 7890 8812 7896
rect 8956 7886 8984 11494
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8680 7274 8708 7482
rect 8668 7268 8720 7274
rect 8668 7210 8720 7216
rect 8392 6928 8444 6934
rect 8392 6870 8444 6876
rect 8208 6724 8260 6730
rect 8208 6666 8260 6672
rect 8404 6118 8432 6870
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8404 5846 8432 6054
rect 8116 5840 8168 5846
rect 8116 5782 8168 5788
rect 8392 5840 8444 5846
rect 8392 5782 8444 5788
rect 8574 5808 8630 5817
rect 8024 5568 8076 5574
rect 8024 5510 8076 5516
rect 7622 5468 7918 5488
rect 7678 5466 7702 5468
rect 7758 5466 7782 5468
rect 7838 5466 7862 5468
rect 7700 5414 7702 5466
rect 7764 5414 7776 5466
rect 7838 5414 7840 5466
rect 7678 5412 7702 5414
rect 7758 5412 7782 5414
rect 7838 5412 7862 5414
rect 7622 5392 7918 5412
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7484 4486 7512 5170
rect 8036 4826 8064 5510
rect 8404 5370 8432 5782
rect 8574 5743 8630 5752
rect 8392 5364 8444 5370
rect 8392 5306 8444 5312
rect 8024 4820 8076 4826
rect 8024 4762 8076 4768
rect 8588 4690 8616 5743
rect 9048 5574 9076 12038
rect 9600 11762 9628 12242
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 9312 11688 9364 11694
rect 9312 11630 9364 11636
rect 9140 10577 9168 11630
rect 9126 10568 9182 10577
rect 9126 10503 9182 10512
rect 9324 9217 9352 11630
rect 9876 11218 9904 11698
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 9588 11212 9640 11218
rect 9588 11154 9640 11160
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 9600 10810 9628 11154
rect 10232 11076 10284 11082
rect 10232 11018 10284 11024
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 9310 9208 9366 9217
rect 9310 9143 9366 9152
rect 9692 8090 9720 10950
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9784 10198 9812 10406
rect 9772 10192 9824 10198
rect 9772 10134 9824 10140
rect 9864 10192 9916 10198
rect 9864 10134 9916 10140
rect 9784 9722 9812 10134
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9876 9654 9904 10134
rect 10048 10056 10100 10062
rect 10048 9998 10100 10004
rect 9864 9648 9916 9654
rect 9864 9590 9916 9596
rect 10060 9450 10088 9998
rect 10244 9722 10272 11018
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 10048 9444 10100 9450
rect 10048 9386 10100 9392
rect 9864 9104 9916 9110
rect 9864 9046 9916 9052
rect 9876 8634 9904 9046
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9876 8294 9904 8570
rect 10048 8356 10100 8362
rect 10048 8298 10100 8304
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 9140 7002 9168 7346
rect 9312 7268 9364 7274
rect 9312 7210 9364 7216
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 9324 6186 9352 7210
rect 9692 7002 9720 8026
rect 9864 8016 9916 8022
rect 9864 7958 9916 7964
rect 9876 7886 9904 7958
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9876 7206 9904 7822
rect 10060 7750 10088 8298
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9876 7002 9904 7142
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9312 6180 9364 6186
rect 9312 6122 9364 6128
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 9036 5568 9088 5574
rect 9036 5510 9088 5516
rect 9128 5296 9180 5302
rect 9128 5238 9180 5244
rect 9140 5098 9168 5238
rect 9036 5092 9088 5098
rect 9036 5034 9088 5040
rect 9128 5092 9180 5098
rect 9128 5034 9180 5040
rect 8392 4684 8444 4690
rect 8576 4684 8628 4690
rect 8444 4644 8524 4672
rect 8392 4626 8444 4632
rect 8024 4548 8076 4554
rect 8024 4490 8076 4496
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 7380 3460 7432 3466
rect 7380 3402 7432 3408
rect 7392 2990 7420 3402
rect 7484 3058 7512 4422
rect 7622 4380 7918 4400
rect 7678 4378 7702 4380
rect 7758 4378 7782 4380
rect 7838 4378 7862 4380
rect 7700 4326 7702 4378
rect 7764 4326 7776 4378
rect 7838 4326 7840 4378
rect 7678 4324 7702 4326
rect 7758 4324 7782 4326
rect 7838 4324 7862 4326
rect 7622 4304 7918 4324
rect 8036 4146 8064 4490
rect 8116 4276 8168 4282
rect 8116 4218 8168 4224
rect 8024 4140 8076 4146
rect 8024 4082 8076 4088
rect 8128 3738 8156 4218
rect 8496 4078 8524 4644
rect 8576 4626 8628 4632
rect 8588 4282 8616 4626
rect 9048 4622 9076 5034
rect 9232 4758 9260 6054
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9324 5234 9352 5646
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 9324 4826 9352 5170
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 9220 4752 9272 4758
rect 9126 4720 9182 4729
rect 9220 4694 9272 4700
rect 9126 4655 9182 4664
rect 9036 4616 9088 4622
rect 9036 4558 9088 4564
rect 8576 4276 8628 4282
rect 8576 4218 8628 4224
rect 8484 4072 8536 4078
rect 8482 4040 8484 4049
rect 8536 4040 8538 4049
rect 8404 3998 8482 4026
rect 8116 3732 8168 3738
rect 8116 3674 8168 3680
rect 8404 3670 8432 3998
rect 8482 3975 8538 3984
rect 8496 3949 8524 3975
rect 8668 3936 8720 3942
rect 8668 3878 8720 3884
rect 8392 3664 8444 3670
rect 8392 3606 8444 3612
rect 8116 3596 8168 3602
rect 8116 3538 8168 3544
rect 7622 3292 7918 3312
rect 7678 3290 7702 3292
rect 7758 3290 7782 3292
rect 7838 3290 7862 3292
rect 7700 3238 7702 3290
rect 7764 3238 7776 3290
rect 7838 3238 7840 3290
rect 7678 3236 7702 3238
rect 7758 3236 7782 3238
rect 7838 3236 7862 3238
rect 7622 3216 7918 3236
rect 8128 3194 8156 3538
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 7380 2984 7432 2990
rect 7380 2926 7432 2932
rect 8128 2582 8156 3130
rect 8576 2984 8628 2990
rect 8496 2944 8576 2972
rect 8496 2854 8524 2944
rect 8576 2926 8628 2932
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 8116 2576 8168 2582
rect 8116 2518 8168 2524
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 6644 2508 6696 2514
rect 6644 2450 6696 2456
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 7380 2508 7432 2514
rect 7380 2450 7432 2456
rect 6012 2106 6040 2450
rect 6656 2310 6684 2450
rect 6276 2304 6328 2310
rect 6276 2246 6328 2252
rect 6644 2304 6696 2310
rect 6644 2246 6696 2252
rect 6000 2100 6052 2106
rect 6000 2042 6052 2048
rect 6288 2038 6316 2246
rect 6276 2032 6328 2038
rect 6276 1974 6328 1980
rect 6288 1601 6316 1974
rect 6274 1592 6330 1601
rect 6274 1527 6330 1536
rect 6656 1057 6684 2246
rect 7392 2038 7420 2450
rect 7622 2204 7918 2224
rect 7678 2202 7702 2204
rect 7758 2202 7782 2204
rect 7838 2202 7862 2204
rect 7700 2150 7702 2202
rect 7764 2150 7776 2202
rect 7838 2150 7840 2202
rect 7678 2148 7702 2150
rect 7758 2148 7782 2150
rect 7838 2148 7862 2150
rect 7622 2128 7918 2148
rect 7380 2032 7432 2038
rect 7380 1974 7432 1980
rect 8496 1601 8524 2790
rect 8680 2038 8708 3878
rect 9140 3058 9168 4655
rect 9968 4593 9996 7142
rect 10060 6322 10088 7686
rect 10336 7002 10364 11494
rect 10416 8560 10468 8566
rect 10416 8502 10468 8508
rect 10428 8022 10456 8502
rect 10416 8016 10468 8022
rect 10416 7958 10468 7964
rect 10324 6996 10376 7002
rect 10324 6938 10376 6944
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 10232 6180 10284 6186
rect 10232 6122 10284 6128
rect 10140 5840 10192 5846
rect 10140 5782 10192 5788
rect 10152 5370 10180 5782
rect 10140 5364 10192 5370
rect 10140 5306 10192 5312
rect 10244 5098 10272 6122
rect 10336 5914 10364 6938
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 10520 5710 10548 12038
rect 10796 11558 10824 12242
rect 11796 11688 11848 11694
rect 12544 11665 12572 15558
rect 12622 15520 12678 15558
rect 16302 15586 16358 16000
rect 19890 15586 19946 16000
rect 16302 15558 16620 15586
rect 16302 15520 16358 15558
rect 14289 13628 14585 13648
rect 14345 13626 14369 13628
rect 14425 13626 14449 13628
rect 14505 13626 14529 13628
rect 14367 13574 14369 13626
rect 14431 13574 14443 13626
rect 14505 13574 14507 13626
rect 14345 13572 14369 13574
rect 14425 13572 14449 13574
rect 14505 13572 14529 13574
rect 14289 13552 14585 13572
rect 12900 12708 12952 12714
rect 12900 12650 12952 12656
rect 11796 11630 11848 11636
rect 12530 11656 12586 11665
rect 11808 11558 11836 11630
rect 12530 11591 12586 11600
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 10796 10470 10824 11494
rect 10968 11212 11020 11218
rect 10968 11154 11020 11160
rect 10980 10810 11008 11154
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 10980 10606 11008 10746
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10704 7206 10732 8434
rect 10796 7449 10824 10406
rect 10980 10266 11008 10542
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10888 7857 10916 9318
rect 11072 8974 11100 10406
rect 11808 9625 11836 11494
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11900 10742 11928 10950
rect 11888 10736 11940 10742
rect 11886 10704 11888 10713
rect 11940 10704 11942 10713
rect 11886 10639 11942 10648
rect 11900 10606 11928 10639
rect 12268 10606 12296 11086
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 11888 10600 11940 10606
rect 11888 10542 11940 10548
rect 12256 10600 12308 10606
rect 12256 10542 12308 10548
rect 12268 9994 12296 10542
rect 12452 10266 12480 10950
rect 12636 10606 12664 10950
rect 12624 10600 12676 10606
rect 12544 10560 12624 10588
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 12256 9988 12308 9994
rect 12256 9930 12308 9936
rect 11794 9616 11850 9625
rect 11794 9551 11850 9560
rect 11808 9518 11836 9551
rect 11796 9512 11848 9518
rect 11796 9454 11848 9460
rect 11704 9376 11756 9382
rect 11704 9318 11756 9324
rect 11716 9110 11744 9318
rect 11704 9104 11756 9110
rect 11704 9046 11756 9052
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11072 8634 11100 8910
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 11164 8566 11192 8910
rect 11716 8634 11744 9046
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11152 8560 11204 8566
rect 11152 8502 11204 8508
rect 12268 8401 12296 9930
rect 12360 9722 12388 10066
rect 12348 9716 12400 9722
rect 12348 9658 12400 9664
rect 12360 9489 12388 9658
rect 12452 9654 12480 10202
rect 12544 10130 12572 10560
rect 12624 10542 12676 10548
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12346 9480 12402 9489
rect 12346 9415 12402 9424
rect 12544 9382 12572 10066
rect 12716 9648 12768 9654
rect 12716 9590 12768 9596
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12624 8424 12676 8430
rect 12254 8392 12310 8401
rect 12624 8366 12676 8372
rect 12254 8327 12310 8336
rect 11336 8084 11388 8090
rect 11336 8026 11388 8032
rect 10874 7848 10930 7857
rect 10874 7783 10930 7792
rect 10782 7440 10838 7449
rect 11348 7410 11376 8026
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11716 7546 11744 7890
rect 12072 7880 12124 7886
rect 12072 7822 12124 7828
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 10782 7375 10838 7384
rect 11336 7404 11388 7410
rect 11336 7346 11388 7352
rect 11716 7342 11744 7482
rect 11704 7336 11756 7342
rect 11704 7278 11756 7284
rect 10692 7200 10744 7206
rect 10692 7142 10744 7148
rect 10692 6928 10744 6934
rect 10692 6870 10744 6876
rect 10704 6118 10732 6870
rect 11716 6458 11744 7278
rect 12084 7206 12112 7822
rect 12636 7750 12664 8366
rect 12728 7954 12756 9590
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12820 8906 12848 9522
rect 12808 8900 12860 8906
rect 12808 8842 12860 8848
rect 12716 7948 12768 7954
rect 12716 7890 12768 7896
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10704 5846 10732 6054
rect 11808 5914 11836 6734
rect 11992 6118 12020 6802
rect 11980 6112 12032 6118
rect 11980 6054 12032 6060
rect 11796 5908 11848 5914
rect 11796 5850 11848 5856
rect 10692 5840 10744 5846
rect 10692 5782 10744 5788
rect 11808 5710 11836 5850
rect 11992 5817 12020 6054
rect 11978 5808 12034 5817
rect 11978 5743 12034 5752
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11888 5568 11940 5574
rect 11888 5510 11940 5516
rect 10232 5092 10284 5098
rect 10232 5034 10284 5040
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 10232 4820 10284 4826
rect 10232 4762 10284 4768
rect 10244 4729 10272 4762
rect 11532 4758 11560 4966
rect 11520 4752 11572 4758
rect 10230 4720 10286 4729
rect 10048 4684 10100 4690
rect 11520 4694 11572 4700
rect 10230 4655 10286 4664
rect 10048 4626 10100 4632
rect 9954 4584 10010 4593
rect 9954 4519 10010 4528
rect 9864 4004 9916 4010
rect 9864 3946 9916 3952
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9312 3120 9364 3126
rect 9312 3062 9364 3068
rect 9128 3052 9180 3058
rect 9128 2994 9180 3000
rect 8760 2848 8812 2854
rect 8760 2790 8812 2796
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 8772 2446 8800 2790
rect 9048 2582 9076 2790
rect 9036 2576 9088 2582
rect 9036 2518 9088 2524
rect 9220 2508 9272 2514
rect 9220 2450 9272 2456
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 9232 2310 9260 2450
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 8668 2032 8720 2038
rect 9048 2009 9076 2246
rect 8668 1974 8720 1980
rect 9034 2000 9090 2009
rect 9034 1935 9090 1944
rect 8482 1592 8538 1601
rect 8482 1527 8538 1536
rect 6642 1048 6698 1057
rect 6642 983 6698 992
rect 4250 54 4476 82
rect 7102 128 7158 480
rect 8496 134 8524 1527
rect 9232 1329 9260 2246
rect 9324 1737 9352 3062
rect 9784 3058 9812 3538
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 9876 2990 9904 3946
rect 9968 3738 9996 4519
rect 10060 3942 10088 4626
rect 10784 4480 10836 4486
rect 10784 4422 10836 4428
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 10140 4072 10192 4078
rect 10140 4014 10192 4020
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 10060 3534 10088 3878
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 10152 3058 10180 4014
rect 10244 3942 10272 4082
rect 10796 4078 10824 4422
rect 11796 4208 11848 4214
rect 11796 4150 11848 4156
rect 10508 4072 10560 4078
rect 10508 4014 10560 4020
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 10244 3126 10272 3878
rect 10520 3670 10548 4014
rect 11808 4010 11836 4150
rect 11244 4004 11296 4010
rect 11244 3946 11296 3952
rect 11796 4004 11848 4010
rect 11796 3946 11848 3952
rect 10876 3936 10928 3942
rect 10876 3878 10928 3884
rect 10508 3664 10560 3670
rect 10508 3606 10560 3612
rect 10888 3602 10916 3878
rect 11256 3738 11284 3946
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 10876 3596 10928 3602
rect 10876 3538 10928 3544
rect 10324 3392 10376 3398
rect 10324 3334 10376 3340
rect 10232 3120 10284 3126
rect 10232 3062 10284 3068
rect 10140 3052 10192 3058
rect 10140 2994 10192 3000
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 9772 2916 9824 2922
rect 9772 2858 9824 2864
rect 9310 1728 9366 1737
rect 9310 1663 9366 1672
rect 9218 1320 9274 1329
rect 9218 1255 9274 1264
rect 7102 76 7104 128
rect 7156 76 7158 128
rect 4250 0 4306 54
rect 7102 0 7158 76
rect 8484 128 8536 134
rect 8484 70 8536 76
rect 9784 82 9812 2858
rect 9876 2650 9904 2926
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 10244 2310 10272 3062
rect 10140 2304 10192 2310
rect 10140 2246 10192 2252
rect 10232 2304 10284 2310
rect 10232 2246 10284 2252
rect 10152 2038 10180 2246
rect 10140 2032 10192 2038
rect 10140 1974 10192 1980
rect 9954 82 10010 480
rect 10336 134 10364 3334
rect 10888 3194 10916 3538
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 11256 2990 11284 3674
rect 11244 2984 11296 2990
rect 11244 2926 11296 2932
rect 11808 2582 11836 3946
rect 11900 3194 11928 5510
rect 12084 4729 12112 7142
rect 12636 6934 12664 7686
rect 12624 6928 12676 6934
rect 12624 6870 12676 6876
rect 12728 6866 12756 7890
rect 12716 6860 12768 6866
rect 12716 6802 12768 6808
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12820 6254 12848 6598
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 12164 5840 12216 5846
rect 12164 5782 12216 5788
rect 12176 5302 12204 5782
rect 12348 5704 12400 5710
rect 12348 5646 12400 5652
rect 12164 5296 12216 5302
rect 12164 5238 12216 5244
rect 12070 4720 12126 4729
rect 12070 4655 12126 4664
rect 12360 4622 12388 5646
rect 12544 5370 12572 6054
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 12348 4616 12400 4622
rect 12348 4558 12400 4564
rect 12716 4480 12768 4486
rect 12716 4422 12768 4428
rect 12728 4078 12756 4422
rect 12716 4072 12768 4078
rect 12716 4014 12768 4020
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 12268 3398 12296 3538
rect 12440 3460 12492 3466
rect 12440 3402 12492 3408
rect 12256 3392 12308 3398
rect 12256 3334 12308 3340
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 12268 2990 12296 3334
rect 12256 2984 12308 2990
rect 12256 2926 12308 2932
rect 11796 2576 11848 2582
rect 11796 2518 11848 2524
rect 12452 2514 12480 3402
rect 12636 3398 12664 3878
rect 12728 3602 12756 4014
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 12532 2984 12584 2990
rect 12532 2926 12584 2932
rect 12544 2582 12572 2926
rect 12532 2576 12584 2582
rect 12532 2518 12584 2524
rect 12636 2514 12664 3334
rect 12728 3126 12756 3538
rect 12716 3120 12768 3126
rect 12716 3062 12768 3068
rect 12808 2984 12860 2990
rect 12728 2944 12808 2972
rect 12728 2650 12756 2944
rect 12808 2926 12860 2932
rect 12716 2644 12768 2650
rect 12716 2586 12768 2592
rect 12912 2582 12940 12650
rect 14289 12540 14585 12560
rect 14345 12538 14369 12540
rect 14425 12538 14449 12540
rect 14505 12538 14529 12540
rect 14367 12486 14369 12538
rect 14431 12486 14443 12538
rect 14505 12486 14507 12538
rect 14345 12484 14369 12486
rect 14425 12484 14449 12486
rect 14505 12484 14529 12486
rect 14289 12464 14585 12484
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 15672 11762 15700 12242
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 14188 11552 14240 11558
rect 14188 11494 14240 11500
rect 14832 11552 14884 11558
rect 14832 11494 14884 11500
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 13544 11008 13596 11014
rect 13544 10950 13596 10956
rect 13268 10532 13320 10538
rect 13268 10474 13320 10480
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 12992 9444 13044 9450
rect 12992 9386 13044 9392
rect 13004 9110 13032 9386
rect 12992 9104 13044 9110
rect 12992 9046 13044 9052
rect 13004 8838 13032 9046
rect 12992 8832 13044 8838
rect 12992 8774 13044 8780
rect 13004 8634 13032 8774
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 12992 6248 13044 6254
rect 13096 6236 13124 9862
rect 13280 6866 13308 10474
rect 13360 10056 13412 10062
rect 13360 9998 13412 10004
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13372 7342 13400 9998
rect 13464 9625 13492 9998
rect 13450 9616 13506 9625
rect 13450 9551 13506 9560
rect 13360 7336 13412 7342
rect 13360 7278 13412 7284
rect 13268 6860 13320 6866
rect 13268 6802 13320 6808
rect 13280 6458 13308 6802
rect 13268 6452 13320 6458
rect 13268 6394 13320 6400
rect 13044 6208 13124 6236
rect 12992 6190 13044 6196
rect 13004 5574 13032 6190
rect 13084 6112 13136 6118
rect 13084 6054 13136 6060
rect 13176 6112 13228 6118
rect 13176 6054 13228 6060
rect 12992 5568 13044 5574
rect 12992 5510 13044 5516
rect 13096 4690 13124 6054
rect 13188 5030 13216 6054
rect 13360 5568 13412 5574
rect 13360 5510 13412 5516
rect 13372 5234 13400 5510
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13176 5024 13228 5030
rect 13176 4966 13228 4972
rect 13084 4684 13136 4690
rect 13084 4626 13136 4632
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 13004 2650 13032 4558
rect 13096 4214 13124 4626
rect 13372 4622 13400 5170
rect 13464 4690 13492 9551
rect 13556 7886 13584 10950
rect 13924 10742 13952 11154
rect 13912 10736 13964 10742
rect 13912 10678 13964 10684
rect 13636 10668 13688 10674
rect 13636 10610 13688 10616
rect 13648 8498 13676 10610
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13740 9042 13768 10202
rect 13832 10130 13860 10406
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 13740 8090 13768 8978
rect 13832 8276 13860 9114
rect 13924 8945 13952 10678
rect 14096 10600 14148 10606
rect 14016 10560 14096 10588
rect 14016 9926 14044 10560
rect 14096 10542 14148 10548
rect 14096 10124 14148 10130
rect 14096 10066 14148 10072
rect 14004 9920 14056 9926
rect 14004 9862 14056 9868
rect 14108 9654 14136 10066
rect 14096 9648 14148 9654
rect 14096 9590 14148 9596
rect 13910 8936 13966 8945
rect 13910 8871 13966 8880
rect 13912 8288 13964 8294
rect 13832 8248 13912 8276
rect 13912 8230 13964 8236
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13820 8016 13872 8022
rect 13820 7958 13872 7964
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13556 7002 13584 7822
rect 13832 7410 13860 7958
rect 13924 7478 13952 8230
rect 13912 7472 13964 7478
rect 13912 7414 13964 7420
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13774 7268 13826 7274
rect 13924 7256 13952 7414
rect 13826 7228 13952 7256
rect 13774 7210 13826 7216
rect 13544 6996 13596 7002
rect 13544 6938 13596 6944
rect 13924 6934 13952 7228
rect 14200 6934 14228 11494
rect 14289 11452 14585 11472
rect 14345 11450 14369 11452
rect 14425 11450 14449 11452
rect 14505 11450 14529 11452
rect 14367 11398 14369 11450
rect 14431 11398 14443 11450
rect 14505 11398 14507 11450
rect 14345 11396 14369 11398
rect 14425 11396 14449 11398
rect 14505 11396 14529 11398
rect 14289 11376 14585 11396
rect 14648 11280 14700 11286
rect 14648 11222 14700 11228
rect 14660 10606 14688 11222
rect 14648 10600 14700 10606
rect 14648 10542 14700 10548
rect 14289 10364 14585 10384
rect 14345 10362 14369 10364
rect 14425 10362 14449 10364
rect 14505 10362 14529 10364
rect 14367 10310 14369 10362
rect 14431 10310 14443 10362
rect 14505 10310 14507 10362
rect 14345 10308 14369 10310
rect 14425 10308 14449 10310
rect 14505 10308 14529 10310
rect 14289 10288 14585 10308
rect 14660 10130 14688 10542
rect 14738 10160 14794 10169
rect 14648 10124 14700 10130
rect 14738 10095 14794 10104
rect 14648 10066 14700 10072
rect 14752 10062 14780 10095
rect 14844 10062 14872 11494
rect 15844 11212 15896 11218
rect 15844 11154 15896 11160
rect 16488 11212 16540 11218
rect 16488 11154 16540 11160
rect 15856 10470 15884 11154
rect 16396 11076 16448 11082
rect 16396 11018 16448 11024
rect 16028 11008 16080 11014
rect 16028 10950 16080 10956
rect 16040 10742 16068 10950
rect 16028 10736 16080 10742
rect 16028 10678 16080 10684
rect 16304 10736 16356 10742
rect 16304 10678 16356 10684
rect 16028 10532 16080 10538
rect 16028 10474 16080 10480
rect 14924 10464 14976 10470
rect 14924 10406 14976 10412
rect 15844 10464 15896 10470
rect 15844 10406 15896 10412
rect 14740 10056 14792 10062
rect 14740 9998 14792 10004
rect 14832 10056 14884 10062
rect 14832 9998 14884 10004
rect 14740 9648 14792 9654
rect 14740 9590 14792 9596
rect 14648 9512 14700 9518
rect 14648 9454 14700 9460
rect 14289 9276 14585 9296
rect 14345 9274 14369 9276
rect 14425 9274 14449 9276
rect 14505 9274 14529 9276
rect 14367 9222 14369 9274
rect 14431 9222 14443 9274
rect 14505 9222 14507 9274
rect 14345 9220 14369 9222
rect 14425 9220 14449 9222
rect 14505 9220 14529 9222
rect 14289 9200 14585 9220
rect 14660 9110 14688 9454
rect 14648 9104 14700 9110
rect 14648 9046 14700 9052
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14289 8188 14585 8208
rect 14345 8186 14369 8188
rect 14425 8186 14449 8188
rect 14505 8186 14529 8188
rect 14367 8134 14369 8186
rect 14431 8134 14443 8186
rect 14505 8134 14507 8186
rect 14345 8132 14369 8134
rect 14425 8132 14449 8134
rect 14505 8132 14529 8134
rect 14289 8112 14585 8132
rect 14660 8090 14688 8434
rect 14752 8294 14780 9590
rect 14844 9178 14872 9998
rect 14832 9172 14884 9178
rect 14832 9114 14884 9120
rect 14740 8288 14792 8294
rect 14740 8230 14792 8236
rect 14648 8084 14700 8090
rect 14648 8026 14700 8032
rect 14648 7880 14700 7886
rect 14648 7822 14700 7828
rect 14289 7100 14585 7120
rect 14345 7098 14369 7100
rect 14425 7098 14449 7100
rect 14505 7098 14529 7100
rect 14367 7046 14369 7098
rect 14431 7046 14443 7098
rect 14505 7046 14507 7098
rect 14345 7044 14369 7046
rect 14425 7044 14449 7046
rect 14505 7044 14529 7046
rect 14289 7024 14585 7044
rect 14660 7002 14688 7822
rect 14648 6996 14700 7002
rect 14648 6938 14700 6944
rect 13912 6928 13964 6934
rect 13912 6870 13964 6876
rect 14188 6928 14240 6934
rect 14188 6870 14240 6876
rect 14936 6798 14964 10406
rect 15198 10296 15254 10305
rect 15198 10231 15254 10240
rect 15016 9648 15068 9654
rect 15016 9590 15068 9596
rect 15028 9450 15056 9590
rect 15016 9444 15068 9450
rect 15016 9386 15068 9392
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 15016 8900 15068 8906
rect 15016 8842 15068 8848
rect 15028 8022 15056 8842
rect 15120 8090 15148 8910
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15016 8016 15068 8022
rect 15016 7958 15068 7964
rect 15028 7546 15056 7958
rect 15016 7540 15068 7546
rect 15016 7482 15068 7488
rect 15016 6928 15068 6934
rect 15016 6870 15068 6876
rect 14188 6792 14240 6798
rect 14188 6734 14240 6740
rect 14924 6792 14976 6798
rect 14924 6734 14976 6740
rect 13912 5772 13964 5778
rect 13912 5714 13964 5720
rect 14096 5772 14148 5778
rect 14096 5714 14148 5720
rect 13924 5681 13952 5714
rect 13910 5672 13966 5681
rect 13910 5607 13966 5616
rect 13924 5001 13952 5607
rect 14108 5370 14136 5714
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 13910 4992 13966 5001
rect 13910 4927 13966 4936
rect 13924 4826 13952 4927
rect 13912 4820 13964 4826
rect 13912 4762 13964 4768
rect 13452 4684 13504 4690
rect 13452 4626 13504 4632
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13084 4208 13136 4214
rect 13084 4150 13136 4156
rect 13096 4049 13124 4150
rect 14200 4146 14228 6734
rect 14648 6248 14700 6254
rect 14648 6190 14700 6196
rect 14289 6012 14585 6032
rect 14345 6010 14369 6012
rect 14425 6010 14449 6012
rect 14505 6010 14529 6012
rect 14367 5958 14369 6010
rect 14431 5958 14443 6010
rect 14505 5958 14507 6010
rect 14345 5956 14369 5958
rect 14425 5956 14449 5958
rect 14505 5956 14529 5958
rect 14289 5936 14585 5956
rect 14660 5710 14688 6190
rect 15028 5914 15056 6870
rect 15016 5908 15068 5914
rect 15016 5850 15068 5856
rect 14648 5704 14700 5710
rect 14648 5646 14700 5652
rect 14646 5536 14702 5545
rect 14646 5471 14702 5480
rect 14660 5098 14688 5471
rect 15212 5098 15240 10231
rect 15384 10192 15436 10198
rect 15384 10134 15436 10140
rect 15396 9722 15424 10134
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 15396 7886 15424 9522
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15476 9104 15528 9110
rect 15476 9046 15528 9052
rect 15488 8634 15516 9046
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 15290 7440 15346 7449
rect 15396 7410 15424 7822
rect 15290 7375 15346 7384
rect 15384 7404 15436 7410
rect 15304 6338 15332 7375
rect 15384 7346 15436 7352
rect 15304 6310 15424 6338
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 15304 5234 15332 5510
rect 15292 5228 15344 5234
rect 15292 5170 15344 5176
rect 14648 5092 14700 5098
rect 14648 5034 14700 5040
rect 15200 5092 15252 5098
rect 15200 5034 15252 5040
rect 14289 4924 14585 4944
rect 14345 4922 14369 4924
rect 14425 4922 14449 4924
rect 14505 4922 14529 4924
rect 14367 4870 14369 4922
rect 14431 4870 14443 4922
rect 14505 4870 14507 4922
rect 14345 4868 14369 4870
rect 14425 4868 14449 4870
rect 14505 4868 14529 4870
rect 14289 4848 14585 4868
rect 14660 4826 14688 5034
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 15016 4684 15068 4690
rect 15016 4626 15068 4632
rect 15028 4486 15056 4626
rect 15292 4616 15344 4622
rect 15292 4558 15344 4564
rect 15016 4480 15068 4486
rect 15016 4422 15068 4428
rect 14832 4276 14884 4282
rect 14832 4218 14884 4224
rect 14188 4140 14240 4146
rect 14188 4082 14240 4088
rect 13082 4040 13138 4049
rect 13082 3975 13138 3984
rect 13912 3596 13964 3602
rect 13912 3538 13964 3544
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 12992 2644 13044 2650
rect 12992 2586 13044 2592
rect 12900 2576 12952 2582
rect 12900 2518 12952 2524
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 13648 2310 13676 3334
rect 13924 3058 13952 3538
rect 14096 3460 14148 3466
rect 14096 3402 14148 3408
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 14108 2310 14136 3402
rect 14200 2446 14228 4082
rect 14844 4078 14872 4218
rect 15028 4185 15056 4422
rect 15014 4176 15070 4185
rect 15014 4111 15070 4120
rect 14832 4072 14884 4078
rect 14832 4014 14884 4020
rect 14924 4072 14976 4078
rect 14924 4014 14976 4020
rect 14936 3942 14964 4014
rect 14924 3936 14976 3942
rect 14924 3878 14976 3884
rect 14289 3836 14585 3856
rect 14345 3834 14369 3836
rect 14425 3834 14449 3836
rect 14505 3834 14529 3836
rect 14367 3782 14369 3834
rect 14431 3782 14443 3834
rect 14505 3782 14507 3834
rect 14345 3780 14369 3782
rect 14425 3780 14449 3782
rect 14505 3780 14529 3782
rect 14289 3760 14585 3780
rect 14936 3126 14964 3878
rect 15304 3670 15332 4558
rect 15292 3664 15344 3670
rect 15292 3606 15344 3612
rect 15200 3596 15252 3602
rect 15200 3538 15252 3544
rect 15212 3398 15240 3538
rect 15200 3392 15252 3398
rect 15200 3334 15252 3340
rect 14924 3120 14976 3126
rect 14924 3062 14976 3068
rect 15108 2848 15160 2854
rect 15108 2790 15160 2796
rect 14289 2748 14585 2768
rect 14345 2746 14369 2748
rect 14425 2746 14449 2748
rect 14505 2746 14529 2748
rect 14367 2694 14369 2746
rect 14431 2694 14443 2746
rect 14505 2694 14507 2746
rect 14345 2692 14369 2694
rect 14425 2692 14449 2694
rect 14505 2692 14529 2694
rect 14289 2672 14585 2692
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 13636 2304 13688 2310
rect 13636 2246 13688 2252
rect 14096 2304 14148 2310
rect 14096 2246 14148 2252
rect 13648 2106 13676 2246
rect 13636 2100 13688 2106
rect 13636 2042 13688 2048
rect 14108 2038 14136 2246
rect 14096 2032 14148 2038
rect 14096 1974 14148 1980
rect 15120 1601 15148 2790
rect 15304 2650 15332 3606
rect 15292 2644 15344 2650
rect 15292 2586 15344 2592
rect 15200 2304 15252 2310
rect 15200 2246 15252 2252
rect 15212 2009 15240 2246
rect 15198 2000 15254 2009
rect 15198 1935 15254 1944
rect 15106 1592 15162 1601
rect 15106 1527 15162 1536
rect 9784 54 10010 82
rect 10324 128 10376 134
rect 10324 70 10376 76
rect 12806 128 12862 480
rect 12806 76 12808 128
rect 12860 76 12862 128
rect 9954 0 10010 54
rect 12806 0 12862 76
rect 15396 82 15424 6310
rect 15580 5914 15608 9318
rect 15660 7336 15712 7342
rect 15660 7278 15712 7284
rect 15672 6934 15700 7278
rect 15752 7200 15804 7206
rect 15752 7142 15804 7148
rect 15660 6928 15712 6934
rect 15660 6870 15712 6876
rect 15672 6390 15700 6870
rect 15764 6458 15792 7142
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15660 6384 15712 6390
rect 15660 6326 15712 6332
rect 15568 5908 15620 5914
rect 15488 5868 15568 5896
rect 15488 5778 15516 5868
rect 15568 5850 15620 5856
rect 15476 5772 15528 5778
rect 15476 5714 15528 5720
rect 15568 5772 15620 5778
rect 15568 5714 15620 5720
rect 15476 5636 15528 5642
rect 15476 5578 15528 5584
rect 15488 3738 15516 5578
rect 15580 5030 15608 5714
rect 15568 5024 15620 5030
rect 15568 4966 15620 4972
rect 15580 4146 15608 4966
rect 15856 4826 15884 10406
rect 16040 10062 16068 10474
rect 16120 10464 16172 10470
rect 16120 10406 16172 10412
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 15934 9616 15990 9625
rect 15934 9551 15990 9560
rect 15948 8537 15976 9551
rect 16040 8974 16068 9998
rect 16028 8968 16080 8974
rect 16028 8910 16080 8916
rect 15934 8528 15990 8537
rect 15934 8463 15990 8472
rect 15936 8288 15988 8294
rect 15936 8230 15988 8236
rect 15948 5642 15976 8230
rect 16040 8022 16068 8910
rect 16028 8016 16080 8022
rect 16028 7958 16080 7964
rect 16028 7404 16080 7410
rect 16028 7346 16080 7352
rect 16040 7002 16068 7346
rect 16028 6996 16080 7002
rect 16028 6938 16080 6944
rect 16028 6180 16080 6186
rect 16028 6122 16080 6128
rect 15936 5636 15988 5642
rect 15936 5578 15988 5584
rect 16040 5098 16068 6122
rect 16028 5092 16080 5098
rect 16028 5034 16080 5040
rect 15844 4820 15896 4826
rect 15844 4762 15896 4768
rect 15936 4752 15988 4758
rect 15936 4694 15988 4700
rect 15660 4208 15712 4214
rect 15660 4150 15712 4156
rect 15568 4140 15620 4146
rect 15568 4082 15620 4088
rect 15672 3738 15700 4150
rect 15948 3942 15976 4694
rect 15936 3936 15988 3942
rect 15936 3878 15988 3884
rect 15476 3732 15528 3738
rect 15476 3674 15528 3680
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 15568 3460 15620 3466
rect 15568 3402 15620 3408
rect 15580 3126 15608 3402
rect 15568 3120 15620 3126
rect 15568 3062 15620 3068
rect 15672 2922 15700 3470
rect 15752 3392 15804 3398
rect 15752 3334 15804 3340
rect 15844 3392 15896 3398
rect 15844 3334 15896 3340
rect 15660 2916 15712 2922
rect 15660 2858 15712 2864
rect 15764 2145 15792 3334
rect 15856 2514 15884 3334
rect 15948 2514 15976 3878
rect 15844 2508 15896 2514
rect 15844 2450 15896 2456
rect 15936 2508 15988 2514
rect 15936 2450 15988 2456
rect 16132 2378 16160 10406
rect 16212 6656 16264 6662
rect 16212 6598 16264 6604
rect 16224 6254 16252 6598
rect 16212 6248 16264 6254
rect 16212 6190 16264 6196
rect 16224 5846 16252 6190
rect 16212 5840 16264 5846
rect 16212 5782 16264 5788
rect 16316 5574 16344 10678
rect 16408 9110 16436 11018
rect 16500 10538 16528 11154
rect 16488 10532 16540 10538
rect 16488 10474 16540 10480
rect 16592 10266 16620 15558
rect 19628 15558 19946 15586
rect 19628 12986 19656 15558
rect 19890 15520 19946 15558
rect 23570 15586 23626 16000
rect 27158 15586 27214 16000
rect 23570 15558 23704 15586
rect 23570 15520 23626 15558
rect 23676 13814 23704 15558
rect 23584 13786 23704 13814
rect 26988 15558 27214 15586
rect 20956 13084 21252 13104
rect 21012 13082 21036 13084
rect 21092 13082 21116 13084
rect 21172 13082 21196 13084
rect 21034 13030 21036 13082
rect 21098 13030 21110 13082
rect 21172 13030 21174 13082
rect 21012 13028 21036 13030
rect 21092 13028 21116 13030
rect 21172 13028 21196 13030
rect 20956 13008 21252 13028
rect 19616 12980 19668 12986
rect 19616 12922 19668 12928
rect 16856 12708 16908 12714
rect 16856 12650 16908 12656
rect 16764 12096 16816 12102
rect 16764 12038 16816 12044
rect 16672 10668 16724 10674
rect 16672 10610 16724 10616
rect 16684 10470 16712 10610
rect 16672 10464 16724 10470
rect 16672 10406 16724 10412
rect 16580 10260 16632 10266
rect 16580 10202 16632 10208
rect 16488 9512 16540 9518
rect 16488 9454 16540 9460
rect 16396 9104 16448 9110
rect 16396 9046 16448 9052
rect 16408 8566 16436 9046
rect 16396 8560 16448 8566
rect 16396 8502 16448 8508
rect 16500 7993 16528 9454
rect 16580 8356 16632 8362
rect 16580 8298 16632 8304
rect 16592 8090 16620 8298
rect 16580 8084 16632 8090
rect 16580 8026 16632 8032
rect 16486 7984 16542 7993
rect 16486 7919 16542 7928
rect 16500 7818 16528 7919
rect 16488 7812 16540 7818
rect 16488 7754 16540 7760
rect 16304 5568 16356 5574
rect 16304 5510 16356 5516
rect 16304 4616 16356 4622
rect 16304 4558 16356 4564
rect 16316 4154 16344 4558
rect 16580 4276 16632 4282
rect 16684 4264 16712 10406
rect 16776 7002 16804 12038
rect 16868 11354 16896 12650
rect 19248 12640 19300 12646
rect 19248 12582 19300 12588
rect 19260 12306 19288 12582
rect 17040 12300 17092 12306
rect 17040 12242 17092 12248
rect 19248 12300 19300 12306
rect 19248 12242 19300 12248
rect 19708 12300 19760 12306
rect 19708 12242 19760 12248
rect 23480 12300 23532 12306
rect 23480 12242 23532 12248
rect 17052 11898 17080 12242
rect 18144 12232 18196 12238
rect 18144 12174 18196 12180
rect 17040 11892 17092 11898
rect 17040 11834 17092 11840
rect 17590 11792 17646 11801
rect 17590 11727 17646 11736
rect 17224 11620 17276 11626
rect 17224 11562 17276 11568
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 17236 10130 17264 11562
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 17236 9722 17264 10066
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 16948 9444 17000 9450
rect 16948 9386 17000 9392
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16868 8294 16896 8978
rect 16856 8288 16908 8294
rect 16856 8230 16908 8236
rect 16960 7954 16988 9386
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 17040 8016 17092 8022
rect 17040 7958 17092 7964
rect 16948 7948 17000 7954
rect 16948 7890 17000 7896
rect 16960 7546 16988 7890
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 17052 7478 17080 7958
rect 17040 7472 17092 7478
rect 17040 7414 17092 7420
rect 16764 6996 16816 7002
rect 16764 6938 16816 6944
rect 17052 6186 17080 7414
rect 17144 7410 17172 8434
rect 17132 7404 17184 7410
rect 17132 7346 17184 7352
rect 17316 7268 17368 7274
rect 17316 7210 17368 7216
rect 17132 6928 17184 6934
rect 17132 6870 17184 6876
rect 17144 6798 17172 6870
rect 17132 6792 17184 6798
rect 17132 6734 17184 6740
rect 17144 6440 17172 6734
rect 17224 6452 17276 6458
rect 17144 6412 17224 6440
rect 17224 6394 17276 6400
rect 17040 6180 17092 6186
rect 17040 6122 17092 6128
rect 17328 6118 17356 7210
rect 17420 6322 17448 11494
rect 17604 11286 17632 11727
rect 17960 11552 18012 11558
rect 17960 11494 18012 11500
rect 17500 11280 17552 11286
rect 17500 11222 17552 11228
rect 17592 11280 17644 11286
rect 17592 11222 17644 11228
rect 17512 9042 17540 11222
rect 17776 11008 17828 11014
rect 17776 10950 17828 10956
rect 17788 10470 17816 10950
rect 17776 10464 17828 10470
rect 17776 10406 17828 10412
rect 17788 9994 17816 10406
rect 17972 10266 18000 11494
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 17776 9988 17828 9994
rect 17776 9930 17828 9936
rect 17868 9648 17920 9654
rect 17868 9590 17920 9596
rect 17880 9450 17908 9590
rect 17972 9586 18000 10202
rect 18156 10062 18184 12174
rect 18604 12164 18656 12170
rect 18604 12106 18656 12112
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 18236 11688 18288 11694
rect 18236 11630 18288 11636
rect 18248 11014 18276 11630
rect 18236 11008 18288 11014
rect 18236 10950 18288 10956
rect 18248 10305 18276 10950
rect 18234 10296 18290 10305
rect 18234 10231 18290 10240
rect 18236 10192 18288 10198
rect 18236 10134 18288 10140
rect 18144 10056 18196 10062
rect 18144 9998 18196 10004
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 17868 9444 17920 9450
rect 17868 9386 17920 9392
rect 17500 9036 17552 9042
rect 17500 8978 17552 8984
rect 17512 8634 17540 8978
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 17776 8084 17828 8090
rect 17776 8026 17828 8032
rect 17788 7546 17816 8026
rect 17880 8022 17908 9386
rect 18156 9178 18184 9998
rect 18248 9518 18276 10134
rect 18236 9512 18288 9518
rect 18236 9454 18288 9460
rect 18248 9178 18276 9454
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 18236 9172 18288 9178
rect 18236 9114 18288 9120
rect 18432 8090 18460 12038
rect 18420 8084 18472 8090
rect 18420 8026 18472 8032
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17776 7540 17828 7546
rect 17776 7482 17828 7488
rect 17788 7206 17816 7482
rect 17960 7472 18012 7478
rect 17960 7414 18012 7420
rect 17776 7200 17828 7206
rect 17776 7142 17828 7148
rect 17972 6730 18000 7414
rect 18432 7410 18460 8026
rect 18420 7404 18472 7410
rect 18420 7346 18472 7352
rect 18616 6798 18644 12106
rect 18696 11688 18748 11694
rect 18696 11630 18748 11636
rect 19062 11656 19118 11665
rect 18708 11150 18736 11630
rect 19062 11591 19118 11600
rect 19076 11558 19104 11591
rect 19260 11558 19288 12242
rect 19720 11830 19748 12242
rect 19800 12096 19852 12102
rect 19800 12038 19852 12044
rect 19708 11824 19760 11830
rect 19708 11766 19760 11772
rect 19064 11552 19116 11558
rect 19248 11552 19300 11558
rect 19064 11494 19116 11500
rect 19168 11512 19248 11540
rect 19064 11348 19116 11354
rect 19064 11290 19116 11296
rect 18696 11144 18748 11150
rect 18696 11086 18748 11092
rect 18880 10600 18932 10606
rect 18880 10542 18932 10548
rect 18694 9480 18750 9489
rect 18694 9415 18750 9424
rect 18708 8430 18736 9415
rect 18788 9376 18840 9382
rect 18788 9318 18840 9324
rect 18696 8424 18748 8430
rect 18696 8366 18748 8372
rect 18708 7954 18736 8366
rect 18696 7948 18748 7954
rect 18696 7890 18748 7896
rect 18604 6792 18656 6798
rect 18050 6760 18106 6769
rect 17960 6724 18012 6730
rect 18604 6734 18656 6740
rect 18050 6695 18106 6704
rect 17960 6666 18012 6672
rect 17972 6322 18000 6666
rect 17408 6316 17460 6322
rect 17408 6258 17460 6264
rect 17960 6316 18012 6322
rect 17960 6258 18012 6264
rect 17316 6112 17368 6118
rect 17316 6054 17368 6060
rect 17040 5840 17092 5846
rect 17040 5782 17092 5788
rect 16764 5568 16816 5574
rect 16764 5510 16816 5516
rect 16776 5030 16804 5510
rect 17052 5370 17080 5782
rect 17224 5636 17276 5642
rect 17328 5624 17356 6054
rect 17420 5914 17448 6258
rect 18064 5914 18092 6695
rect 18236 6656 18288 6662
rect 18236 6598 18288 6604
rect 18248 6390 18276 6598
rect 18236 6384 18288 6390
rect 18236 6326 18288 6332
rect 18248 6186 18276 6326
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 18236 6180 18288 6186
rect 18236 6122 18288 6128
rect 18524 5914 18552 6258
rect 18616 5914 18644 6734
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 18512 5908 18564 5914
rect 18512 5850 18564 5856
rect 18604 5908 18656 5914
rect 18604 5850 18656 5856
rect 17408 5636 17460 5642
rect 17328 5596 17408 5624
rect 17224 5578 17276 5584
rect 17408 5578 17460 5584
rect 17040 5364 17092 5370
rect 17040 5306 17092 5312
rect 17236 5234 17264 5578
rect 17420 5273 17448 5578
rect 17406 5264 17462 5273
rect 17224 5228 17276 5234
rect 17406 5199 17462 5208
rect 17224 5170 17276 5176
rect 18064 5166 18092 5850
rect 18144 5704 18196 5710
rect 18144 5646 18196 5652
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 18156 5030 18184 5646
rect 16764 5024 16816 5030
rect 16764 4966 16816 4972
rect 18144 5024 18196 5030
rect 18144 4966 18196 4972
rect 16776 4554 16804 4966
rect 16948 4684 17000 4690
rect 16948 4626 17000 4632
rect 16764 4548 16816 4554
rect 16764 4490 16816 4496
rect 16776 4282 16804 4490
rect 16632 4236 16712 4264
rect 16580 4218 16632 4224
rect 16486 4176 16542 4185
rect 16316 4126 16436 4154
rect 16408 4078 16436 4126
rect 16486 4111 16542 4120
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16500 2582 16528 4111
rect 16580 4072 16632 4078
rect 16580 4014 16632 4020
rect 16592 3670 16620 4014
rect 16580 3664 16632 3670
rect 16580 3606 16632 3612
rect 16592 2854 16620 3606
rect 16684 3466 16712 4236
rect 16764 4276 16816 4282
rect 16764 4218 16816 4224
rect 16776 3602 16804 4218
rect 16856 4140 16908 4146
rect 16856 4082 16908 4088
rect 16764 3596 16816 3602
rect 16764 3538 16816 3544
rect 16672 3460 16724 3466
rect 16672 3402 16724 3408
rect 16684 2922 16712 3402
rect 16868 3126 16896 4082
rect 16960 3942 16988 4626
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17420 3942 17448 4558
rect 18144 4480 18196 4486
rect 18144 4422 18196 4428
rect 18156 4078 18184 4422
rect 18800 4214 18828 9318
rect 18892 9217 18920 10542
rect 18878 9208 18934 9217
rect 18878 9143 18934 9152
rect 19076 9042 19104 11290
rect 19064 9036 19116 9042
rect 19064 8978 19116 8984
rect 18972 8832 19024 8838
rect 18972 8774 19024 8780
rect 18984 8498 19012 8774
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 18972 8492 19024 8498
rect 18972 8434 19024 8440
rect 18892 6798 18920 8434
rect 18984 8090 19012 8434
rect 18972 8084 19024 8090
rect 18972 8026 19024 8032
rect 18972 7948 19024 7954
rect 18972 7890 19024 7896
rect 18984 7546 19012 7890
rect 19076 7886 19104 8978
rect 19168 8634 19196 11512
rect 19248 11494 19300 11500
rect 19340 11212 19392 11218
rect 19340 11154 19392 11160
rect 19248 10532 19300 10538
rect 19248 10474 19300 10480
rect 19260 9586 19288 10474
rect 19352 10470 19380 11154
rect 19432 10600 19484 10606
rect 19432 10542 19484 10548
rect 19340 10464 19392 10470
rect 19340 10406 19392 10412
rect 19248 9580 19300 9586
rect 19248 9522 19300 9528
rect 19246 9208 19302 9217
rect 19246 9143 19302 9152
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 18972 7540 19024 7546
rect 18972 7482 19024 7488
rect 18880 6792 18932 6798
rect 18880 6734 18932 6740
rect 19260 5778 19288 9143
rect 19352 6322 19380 10406
rect 19444 7954 19472 10542
rect 19524 10124 19576 10130
rect 19524 10066 19576 10072
rect 19536 9382 19564 10066
rect 19524 9376 19576 9382
rect 19524 9318 19576 9324
rect 19524 8356 19576 8362
rect 19524 8298 19576 8304
rect 19536 8090 19564 8298
rect 19524 8084 19576 8090
rect 19524 8026 19576 8032
rect 19432 7948 19484 7954
rect 19432 7890 19484 7896
rect 19444 7546 19472 7890
rect 19432 7540 19484 7546
rect 19432 7482 19484 7488
rect 19340 6316 19392 6322
rect 19340 6258 19392 6264
rect 19248 5772 19300 5778
rect 19248 5714 19300 5720
rect 19260 5681 19288 5714
rect 19246 5672 19302 5681
rect 19246 5607 19302 5616
rect 19260 5370 19288 5607
rect 19248 5364 19300 5370
rect 19248 5306 19300 5312
rect 18880 4684 18932 4690
rect 18880 4626 18932 4632
rect 19156 4684 19208 4690
rect 19156 4626 19208 4632
rect 18788 4208 18840 4214
rect 18788 4150 18840 4156
rect 18892 4078 18920 4626
rect 17960 4072 18012 4078
rect 17960 4014 18012 4020
rect 18144 4072 18196 4078
rect 18144 4014 18196 4020
rect 18880 4072 18932 4078
rect 18880 4014 18932 4020
rect 16948 3936 17000 3942
rect 16948 3878 17000 3884
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 16960 3602 16988 3878
rect 17420 3670 17448 3878
rect 17408 3664 17460 3670
rect 17408 3606 17460 3612
rect 16948 3596 17000 3602
rect 16948 3538 17000 3544
rect 17224 3528 17276 3534
rect 17224 3470 17276 3476
rect 17236 3194 17264 3470
rect 17420 3398 17448 3606
rect 17972 3602 18000 4014
rect 18156 3602 18184 4014
rect 17960 3596 18012 3602
rect 17960 3538 18012 3544
rect 18144 3596 18196 3602
rect 18144 3538 18196 3544
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 17972 3194 18000 3538
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 16856 3120 16908 3126
rect 16856 3062 16908 3068
rect 18156 3058 18184 3538
rect 18788 3460 18840 3466
rect 18788 3402 18840 3408
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 18800 2990 18828 3402
rect 18892 3398 18920 4014
rect 19168 3942 19196 4626
rect 19248 4548 19300 4554
rect 19248 4490 19300 4496
rect 19260 4128 19288 4490
rect 19340 4140 19392 4146
rect 19260 4100 19340 4128
rect 19340 4082 19392 4088
rect 19156 3936 19208 3942
rect 19156 3878 19208 3884
rect 18972 3732 19024 3738
rect 18972 3674 19024 3680
rect 18880 3392 18932 3398
rect 18880 3334 18932 3340
rect 18788 2984 18840 2990
rect 18788 2926 18840 2932
rect 16672 2916 16724 2922
rect 16672 2858 16724 2864
rect 17224 2916 17276 2922
rect 17224 2858 17276 2864
rect 16580 2848 16632 2854
rect 16580 2790 16632 2796
rect 17236 2582 17264 2858
rect 18604 2848 18656 2854
rect 18604 2790 18656 2796
rect 16488 2576 16540 2582
rect 16488 2518 16540 2524
rect 17224 2576 17276 2582
rect 17224 2518 17276 2524
rect 17776 2576 17828 2582
rect 17776 2518 17828 2524
rect 16396 2508 16448 2514
rect 16396 2450 16448 2456
rect 16120 2372 16172 2378
rect 16120 2314 16172 2320
rect 16408 2310 16436 2450
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 16396 2304 16448 2310
rect 16396 2246 16448 2252
rect 15750 2136 15806 2145
rect 15750 2071 15806 2080
rect 16960 1329 16988 2382
rect 17788 1737 17816 2518
rect 18616 2514 18644 2790
rect 18984 2650 19012 3674
rect 19168 3126 19196 3878
rect 19522 3496 19578 3505
rect 19522 3431 19578 3440
rect 19156 3120 19208 3126
rect 19156 3062 19208 3068
rect 19536 3058 19564 3431
rect 19720 3058 19748 11766
rect 19812 11218 19840 12038
rect 20956 11996 21252 12016
rect 21012 11994 21036 11996
rect 21092 11994 21116 11996
rect 21172 11994 21196 11996
rect 21034 11942 21036 11994
rect 21098 11942 21110 11994
rect 21172 11942 21174 11994
rect 21012 11940 21036 11942
rect 21092 11940 21116 11942
rect 21172 11940 21196 11942
rect 20956 11920 21252 11940
rect 23020 11892 23072 11898
rect 23020 11834 23072 11840
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 19984 11552 20036 11558
rect 19984 11494 20036 11500
rect 19996 11218 20024 11494
rect 19800 11212 19852 11218
rect 19800 11154 19852 11160
rect 19984 11212 20036 11218
rect 19984 11154 20036 11160
rect 19812 10742 19840 11154
rect 20168 11008 20220 11014
rect 20168 10950 20220 10956
rect 19800 10736 19852 10742
rect 19800 10678 19852 10684
rect 20180 10674 20208 10950
rect 20168 10668 20220 10674
rect 20168 10610 20220 10616
rect 20168 10532 20220 10538
rect 20168 10474 20220 10480
rect 20180 9926 20208 10474
rect 19892 9920 19944 9926
rect 19892 9862 19944 9868
rect 20168 9920 20220 9926
rect 20168 9862 20220 9868
rect 19904 8566 19932 9862
rect 20180 9654 20208 9862
rect 20168 9648 20220 9654
rect 20168 9590 20220 9596
rect 20076 9444 20128 9450
rect 20076 9386 20128 9392
rect 19984 9376 20036 9382
rect 19984 9318 20036 9324
rect 19892 8560 19944 8566
rect 19892 8502 19944 8508
rect 19890 8392 19946 8401
rect 19996 8378 20024 9318
rect 20088 9178 20116 9386
rect 20076 9172 20128 9178
rect 20076 9114 20128 9120
rect 19946 8350 20024 8378
rect 20088 8362 20116 9114
rect 20180 8634 20208 9590
rect 20260 9580 20312 9586
rect 20260 9522 20312 9528
rect 20272 9178 20300 9522
rect 20260 9172 20312 9178
rect 20260 9114 20312 9120
rect 20168 8628 20220 8634
rect 20168 8570 20220 8576
rect 20076 8356 20128 8362
rect 19890 8327 19946 8336
rect 19904 7546 19932 8327
rect 20076 8298 20128 8304
rect 20088 7750 20116 8298
rect 20076 7744 20128 7750
rect 20076 7686 20128 7692
rect 19892 7540 19944 7546
rect 19892 7482 19944 7488
rect 19904 7342 19932 7482
rect 19892 7336 19944 7342
rect 19892 7278 19944 7284
rect 20168 7336 20220 7342
rect 20168 7278 20220 7284
rect 20180 7002 20208 7278
rect 20168 6996 20220 7002
rect 20168 6938 20220 6944
rect 20180 6458 20208 6938
rect 20364 6866 20392 11698
rect 22376 11688 22428 11694
rect 22376 11630 22428 11636
rect 21640 11620 21692 11626
rect 21640 11562 21692 11568
rect 21272 11076 21324 11082
rect 21272 11018 21324 11024
rect 20956 10908 21252 10928
rect 21012 10906 21036 10908
rect 21092 10906 21116 10908
rect 21172 10906 21196 10908
rect 21034 10854 21036 10906
rect 21098 10854 21110 10906
rect 21172 10854 21174 10906
rect 21012 10852 21036 10854
rect 21092 10852 21116 10854
rect 21172 10852 21196 10854
rect 20956 10832 21252 10852
rect 21284 10810 21312 11018
rect 21272 10804 21324 10810
rect 21272 10746 21324 10752
rect 20812 10532 20864 10538
rect 20812 10474 20864 10480
rect 20824 10062 20852 10474
rect 21272 10192 21324 10198
rect 21272 10134 21324 10140
rect 20812 10056 20864 10062
rect 20812 9998 20864 10004
rect 20824 9178 20852 9998
rect 20956 9820 21252 9840
rect 21012 9818 21036 9820
rect 21092 9818 21116 9820
rect 21172 9818 21196 9820
rect 21034 9766 21036 9818
rect 21098 9766 21110 9818
rect 21172 9766 21174 9818
rect 21012 9764 21036 9766
rect 21092 9764 21116 9766
rect 21172 9764 21196 9766
rect 20956 9744 21252 9764
rect 21284 9722 21312 10134
rect 21548 9988 21600 9994
rect 21548 9930 21600 9936
rect 21272 9716 21324 9722
rect 21272 9658 21324 9664
rect 20812 9172 20864 9178
rect 20812 9114 20864 9120
rect 20720 8968 20772 8974
rect 20720 8910 20772 8916
rect 20732 8022 20760 8910
rect 21560 8906 21588 9930
rect 21652 9586 21680 11562
rect 22388 10606 22416 11630
rect 22928 11552 22980 11558
rect 22928 11494 22980 11500
rect 22940 11354 22968 11494
rect 22928 11348 22980 11354
rect 22928 11290 22980 11296
rect 23032 11286 23060 11834
rect 23492 11558 23520 12242
rect 23480 11552 23532 11558
rect 23480 11494 23532 11500
rect 23020 11280 23072 11286
rect 23020 11222 23072 11228
rect 23492 11218 23520 11494
rect 23480 11212 23532 11218
rect 23480 11154 23532 11160
rect 23020 11144 23072 11150
rect 23020 11086 23072 11092
rect 22836 10736 22888 10742
rect 22836 10678 22888 10684
rect 22376 10600 22428 10606
rect 22376 10542 22428 10548
rect 22560 10600 22612 10606
rect 22560 10542 22612 10548
rect 22468 10532 22520 10538
rect 22468 10474 22520 10480
rect 22480 10130 22508 10474
rect 22468 10124 22520 10130
rect 22468 10066 22520 10072
rect 21732 9648 21784 9654
rect 21732 9590 21784 9596
rect 21640 9580 21692 9586
rect 21640 9522 21692 9528
rect 21652 9178 21680 9522
rect 21744 9450 21772 9590
rect 21916 9580 21968 9586
rect 21916 9522 21968 9528
rect 21928 9489 21956 9522
rect 21914 9480 21970 9489
rect 21732 9444 21784 9450
rect 21914 9415 21970 9424
rect 21732 9386 21784 9392
rect 21640 9172 21692 9178
rect 21640 9114 21692 9120
rect 21928 8974 21956 9415
rect 22480 9382 22508 10066
rect 22468 9376 22520 9382
rect 22468 9318 22520 9324
rect 22100 9104 22152 9110
rect 22100 9046 22152 9052
rect 21916 8968 21968 8974
rect 21916 8910 21968 8916
rect 21548 8900 21600 8906
rect 21548 8842 21600 8848
rect 21272 8832 21324 8838
rect 21272 8774 21324 8780
rect 20956 8732 21252 8752
rect 21012 8730 21036 8732
rect 21092 8730 21116 8732
rect 21172 8730 21196 8732
rect 21034 8678 21036 8730
rect 21098 8678 21110 8730
rect 21172 8678 21174 8730
rect 21012 8676 21036 8678
rect 21092 8676 21116 8678
rect 21172 8676 21196 8678
rect 20956 8656 21252 8676
rect 21284 8430 21312 8774
rect 22112 8634 22140 9046
rect 22100 8628 22152 8634
rect 22100 8570 22152 8576
rect 21364 8492 21416 8498
rect 21364 8434 21416 8440
rect 21272 8424 21324 8430
rect 21272 8366 21324 8372
rect 20720 8016 20772 8022
rect 20720 7958 20772 7964
rect 21376 7954 21404 8434
rect 21824 8356 21876 8362
rect 21824 8298 21876 8304
rect 21364 7948 21416 7954
rect 21364 7890 21416 7896
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 20956 7644 21252 7664
rect 21012 7642 21036 7644
rect 21092 7642 21116 7644
rect 21172 7642 21196 7644
rect 21034 7590 21036 7642
rect 21098 7590 21110 7642
rect 21172 7590 21174 7642
rect 21012 7588 21036 7590
rect 21092 7588 21116 7590
rect 21172 7588 21196 7590
rect 20956 7568 21252 7588
rect 21180 7404 21232 7410
rect 21284 7392 21312 7822
rect 21232 7364 21312 7392
rect 21180 7346 21232 7352
rect 21192 7313 21220 7346
rect 21376 7342 21404 7890
rect 21640 7880 21692 7886
rect 21640 7822 21692 7828
rect 21548 7744 21600 7750
rect 21548 7686 21600 7692
rect 21364 7336 21416 7342
rect 21178 7304 21234 7313
rect 20812 7268 20864 7274
rect 21364 7278 21416 7284
rect 21560 7274 21588 7686
rect 21652 7410 21680 7822
rect 21640 7404 21692 7410
rect 21640 7346 21692 7352
rect 21178 7239 21234 7248
rect 21548 7268 21600 7274
rect 20812 7210 20864 7216
rect 21548 7210 21600 7216
rect 20824 7002 20852 7210
rect 20812 6996 20864 7002
rect 20812 6938 20864 6944
rect 21732 6996 21784 7002
rect 21732 6938 21784 6944
rect 20352 6860 20404 6866
rect 20352 6802 20404 6808
rect 21364 6860 21416 6866
rect 21364 6802 21416 6808
rect 20956 6556 21252 6576
rect 21012 6554 21036 6556
rect 21092 6554 21116 6556
rect 21172 6554 21196 6556
rect 21034 6502 21036 6554
rect 21098 6502 21110 6554
rect 21172 6502 21174 6554
rect 21012 6500 21036 6502
rect 21092 6500 21116 6502
rect 21172 6500 21196 6502
rect 20956 6480 21252 6500
rect 19800 6452 19852 6458
rect 19800 6394 19852 6400
rect 20168 6452 20220 6458
rect 20168 6394 20220 6400
rect 19812 5778 19840 6394
rect 20166 6352 20222 6361
rect 20166 6287 20222 6296
rect 20180 6254 20208 6287
rect 20168 6248 20220 6254
rect 20168 6190 20220 6196
rect 21376 6118 21404 6802
rect 21744 6322 21772 6938
rect 21836 6866 21864 8298
rect 21824 6860 21876 6866
rect 21824 6802 21876 6808
rect 22468 6860 22520 6866
rect 22468 6802 22520 6808
rect 21732 6316 21784 6322
rect 21732 6258 21784 6264
rect 22376 6248 22428 6254
rect 22376 6190 22428 6196
rect 21456 6180 21508 6186
rect 21456 6122 21508 6128
rect 21916 6180 21968 6186
rect 21916 6122 21968 6128
rect 21364 6112 21416 6118
rect 21364 6054 21416 6060
rect 19800 5772 19852 5778
rect 19800 5714 19852 5720
rect 19812 5166 19840 5714
rect 21468 5710 21496 6122
rect 21824 6112 21876 6118
rect 21824 6054 21876 6060
rect 21272 5704 21324 5710
rect 21272 5646 21324 5652
rect 21456 5704 21508 5710
rect 21456 5646 21508 5652
rect 20956 5468 21252 5488
rect 21012 5466 21036 5468
rect 21092 5466 21116 5468
rect 21172 5466 21196 5468
rect 21034 5414 21036 5466
rect 21098 5414 21110 5466
rect 21172 5414 21174 5466
rect 21012 5412 21036 5414
rect 21092 5412 21116 5414
rect 21172 5412 21196 5414
rect 20956 5392 21252 5412
rect 21284 5234 21312 5646
rect 21468 5302 21496 5646
rect 21456 5296 21508 5302
rect 21456 5238 21508 5244
rect 21272 5228 21324 5234
rect 21272 5170 21324 5176
rect 19800 5160 19852 5166
rect 19800 5102 19852 5108
rect 19812 4826 19840 5102
rect 20444 5092 20496 5098
rect 20444 5034 20496 5040
rect 19800 4820 19852 4826
rect 19800 4762 19852 4768
rect 20456 4622 20484 5034
rect 21548 5024 21600 5030
rect 21548 4966 21600 4972
rect 21560 4826 21588 4966
rect 21548 4820 21600 4826
rect 21548 4762 21600 4768
rect 20444 4616 20496 4622
rect 20444 4558 20496 4564
rect 21640 4616 21692 4622
rect 21640 4558 21692 4564
rect 20956 4380 21252 4400
rect 21012 4378 21036 4380
rect 21092 4378 21116 4380
rect 21172 4378 21196 4380
rect 21034 4326 21036 4378
rect 21098 4326 21110 4378
rect 21172 4326 21174 4378
rect 21012 4324 21036 4326
rect 21092 4324 21116 4326
rect 21172 4324 21196 4326
rect 20956 4304 21252 4324
rect 21652 4214 21680 4558
rect 21640 4208 21692 4214
rect 21640 4150 21692 4156
rect 20352 4140 20404 4146
rect 20352 4082 20404 4088
rect 20364 3738 20392 4082
rect 21088 4072 21140 4078
rect 21088 4014 21140 4020
rect 21100 3738 21128 4014
rect 20352 3732 20404 3738
rect 20352 3674 20404 3680
rect 21088 3732 21140 3738
rect 21088 3674 21140 3680
rect 19800 3460 19852 3466
rect 19800 3402 19852 3408
rect 19524 3052 19576 3058
rect 19524 2994 19576 3000
rect 19708 3052 19760 3058
rect 19708 2994 19760 3000
rect 19812 2990 19840 3402
rect 20364 3126 20392 3674
rect 20628 3392 20680 3398
rect 20628 3334 20680 3340
rect 20352 3120 20404 3126
rect 20352 3062 20404 3068
rect 19800 2984 19852 2990
rect 19800 2926 19852 2932
rect 20352 2984 20404 2990
rect 20352 2926 20404 2932
rect 19984 2916 20036 2922
rect 19984 2858 20036 2864
rect 18972 2644 19024 2650
rect 18972 2586 19024 2592
rect 19996 2582 20024 2858
rect 20364 2854 20392 2926
rect 20536 2916 20588 2922
rect 20536 2858 20588 2864
rect 20352 2848 20404 2854
rect 20352 2790 20404 2796
rect 20548 2650 20576 2858
rect 20640 2650 20668 3334
rect 20956 3292 21252 3312
rect 21012 3290 21036 3292
rect 21092 3290 21116 3292
rect 21172 3290 21196 3292
rect 21034 3238 21036 3290
rect 21098 3238 21110 3290
rect 21172 3238 21174 3290
rect 21012 3236 21036 3238
rect 21092 3236 21116 3238
rect 21172 3236 21196 3238
rect 20956 3216 21252 3236
rect 20536 2644 20588 2650
rect 20536 2586 20588 2592
rect 20628 2644 20680 2650
rect 20628 2586 20680 2592
rect 21088 2644 21140 2650
rect 21088 2586 21140 2592
rect 19984 2576 20036 2582
rect 19984 2518 20036 2524
rect 18328 2508 18380 2514
rect 18328 2450 18380 2456
rect 18420 2508 18472 2514
rect 18420 2450 18472 2456
rect 18604 2508 18656 2514
rect 18604 2450 18656 2456
rect 18340 2310 18368 2450
rect 18432 2417 18460 2450
rect 18418 2408 18474 2417
rect 18418 2343 18474 2352
rect 18616 2310 18644 2450
rect 20548 2446 20576 2586
rect 21100 2514 21128 2586
rect 21088 2508 21140 2514
rect 21088 2450 21140 2456
rect 20536 2440 20588 2446
rect 20536 2382 20588 2388
rect 18328 2304 18380 2310
rect 18328 2246 18380 2252
rect 18604 2304 18656 2310
rect 18604 2246 18656 2252
rect 17774 1728 17830 1737
rect 17774 1663 17830 1672
rect 16946 1320 17002 1329
rect 16946 1255 17002 1264
rect 15658 82 15714 480
rect 18340 241 18368 2246
rect 20956 2204 21252 2224
rect 21012 2202 21036 2204
rect 21092 2202 21116 2204
rect 21172 2202 21196 2204
rect 21034 2150 21036 2202
rect 21098 2150 21110 2202
rect 21172 2150 21174 2202
rect 21012 2148 21036 2150
rect 21092 2148 21116 2150
rect 21172 2148 21196 2150
rect 20956 2128 21252 2148
rect 18786 1864 18842 1873
rect 18786 1799 18842 1808
rect 18326 232 18382 241
rect 18326 167 18382 176
rect 15396 54 15714 82
rect 15658 0 15714 54
rect 18510 82 18566 480
rect 18800 82 18828 1799
rect 21836 1465 21864 6054
rect 21928 5846 21956 6122
rect 22388 5914 22416 6190
rect 22480 5914 22508 6802
rect 22376 5908 22428 5914
rect 22376 5850 22428 5856
rect 22468 5908 22520 5914
rect 22468 5850 22520 5856
rect 21916 5840 21968 5846
rect 21916 5782 21968 5788
rect 21928 5030 21956 5782
rect 21916 5024 21968 5030
rect 21968 4984 22048 5012
rect 21916 4966 21968 4972
rect 22020 4826 22048 4984
rect 22008 4820 22060 4826
rect 22008 4762 22060 4768
rect 22020 4146 22048 4762
rect 22572 4154 22600 10542
rect 22744 10260 22796 10266
rect 22744 10202 22796 10208
rect 22652 8084 22704 8090
rect 22652 8026 22704 8032
rect 22664 7410 22692 8026
rect 22756 7954 22784 10202
rect 22848 10130 22876 10678
rect 22928 10464 22980 10470
rect 22928 10406 22980 10412
rect 22836 10124 22888 10130
rect 22836 10066 22888 10072
rect 22848 9382 22876 10066
rect 22836 9376 22888 9382
rect 22836 9318 22888 9324
rect 22836 8016 22888 8022
rect 22836 7958 22888 7964
rect 22744 7948 22796 7954
rect 22744 7890 22796 7896
rect 22756 7546 22784 7890
rect 22744 7540 22796 7546
rect 22744 7482 22796 7488
rect 22848 7478 22876 7958
rect 22940 7478 22968 10406
rect 22836 7472 22888 7478
rect 22836 7414 22888 7420
rect 22928 7472 22980 7478
rect 22928 7414 22980 7420
rect 22652 7404 22704 7410
rect 22652 7346 22704 7352
rect 22848 7274 22876 7414
rect 22836 7268 22888 7274
rect 22836 7210 22888 7216
rect 22848 6934 22876 7210
rect 22836 6928 22888 6934
rect 22836 6870 22888 6876
rect 22848 6390 22876 6870
rect 22836 6384 22888 6390
rect 22836 6326 22888 6332
rect 22848 6186 22876 6326
rect 22836 6180 22888 6186
rect 22836 6122 22888 6128
rect 23032 5234 23060 11086
rect 23296 11008 23348 11014
rect 23296 10950 23348 10956
rect 23204 10056 23256 10062
rect 23204 9998 23256 10004
rect 23216 9625 23244 9998
rect 23202 9616 23258 9625
rect 23202 9551 23258 9560
rect 23204 9376 23256 9382
rect 23204 9318 23256 9324
rect 23216 8974 23244 9318
rect 23112 8968 23164 8974
rect 23112 8910 23164 8916
rect 23204 8968 23256 8974
rect 23204 8910 23256 8916
rect 23124 8634 23152 8910
rect 23112 8628 23164 8634
rect 23112 8570 23164 8576
rect 23308 8090 23336 10950
rect 23492 10470 23520 11154
rect 23480 10464 23532 10470
rect 23584 10441 23612 13786
rect 25136 12300 25188 12306
rect 25136 12242 25188 12248
rect 24124 12096 24176 12102
rect 24124 12038 24176 12044
rect 24676 12096 24728 12102
rect 24676 12038 24728 12044
rect 23848 11348 23900 11354
rect 23848 11290 23900 11296
rect 23860 10674 23888 11290
rect 23848 10668 23900 10674
rect 23848 10610 23900 10616
rect 23940 10532 23992 10538
rect 23940 10474 23992 10480
rect 23480 10406 23532 10412
rect 23570 10432 23626 10441
rect 23492 9994 23520 10406
rect 23570 10367 23626 10376
rect 23952 10198 23980 10474
rect 23940 10192 23992 10198
rect 23940 10134 23992 10140
rect 23480 9988 23532 9994
rect 23480 9930 23532 9936
rect 23952 9926 23980 10134
rect 23388 9920 23440 9926
rect 23388 9862 23440 9868
rect 23940 9920 23992 9926
rect 23940 9862 23992 9868
rect 23400 9654 23428 9862
rect 23388 9648 23440 9654
rect 23388 9590 23440 9596
rect 23400 8906 23428 9590
rect 24136 9450 24164 12038
rect 24400 11824 24452 11830
rect 24400 11766 24452 11772
rect 24308 11552 24360 11558
rect 24308 11494 24360 11500
rect 24216 11076 24268 11082
rect 24216 11018 24268 11024
rect 24228 10130 24256 11018
rect 24320 10305 24348 11494
rect 24306 10296 24362 10305
rect 24306 10231 24362 10240
rect 24216 10124 24268 10130
rect 24216 10066 24268 10072
rect 24228 9586 24256 10066
rect 24216 9580 24268 9586
rect 24216 9522 24268 9528
rect 24124 9444 24176 9450
rect 24124 9386 24176 9392
rect 23664 9376 23716 9382
rect 23664 9318 23716 9324
rect 23480 9172 23532 9178
rect 23480 9114 23532 9120
rect 23388 8900 23440 8906
rect 23388 8842 23440 8848
rect 23492 8294 23520 9114
rect 23480 8288 23532 8294
rect 23480 8230 23532 8236
rect 23296 8084 23348 8090
rect 23296 8026 23348 8032
rect 23492 8022 23520 8230
rect 23480 8016 23532 8022
rect 23480 7958 23532 7964
rect 23676 7954 23704 9318
rect 23754 8936 23810 8945
rect 23754 8871 23810 8880
rect 23768 8430 23796 8871
rect 23756 8424 23808 8430
rect 23756 8366 23808 8372
rect 23664 7948 23716 7954
rect 23664 7890 23716 7896
rect 24122 7848 24178 7857
rect 24320 7818 24348 10231
rect 24412 10062 24440 11766
rect 24490 11656 24546 11665
rect 24490 11591 24546 11600
rect 24504 11354 24532 11591
rect 24492 11348 24544 11354
rect 24492 11290 24544 11296
rect 24688 10674 24716 12038
rect 25148 11558 25176 12242
rect 26332 11756 26384 11762
rect 26332 11698 26384 11704
rect 25136 11552 25188 11558
rect 25136 11494 25188 11500
rect 24860 11212 24912 11218
rect 24860 11154 24912 11160
rect 24676 10668 24728 10674
rect 24676 10610 24728 10616
rect 24584 10532 24636 10538
rect 24584 10474 24636 10480
rect 24400 10056 24452 10062
rect 24400 9998 24452 10004
rect 24492 10056 24544 10062
rect 24492 9998 24544 10004
rect 24412 9178 24440 9998
rect 24504 9625 24532 9998
rect 24490 9616 24546 9625
rect 24596 9586 24624 10474
rect 24490 9551 24492 9560
rect 24544 9551 24546 9560
rect 24584 9580 24636 9586
rect 24492 9522 24544 9528
rect 24584 9522 24636 9528
rect 24504 9491 24532 9522
rect 24596 9489 24624 9522
rect 24582 9480 24638 9489
rect 24582 9415 24638 9424
rect 24400 9172 24452 9178
rect 24400 9114 24452 9120
rect 24688 8838 24716 10610
rect 24872 10606 24900 11154
rect 24860 10600 24912 10606
rect 24860 10542 24912 10548
rect 24768 10464 24820 10470
rect 24768 10406 24820 10412
rect 24676 8832 24728 8838
rect 24676 8774 24728 8780
rect 24780 8650 24808 10406
rect 24504 8622 24808 8650
rect 24122 7783 24178 7792
rect 24308 7812 24360 7818
rect 23756 7200 23808 7206
rect 23756 7142 23808 7148
rect 23768 7002 23796 7142
rect 23756 6996 23808 7002
rect 23756 6938 23808 6944
rect 23296 6384 23348 6390
rect 23296 6326 23348 6332
rect 23112 6180 23164 6186
rect 23112 6122 23164 6128
rect 23124 5914 23152 6122
rect 23112 5908 23164 5914
rect 23112 5850 23164 5856
rect 23308 5710 23336 6326
rect 23388 5840 23440 5846
rect 23388 5782 23440 5788
rect 23296 5704 23348 5710
rect 23296 5646 23348 5652
rect 23020 5228 23072 5234
rect 23020 5170 23072 5176
rect 23308 4758 23336 5646
rect 23400 5370 23428 5782
rect 24136 5681 24164 7783
rect 24308 7754 24360 7760
rect 24216 6928 24268 6934
rect 24216 6870 24268 6876
rect 24400 6928 24452 6934
rect 24400 6870 24452 6876
rect 24228 6458 24256 6870
rect 24308 6792 24360 6798
rect 24308 6734 24360 6740
rect 24216 6452 24268 6458
rect 24216 6394 24268 6400
rect 24122 5672 24178 5681
rect 24122 5607 24178 5616
rect 23388 5364 23440 5370
rect 23388 5306 23440 5312
rect 23296 4752 23348 4758
rect 23480 4752 23532 4758
rect 23296 4694 23348 4700
rect 23400 4712 23480 4740
rect 23400 4282 23428 4712
rect 23480 4694 23532 4700
rect 23480 4616 23532 4622
rect 23480 4558 23532 4564
rect 23940 4616 23992 4622
rect 23940 4558 23992 4564
rect 23112 4276 23164 4282
rect 23112 4218 23164 4224
rect 23388 4276 23440 4282
rect 23388 4218 23440 4224
rect 22008 4140 22060 4146
rect 22572 4126 22692 4154
rect 22008 4082 22060 4088
rect 22020 3670 22048 4082
rect 22008 3664 22060 3670
rect 22008 3606 22060 3612
rect 22020 3194 22048 3606
rect 22008 3188 22060 3194
rect 22008 3130 22060 3136
rect 22664 2514 22692 4126
rect 23124 3194 23152 4218
rect 23388 4004 23440 4010
rect 23388 3946 23440 3952
rect 23112 3188 23164 3194
rect 23112 3130 23164 3136
rect 23124 2990 23152 3130
rect 23400 3058 23428 3946
rect 23492 3738 23520 4558
rect 23952 4146 23980 4558
rect 23940 4140 23992 4146
rect 23940 4082 23992 4088
rect 23480 3732 23532 3738
rect 23480 3674 23532 3680
rect 23388 3052 23440 3058
rect 23388 2994 23440 3000
rect 23112 2984 23164 2990
rect 23112 2926 23164 2932
rect 23492 2650 23520 3674
rect 23952 3670 23980 4082
rect 23940 3664 23992 3670
rect 23940 3606 23992 3612
rect 24032 2848 24084 2854
rect 24032 2790 24084 2796
rect 23480 2644 23532 2650
rect 23480 2586 23532 2592
rect 24044 2582 24072 2790
rect 24032 2576 24084 2582
rect 24032 2518 24084 2524
rect 22652 2508 22704 2514
rect 22652 2450 22704 2456
rect 21822 1456 21878 1465
rect 21822 1391 21878 1400
rect 18510 54 18828 82
rect 21362 128 21418 480
rect 21362 76 21364 128
rect 21416 76 21418 128
rect 18510 0 18566 54
rect 21362 0 21418 76
rect 24136 82 24164 5607
rect 24320 5574 24348 6734
rect 24412 6730 24440 6870
rect 24400 6724 24452 6730
rect 24400 6666 24452 6672
rect 24400 6180 24452 6186
rect 24400 6122 24452 6128
rect 24412 5710 24440 6122
rect 24400 5704 24452 5710
rect 24400 5646 24452 5652
rect 24216 5568 24268 5574
rect 24216 5510 24268 5516
rect 24308 5568 24360 5574
rect 24308 5510 24360 5516
rect 24228 5098 24256 5510
rect 24412 5098 24440 5646
rect 24216 5092 24268 5098
rect 24216 5034 24268 5040
rect 24400 5092 24452 5098
rect 24400 5034 24452 5040
rect 24228 4826 24256 5034
rect 24216 4820 24268 4826
rect 24216 4762 24268 4768
rect 24216 3664 24268 3670
rect 24216 3606 24268 3612
rect 24228 3466 24256 3606
rect 24216 3460 24268 3466
rect 24216 3402 24268 3408
rect 24228 2514 24256 3402
rect 24216 2508 24268 2514
rect 24216 2450 24268 2456
rect 24214 82 24270 480
rect 24504 134 24532 8622
rect 24584 8424 24636 8430
rect 24584 8366 24636 8372
rect 24860 8424 24912 8430
rect 24860 8366 24912 8372
rect 24596 4185 24624 8366
rect 24768 8016 24820 8022
rect 24768 7958 24820 7964
rect 24676 7880 24728 7886
rect 24676 7822 24728 7828
rect 24688 7342 24716 7822
rect 24780 7546 24808 7958
rect 24872 7750 24900 8366
rect 24952 8356 25004 8362
rect 24952 8298 25004 8304
rect 24860 7744 24912 7750
rect 24860 7686 24912 7692
rect 24768 7540 24820 7546
rect 24768 7482 24820 7488
rect 24676 7336 24728 7342
rect 24676 7278 24728 7284
rect 24688 6780 24716 7278
rect 24780 7002 24808 7482
rect 24768 6996 24820 7002
rect 24768 6938 24820 6944
rect 24768 6792 24820 6798
rect 24688 6752 24768 6780
rect 24768 6734 24820 6740
rect 24780 6390 24808 6734
rect 24768 6384 24820 6390
rect 24768 6326 24820 6332
rect 24872 5914 24900 7686
rect 24964 6934 24992 8298
rect 24952 6928 25004 6934
rect 24952 6870 25004 6876
rect 24860 5908 24912 5914
rect 24860 5850 24912 5856
rect 25148 5846 25176 11494
rect 25228 11212 25280 11218
rect 25228 11154 25280 11160
rect 25240 10470 25268 11154
rect 25872 11008 25924 11014
rect 25872 10950 25924 10956
rect 25884 10606 25912 10950
rect 26344 10656 26372 11698
rect 26424 11212 26476 11218
rect 26424 11154 26476 11160
rect 26436 10810 26464 11154
rect 26988 11150 27016 15558
rect 27158 15520 27214 15558
rect 30838 15586 30894 16000
rect 34426 15586 34482 16000
rect 38106 15586 38162 16000
rect 30838 15558 30972 15586
rect 30838 15520 30894 15558
rect 27622 13628 27918 13648
rect 27678 13626 27702 13628
rect 27758 13626 27782 13628
rect 27838 13626 27862 13628
rect 27700 13574 27702 13626
rect 27764 13574 27776 13626
rect 27838 13574 27840 13626
rect 27678 13572 27702 13574
rect 27758 13572 27782 13574
rect 27838 13572 27862 13574
rect 27622 13552 27918 13572
rect 28264 13184 28316 13190
rect 28264 13126 28316 13132
rect 28276 12986 28304 13126
rect 28264 12980 28316 12986
rect 28264 12922 28316 12928
rect 28724 12776 28776 12782
rect 28724 12718 28776 12724
rect 28736 12646 28764 12718
rect 28724 12640 28776 12646
rect 28724 12582 28776 12588
rect 27622 12540 27918 12560
rect 27678 12538 27702 12540
rect 27758 12538 27782 12540
rect 27838 12538 27862 12540
rect 27700 12486 27702 12538
rect 27764 12486 27776 12538
rect 27838 12486 27840 12538
rect 27678 12484 27702 12486
rect 27758 12484 27782 12486
rect 27838 12484 27862 12486
rect 27622 12464 27918 12484
rect 28080 12300 28132 12306
rect 28080 12242 28132 12248
rect 27528 12096 27580 12102
rect 27528 12038 27580 12044
rect 27344 11552 27396 11558
rect 27344 11494 27396 11500
rect 26976 11144 27028 11150
rect 26976 11086 27028 11092
rect 27068 11008 27120 11014
rect 27068 10950 27120 10956
rect 26424 10804 26476 10810
rect 26424 10746 26476 10752
rect 26344 10628 26464 10656
rect 25412 10600 25464 10606
rect 25412 10542 25464 10548
rect 25504 10600 25556 10606
rect 25504 10542 25556 10548
rect 25872 10600 25924 10606
rect 26056 10600 26108 10606
rect 25924 10560 26004 10588
rect 25872 10542 25924 10548
rect 25228 10464 25280 10470
rect 25228 10406 25280 10412
rect 25320 9444 25372 9450
rect 25320 9386 25372 9392
rect 25332 9178 25360 9386
rect 25320 9172 25372 9178
rect 25320 9114 25372 9120
rect 25320 6996 25372 7002
rect 25320 6938 25372 6944
rect 25332 6322 25360 6938
rect 25320 6316 25372 6322
rect 25320 6258 25372 6264
rect 25136 5840 25188 5846
rect 24766 5808 24822 5817
rect 25136 5782 25188 5788
rect 24766 5743 24768 5752
rect 24820 5743 24822 5752
rect 25228 5772 25280 5778
rect 24768 5714 24820 5720
rect 25228 5714 25280 5720
rect 24780 5030 24808 5714
rect 25044 5568 25096 5574
rect 25044 5510 25096 5516
rect 24858 5128 24914 5137
rect 24858 5063 24914 5072
rect 24952 5092 25004 5098
rect 24768 5024 24820 5030
rect 24768 4966 24820 4972
rect 24872 4758 24900 5063
rect 24952 5034 25004 5040
rect 24860 4752 24912 4758
rect 24860 4694 24912 4700
rect 24964 4690 24992 5034
rect 24952 4684 25004 4690
rect 24952 4626 25004 4632
rect 24768 4208 24820 4214
rect 24582 4176 24638 4185
rect 24768 4150 24820 4156
rect 24582 4111 24638 4120
rect 24780 3942 24808 4150
rect 24768 3936 24820 3942
rect 24768 3878 24820 3884
rect 24780 3534 24808 3878
rect 24964 3738 24992 4626
rect 25056 3738 25084 5510
rect 25240 5370 25268 5714
rect 25228 5364 25280 5370
rect 25228 5306 25280 5312
rect 25228 5024 25280 5030
rect 25228 4966 25280 4972
rect 25240 4758 25268 4966
rect 25228 4752 25280 4758
rect 25228 4694 25280 4700
rect 24952 3732 25004 3738
rect 24952 3674 25004 3680
rect 25044 3732 25096 3738
rect 25044 3674 25096 3680
rect 25424 3602 25452 10542
rect 25516 10169 25544 10542
rect 25594 10432 25650 10441
rect 25594 10367 25650 10376
rect 25502 10160 25558 10169
rect 25502 10095 25558 10104
rect 25504 9104 25556 9110
rect 25504 9046 25556 9052
rect 25516 7750 25544 9046
rect 25608 8514 25636 10367
rect 25688 9444 25740 9450
rect 25688 9386 25740 9392
rect 25700 8634 25728 9386
rect 25688 8628 25740 8634
rect 25688 8570 25740 8576
rect 25608 8486 25728 8514
rect 25504 7744 25556 7750
rect 25504 7686 25556 7692
rect 25516 7313 25544 7686
rect 25596 7404 25648 7410
rect 25596 7346 25648 7352
rect 25502 7304 25558 7313
rect 25502 7239 25558 7248
rect 25504 7200 25556 7206
rect 25504 7142 25556 7148
rect 25412 3596 25464 3602
rect 25412 3538 25464 3544
rect 24584 3528 24636 3534
rect 24584 3470 24636 3476
rect 24768 3528 24820 3534
rect 24768 3470 24820 3476
rect 24596 3126 24624 3470
rect 24584 3120 24636 3126
rect 24584 3062 24636 3068
rect 24596 2650 24624 3062
rect 25424 2854 25452 3538
rect 25516 3126 25544 7142
rect 25608 7002 25636 7346
rect 25596 6996 25648 7002
rect 25596 6938 25648 6944
rect 25700 6882 25728 8486
rect 25608 6854 25728 6882
rect 25504 3120 25556 3126
rect 25504 3062 25556 3068
rect 25412 2848 25464 2854
rect 25412 2790 25464 2796
rect 24584 2644 24636 2650
rect 24584 2586 24636 2592
rect 25424 1873 25452 2790
rect 25608 2514 25636 6854
rect 25872 5160 25924 5166
rect 25872 5102 25924 5108
rect 25688 5024 25740 5030
rect 25688 4966 25740 4972
rect 25700 4010 25728 4966
rect 25884 4486 25912 5102
rect 25976 4690 26004 10560
rect 26056 10542 26108 10548
rect 26068 9926 26096 10542
rect 26332 10532 26384 10538
rect 26332 10474 26384 10480
rect 26240 10124 26292 10130
rect 26240 10066 26292 10072
rect 26056 9920 26108 9926
rect 26056 9862 26108 9868
rect 26252 9382 26280 10066
rect 26240 9376 26292 9382
rect 26240 9318 26292 9324
rect 26252 8537 26280 9318
rect 26238 8528 26294 8537
rect 26344 8498 26372 10474
rect 26238 8463 26294 8472
rect 26332 8492 26384 8498
rect 26252 7206 26280 8463
rect 26332 8434 26384 8440
rect 26436 7954 26464 10628
rect 27080 10266 27108 10950
rect 27068 10260 27120 10266
rect 27068 10202 27120 10208
rect 26608 9920 26660 9926
rect 26608 9862 26660 9868
rect 26792 9920 26844 9926
rect 26792 9862 26844 9868
rect 26516 8968 26568 8974
rect 26516 8910 26568 8916
rect 26528 8090 26556 8910
rect 26516 8084 26568 8090
rect 26516 8026 26568 8032
rect 26620 7954 26648 9862
rect 26804 9217 26832 9862
rect 27080 9586 27108 10202
rect 27356 10198 27384 11494
rect 27540 10606 27568 12038
rect 28092 11558 28120 12242
rect 28080 11552 28132 11558
rect 28080 11494 28132 11500
rect 27622 11452 27918 11472
rect 27678 11450 27702 11452
rect 27758 11450 27782 11452
rect 27838 11450 27862 11452
rect 27700 11398 27702 11450
rect 27764 11398 27776 11450
rect 27838 11398 27840 11450
rect 27678 11396 27702 11398
rect 27758 11396 27782 11398
rect 27838 11396 27862 11398
rect 27622 11376 27918 11396
rect 27712 11008 27764 11014
rect 27712 10950 27764 10956
rect 27724 10606 27752 10950
rect 27528 10600 27580 10606
rect 27528 10542 27580 10548
rect 27712 10600 27764 10606
rect 27712 10542 27764 10548
rect 27622 10364 27918 10384
rect 27678 10362 27702 10364
rect 27758 10362 27782 10364
rect 27838 10362 27862 10364
rect 27700 10310 27702 10362
rect 27764 10310 27776 10362
rect 27838 10310 27840 10362
rect 27678 10308 27702 10310
rect 27758 10308 27782 10310
rect 27838 10308 27862 10310
rect 27622 10288 27918 10308
rect 27344 10192 27396 10198
rect 27344 10134 27396 10140
rect 27712 10192 27764 10198
rect 27712 10134 27764 10140
rect 27724 9722 27752 10134
rect 27712 9716 27764 9722
rect 27712 9658 27764 9664
rect 27160 9648 27212 9654
rect 27160 9590 27212 9596
rect 27068 9580 27120 9586
rect 27068 9522 27120 9528
rect 27172 9450 27200 9590
rect 27160 9444 27212 9450
rect 27160 9386 27212 9392
rect 27622 9276 27918 9296
rect 27678 9274 27702 9276
rect 27758 9274 27782 9276
rect 27838 9274 27862 9276
rect 27700 9222 27702 9274
rect 27764 9222 27776 9274
rect 27838 9222 27840 9274
rect 27678 9220 27702 9222
rect 27758 9220 27782 9222
rect 27838 9220 27862 9222
rect 26790 9208 26846 9217
rect 27622 9200 27918 9220
rect 26846 9166 26924 9194
rect 26790 9143 26846 9152
rect 26424 7948 26476 7954
rect 26608 7948 26660 7954
rect 26424 7890 26476 7896
rect 26528 7908 26608 7936
rect 26436 7342 26464 7890
rect 26424 7336 26476 7342
rect 26424 7278 26476 7284
rect 26528 7206 26556 7908
rect 26608 7890 26660 7896
rect 26896 7546 26924 9166
rect 26976 9104 27028 9110
rect 26976 9046 27028 9052
rect 26988 8362 27016 9046
rect 26976 8356 27028 8362
rect 26976 8298 27028 8304
rect 26988 8090 27016 8298
rect 27622 8188 27918 8208
rect 27678 8186 27702 8188
rect 27758 8186 27782 8188
rect 27838 8186 27862 8188
rect 27700 8134 27702 8186
rect 27764 8134 27776 8186
rect 27838 8134 27840 8186
rect 27678 8132 27702 8134
rect 27758 8132 27782 8134
rect 27838 8132 27862 8134
rect 27622 8112 27918 8132
rect 26976 8084 27028 8090
rect 26976 8026 27028 8032
rect 27528 7744 27580 7750
rect 27528 7686 27580 7692
rect 27712 7744 27764 7750
rect 27712 7686 27764 7692
rect 27540 7546 27568 7686
rect 26792 7540 26844 7546
rect 26792 7482 26844 7488
rect 26884 7540 26936 7546
rect 26884 7482 26936 7488
rect 27528 7540 27580 7546
rect 27528 7482 27580 7488
rect 26700 7268 26752 7274
rect 26700 7210 26752 7216
rect 26240 7200 26292 7206
rect 26240 7142 26292 7148
rect 26516 7200 26568 7206
rect 26516 7142 26568 7148
rect 26528 5370 26556 7142
rect 26608 6928 26660 6934
rect 26608 6870 26660 6876
rect 26620 6458 26648 6870
rect 26712 6798 26740 7210
rect 26804 6934 26832 7482
rect 27724 7342 27752 7686
rect 27712 7336 27764 7342
rect 27712 7278 27764 7284
rect 26884 7200 26936 7206
rect 26884 7142 26936 7148
rect 26792 6928 26844 6934
rect 26792 6870 26844 6876
rect 26700 6792 26752 6798
rect 26700 6734 26752 6740
rect 26608 6452 26660 6458
rect 26608 6394 26660 6400
rect 26712 6322 26740 6734
rect 26804 6390 26832 6870
rect 26792 6384 26844 6390
rect 26792 6326 26844 6332
rect 26700 6316 26752 6322
rect 26700 6258 26752 6264
rect 26516 5364 26568 5370
rect 26516 5306 26568 5312
rect 26896 5166 26924 7142
rect 27622 7100 27918 7120
rect 27678 7098 27702 7100
rect 27758 7098 27782 7100
rect 27838 7098 27862 7100
rect 27700 7046 27702 7098
rect 27764 7046 27776 7098
rect 27838 7046 27840 7098
rect 27678 7044 27702 7046
rect 27758 7044 27782 7046
rect 27838 7044 27862 7046
rect 27622 7024 27918 7044
rect 27344 6452 27396 6458
rect 27344 6394 27396 6400
rect 27356 6361 27384 6394
rect 27342 6352 27398 6361
rect 27342 6287 27398 6296
rect 27356 6254 27384 6287
rect 27344 6248 27396 6254
rect 27344 6190 27396 6196
rect 27068 6180 27120 6186
rect 27068 6122 27120 6128
rect 26884 5160 26936 5166
rect 26884 5102 26936 5108
rect 25964 4684 26016 4690
rect 25964 4626 26016 4632
rect 26792 4684 26844 4690
rect 26792 4626 26844 4632
rect 25872 4480 25924 4486
rect 25872 4422 25924 4428
rect 25780 4072 25832 4078
rect 25884 4049 25912 4422
rect 26804 4214 26832 4626
rect 26792 4208 26844 4214
rect 26792 4150 26844 4156
rect 25780 4014 25832 4020
rect 25870 4040 25926 4049
rect 25688 4004 25740 4010
rect 25688 3946 25740 3952
rect 25792 2854 25820 4014
rect 25870 3975 25926 3984
rect 25964 3732 26016 3738
rect 25964 3674 26016 3680
rect 25976 2990 26004 3674
rect 26804 3602 26832 4150
rect 26896 3738 26924 5102
rect 27080 4570 27108 6122
rect 27252 5840 27304 5846
rect 27252 5782 27304 5788
rect 27160 5704 27212 5710
rect 27160 5646 27212 5652
rect 27172 5370 27200 5646
rect 27160 5364 27212 5370
rect 27160 5306 27212 5312
rect 27264 5234 27292 5782
rect 27252 5228 27304 5234
rect 27252 5170 27304 5176
rect 27356 4826 27384 6190
rect 27622 6012 27918 6032
rect 27678 6010 27702 6012
rect 27758 6010 27782 6012
rect 27838 6010 27862 6012
rect 27700 5958 27702 6010
rect 27764 5958 27776 6010
rect 27838 5958 27840 6010
rect 27678 5956 27702 5958
rect 27758 5956 27782 5958
rect 27838 5956 27862 5958
rect 27622 5936 27918 5956
rect 27528 5160 27580 5166
rect 27528 5102 27580 5108
rect 27344 4820 27396 4826
rect 27344 4762 27396 4768
rect 27540 4706 27568 5102
rect 27622 4924 27918 4944
rect 27678 4922 27702 4924
rect 27758 4922 27782 4924
rect 27838 4922 27862 4924
rect 27700 4870 27702 4922
rect 27764 4870 27776 4922
rect 27838 4870 27840 4922
rect 27678 4868 27702 4870
rect 27758 4868 27782 4870
rect 27838 4868 27862 4870
rect 27622 4848 27918 4868
rect 28092 4729 28120 11494
rect 28632 11212 28684 11218
rect 28632 11154 28684 11160
rect 28540 11144 28592 11150
rect 28540 11086 28592 11092
rect 28172 10192 28224 10198
rect 28224 10152 28304 10180
rect 28172 10134 28224 10140
rect 28276 9382 28304 10152
rect 28552 9926 28580 11086
rect 28644 10470 28672 11154
rect 28632 10464 28684 10470
rect 28632 10406 28684 10412
rect 28632 10124 28684 10130
rect 28632 10066 28684 10072
rect 28540 9920 28592 9926
rect 28540 9862 28592 9868
rect 28356 9444 28408 9450
rect 28356 9386 28408 9392
rect 28264 9376 28316 9382
rect 28264 9318 28316 9324
rect 28276 9178 28304 9318
rect 28264 9172 28316 9178
rect 28264 9114 28316 9120
rect 28368 8974 28396 9386
rect 28448 9104 28500 9110
rect 28448 9046 28500 9052
rect 28356 8968 28408 8974
rect 28356 8910 28408 8916
rect 28368 8498 28396 8910
rect 28460 8634 28488 9046
rect 28448 8628 28500 8634
rect 28448 8570 28500 8576
rect 28356 8492 28408 8498
rect 28356 8434 28408 8440
rect 28448 7200 28500 7206
rect 28448 7142 28500 7148
rect 28460 7002 28488 7142
rect 28448 6996 28500 7002
rect 28448 6938 28500 6944
rect 28460 6254 28488 6938
rect 28448 6248 28500 6254
rect 28448 6190 28500 6196
rect 28552 6186 28580 9862
rect 28644 9518 28672 10066
rect 28736 9518 28764 12582
rect 30944 11626 30972 15558
rect 34072 15558 34482 15586
rect 34072 12986 34100 15558
rect 34426 15520 34482 15558
rect 37752 15558 38162 15586
rect 35622 14104 35678 14113
rect 35622 14039 35678 14048
rect 34289 13084 34585 13104
rect 34345 13082 34369 13084
rect 34425 13082 34449 13084
rect 34505 13082 34529 13084
rect 34367 13030 34369 13082
rect 34431 13030 34443 13082
rect 34505 13030 34507 13082
rect 34345 13028 34369 13030
rect 34425 13028 34449 13030
rect 34505 13028 34529 13030
rect 34289 13008 34585 13028
rect 35636 12986 35664 14039
rect 34060 12980 34112 12986
rect 34060 12922 34112 12928
rect 35624 12980 35676 12986
rect 35624 12922 35676 12928
rect 31392 12776 31444 12782
rect 31392 12718 31444 12724
rect 34796 12776 34848 12782
rect 34796 12718 34848 12724
rect 30932 11620 30984 11626
rect 30932 11562 30984 11568
rect 30944 11218 30972 11562
rect 30932 11212 30984 11218
rect 30932 11154 30984 11160
rect 28908 11144 28960 11150
rect 28908 11086 28960 11092
rect 28816 10736 28868 10742
rect 28816 10678 28868 10684
rect 28828 10606 28856 10678
rect 28816 10600 28868 10606
rect 28816 10542 28868 10548
rect 28632 9512 28684 9518
rect 28632 9454 28684 9460
rect 28724 9512 28776 9518
rect 28724 9454 28776 9460
rect 28724 9376 28776 9382
rect 28724 9318 28776 9324
rect 28736 8022 28764 9318
rect 28724 8016 28776 8022
rect 28724 7958 28776 7964
rect 28828 7954 28856 10542
rect 28920 9178 28948 11086
rect 29276 11008 29328 11014
rect 29276 10950 29328 10956
rect 29288 10742 29316 10950
rect 30944 10742 30972 11154
rect 29276 10736 29328 10742
rect 29276 10678 29328 10684
rect 30932 10736 30984 10742
rect 30932 10678 30984 10684
rect 29828 10532 29880 10538
rect 29828 10474 29880 10480
rect 30012 10532 30064 10538
rect 30012 10474 30064 10480
rect 29644 10464 29696 10470
rect 29644 10406 29696 10412
rect 29656 10130 29684 10406
rect 29644 10124 29696 10130
rect 29644 10066 29696 10072
rect 29000 10056 29052 10062
rect 29000 9998 29052 10004
rect 29012 9489 29040 9998
rect 28998 9480 29054 9489
rect 28998 9415 29054 9424
rect 28908 9172 28960 9178
rect 28908 9114 28960 9120
rect 29012 9110 29040 9415
rect 29656 9382 29684 10066
rect 29644 9376 29696 9382
rect 29644 9318 29696 9324
rect 29552 9172 29604 9178
rect 29552 9114 29604 9120
rect 29000 9104 29052 9110
rect 29000 9046 29052 9052
rect 29564 8498 29592 9114
rect 29552 8492 29604 8498
rect 29552 8434 29604 8440
rect 28816 7948 28868 7954
rect 28816 7890 28868 7896
rect 28828 7206 28856 7890
rect 29460 7336 29512 7342
rect 29460 7278 29512 7284
rect 29736 7336 29788 7342
rect 29736 7278 29788 7284
rect 28816 7200 28868 7206
rect 28816 7142 28868 7148
rect 28908 6928 28960 6934
rect 28908 6870 28960 6876
rect 28632 6792 28684 6798
rect 28632 6734 28684 6740
rect 28540 6180 28592 6186
rect 28540 6122 28592 6128
rect 28644 5574 28672 6734
rect 28920 6458 28948 6870
rect 29472 6458 29500 7278
rect 29748 7206 29776 7278
rect 29736 7200 29788 7206
rect 29736 7142 29788 7148
rect 29644 6792 29696 6798
rect 29644 6734 29696 6740
rect 28908 6452 28960 6458
rect 28908 6394 28960 6400
rect 29460 6452 29512 6458
rect 29460 6394 29512 6400
rect 28920 5846 28948 6394
rect 28908 5840 28960 5846
rect 28908 5782 28960 5788
rect 28724 5704 28776 5710
rect 28724 5646 28776 5652
rect 28816 5704 28868 5710
rect 28816 5646 28868 5652
rect 28632 5568 28684 5574
rect 28632 5510 28684 5516
rect 28540 5364 28592 5370
rect 28540 5306 28592 5312
rect 28448 4752 28500 4758
rect 27618 4720 27674 4729
rect 27540 4678 27618 4706
rect 27618 4655 27674 4664
rect 28078 4720 28134 4729
rect 28448 4694 28500 4700
rect 28078 4655 28134 4664
rect 27632 4622 27660 4655
rect 27620 4616 27672 4622
rect 27158 4584 27214 4593
rect 27080 4542 27158 4570
rect 27620 4558 27672 4564
rect 27988 4616 28040 4622
rect 27988 4558 28040 4564
rect 27158 4519 27214 4528
rect 27172 4154 27200 4519
rect 27252 4480 27304 4486
rect 27252 4422 27304 4428
rect 27264 4282 27292 4422
rect 27252 4276 27304 4282
rect 27252 4218 27304 4224
rect 27528 4276 27580 4282
rect 27528 4218 27580 4224
rect 27172 4126 27292 4154
rect 26884 3732 26936 3738
rect 26884 3674 26936 3680
rect 26792 3596 26844 3602
rect 26792 3538 26844 3544
rect 27068 3596 27120 3602
rect 27068 3538 27120 3544
rect 26056 3392 26108 3398
rect 26056 3334 26108 3340
rect 26068 2990 26096 3334
rect 25964 2984 26016 2990
rect 25964 2926 26016 2932
rect 26056 2984 26108 2990
rect 26056 2926 26108 2932
rect 25780 2848 25832 2854
rect 25780 2790 25832 2796
rect 26804 2650 26832 3538
rect 27080 3058 27108 3538
rect 27068 3052 27120 3058
rect 27068 2994 27120 3000
rect 26792 2644 26844 2650
rect 26792 2586 26844 2592
rect 27264 2514 27292 4126
rect 27540 4010 27568 4218
rect 27528 4004 27580 4010
rect 27528 3946 27580 3952
rect 27622 3836 27918 3856
rect 27678 3834 27702 3836
rect 27758 3834 27782 3836
rect 27838 3834 27862 3836
rect 27700 3782 27702 3834
rect 27764 3782 27776 3834
rect 27838 3782 27840 3834
rect 27678 3780 27702 3782
rect 27758 3780 27782 3782
rect 27838 3780 27862 3782
rect 27622 3760 27918 3780
rect 28000 3738 28028 4558
rect 27988 3732 28040 3738
rect 27988 3674 28040 3680
rect 28000 3058 28028 3674
rect 27988 3052 28040 3058
rect 27988 2994 28040 3000
rect 28092 2990 28120 4655
rect 28460 4282 28488 4694
rect 28448 4276 28500 4282
rect 28448 4218 28500 4224
rect 28356 3596 28408 3602
rect 28356 3538 28408 3544
rect 27344 2984 27396 2990
rect 27344 2926 27396 2932
rect 28080 2984 28132 2990
rect 28080 2926 28132 2932
rect 27356 2650 27384 2926
rect 28368 2854 28396 3538
rect 28356 2848 28408 2854
rect 28356 2790 28408 2796
rect 27622 2748 27918 2768
rect 27678 2746 27702 2748
rect 27758 2746 27782 2748
rect 27838 2746 27862 2748
rect 27700 2694 27702 2746
rect 27764 2694 27776 2746
rect 27838 2694 27840 2746
rect 27678 2692 27702 2694
rect 27758 2692 27782 2694
rect 27838 2692 27862 2694
rect 27622 2672 27918 2692
rect 27344 2644 27396 2650
rect 27344 2586 27396 2592
rect 25596 2508 25648 2514
rect 25596 2450 25648 2456
rect 27252 2508 27304 2514
rect 27252 2450 27304 2456
rect 28448 2508 28500 2514
rect 28448 2450 28500 2456
rect 28460 2378 28488 2450
rect 28552 2378 28580 5306
rect 28644 3738 28672 5510
rect 28736 4826 28764 5646
rect 28828 5030 28856 5646
rect 29184 5160 29236 5166
rect 29184 5102 29236 5108
rect 28816 5024 28868 5030
rect 28816 4966 28868 4972
rect 28724 4820 28776 4826
rect 28724 4762 28776 4768
rect 28724 4480 28776 4486
rect 28724 4422 28776 4428
rect 28736 4010 28764 4422
rect 28724 4004 28776 4010
rect 28724 3946 28776 3952
rect 28632 3732 28684 3738
rect 28632 3674 28684 3680
rect 28724 3528 28776 3534
rect 28724 3470 28776 3476
rect 28736 3194 28764 3470
rect 28724 3188 28776 3194
rect 28724 3130 28776 3136
rect 28828 2582 28856 4966
rect 29092 4616 29144 4622
rect 29092 4558 29144 4564
rect 29104 4282 29132 4558
rect 29196 4554 29224 5102
rect 29368 4820 29420 4826
rect 29368 4762 29420 4768
rect 29184 4548 29236 4554
rect 29184 4490 29236 4496
rect 29092 4276 29144 4282
rect 29092 4218 29144 4224
rect 29104 4154 29132 4218
rect 28920 4126 29132 4154
rect 29380 4146 29408 4762
rect 29656 4554 29684 6734
rect 29748 4826 29776 7142
rect 29840 6866 29868 10474
rect 30024 8498 30052 10474
rect 30564 9988 30616 9994
rect 30564 9930 30616 9936
rect 30104 9376 30156 9382
rect 30104 9318 30156 9324
rect 30116 8906 30144 9318
rect 30576 9110 30604 9930
rect 30656 9920 30708 9926
rect 30656 9862 30708 9868
rect 30668 9586 30696 9862
rect 30748 9716 30800 9722
rect 30748 9658 30800 9664
rect 30656 9580 30708 9586
rect 30656 9522 30708 9528
rect 30760 9450 30788 9658
rect 30932 9580 30984 9586
rect 30932 9522 30984 9528
rect 30748 9444 30800 9450
rect 30748 9386 30800 9392
rect 30564 9104 30616 9110
rect 30564 9046 30616 9052
rect 30104 8900 30156 8906
rect 30104 8842 30156 8848
rect 30576 8634 30604 9046
rect 30564 8628 30616 8634
rect 30564 8570 30616 8576
rect 30012 8492 30064 8498
rect 30012 8434 30064 8440
rect 30760 8430 30788 9386
rect 30840 9104 30892 9110
rect 30840 9046 30892 9052
rect 30852 8566 30880 9046
rect 30944 8974 30972 9522
rect 30932 8968 30984 8974
rect 30932 8910 30984 8916
rect 30840 8560 30892 8566
rect 30840 8502 30892 8508
rect 30748 8424 30800 8430
rect 30748 8366 30800 8372
rect 29920 8288 29972 8294
rect 29920 8230 29972 8236
rect 29932 8090 29960 8230
rect 30852 8090 30880 8502
rect 29920 8084 29972 8090
rect 29920 8026 29972 8032
rect 30656 8084 30708 8090
rect 30656 8026 30708 8032
rect 30840 8084 30892 8090
rect 30840 8026 30892 8032
rect 29920 7880 29972 7886
rect 29920 7822 29972 7828
rect 29932 7342 29960 7822
rect 30380 7812 30432 7818
rect 30380 7754 30432 7760
rect 29920 7336 29972 7342
rect 29920 7278 29972 7284
rect 29828 6860 29880 6866
rect 29828 6802 29880 6808
rect 29828 6112 29880 6118
rect 29828 6054 29880 6060
rect 29840 5914 29868 6054
rect 29828 5908 29880 5914
rect 29828 5850 29880 5856
rect 29840 5030 29868 5850
rect 29932 5234 29960 7278
rect 30196 6656 30248 6662
rect 30196 6598 30248 6604
rect 30208 6390 30236 6598
rect 30196 6384 30248 6390
rect 30196 6326 30248 6332
rect 29920 5228 29972 5234
rect 29920 5170 29972 5176
rect 29828 5024 29880 5030
rect 29828 4966 29880 4972
rect 29736 4820 29788 4826
rect 29736 4762 29788 4768
rect 29840 4758 29868 4966
rect 29828 4752 29880 4758
rect 29828 4694 29880 4700
rect 29644 4548 29696 4554
rect 29644 4490 29696 4496
rect 29368 4140 29420 4146
rect 28920 3670 28948 4126
rect 29368 4082 29420 4088
rect 29368 4004 29420 4010
rect 29368 3946 29420 3952
rect 29380 3738 29408 3946
rect 29368 3732 29420 3738
rect 29368 3674 29420 3680
rect 28908 3664 28960 3670
rect 28908 3606 28960 3612
rect 29656 3534 29684 4490
rect 29840 4282 29868 4694
rect 29828 4276 29880 4282
rect 29828 4218 29880 4224
rect 30392 4154 30420 7754
rect 30668 7206 30696 8026
rect 31404 7426 31432 12718
rect 34289 11996 34585 12016
rect 34345 11994 34369 11996
rect 34425 11994 34449 11996
rect 34505 11994 34529 11996
rect 34367 11942 34369 11994
rect 34431 11942 34443 11994
rect 34505 11942 34507 11994
rect 34345 11940 34369 11942
rect 34425 11940 34449 11942
rect 34505 11940 34529 11942
rect 34289 11920 34585 11940
rect 32588 11212 32640 11218
rect 32588 11154 32640 11160
rect 32680 11212 32732 11218
rect 32680 11154 32732 11160
rect 31576 11008 31628 11014
rect 31576 10950 31628 10956
rect 31668 11008 31720 11014
rect 31668 10950 31720 10956
rect 31484 10532 31536 10538
rect 31484 10474 31536 10480
rect 31496 9110 31524 10474
rect 31588 10198 31616 10950
rect 31680 10674 31708 10950
rect 32600 10810 32628 11154
rect 32588 10804 32640 10810
rect 32588 10746 32640 10752
rect 32692 10674 32720 11154
rect 34289 10908 34585 10928
rect 34345 10906 34369 10908
rect 34425 10906 34449 10908
rect 34505 10906 34529 10908
rect 34367 10854 34369 10906
rect 34431 10854 34443 10906
rect 34505 10854 34507 10906
rect 34345 10852 34369 10854
rect 34425 10852 34449 10854
rect 34505 10852 34529 10854
rect 34289 10832 34585 10852
rect 31668 10668 31720 10674
rect 31668 10610 31720 10616
rect 32680 10668 32732 10674
rect 32680 10610 32732 10616
rect 31680 10266 31708 10610
rect 32496 10532 32548 10538
rect 32496 10474 32548 10480
rect 31668 10260 31720 10266
rect 31668 10202 31720 10208
rect 31576 10192 31628 10198
rect 31576 10134 31628 10140
rect 32312 10192 32364 10198
rect 32312 10134 32364 10140
rect 31588 9178 31616 10134
rect 31760 10124 31812 10130
rect 31760 10066 31812 10072
rect 31772 9382 31800 10066
rect 32036 10056 32088 10062
rect 32036 9998 32088 10004
rect 31760 9376 31812 9382
rect 31760 9318 31812 9324
rect 31576 9172 31628 9178
rect 31576 9114 31628 9120
rect 31484 9104 31536 9110
rect 31484 9046 31536 9052
rect 31668 8492 31720 8498
rect 31668 8434 31720 8440
rect 31680 8090 31708 8434
rect 31668 8084 31720 8090
rect 31668 8026 31720 8032
rect 31772 7818 31800 9318
rect 32048 9042 32076 9998
rect 32324 9722 32352 10134
rect 32508 10062 32536 10474
rect 32496 10056 32548 10062
rect 32496 9998 32548 10004
rect 32312 9716 32364 9722
rect 32312 9658 32364 9664
rect 32508 9586 32536 9998
rect 32692 9586 32720 10610
rect 33508 10464 33560 10470
rect 33508 10406 33560 10412
rect 33520 10062 33548 10406
rect 33876 10192 33928 10198
rect 33876 10134 33928 10140
rect 33508 10056 33560 10062
rect 33508 9998 33560 10004
rect 33520 9654 33548 9998
rect 33888 9722 33916 10134
rect 34289 9820 34585 9840
rect 34345 9818 34369 9820
rect 34425 9818 34449 9820
rect 34505 9818 34529 9820
rect 34367 9766 34369 9818
rect 34431 9766 34443 9818
rect 34505 9766 34507 9818
rect 34345 9764 34369 9766
rect 34425 9764 34449 9766
rect 34505 9764 34529 9766
rect 34289 9744 34585 9764
rect 33876 9716 33928 9722
rect 33876 9658 33928 9664
rect 33508 9648 33560 9654
rect 33508 9590 33560 9596
rect 32496 9580 32548 9586
rect 32496 9522 32548 9528
rect 32680 9580 32732 9586
rect 32680 9522 32732 9528
rect 32692 9489 32720 9522
rect 32678 9480 32734 9489
rect 32678 9415 32734 9424
rect 33140 9376 33192 9382
rect 33140 9318 33192 9324
rect 33152 9178 33180 9318
rect 32496 9172 32548 9178
rect 32496 9114 32548 9120
rect 33140 9172 33192 9178
rect 33140 9114 33192 9120
rect 32036 9036 32088 9042
rect 32036 8978 32088 8984
rect 32508 8294 32536 9114
rect 34612 9104 34664 9110
rect 34150 9072 34206 9081
rect 33232 9036 33284 9042
rect 34612 9046 34664 9052
rect 34150 9007 34206 9016
rect 33232 8978 33284 8984
rect 33244 8634 33272 8978
rect 33232 8628 33284 8634
rect 33232 8570 33284 8576
rect 34164 8430 34192 9007
rect 34289 8732 34585 8752
rect 34345 8730 34369 8732
rect 34425 8730 34449 8732
rect 34505 8730 34529 8732
rect 34367 8678 34369 8730
rect 34431 8678 34443 8730
rect 34505 8678 34507 8730
rect 34345 8676 34369 8678
rect 34425 8676 34449 8678
rect 34505 8676 34529 8678
rect 34289 8656 34585 8676
rect 34624 8498 34652 9046
rect 34704 8968 34756 8974
rect 34704 8910 34756 8916
rect 34716 8634 34744 8910
rect 34704 8628 34756 8634
rect 34704 8570 34756 8576
rect 34612 8492 34664 8498
rect 34612 8434 34664 8440
rect 34152 8424 34204 8430
rect 34152 8366 34204 8372
rect 32496 8288 32548 8294
rect 32496 8230 32548 8236
rect 34152 8288 34204 8294
rect 34152 8230 34204 8236
rect 32508 8090 32536 8230
rect 32496 8084 32548 8090
rect 32496 8026 32548 8032
rect 31852 7948 31904 7954
rect 31852 7890 31904 7896
rect 31760 7812 31812 7818
rect 31760 7754 31812 7760
rect 31482 7440 31538 7449
rect 31404 7398 31482 7426
rect 31482 7375 31538 7384
rect 30656 7200 30708 7206
rect 30656 7142 30708 7148
rect 30668 7002 30696 7142
rect 30656 6996 30708 7002
rect 30656 6938 30708 6944
rect 30472 6656 30524 6662
rect 30472 6598 30524 6604
rect 30484 6322 30512 6598
rect 30472 6316 30524 6322
rect 30472 6258 30524 6264
rect 30668 6118 30696 6938
rect 31116 6860 31168 6866
rect 31116 6802 31168 6808
rect 30932 6316 30984 6322
rect 30932 6258 30984 6264
rect 30748 6180 30800 6186
rect 30748 6122 30800 6128
rect 30656 6112 30708 6118
rect 30656 6054 30708 6060
rect 30760 5778 30788 6122
rect 30748 5772 30800 5778
rect 30748 5714 30800 5720
rect 30944 5642 30972 6258
rect 31128 5914 31156 6802
rect 31116 5908 31168 5914
rect 31116 5850 31168 5856
rect 30932 5636 30984 5642
rect 30932 5578 30984 5584
rect 30944 5234 30972 5578
rect 30932 5228 30984 5234
rect 30932 5170 30984 5176
rect 30656 5160 30708 5166
rect 30656 5102 30708 5108
rect 30668 4826 30696 5102
rect 30656 4820 30708 4826
rect 30708 4780 30788 4808
rect 30656 4762 30708 4768
rect 30656 4684 30708 4690
rect 30656 4626 30708 4632
rect 30472 4480 30524 4486
rect 30472 4422 30524 4428
rect 30208 4126 30420 4154
rect 29644 3528 29696 3534
rect 29644 3470 29696 3476
rect 29276 2984 29328 2990
rect 29276 2926 29328 2932
rect 29920 2984 29972 2990
rect 29920 2926 29972 2932
rect 29288 2650 29316 2926
rect 29932 2650 29960 2926
rect 30208 2854 30236 4126
rect 30288 4072 30340 4078
rect 30288 4014 30340 4020
rect 30300 3602 30328 4014
rect 30484 3670 30512 4422
rect 30668 4214 30696 4626
rect 30656 4208 30708 4214
rect 30656 4150 30708 4156
rect 30668 4078 30696 4150
rect 30656 4072 30708 4078
rect 30656 4014 30708 4020
rect 30472 3664 30524 3670
rect 30472 3606 30524 3612
rect 30288 3596 30340 3602
rect 30288 3538 30340 3544
rect 30484 3194 30512 3606
rect 30472 3188 30524 3194
rect 30472 3130 30524 3136
rect 30760 3058 30788 4780
rect 31496 4078 31524 7375
rect 31760 7336 31812 7342
rect 31760 7278 31812 7284
rect 31772 6662 31800 7278
rect 31760 6656 31812 6662
rect 31760 6598 31812 6604
rect 31864 6322 31892 7890
rect 32128 7880 32180 7886
rect 32128 7822 32180 7828
rect 32140 7410 32168 7822
rect 32128 7404 32180 7410
rect 32128 7346 32180 7352
rect 32404 7336 32456 7342
rect 32404 7278 32456 7284
rect 31944 7268 31996 7274
rect 31944 7210 31996 7216
rect 31956 6866 31984 7210
rect 31944 6860 31996 6866
rect 31944 6802 31996 6808
rect 31956 6458 31984 6802
rect 31944 6452 31996 6458
rect 31944 6394 31996 6400
rect 31852 6316 31904 6322
rect 31852 6258 31904 6264
rect 31944 5840 31996 5846
rect 31944 5782 31996 5788
rect 31956 5370 31984 5782
rect 32416 5681 32444 7278
rect 32508 7274 32536 8026
rect 34164 8022 34192 8230
rect 34716 8090 34744 8570
rect 34704 8084 34756 8090
rect 34704 8026 34756 8032
rect 34152 8016 34204 8022
rect 34152 7958 34204 7964
rect 34520 8016 34572 8022
rect 34520 7958 34572 7964
rect 33692 7880 33744 7886
rect 33692 7822 33744 7828
rect 33704 7750 33732 7822
rect 33692 7744 33744 7750
rect 33692 7686 33744 7692
rect 33704 7546 33732 7686
rect 33692 7540 33744 7546
rect 33692 7482 33744 7488
rect 33968 7404 34020 7410
rect 33968 7346 34020 7352
rect 32496 7268 32548 7274
rect 32496 7210 32548 7216
rect 32508 6934 32536 7210
rect 32680 7200 32732 7206
rect 32680 7142 32732 7148
rect 32692 6934 32720 7142
rect 33980 7002 34008 7346
rect 34164 7002 34192 7958
rect 34532 7886 34560 7958
rect 34520 7880 34572 7886
rect 34520 7822 34572 7828
rect 34289 7644 34585 7664
rect 34345 7642 34369 7644
rect 34425 7642 34449 7644
rect 34505 7642 34529 7644
rect 34367 7590 34369 7642
rect 34431 7590 34443 7642
rect 34505 7590 34507 7642
rect 34345 7588 34369 7590
rect 34425 7588 34449 7590
rect 34505 7588 34529 7590
rect 34289 7568 34585 7588
rect 34808 7546 34836 12718
rect 35622 12608 35678 12617
rect 35622 12543 35678 12552
rect 35636 11898 35664 12543
rect 35624 11892 35676 11898
rect 35624 11834 35676 11840
rect 35440 11688 35492 11694
rect 35440 11630 35492 11636
rect 35452 10810 35480 11630
rect 37752 11354 37780 15558
rect 38106 15520 38162 15558
rect 39578 15464 39634 15473
rect 39578 15399 39634 15408
rect 39592 12714 39620 15399
rect 39580 12708 39632 12714
rect 39580 12650 39632 12656
rect 37740 11348 37792 11354
rect 37740 11290 37792 11296
rect 35440 10804 35492 10810
rect 35440 10746 35492 10752
rect 35256 10736 35308 10742
rect 35256 10678 35308 10684
rect 35268 10130 35296 10678
rect 35256 10124 35308 10130
rect 35256 10066 35308 10072
rect 34980 9920 35032 9926
rect 34980 9862 35032 9868
rect 34992 8498 35020 9862
rect 35268 9722 35296 10066
rect 35256 9716 35308 9722
rect 35256 9658 35308 9664
rect 35268 9518 35296 9658
rect 35256 9512 35308 9518
rect 35256 9454 35308 9460
rect 35452 8498 35480 10746
rect 35900 10600 35952 10606
rect 35900 10542 35952 10548
rect 35622 9752 35678 9761
rect 35622 9687 35678 9696
rect 35636 9654 35664 9687
rect 35624 9648 35676 9654
rect 35624 9590 35676 9596
rect 35912 9042 35940 10542
rect 37002 10296 37058 10305
rect 37002 10231 37058 10240
rect 37016 9081 37044 10231
rect 37002 9072 37058 9081
rect 35900 9036 35952 9042
rect 37002 9007 37058 9016
rect 35900 8978 35952 8984
rect 35912 8566 35940 8978
rect 36268 8968 36320 8974
rect 36268 8910 36320 8916
rect 35900 8560 35952 8566
rect 35900 8502 35952 8508
rect 34980 8492 35032 8498
rect 34980 8434 35032 8440
rect 35256 8492 35308 8498
rect 35256 8434 35308 8440
rect 35440 8492 35492 8498
rect 35440 8434 35492 8440
rect 34992 8090 35020 8434
rect 34980 8084 35032 8090
rect 34980 8026 35032 8032
rect 35268 8022 35296 8434
rect 35256 8016 35308 8022
rect 35256 7958 35308 7964
rect 34796 7540 34848 7546
rect 34796 7482 34848 7488
rect 35268 7410 35296 7958
rect 35912 7478 35940 8502
rect 35992 8288 36044 8294
rect 35992 8230 36044 8236
rect 36004 8022 36032 8230
rect 35992 8016 36044 8022
rect 35992 7958 36044 7964
rect 36084 8016 36136 8022
rect 36084 7958 36136 7964
rect 36004 7546 36032 7958
rect 36096 7886 36124 7958
rect 36280 7886 36308 8910
rect 36636 8900 36688 8906
rect 36636 8842 36688 8848
rect 36648 8430 36676 8842
rect 36636 8424 36688 8430
rect 36636 8366 36688 8372
rect 36084 7880 36136 7886
rect 36084 7822 36136 7828
rect 36268 7880 36320 7886
rect 36268 7822 36320 7828
rect 35992 7540 36044 7546
rect 35992 7482 36044 7488
rect 35900 7472 35952 7478
rect 35820 7432 35900 7460
rect 35072 7404 35124 7410
rect 35072 7346 35124 7352
rect 35256 7404 35308 7410
rect 35256 7346 35308 7352
rect 35084 7274 35112 7346
rect 34980 7268 35032 7274
rect 34980 7210 35032 7216
rect 35072 7268 35124 7274
rect 35072 7210 35124 7216
rect 34992 7002 35020 7210
rect 33968 6996 34020 7002
rect 33968 6938 34020 6944
rect 34152 6996 34204 7002
rect 34152 6938 34204 6944
rect 34980 6996 35032 7002
rect 34980 6938 35032 6944
rect 35084 6934 35112 7210
rect 32496 6928 32548 6934
rect 32496 6870 32548 6876
rect 32680 6928 32732 6934
rect 32680 6870 32732 6876
rect 34060 6928 34112 6934
rect 34060 6870 34112 6876
rect 35072 6928 35124 6934
rect 35072 6870 35124 6876
rect 34072 6458 34100 6870
rect 34888 6724 34940 6730
rect 34888 6666 34940 6672
rect 34612 6656 34664 6662
rect 34612 6598 34664 6604
rect 34289 6556 34585 6576
rect 34345 6554 34369 6556
rect 34425 6554 34449 6556
rect 34505 6554 34529 6556
rect 34367 6502 34369 6554
rect 34431 6502 34443 6554
rect 34505 6502 34507 6554
rect 34345 6500 34369 6502
rect 34425 6500 34449 6502
rect 34505 6500 34529 6502
rect 34289 6480 34585 6500
rect 34624 6458 34652 6598
rect 34060 6452 34112 6458
rect 34060 6394 34112 6400
rect 34612 6452 34664 6458
rect 34612 6394 34664 6400
rect 34624 6118 34652 6394
rect 33048 6112 33100 6118
rect 33048 6054 33100 6060
rect 34612 6112 34664 6118
rect 34612 6054 34664 6060
rect 33060 5846 33088 6054
rect 34900 5914 34928 6666
rect 35268 6322 35296 7346
rect 35348 6792 35400 6798
rect 35348 6734 35400 6740
rect 35360 6322 35388 6734
rect 35256 6316 35308 6322
rect 35256 6258 35308 6264
rect 35348 6316 35400 6322
rect 35348 6258 35400 6264
rect 35268 5914 35296 6258
rect 34888 5908 34940 5914
rect 34888 5850 34940 5856
rect 35256 5908 35308 5914
rect 35256 5850 35308 5856
rect 35360 5846 35388 6258
rect 33048 5840 33100 5846
rect 33048 5782 33100 5788
rect 33968 5840 34020 5846
rect 33968 5782 34020 5788
rect 35348 5840 35400 5846
rect 35348 5782 35400 5788
rect 33416 5704 33468 5710
rect 32402 5672 32458 5681
rect 33416 5646 33468 5652
rect 33876 5704 33928 5710
rect 33876 5646 33928 5652
rect 32402 5607 32458 5616
rect 32772 5636 32824 5642
rect 31944 5364 31996 5370
rect 31944 5306 31996 5312
rect 32312 5160 32364 5166
rect 32312 5102 32364 5108
rect 32324 5030 32352 5102
rect 32312 5024 32364 5030
rect 32312 4966 32364 4972
rect 32324 4758 32352 4966
rect 32312 4752 32364 4758
rect 32312 4694 32364 4700
rect 32324 4282 32352 4694
rect 32312 4276 32364 4282
rect 32312 4218 32364 4224
rect 31300 4072 31352 4078
rect 30930 4040 30986 4049
rect 31300 4014 31352 4020
rect 31484 4072 31536 4078
rect 31484 4014 31536 4020
rect 30930 3975 30986 3984
rect 30944 3942 30972 3975
rect 30932 3936 30984 3942
rect 30932 3878 30984 3884
rect 31312 3670 31340 4014
rect 31300 3664 31352 3670
rect 31300 3606 31352 3612
rect 30748 3052 30800 3058
rect 30748 2994 30800 3000
rect 31312 2990 31340 3606
rect 32416 3126 32444 5607
rect 32772 5578 32824 5584
rect 32496 5092 32548 5098
rect 32496 5034 32548 5040
rect 32508 4486 32536 5034
rect 32784 4554 32812 5578
rect 33428 5370 33456 5646
rect 33888 5370 33916 5646
rect 33980 5370 34008 5782
rect 34289 5468 34585 5488
rect 34345 5466 34369 5468
rect 34425 5466 34449 5468
rect 34505 5466 34529 5468
rect 34367 5414 34369 5466
rect 34431 5414 34443 5466
rect 34505 5414 34507 5466
rect 34345 5412 34369 5414
rect 34425 5412 34449 5414
rect 34505 5412 34529 5414
rect 34289 5392 34585 5412
rect 33416 5364 33468 5370
rect 33416 5306 33468 5312
rect 33876 5364 33928 5370
rect 33876 5306 33928 5312
rect 33968 5364 34020 5370
rect 33968 5306 34020 5312
rect 32864 4616 32916 4622
rect 32864 4558 32916 4564
rect 32772 4548 32824 4554
rect 32772 4490 32824 4496
rect 32496 4480 32548 4486
rect 32496 4422 32548 4428
rect 32508 3194 32536 4422
rect 32876 4282 32904 4558
rect 32864 4276 32916 4282
rect 32864 4218 32916 4224
rect 33428 4214 33456 5306
rect 35360 5166 35388 5782
rect 35348 5160 35400 5166
rect 35348 5102 35400 5108
rect 35820 4690 35848 7432
rect 35900 7414 35952 7420
rect 36096 7410 36124 7822
rect 36084 7404 36136 7410
rect 36084 7346 36136 7352
rect 36280 6934 36308 7822
rect 36452 7812 36504 7818
rect 36452 7754 36504 7760
rect 36464 7342 36492 7754
rect 36634 7712 36690 7721
rect 36634 7647 36690 7656
rect 36648 7546 36676 7647
rect 36636 7540 36688 7546
rect 36636 7482 36688 7488
rect 36452 7336 36504 7342
rect 36452 7278 36504 7284
rect 35900 6928 35952 6934
rect 35900 6870 35952 6876
rect 36268 6928 36320 6934
rect 36268 6870 36320 6876
rect 35912 6458 35940 6870
rect 36280 6730 36308 6870
rect 36360 6792 36412 6798
rect 36360 6734 36412 6740
rect 36268 6724 36320 6730
rect 36268 6666 36320 6672
rect 36372 6458 36400 6734
rect 37016 6458 37044 9007
rect 39580 8832 39632 8838
rect 39580 8774 39632 8780
rect 39592 8673 39620 8774
rect 39578 8664 39634 8673
rect 39578 8599 39634 8608
rect 38108 8288 38160 8294
rect 38108 8230 38160 8236
rect 37096 7200 37148 7206
rect 37096 7142 37148 7148
rect 37108 6798 37136 7142
rect 38120 6905 38148 8230
rect 38106 6896 38162 6905
rect 38106 6831 38162 6840
rect 37096 6792 37148 6798
rect 37096 6734 37148 6740
rect 35900 6452 35952 6458
rect 35900 6394 35952 6400
rect 36360 6452 36412 6458
rect 36360 6394 36412 6400
rect 37004 6452 37056 6458
rect 37004 6394 37056 6400
rect 37016 6254 37044 6394
rect 37004 6248 37056 6254
rect 37004 6190 37056 6196
rect 34152 4684 34204 4690
rect 34152 4626 34204 4632
rect 35348 4684 35400 4690
rect 35348 4626 35400 4632
rect 35808 4684 35860 4690
rect 35808 4626 35860 4632
rect 33968 4480 34020 4486
rect 33968 4422 34020 4428
rect 33980 4282 34008 4422
rect 33968 4276 34020 4282
rect 33968 4218 34020 4224
rect 33416 4208 33468 4214
rect 33416 4150 33468 4156
rect 34164 3942 34192 4626
rect 34289 4380 34585 4400
rect 34345 4378 34369 4380
rect 34425 4378 34449 4380
rect 34505 4378 34529 4380
rect 34367 4326 34369 4378
rect 34431 4326 34443 4378
rect 34505 4326 34507 4378
rect 34345 4324 34369 4326
rect 34425 4324 34449 4326
rect 34505 4324 34529 4326
rect 34289 4304 34585 4324
rect 35360 3942 35388 4626
rect 34152 3936 34204 3942
rect 34152 3878 34204 3884
rect 35348 3936 35400 3942
rect 35348 3878 35400 3884
rect 32680 3596 32732 3602
rect 32680 3538 32732 3544
rect 33232 3596 33284 3602
rect 33232 3538 33284 3544
rect 32692 3194 32720 3538
rect 33244 3194 33272 3538
rect 34164 3505 34192 3878
rect 34150 3496 34206 3505
rect 34150 3431 34206 3440
rect 34289 3292 34585 3312
rect 34345 3290 34369 3292
rect 34425 3290 34449 3292
rect 34505 3290 34529 3292
rect 34367 3238 34369 3290
rect 34431 3238 34443 3290
rect 34505 3238 34507 3290
rect 34345 3236 34369 3238
rect 34425 3236 34449 3238
rect 34505 3236 34529 3238
rect 34289 3216 34585 3236
rect 32496 3188 32548 3194
rect 32496 3130 32548 3136
rect 32680 3188 32732 3194
rect 32680 3130 32732 3136
rect 33232 3188 33284 3194
rect 33232 3130 33284 3136
rect 32404 3120 32456 3126
rect 32404 3062 32456 3068
rect 31300 2984 31352 2990
rect 31300 2926 31352 2932
rect 30196 2848 30248 2854
rect 30196 2790 30248 2796
rect 30208 2650 30236 2790
rect 29276 2644 29328 2650
rect 29276 2586 29328 2592
rect 29920 2644 29972 2650
rect 29920 2586 29972 2592
rect 30196 2644 30248 2650
rect 30196 2586 30248 2592
rect 32404 2644 32456 2650
rect 32404 2586 32456 2592
rect 28816 2576 28868 2582
rect 28816 2518 28868 2524
rect 26792 2372 26844 2378
rect 26792 2314 26844 2320
rect 28448 2372 28500 2378
rect 28448 2314 28500 2320
rect 28540 2372 28592 2378
rect 28540 2314 28592 2320
rect 25410 1864 25466 1873
rect 25410 1799 25466 1808
rect 24136 54 24270 82
rect 24492 128 24544 134
rect 24492 70 24544 76
rect 26804 82 26832 2314
rect 27252 2304 27304 2310
rect 27252 2246 27304 2252
rect 27264 1329 27292 2246
rect 29642 1456 29698 1465
rect 29642 1391 29698 1400
rect 27250 1320 27306 1329
rect 27250 1255 27306 1264
rect 27066 82 27122 480
rect 26804 54 27122 82
rect 29656 82 29684 1391
rect 29918 82 29974 480
rect 29656 54 29974 82
rect 32416 82 32444 2586
rect 34289 2204 34585 2224
rect 34345 2202 34369 2204
rect 34425 2202 34449 2204
rect 34505 2202 34529 2204
rect 34367 2150 34369 2202
rect 34431 2150 34443 2202
rect 34505 2150 34507 2202
rect 34345 2148 34369 2150
rect 34425 2148 34449 2150
rect 34505 2148 34529 2150
rect 34289 2128 34585 2148
rect 32770 82 32826 480
rect 32416 54 32826 82
rect 35360 82 35388 3878
rect 38120 3602 38148 6831
rect 39580 5092 39632 5098
rect 39580 5034 39632 5040
rect 39592 4049 39620 5034
rect 39578 4040 39634 4049
rect 39578 3975 39634 3984
rect 38108 3596 38160 3602
rect 38108 3538 38160 3544
rect 39580 3460 39632 3466
rect 39580 3402 39632 3408
rect 39592 2825 39620 3402
rect 39578 2816 39634 2825
rect 39578 2751 39634 2760
rect 38566 1320 38622 1329
rect 38566 1255 38622 1264
rect 35622 82 35678 480
rect 35360 54 35678 82
rect 24214 0 24270 54
rect 27066 0 27122 54
rect 29918 0 29974 54
rect 32770 0 32826 54
rect 35622 0 35678 54
rect 38474 82 38530 480
rect 38580 82 38608 1255
rect 38474 54 38608 82
rect 38474 0 38530 54
<< via2 >>
rect 1122 15000 1178 15056
rect 110 13640 166 13696
rect 1582 12416 1638 12472
rect 110 11736 166 11792
rect 1398 10240 1454 10296
rect 110 9832 166 9888
rect 110 8880 166 8936
rect 18 7928 74 7984
rect 1766 10648 1822 10704
rect 1490 5752 1546 5808
rect 1950 14184 2006 14240
rect 2042 11600 2098 11656
rect 1950 9560 2006 9616
rect 2962 10240 3018 10296
rect 1674 4936 1730 4992
rect 2778 6704 2834 6760
rect 4526 10240 4582 10296
rect 2962 5616 3018 5672
rect 3698 9152 3754 9208
rect 3606 6704 3662 6760
rect 3974 7384 4030 7440
rect 110 3168 166 3224
rect 110 2216 166 2272
rect 2502 1672 2558 1728
rect 7622 13082 7678 13084
rect 7702 13082 7758 13084
rect 7782 13082 7838 13084
rect 7862 13082 7918 13084
rect 7622 13030 7648 13082
rect 7648 13030 7678 13082
rect 7702 13030 7712 13082
rect 7712 13030 7758 13082
rect 7782 13030 7828 13082
rect 7828 13030 7838 13082
rect 7862 13030 7892 13082
rect 7892 13030 7918 13082
rect 7622 13028 7678 13030
rect 7702 13028 7758 13030
rect 7782 13028 7838 13030
rect 7862 13028 7918 13030
rect 5630 11736 5686 11792
rect 7622 11994 7678 11996
rect 7702 11994 7758 11996
rect 7782 11994 7838 11996
rect 7862 11994 7918 11996
rect 7622 11942 7648 11994
rect 7648 11942 7678 11994
rect 7702 11942 7712 11994
rect 7712 11942 7758 11994
rect 7782 11942 7828 11994
rect 7828 11942 7838 11994
rect 7862 11942 7892 11994
rect 7892 11942 7918 11994
rect 7622 11940 7678 11942
rect 7702 11940 7758 11942
rect 7782 11940 7838 11942
rect 7862 11940 7918 11942
rect 5078 5208 5134 5264
rect 5446 5616 5502 5672
rect 5998 9716 6054 9752
rect 5998 9696 6000 9716
rect 6000 9696 6052 9716
rect 6052 9696 6054 9716
rect 6366 9424 6422 9480
rect 7622 10906 7678 10908
rect 7702 10906 7758 10908
rect 7782 10906 7838 10908
rect 7862 10906 7918 10908
rect 7622 10854 7648 10906
rect 7648 10854 7678 10906
rect 7702 10854 7712 10906
rect 7712 10854 7758 10906
rect 7782 10854 7828 10906
rect 7828 10854 7838 10906
rect 7862 10854 7892 10906
rect 7892 10854 7918 10906
rect 7622 10852 7678 10854
rect 7702 10852 7758 10854
rect 7782 10852 7838 10854
rect 7862 10852 7918 10854
rect 7622 9818 7678 9820
rect 7702 9818 7758 9820
rect 7782 9818 7838 9820
rect 7862 9818 7918 9820
rect 7622 9766 7648 9818
rect 7648 9766 7678 9818
rect 7702 9766 7712 9818
rect 7712 9766 7758 9818
rect 7782 9766 7828 9818
rect 7828 9766 7838 9818
rect 7862 9766 7892 9818
rect 7892 9766 7918 9818
rect 7622 9764 7678 9766
rect 7702 9764 7758 9766
rect 7782 9764 7838 9766
rect 7862 9764 7918 9766
rect 7622 8730 7678 8732
rect 7702 8730 7758 8732
rect 7782 8730 7838 8732
rect 7862 8730 7918 8732
rect 7622 8678 7648 8730
rect 7648 8678 7678 8730
rect 7702 8678 7712 8730
rect 7712 8678 7758 8730
rect 7782 8678 7828 8730
rect 7828 8678 7838 8730
rect 7862 8678 7892 8730
rect 7892 8678 7918 8730
rect 7622 8676 7678 8678
rect 7702 8676 7758 8678
rect 7782 8676 7838 8678
rect 7862 8676 7918 8678
rect 7102 7928 7158 7984
rect 5906 4120 5962 4176
rect 7622 7642 7678 7644
rect 7702 7642 7758 7644
rect 7782 7642 7838 7644
rect 7862 7642 7918 7644
rect 7622 7590 7648 7642
rect 7648 7590 7678 7642
rect 7702 7590 7712 7642
rect 7712 7590 7758 7642
rect 7782 7590 7828 7642
rect 7828 7590 7838 7642
rect 7862 7590 7892 7642
rect 7892 7590 7918 7642
rect 7622 7588 7678 7590
rect 7702 7588 7758 7590
rect 7782 7588 7838 7590
rect 7862 7588 7918 7590
rect 8114 9036 8170 9072
rect 8114 9016 8116 9036
rect 8116 9016 8168 9036
rect 8168 9016 8170 9036
rect 7622 6554 7678 6556
rect 7702 6554 7758 6556
rect 7782 6554 7838 6556
rect 7862 6554 7918 6556
rect 7622 6502 7648 6554
rect 7648 6502 7678 6554
rect 7702 6502 7712 6554
rect 7712 6502 7758 6554
rect 7782 6502 7828 6554
rect 7828 6502 7838 6554
rect 7862 6502 7892 6554
rect 7892 6502 7918 6554
rect 7622 6500 7678 6502
rect 7702 6500 7758 6502
rect 7782 6500 7838 6502
rect 7862 6500 7918 6502
rect 7622 5466 7678 5468
rect 7702 5466 7758 5468
rect 7782 5466 7838 5468
rect 7862 5466 7918 5468
rect 7622 5414 7648 5466
rect 7648 5414 7678 5466
rect 7702 5414 7712 5466
rect 7712 5414 7758 5466
rect 7782 5414 7828 5466
rect 7828 5414 7838 5466
rect 7862 5414 7892 5466
rect 7892 5414 7918 5466
rect 7622 5412 7678 5414
rect 7702 5412 7758 5414
rect 7782 5412 7838 5414
rect 7862 5412 7918 5414
rect 8574 5752 8630 5808
rect 9126 10512 9182 10568
rect 9310 9152 9366 9208
rect 7622 4378 7678 4380
rect 7702 4378 7758 4380
rect 7782 4378 7838 4380
rect 7862 4378 7918 4380
rect 7622 4326 7648 4378
rect 7648 4326 7678 4378
rect 7702 4326 7712 4378
rect 7712 4326 7758 4378
rect 7782 4326 7828 4378
rect 7828 4326 7838 4378
rect 7862 4326 7892 4378
rect 7892 4326 7918 4378
rect 7622 4324 7678 4326
rect 7702 4324 7758 4326
rect 7782 4324 7838 4326
rect 7862 4324 7918 4326
rect 9126 4664 9182 4720
rect 8482 4020 8484 4040
rect 8484 4020 8536 4040
rect 8536 4020 8538 4040
rect 8482 3984 8538 4020
rect 7622 3290 7678 3292
rect 7702 3290 7758 3292
rect 7782 3290 7838 3292
rect 7862 3290 7918 3292
rect 7622 3238 7648 3290
rect 7648 3238 7678 3290
rect 7702 3238 7712 3290
rect 7712 3238 7758 3290
rect 7782 3238 7828 3290
rect 7828 3238 7838 3290
rect 7862 3238 7892 3290
rect 7892 3238 7918 3290
rect 7622 3236 7678 3238
rect 7702 3236 7758 3238
rect 7782 3236 7838 3238
rect 7862 3236 7918 3238
rect 6274 1536 6330 1592
rect 7622 2202 7678 2204
rect 7702 2202 7758 2204
rect 7782 2202 7838 2204
rect 7862 2202 7918 2204
rect 7622 2150 7648 2202
rect 7648 2150 7678 2202
rect 7702 2150 7712 2202
rect 7712 2150 7758 2202
rect 7782 2150 7828 2202
rect 7828 2150 7838 2202
rect 7862 2150 7892 2202
rect 7892 2150 7918 2202
rect 7622 2148 7678 2150
rect 7702 2148 7758 2150
rect 7782 2148 7838 2150
rect 7862 2148 7918 2150
rect 14289 13626 14345 13628
rect 14369 13626 14425 13628
rect 14449 13626 14505 13628
rect 14529 13626 14585 13628
rect 14289 13574 14315 13626
rect 14315 13574 14345 13626
rect 14369 13574 14379 13626
rect 14379 13574 14425 13626
rect 14449 13574 14495 13626
rect 14495 13574 14505 13626
rect 14529 13574 14559 13626
rect 14559 13574 14585 13626
rect 14289 13572 14345 13574
rect 14369 13572 14425 13574
rect 14449 13572 14505 13574
rect 14529 13572 14585 13574
rect 12530 11600 12586 11656
rect 11886 10684 11888 10704
rect 11888 10684 11940 10704
rect 11940 10684 11942 10704
rect 11886 10648 11942 10684
rect 11794 9560 11850 9616
rect 12346 9424 12402 9480
rect 12254 8336 12310 8392
rect 10874 7792 10930 7848
rect 10782 7384 10838 7440
rect 11978 5752 12034 5808
rect 10230 4664 10286 4720
rect 9954 4528 10010 4584
rect 9034 1944 9090 2000
rect 8482 1536 8538 1592
rect 6642 992 6698 1048
rect 9310 1672 9366 1728
rect 9218 1264 9274 1320
rect 12070 4664 12126 4720
rect 14289 12538 14345 12540
rect 14369 12538 14425 12540
rect 14449 12538 14505 12540
rect 14529 12538 14585 12540
rect 14289 12486 14315 12538
rect 14315 12486 14345 12538
rect 14369 12486 14379 12538
rect 14379 12486 14425 12538
rect 14449 12486 14495 12538
rect 14495 12486 14505 12538
rect 14529 12486 14559 12538
rect 14559 12486 14585 12538
rect 14289 12484 14345 12486
rect 14369 12484 14425 12486
rect 14449 12484 14505 12486
rect 14529 12484 14585 12486
rect 13450 9560 13506 9616
rect 13910 8880 13966 8936
rect 14289 11450 14345 11452
rect 14369 11450 14425 11452
rect 14449 11450 14505 11452
rect 14529 11450 14585 11452
rect 14289 11398 14315 11450
rect 14315 11398 14345 11450
rect 14369 11398 14379 11450
rect 14379 11398 14425 11450
rect 14449 11398 14495 11450
rect 14495 11398 14505 11450
rect 14529 11398 14559 11450
rect 14559 11398 14585 11450
rect 14289 11396 14345 11398
rect 14369 11396 14425 11398
rect 14449 11396 14505 11398
rect 14529 11396 14585 11398
rect 14289 10362 14345 10364
rect 14369 10362 14425 10364
rect 14449 10362 14505 10364
rect 14529 10362 14585 10364
rect 14289 10310 14315 10362
rect 14315 10310 14345 10362
rect 14369 10310 14379 10362
rect 14379 10310 14425 10362
rect 14449 10310 14495 10362
rect 14495 10310 14505 10362
rect 14529 10310 14559 10362
rect 14559 10310 14585 10362
rect 14289 10308 14345 10310
rect 14369 10308 14425 10310
rect 14449 10308 14505 10310
rect 14529 10308 14585 10310
rect 14738 10104 14794 10160
rect 14289 9274 14345 9276
rect 14369 9274 14425 9276
rect 14449 9274 14505 9276
rect 14529 9274 14585 9276
rect 14289 9222 14315 9274
rect 14315 9222 14345 9274
rect 14369 9222 14379 9274
rect 14379 9222 14425 9274
rect 14449 9222 14495 9274
rect 14495 9222 14505 9274
rect 14529 9222 14559 9274
rect 14559 9222 14585 9274
rect 14289 9220 14345 9222
rect 14369 9220 14425 9222
rect 14449 9220 14505 9222
rect 14529 9220 14585 9222
rect 14289 8186 14345 8188
rect 14369 8186 14425 8188
rect 14449 8186 14505 8188
rect 14529 8186 14585 8188
rect 14289 8134 14315 8186
rect 14315 8134 14345 8186
rect 14369 8134 14379 8186
rect 14379 8134 14425 8186
rect 14449 8134 14495 8186
rect 14495 8134 14505 8186
rect 14529 8134 14559 8186
rect 14559 8134 14585 8186
rect 14289 8132 14345 8134
rect 14369 8132 14425 8134
rect 14449 8132 14505 8134
rect 14529 8132 14585 8134
rect 14289 7098 14345 7100
rect 14369 7098 14425 7100
rect 14449 7098 14505 7100
rect 14529 7098 14585 7100
rect 14289 7046 14315 7098
rect 14315 7046 14345 7098
rect 14369 7046 14379 7098
rect 14379 7046 14425 7098
rect 14449 7046 14495 7098
rect 14495 7046 14505 7098
rect 14529 7046 14559 7098
rect 14559 7046 14585 7098
rect 14289 7044 14345 7046
rect 14369 7044 14425 7046
rect 14449 7044 14505 7046
rect 14529 7044 14585 7046
rect 15198 10240 15254 10296
rect 13910 5616 13966 5672
rect 13910 4936 13966 4992
rect 14289 6010 14345 6012
rect 14369 6010 14425 6012
rect 14449 6010 14505 6012
rect 14529 6010 14585 6012
rect 14289 5958 14315 6010
rect 14315 5958 14345 6010
rect 14369 5958 14379 6010
rect 14379 5958 14425 6010
rect 14449 5958 14495 6010
rect 14495 5958 14505 6010
rect 14529 5958 14559 6010
rect 14559 5958 14585 6010
rect 14289 5956 14345 5958
rect 14369 5956 14425 5958
rect 14449 5956 14505 5958
rect 14529 5956 14585 5958
rect 14646 5480 14702 5536
rect 15290 7384 15346 7440
rect 14289 4922 14345 4924
rect 14369 4922 14425 4924
rect 14449 4922 14505 4924
rect 14529 4922 14585 4924
rect 14289 4870 14315 4922
rect 14315 4870 14345 4922
rect 14369 4870 14379 4922
rect 14379 4870 14425 4922
rect 14449 4870 14495 4922
rect 14495 4870 14505 4922
rect 14529 4870 14559 4922
rect 14559 4870 14585 4922
rect 14289 4868 14345 4870
rect 14369 4868 14425 4870
rect 14449 4868 14505 4870
rect 14529 4868 14585 4870
rect 13082 3984 13138 4040
rect 15014 4120 15070 4176
rect 14289 3834 14345 3836
rect 14369 3834 14425 3836
rect 14449 3834 14505 3836
rect 14529 3834 14585 3836
rect 14289 3782 14315 3834
rect 14315 3782 14345 3834
rect 14369 3782 14379 3834
rect 14379 3782 14425 3834
rect 14449 3782 14495 3834
rect 14495 3782 14505 3834
rect 14529 3782 14559 3834
rect 14559 3782 14585 3834
rect 14289 3780 14345 3782
rect 14369 3780 14425 3782
rect 14449 3780 14505 3782
rect 14529 3780 14585 3782
rect 14289 2746 14345 2748
rect 14369 2746 14425 2748
rect 14449 2746 14505 2748
rect 14529 2746 14585 2748
rect 14289 2694 14315 2746
rect 14315 2694 14345 2746
rect 14369 2694 14379 2746
rect 14379 2694 14425 2746
rect 14449 2694 14495 2746
rect 14495 2694 14505 2746
rect 14529 2694 14559 2746
rect 14559 2694 14585 2746
rect 14289 2692 14345 2694
rect 14369 2692 14425 2694
rect 14449 2692 14505 2694
rect 14529 2692 14585 2694
rect 15198 1944 15254 2000
rect 15106 1536 15162 1592
rect 15934 9560 15990 9616
rect 15934 8472 15990 8528
rect 20956 13082 21012 13084
rect 21036 13082 21092 13084
rect 21116 13082 21172 13084
rect 21196 13082 21252 13084
rect 20956 13030 20982 13082
rect 20982 13030 21012 13082
rect 21036 13030 21046 13082
rect 21046 13030 21092 13082
rect 21116 13030 21162 13082
rect 21162 13030 21172 13082
rect 21196 13030 21226 13082
rect 21226 13030 21252 13082
rect 20956 13028 21012 13030
rect 21036 13028 21092 13030
rect 21116 13028 21172 13030
rect 21196 13028 21252 13030
rect 16486 7928 16542 7984
rect 17590 11736 17646 11792
rect 18234 10240 18290 10296
rect 19062 11600 19118 11656
rect 18694 9424 18750 9480
rect 18050 6704 18106 6760
rect 17406 5208 17462 5264
rect 16486 4120 16542 4176
rect 18878 9152 18934 9208
rect 19246 9152 19302 9208
rect 19246 5616 19302 5672
rect 15750 2080 15806 2136
rect 19522 3440 19578 3496
rect 20956 11994 21012 11996
rect 21036 11994 21092 11996
rect 21116 11994 21172 11996
rect 21196 11994 21252 11996
rect 20956 11942 20982 11994
rect 20982 11942 21012 11994
rect 21036 11942 21046 11994
rect 21046 11942 21092 11994
rect 21116 11942 21162 11994
rect 21162 11942 21172 11994
rect 21196 11942 21226 11994
rect 21226 11942 21252 11994
rect 20956 11940 21012 11942
rect 21036 11940 21092 11942
rect 21116 11940 21172 11942
rect 21196 11940 21252 11942
rect 19890 8336 19946 8392
rect 20956 10906 21012 10908
rect 21036 10906 21092 10908
rect 21116 10906 21172 10908
rect 21196 10906 21252 10908
rect 20956 10854 20982 10906
rect 20982 10854 21012 10906
rect 21036 10854 21046 10906
rect 21046 10854 21092 10906
rect 21116 10854 21162 10906
rect 21162 10854 21172 10906
rect 21196 10854 21226 10906
rect 21226 10854 21252 10906
rect 20956 10852 21012 10854
rect 21036 10852 21092 10854
rect 21116 10852 21172 10854
rect 21196 10852 21252 10854
rect 20956 9818 21012 9820
rect 21036 9818 21092 9820
rect 21116 9818 21172 9820
rect 21196 9818 21252 9820
rect 20956 9766 20982 9818
rect 20982 9766 21012 9818
rect 21036 9766 21046 9818
rect 21046 9766 21092 9818
rect 21116 9766 21162 9818
rect 21162 9766 21172 9818
rect 21196 9766 21226 9818
rect 21226 9766 21252 9818
rect 20956 9764 21012 9766
rect 21036 9764 21092 9766
rect 21116 9764 21172 9766
rect 21196 9764 21252 9766
rect 21914 9424 21970 9480
rect 20956 8730 21012 8732
rect 21036 8730 21092 8732
rect 21116 8730 21172 8732
rect 21196 8730 21252 8732
rect 20956 8678 20982 8730
rect 20982 8678 21012 8730
rect 21036 8678 21046 8730
rect 21046 8678 21092 8730
rect 21116 8678 21162 8730
rect 21162 8678 21172 8730
rect 21196 8678 21226 8730
rect 21226 8678 21252 8730
rect 20956 8676 21012 8678
rect 21036 8676 21092 8678
rect 21116 8676 21172 8678
rect 21196 8676 21252 8678
rect 20956 7642 21012 7644
rect 21036 7642 21092 7644
rect 21116 7642 21172 7644
rect 21196 7642 21252 7644
rect 20956 7590 20982 7642
rect 20982 7590 21012 7642
rect 21036 7590 21046 7642
rect 21046 7590 21092 7642
rect 21116 7590 21162 7642
rect 21162 7590 21172 7642
rect 21196 7590 21226 7642
rect 21226 7590 21252 7642
rect 20956 7588 21012 7590
rect 21036 7588 21092 7590
rect 21116 7588 21172 7590
rect 21196 7588 21252 7590
rect 21178 7248 21234 7304
rect 20956 6554 21012 6556
rect 21036 6554 21092 6556
rect 21116 6554 21172 6556
rect 21196 6554 21252 6556
rect 20956 6502 20982 6554
rect 20982 6502 21012 6554
rect 21036 6502 21046 6554
rect 21046 6502 21092 6554
rect 21116 6502 21162 6554
rect 21162 6502 21172 6554
rect 21196 6502 21226 6554
rect 21226 6502 21252 6554
rect 20956 6500 21012 6502
rect 21036 6500 21092 6502
rect 21116 6500 21172 6502
rect 21196 6500 21252 6502
rect 20166 6296 20222 6352
rect 20956 5466 21012 5468
rect 21036 5466 21092 5468
rect 21116 5466 21172 5468
rect 21196 5466 21252 5468
rect 20956 5414 20982 5466
rect 20982 5414 21012 5466
rect 21036 5414 21046 5466
rect 21046 5414 21092 5466
rect 21116 5414 21162 5466
rect 21162 5414 21172 5466
rect 21196 5414 21226 5466
rect 21226 5414 21252 5466
rect 20956 5412 21012 5414
rect 21036 5412 21092 5414
rect 21116 5412 21172 5414
rect 21196 5412 21252 5414
rect 20956 4378 21012 4380
rect 21036 4378 21092 4380
rect 21116 4378 21172 4380
rect 21196 4378 21252 4380
rect 20956 4326 20982 4378
rect 20982 4326 21012 4378
rect 21036 4326 21046 4378
rect 21046 4326 21092 4378
rect 21116 4326 21162 4378
rect 21162 4326 21172 4378
rect 21196 4326 21226 4378
rect 21226 4326 21252 4378
rect 20956 4324 21012 4326
rect 21036 4324 21092 4326
rect 21116 4324 21172 4326
rect 21196 4324 21252 4326
rect 20956 3290 21012 3292
rect 21036 3290 21092 3292
rect 21116 3290 21172 3292
rect 21196 3290 21252 3292
rect 20956 3238 20982 3290
rect 20982 3238 21012 3290
rect 21036 3238 21046 3290
rect 21046 3238 21092 3290
rect 21116 3238 21162 3290
rect 21162 3238 21172 3290
rect 21196 3238 21226 3290
rect 21226 3238 21252 3290
rect 20956 3236 21012 3238
rect 21036 3236 21092 3238
rect 21116 3236 21172 3238
rect 21196 3236 21252 3238
rect 18418 2352 18474 2408
rect 17774 1672 17830 1728
rect 16946 1264 17002 1320
rect 20956 2202 21012 2204
rect 21036 2202 21092 2204
rect 21116 2202 21172 2204
rect 21196 2202 21252 2204
rect 20956 2150 20982 2202
rect 20982 2150 21012 2202
rect 21036 2150 21046 2202
rect 21046 2150 21092 2202
rect 21116 2150 21162 2202
rect 21162 2150 21172 2202
rect 21196 2150 21226 2202
rect 21226 2150 21252 2202
rect 20956 2148 21012 2150
rect 21036 2148 21092 2150
rect 21116 2148 21172 2150
rect 21196 2148 21252 2150
rect 18786 1808 18842 1864
rect 18326 176 18382 232
rect 23202 9560 23258 9616
rect 23570 10376 23626 10432
rect 24306 10240 24362 10296
rect 23754 8880 23810 8936
rect 24122 7792 24178 7848
rect 24490 11600 24546 11656
rect 24490 9580 24546 9616
rect 24490 9560 24492 9580
rect 24492 9560 24544 9580
rect 24544 9560 24546 9580
rect 24582 9424 24638 9480
rect 24122 5616 24178 5672
rect 21822 1400 21878 1456
rect 27622 13626 27678 13628
rect 27702 13626 27758 13628
rect 27782 13626 27838 13628
rect 27862 13626 27918 13628
rect 27622 13574 27648 13626
rect 27648 13574 27678 13626
rect 27702 13574 27712 13626
rect 27712 13574 27758 13626
rect 27782 13574 27828 13626
rect 27828 13574 27838 13626
rect 27862 13574 27892 13626
rect 27892 13574 27918 13626
rect 27622 13572 27678 13574
rect 27702 13572 27758 13574
rect 27782 13572 27838 13574
rect 27862 13572 27918 13574
rect 27622 12538 27678 12540
rect 27702 12538 27758 12540
rect 27782 12538 27838 12540
rect 27862 12538 27918 12540
rect 27622 12486 27648 12538
rect 27648 12486 27678 12538
rect 27702 12486 27712 12538
rect 27712 12486 27758 12538
rect 27782 12486 27828 12538
rect 27828 12486 27838 12538
rect 27862 12486 27892 12538
rect 27892 12486 27918 12538
rect 27622 12484 27678 12486
rect 27702 12484 27758 12486
rect 27782 12484 27838 12486
rect 27862 12484 27918 12486
rect 24766 5772 24822 5808
rect 24766 5752 24768 5772
rect 24768 5752 24820 5772
rect 24820 5752 24822 5772
rect 24858 5072 24914 5128
rect 24582 4120 24638 4176
rect 25594 10376 25650 10432
rect 25502 10104 25558 10160
rect 25502 7248 25558 7304
rect 26238 8472 26294 8528
rect 27622 11450 27678 11452
rect 27702 11450 27758 11452
rect 27782 11450 27838 11452
rect 27862 11450 27918 11452
rect 27622 11398 27648 11450
rect 27648 11398 27678 11450
rect 27702 11398 27712 11450
rect 27712 11398 27758 11450
rect 27782 11398 27828 11450
rect 27828 11398 27838 11450
rect 27862 11398 27892 11450
rect 27892 11398 27918 11450
rect 27622 11396 27678 11398
rect 27702 11396 27758 11398
rect 27782 11396 27838 11398
rect 27862 11396 27918 11398
rect 27622 10362 27678 10364
rect 27702 10362 27758 10364
rect 27782 10362 27838 10364
rect 27862 10362 27918 10364
rect 27622 10310 27648 10362
rect 27648 10310 27678 10362
rect 27702 10310 27712 10362
rect 27712 10310 27758 10362
rect 27782 10310 27828 10362
rect 27828 10310 27838 10362
rect 27862 10310 27892 10362
rect 27892 10310 27918 10362
rect 27622 10308 27678 10310
rect 27702 10308 27758 10310
rect 27782 10308 27838 10310
rect 27862 10308 27918 10310
rect 27622 9274 27678 9276
rect 27702 9274 27758 9276
rect 27782 9274 27838 9276
rect 27862 9274 27918 9276
rect 27622 9222 27648 9274
rect 27648 9222 27678 9274
rect 27702 9222 27712 9274
rect 27712 9222 27758 9274
rect 27782 9222 27828 9274
rect 27828 9222 27838 9274
rect 27862 9222 27892 9274
rect 27892 9222 27918 9274
rect 27622 9220 27678 9222
rect 27702 9220 27758 9222
rect 27782 9220 27838 9222
rect 27862 9220 27918 9222
rect 26790 9152 26846 9208
rect 27622 8186 27678 8188
rect 27702 8186 27758 8188
rect 27782 8186 27838 8188
rect 27862 8186 27918 8188
rect 27622 8134 27648 8186
rect 27648 8134 27678 8186
rect 27702 8134 27712 8186
rect 27712 8134 27758 8186
rect 27782 8134 27828 8186
rect 27828 8134 27838 8186
rect 27862 8134 27892 8186
rect 27892 8134 27918 8186
rect 27622 8132 27678 8134
rect 27702 8132 27758 8134
rect 27782 8132 27838 8134
rect 27862 8132 27918 8134
rect 27622 7098 27678 7100
rect 27702 7098 27758 7100
rect 27782 7098 27838 7100
rect 27862 7098 27918 7100
rect 27622 7046 27648 7098
rect 27648 7046 27678 7098
rect 27702 7046 27712 7098
rect 27712 7046 27758 7098
rect 27782 7046 27828 7098
rect 27828 7046 27838 7098
rect 27862 7046 27892 7098
rect 27892 7046 27918 7098
rect 27622 7044 27678 7046
rect 27702 7044 27758 7046
rect 27782 7044 27838 7046
rect 27862 7044 27918 7046
rect 27342 6296 27398 6352
rect 25870 3984 25926 4040
rect 27622 6010 27678 6012
rect 27702 6010 27758 6012
rect 27782 6010 27838 6012
rect 27862 6010 27918 6012
rect 27622 5958 27648 6010
rect 27648 5958 27678 6010
rect 27702 5958 27712 6010
rect 27712 5958 27758 6010
rect 27782 5958 27828 6010
rect 27828 5958 27838 6010
rect 27862 5958 27892 6010
rect 27892 5958 27918 6010
rect 27622 5956 27678 5958
rect 27702 5956 27758 5958
rect 27782 5956 27838 5958
rect 27862 5956 27918 5958
rect 27622 4922 27678 4924
rect 27702 4922 27758 4924
rect 27782 4922 27838 4924
rect 27862 4922 27918 4924
rect 27622 4870 27648 4922
rect 27648 4870 27678 4922
rect 27702 4870 27712 4922
rect 27712 4870 27758 4922
rect 27782 4870 27828 4922
rect 27828 4870 27838 4922
rect 27862 4870 27892 4922
rect 27892 4870 27918 4922
rect 27622 4868 27678 4870
rect 27702 4868 27758 4870
rect 27782 4868 27838 4870
rect 27862 4868 27918 4870
rect 35622 14048 35678 14104
rect 34289 13082 34345 13084
rect 34369 13082 34425 13084
rect 34449 13082 34505 13084
rect 34529 13082 34585 13084
rect 34289 13030 34315 13082
rect 34315 13030 34345 13082
rect 34369 13030 34379 13082
rect 34379 13030 34425 13082
rect 34449 13030 34495 13082
rect 34495 13030 34505 13082
rect 34529 13030 34559 13082
rect 34559 13030 34585 13082
rect 34289 13028 34345 13030
rect 34369 13028 34425 13030
rect 34449 13028 34505 13030
rect 34529 13028 34585 13030
rect 28998 9424 29054 9480
rect 27618 4664 27674 4720
rect 28078 4664 28134 4720
rect 27158 4528 27214 4584
rect 27622 3834 27678 3836
rect 27702 3834 27758 3836
rect 27782 3834 27838 3836
rect 27862 3834 27918 3836
rect 27622 3782 27648 3834
rect 27648 3782 27678 3834
rect 27702 3782 27712 3834
rect 27712 3782 27758 3834
rect 27782 3782 27828 3834
rect 27828 3782 27838 3834
rect 27862 3782 27892 3834
rect 27892 3782 27918 3834
rect 27622 3780 27678 3782
rect 27702 3780 27758 3782
rect 27782 3780 27838 3782
rect 27862 3780 27918 3782
rect 27622 2746 27678 2748
rect 27702 2746 27758 2748
rect 27782 2746 27838 2748
rect 27862 2746 27918 2748
rect 27622 2694 27648 2746
rect 27648 2694 27678 2746
rect 27702 2694 27712 2746
rect 27712 2694 27758 2746
rect 27782 2694 27828 2746
rect 27828 2694 27838 2746
rect 27862 2694 27892 2746
rect 27892 2694 27918 2746
rect 27622 2692 27678 2694
rect 27702 2692 27758 2694
rect 27782 2692 27838 2694
rect 27862 2692 27918 2694
rect 34289 11994 34345 11996
rect 34369 11994 34425 11996
rect 34449 11994 34505 11996
rect 34529 11994 34585 11996
rect 34289 11942 34315 11994
rect 34315 11942 34345 11994
rect 34369 11942 34379 11994
rect 34379 11942 34425 11994
rect 34449 11942 34495 11994
rect 34495 11942 34505 11994
rect 34529 11942 34559 11994
rect 34559 11942 34585 11994
rect 34289 11940 34345 11942
rect 34369 11940 34425 11942
rect 34449 11940 34505 11942
rect 34529 11940 34585 11942
rect 34289 10906 34345 10908
rect 34369 10906 34425 10908
rect 34449 10906 34505 10908
rect 34529 10906 34585 10908
rect 34289 10854 34315 10906
rect 34315 10854 34345 10906
rect 34369 10854 34379 10906
rect 34379 10854 34425 10906
rect 34449 10854 34495 10906
rect 34495 10854 34505 10906
rect 34529 10854 34559 10906
rect 34559 10854 34585 10906
rect 34289 10852 34345 10854
rect 34369 10852 34425 10854
rect 34449 10852 34505 10854
rect 34529 10852 34585 10854
rect 34289 9818 34345 9820
rect 34369 9818 34425 9820
rect 34449 9818 34505 9820
rect 34529 9818 34585 9820
rect 34289 9766 34315 9818
rect 34315 9766 34345 9818
rect 34369 9766 34379 9818
rect 34379 9766 34425 9818
rect 34449 9766 34495 9818
rect 34495 9766 34505 9818
rect 34529 9766 34559 9818
rect 34559 9766 34585 9818
rect 34289 9764 34345 9766
rect 34369 9764 34425 9766
rect 34449 9764 34505 9766
rect 34529 9764 34585 9766
rect 32678 9424 32734 9480
rect 34150 9016 34206 9072
rect 34289 8730 34345 8732
rect 34369 8730 34425 8732
rect 34449 8730 34505 8732
rect 34529 8730 34585 8732
rect 34289 8678 34315 8730
rect 34315 8678 34345 8730
rect 34369 8678 34379 8730
rect 34379 8678 34425 8730
rect 34449 8678 34495 8730
rect 34495 8678 34505 8730
rect 34529 8678 34559 8730
rect 34559 8678 34585 8730
rect 34289 8676 34345 8678
rect 34369 8676 34425 8678
rect 34449 8676 34505 8678
rect 34529 8676 34585 8678
rect 31482 7384 31538 7440
rect 34289 7642 34345 7644
rect 34369 7642 34425 7644
rect 34449 7642 34505 7644
rect 34529 7642 34585 7644
rect 34289 7590 34315 7642
rect 34315 7590 34345 7642
rect 34369 7590 34379 7642
rect 34379 7590 34425 7642
rect 34449 7590 34495 7642
rect 34495 7590 34505 7642
rect 34529 7590 34559 7642
rect 34559 7590 34585 7642
rect 34289 7588 34345 7590
rect 34369 7588 34425 7590
rect 34449 7588 34505 7590
rect 34529 7588 34585 7590
rect 35622 12552 35678 12608
rect 39578 15408 39634 15464
rect 35622 9696 35678 9752
rect 37002 10240 37058 10296
rect 37002 9016 37058 9072
rect 34289 6554 34345 6556
rect 34369 6554 34425 6556
rect 34449 6554 34505 6556
rect 34529 6554 34585 6556
rect 34289 6502 34315 6554
rect 34315 6502 34345 6554
rect 34369 6502 34379 6554
rect 34379 6502 34425 6554
rect 34449 6502 34495 6554
rect 34495 6502 34505 6554
rect 34529 6502 34559 6554
rect 34559 6502 34585 6554
rect 34289 6500 34345 6502
rect 34369 6500 34425 6502
rect 34449 6500 34505 6502
rect 34529 6500 34585 6502
rect 32402 5616 32458 5672
rect 30930 3984 30986 4040
rect 34289 5466 34345 5468
rect 34369 5466 34425 5468
rect 34449 5466 34505 5468
rect 34529 5466 34585 5468
rect 34289 5414 34315 5466
rect 34315 5414 34345 5466
rect 34369 5414 34379 5466
rect 34379 5414 34425 5466
rect 34449 5414 34495 5466
rect 34495 5414 34505 5466
rect 34529 5414 34559 5466
rect 34559 5414 34585 5466
rect 34289 5412 34345 5414
rect 34369 5412 34425 5414
rect 34449 5412 34505 5414
rect 34529 5412 34585 5414
rect 36634 7656 36690 7712
rect 39578 8608 39634 8664
rect 38106 6840 38162 6896
rect 34289 4378 34345 4380
rect 34369 4378 34425 4380
rect 34449 4378 34505 4380
rect 34529 4378 34585 4380
rect 34289 4326 34315 4378
rect 34315 4326 34345 4378
rect 34369 4326 34379 4378
rect 34379 4326 34425 4378
rect 34449 4326 34495 4378
rect 34495 4326 34505 4378
rect 34529 4326 34559 4378
rect 34559 4326 34585 4378
rect 34289 4324 34345 4326
rect 34369 4324 34425 4326
rect 34449 4324 34505 4326
rect 34529 4324 34585 4326
rect 34150 3440 34206 3496
rect 34289 3290 34345 3292
rect 34369 3290 34425 3292
rect 34449 3290 34505 3292
rect 34529 3290 34585 3292
rect 34289 3238 34315 3290
rect 34315 3238 34345 3290
rect 34369 3238 34379 3290
rect 34379 3238 34425 3290
rect 34449 3238 34495 3290
rect 34495 3238 34505 3290
rect 34529 3238 34559 3290
rect 34559 3238 34585 3290
rect 34289 3236 34345 3238
rect 34369 3236 34425 3238
rect 34449 3236 34505 3238
rect 34529 3236 34585 3238
rect 25410 1808 25466 1864
rect 29642 1400 29698 1456
rect 27250 1264 27306 1320
rect 34289 2202 34345 2204
rect 34369 2202 34425 2204
rect 34449 2202 34505 2204
rect 34529 2202 34585 2204
rect 34289 2150 34315 2202
rect 34315 2150 34345 2202
rect 34369 2150 34379 2202
rect 34379 2150 34425 2202
rect 34449 2150 34495 2202
rect 34495 2150 34505 2202
rect 34529 2150 34559 2202
rect 34559 2150 34585 2202
rect 34289 2148 34345 2150
rect 34369 2148 34425 2150
rect 34449 2148 34505 2150
rect 34529 2148 34585 2150
rect 39578 3984 39634 4040
rect 39578 2760 39634 2816
rect 38566 1264 38622 1320
<< metal3 >>
rect 0 15512 480 15632
rect 62 15058 122 15512
rect 39520 15466 40000 15496
rect 39492 15464 40000 15466
rect 39492 15408 39578 15464
rect 39634 15408 40000 15464
rect 39492 15406 40000 15408
rect 39520 15376 40000 15406
rect 1117 15058 1183 15061
rect 62 15056 1183 15058
rect 62 15000 1122 15056
rect 1178 15000 1183 15056
rect 62 14998 1183 15000
rect 1117 14995 1183 14998
rect 0 14560 480 14680
rect 62 14242 122 14560
rect 39520 14288 40000 14408
rect 1945 14242 2011 14245
rect 62 14240 2011 14242
rect 62 14184 1950 14240
rect 2006 14184 2011 14240
rect 62 14182 2011 14184
rect 1945 14179 2011 14182
rect 35617 14106 35683 14109
rect 39622 14106 39682 14288
rect 35617 14104 39682 14106
rect 35617 14048 35622 14104
rect 35678 14048 39682 14104
rect 35617 14046 39682 14048
rect 35617 14043 35683 14046
rect 0 13696 480 13728
rect 0 13640 110 13696
rect 166 13640 480 13696
rect 0 13608 480 13640
rect 14277 13632 14597 13633
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 13567 14597 13568
rect 27610 13632 27930 13633
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 13567 27930 13568
rect 7610 13088 7930 13089
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7930 13088
rect 7610 13023 7930 13024
rect 20944 13088 21264 13089
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 13023 21264 13024
rect 34277 13088 34597 13089
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 39520 13064 40000 13184
rect 34277 13023 34597 13024
rect 0 12656 480 12776
rect 62 12474 122 12656
rect 35617 12610 35683 12613
rect 39622 12610 39682 13064
rect 35617 12608 39682 12610
rect 35617 12552 35622 12608
rect 35678 12552 39682 12608
rect 35617 12550 39682 12552
rect 35617 12547 35683 12550
rect 14277 12544 14597 12545
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 12479 14597 12480
rect 27610 12544 27930 12545
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 27610 12479 27930 12480
rect 1577 12474 1643 12477
rect 62 12472 1643 12474
rect 62 12416 1582 12472
rect 1638 12416 1643 12472
rect 62 12414 1643 12416
rect 1577 12411 1643 12414
rect 7610 12000 7930 12001
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7930 12000
rect 7610 11935 7930 11936
rect 20944 12000 21264 12001
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 11935 21264 11936
rect 34277 12000 34597 12001
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 39520 11976 40000 12096
rect 34277 11935 34597 11936
rect 0 11792 480 11824
rect 0 11736 110 11792
rect 166 11736 480 11792
rect 0 11704 480 11736
rect 5625 11794 5691 11797
rect 17585 11794 17651 11797
rect 5625 11792 17651 11794
rect 5625 11736 5630 11792
rect 5686 11736 17590 11792
rect 17646 11736 17651 11792
rect 5625 11734 17651 11736
rect 5625 11731 5691 11734
rect 17585 11731 17651 11734
rect 2037 11658 2103 11661
rect 12525 11658 12591 11661
rect 19057 11658 19123 11661
rect 2037 11656 19123 11658
rect 2037 11600 2042 11656
rect 2098 11600 12530 11656
rect 12586 11600 19062 11656
rect 19118 11600 19123 11656
rect 2037 11598 19123 11600
rect 2037 11595 2103 11598
rect 12525 11595 12591 11598
rect 19057 11595 19123 11598
rect 24485 11658 24551 11661
rect 39622 11658 39682 11976
rect 24485 11656 39682 11658
rect 24485 11600 24490 11656
rect 24546 11600 39682 11656
rect 24485 11598 39682 11600
rect 24485 11595 24551 11598
rect 14277 11456 14597 11457
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 11391 14597 11392
rect 27610 11456 27930 11457
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 27610 11391 27930 11392
rect 7610 10912 7930 10913
rect 0 10752 480 10872
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7930 10912
rect 7610 10847 7930 10848
rect 20944 10912 21264 10913
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 10847 21264 10848
rect 34277 10912 34597 10913
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 34277 10847 34597 10848
rect 39520 10752 40000 10872
rect 62 10298 122 10752
rect 1761 10706 1827 10709
rect 11881 10706 11947 10709
rect 1761 10704 11947 10706
rect 1761 10648 1766 10704
rect 1822 10648 11886 10704
rect 11942 10648 11947 10704
rect 1761 10646 11947 10648
rect 1761 10643 1827 10646
rect 11881 10643 11947 10646
rect 9121 10570 9187 10573
rect 9121 10568 18660 10570
rect 9121 10512 9126 10568
rect 9182 10512 18660 10568
rect 9121 10510 18660 10512
rect 9121 10507 9187 10510
rect 18600 10434 18660 10510
rect 23565 10434 23631 10437
rect 25589 10434 25655 10437
rect 18600 10432 25655 10434
rect 18600 10376 23570 10432
rect 23626 10376 25594 10432
rect 25650 10376 25655 10432
rect 18600 10374 25655 10376
rect 23565 10371 23631 10374
rect 25589 10371 25655 10374
rect 14277 10368 14597 10369
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 10303 14597 10304
rect 27610 10368 27930 10369
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 10303 27930 10304
rect 1393 10298 1459 10301
rect 62 10296 1459 10298
rect 62 10240 1398 10296
rect 1454 10240 1459 10296
rect 62 10238 1459 10240
rect 1393 10235 1459 10238
rect 2957 10298 3023 10301
rect 4521 10298 4587 10301
rect 2957 10296 4587 10298
rect 2957 10240 2962 10296
rect 3018 10240 4526 10296
rect 4582 10240 4587 10296
rect 2957 10238 4587 10240
rect 2957 10235 3023 10238
rect 4521 10235 4587 10238
rect 15193 10298 15259 10301
rect 18229 10298 18295 10301
rect 24301 10298 24367 10301
rect 15193 10296 24367 10298
rect 15193 10240 15198 10296
rect 15254 10240 18234 10296
rect 18290 10240 24306 10296
rect 24362 10240 24367 10296
rect 15193 10238 24367 10240
rect 15193 10235 15259 10238
rect 18229 10235 18295 10238
rect 24301 10235 24367 10238
rect 36997 10298 37063 10301
rect 39622 10298 39682 10752
rect 36997 10296 39682 10298
rect 36997 10240 37002 10296
rect 37058 10240 39682 10296
rect 36997 10238 39682 10240
rect 36997 10235 37063 10238
rect 14733 10162 14799 10165
rect 25497 10162 25563 10165
rect 14733 10160 25563 10162
rect 14733 10104 14738 10160
rect 14794 10104 25502 10160
rect 25558 10104 25563 10160
rect 14733 10102 25563 10104
rect 14733 10099 14799 10102
rect 25497 10099 25563 10102
rect 0 9888 480 9920
rect 0 9832 110 9888
rect 166 9832 480 9888
rect 0 9800 480 9832
rect 7610 9824 7930 9825
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7930 9824
rect 7610 9759 7930 9760
rect 20944 9824 21264 9825
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 9759 21264 9760
rect 34277 9824 34597 9825
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 34277 9759 34597 9760
rect 5993 9752 6059 9757
rect 5993 9696 5998 9752
rect 6054 9696 6059 9752
rect 5993 9691 6059 9696
rect 35617 9754 35683 9757
rect 39520 9754 40000 9784
rect 35617 9752 40000 9754
rect 35617 9696 35622 9752
rect 35678 9696 40000 9752
rect 35617 9694 40000 9696
rect 35617 9691 35683 9694
rect 1945 9618 2011 9621
rect 5996 9618 6056 9691
rect 39520 9664 40000 9694
rect 11789 9618 11855 9621
rect 1945 9616 4170 9618
rect 1945 9560 1950 9616
rect 2006 9560 4170 9616
rect 1945 9558 4170 9560
rect 5996 9616 11855 9618
rect 5996 9560 11794 9616
rect 11850 9560 11855 9616
rect 5996 9558 11855 9560
rect 1945 9555 2011 9558
rect 4110 9482 4170 9558
rect 11789 9555 11855 9558
rect 13445 9618 13511 9621
rect 15929 9618 15995 9621
rect 13445 9616 15995 9618
rect 13445 9560 13450 9616
rect 13506 9560 15934 9616
rect 15990 9560 15995 9616
rect 13445 9558 15995 9560
rect 13445 9555 13511 9558
rect 15929 9555 15995 9558
rect 23197 9618 23263 9621
rect 24485 9618 24551 9621
rect 23197 9616 24551 9618
rect 23197 9560 23202 9616
rect 23258 9560 24490 9616
rect 24546 9560 24551 9616
rect 23197 9558 24551 9560
rect 23197 9555 23263 9558
rect 24485 9555 24551 9558
rect 6361 9482 6427 9485
rect 4110 9480 6427 9482
rect 4110 9424 6366 9480
rect 6422 9424 6427 9480
rect 4110 9422 6427 9424
rect 6361 9419 6427 9422
rect 12341 9482 12407 9485
rect 18689 9482 18755 9485
rect 12341 9480 18755 9482
rect 12341 9424 12346 9480
rect 12402 9424 18694 9480
rect 18750 9424 18755 9480
rect 12341 9422 18755 9424
rect 12341 9419 12407 9422
rect 18689 9419 18755 9422
rect 21909 9482 21975 9485
rect 24577 9482 24643 9485
rect 21909 9480 24643 9482
rect 21909 9424 21914 9480
rect 21970 9424 24582 9480
rect 24638 9424 24643 9480
rect 21909 9422 24643 9424
rect 21909 9419 21975 9422
rect 24577 9419 24643 9422
rect 28993 9482 29059 9485
rect 32673 9482 32739 9485
rect 28993 9480 32739 9482
rect 28993 9424 28998 9480
rect 29054 9424 32678 9480
rect 32734 9424 32739 9480
rect 28993 9422 32739 9424
rect 28993 9419 29059 9422
rect 32673 9419 32739 9422
rect 14277 9280 14597 9281
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 9215 14597 9216
rect 27610 9280 27930 9281
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 27610 9215 27930 9216
rect 3693 9210 3759 9213
rect 9305 9210 9371 9213
rect 3693 9208 9371 9210
rect 3693 9152 3698 9208
rect 3754 9152 9310 9208
rect 9366 9152 9371 9208
rect 3693 9150 9371 9152
rect 3693 9147 3759 9150
rect 9305 9147 9371 9150
rect 18873 9210 18939 9213
rect 19241 9210 19307 9213
rect 26785 9210 26851 9213
rect 18873 9208 26851 9210
rect 18873 9152 18878 9208
rect 18934 9152 19246 9208
rect 19302 9152 26790 9208
rect 26846 9152 26851 9208
rect 18873 9150 26851 9152
rect 18873 9147 18939 9150
rect 19241 9147 19307 9150
rect 26785 9147 26851 9150
rect 8109 9074 8175 9077
rect 34145 9074 34211 9077
rect 36997 9074 37063 9077
rect 8109 9072 37063 9074
rect 8109 9016 8114 9072
rect 8170 9016 34150 9072
rect 34206 9016 37002 9072
rect 37058 9016 37063 9072
rect 8109 9014 37063 9016
rect 8109 9011 8175 9014
rect 34145 9011 34211 9014
rect 36997 9011 37063 9014
rect 0 8936 480 8968
rect 0 8880 110 8936
rect 166 8880 480 8936
rect 0 8848 480 8880
rect 13905 8938 13971 8941
rect 23749 8938 23815 8941
rect 13905 8936 23815 8938
rect 13905 8880 13910 8936
rect 13966 8880 23754 8936
rect 23810 8880 23815 8936
rect 13905 8878 23815 8880
rect 13905 8875 13971 8878
rect 23749 8875 23815 8878
rect 7610 8736 7930 8737
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7930 8736
rect 7610 8671 7930 8672
rect 20944 8736 21264 8737
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 8671 21264 8672
rect 34277 8736 34597 8737
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 8671 34597 8672
rect 39520 8666 40000 8696
rect 39492 8664 40000 8666
rect 39492 8608 39578 8664
rect 39634 8608 40000 8664
rect 39492 8606 40000 8608
rect 39520 8576 40000 8606
rect 15929 8530 15995 8533
rect 26233 8530 26299 8533
rect 15929 8528 26299 8530
rect 15929 8472 15934 8528
rect 15990 8472 26238 8528
rect 26294 8472 26299 8528
rect 15929 8470 26299 8472
rect 15929 8467 15995 8470
rect 26233 8467 26299 8470
rect 12249 8394 12315 8397
rect 19885 8394 19951 8397
rect 12249 8392 19951 8394
rect 12249 8336 12254 8392
rect 12310 8336 19890 8392
rect 19946 8336 19951 8392
rect 12249 8334 19951 8336
rect 12249 8331 12315 8334
rect 19885 8331 19951 8334
rect 14277 8192 14597 8193
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 8127 14597 8128
rect 27610 8192 27930 8193
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 8127 27930 8128
rect 0 7984 480 8016
rect 0 7928 18 7984
rect 74 7928 480 7984
rect 0 7896 480 7928
rect 7097 7986 7163 7989
rect 16481 7986 16547 7989
rect 7097 7984 16547 7986
rect 7097 7928 7102 7984
rect 7158 7928 16486 7984
rect 16542 7928 16547 7984
rect 7097 7926 16547 7928
rect 7097 7923 7163 7926
rect 16481 7923 16547 7926
rect 10869 7850 10935 7853
rect 24117 7850 24183 7853
rect 10869 7848 24183 7850
rect 10869 7792 10874 7848
rect 10930 7792 24122 7848
rect 24178 7792 24183 7848
rect 10869 7790 24183 7792
rect 10869 7787 10935 7790
rect 24117 7787 24183 7790
rect 36629 7714 36695 7717
rect 39614 7714 39620 7716
rect 36629 7712 39620 7714
rect 36629 7656 36634 7712
rect 36690 7656 39620 7712
rect 36629 7654 39620 7656
rect 36629 7651 36695 7654
rect 39614 7652 39620 7654
rect 39684 7652 39690 7716
rect 7610 7648 7930 7649
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7930 7648
rect 7610 7583 7930 7584
rect 20944 7648 21264 7649
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 7583 21264 7584
rect 34277 7648 34597 7649
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 7583 34597 7584
rect 3969 7442 4035 7445
rect 62 7440 4035 7442
rect 62 7384 3974 7440
rect 4030 7384 4035 7440
rect 62 7382 4035 7384
rect 62 7064 122 7382
rect 3969 7379 4035 7382
rect 10777 7442 10843 7445
rect 15285 7442 15351 7445
rect 31477 7442 31543 7445
rect 39520 7444 40000 7472
rect 39520 7442 39620 7444
rect 10777 7440 31543 7442
rect 10777 7384 10782 7440
rect 10838 7384 15290 7440
rect 15346 7384 31482 7440
rect 31538 7384 31543 7440
rect 10777 7382 31543 7384
rect 39492 7382 39620 7442
rect 10777 7379 10843 7382
rect 15285 7379 15351 7382
rect 31477 7379 31543 7382
rect 39520 7380 39620 7382
rect 39684 7380 40000 7444
rect 39520 7352 40000 7380
rect 21173 7306 21239 7309
rect 25497 7306 25563 7309
rect 21173 7304 25563 7306
rect 21173 7248 21178 7304
rect 21234 7248 25502 7304
rect 25558 7248 25563 7304
rect 21173 7246 25563 7248
rect 21173 7243 21239 7246
rect 25497 7243 25563 7246
rect 14277 7104 14597 7105
rect 0 6944 480 7064
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 7039 14597 7040
rect 27610 7104 27930 7105
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 7039 27930 7040
rect 38101 6898 38167 6901
rect 38101 6896 39682 6898
rect 38101 6840 38106 6896
rect 38162 6840 39682 6896
rect 38101 6838 39682 6840
rect 38101 6835 38167 6838
rect 2773 6762 2839 6765
rect 3601 6762 3667 6765
rect 18045 6762 18111 6765
rect 2773 6760 18111 6762
rect 2773 6704 2778 6760
rect 2834 6704 3606 6760
rect 3662 6704 18050 6760
rect 18106 6704 18111 6760
rect 2773 6702 18111 6704
rect 2773 6699 2839 6702
rect 3601 6699 3667 6702
rect 18045 6699 18111 6702
rect 7610 6560 7930 6561
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7930 6560
rect 7610 6495 7930 6496
rect 20944 6560 21264 6561
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 6495 21264 6496
rect 34277 6560 34597 6561
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 34277 6495 34597 6496
rect 39622 6384 39682 6838
rect 20161 6354 20227 6357
rect 27337 6354 27403 6357
rect 20161 6352 27403 6354
rect 20161 6296 20166 6352
rect 20222 6296 27342 6352
rect 27398 6296 27403 6352
rect 20161 6294 27403 6296
rect 20161 6291 20227 6294
rect 27337 6291 27403 6294
rect 39520 6264 40000 6384
rect 0 6084 480 6112
rect 0 6020 60 6084
rect 124 6020 480 6084
rect 0 5992 480 6020
rect 14277 6016 14597 6017
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 5951 14597 5952
rect 27610 6016 27930 6017
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 5951 27930 5952
rect 54 5748 60 5812
rect 124 5810 130 5812
rect 1485 5810 1551 5813
rect 124 5808 1551 5810
rect 124 5752 1490 5808
rect 1546 5752 1551 5808
rect 124 5750 1551 5752
rect 124 5748 130 5750
rect 1485 5747 1551 5750
rect 8569 5810 8635 5813
rect 11973 5810 12039 5813
rect 24761 5810 24827 5813
rect 8569 5808 24827 5810
rect 8569 5752 8574 5808
rect 8630 5752 11978 5808
rect 12034 5752 24766 5808
rect 24822 5752 24827 5808
rect 8569 5750 24827 5752
rect 8569 5747 8635 5750
rect 11973 5747 12039 5750
rect 24761 5747 24827 5750
rect 2957 5674 3023 5677
rect 62 5672 3023 5674
rect 62 5616 2962 5672
rect 3018 5616 3023 5672
rect 62 5614 3023 5616
rect 62 5160 122 5614
rect 2957 5611 3023 5614
rect 5441 5674 5507 5677
rect 13905 5674 13971 5677
rect 19241 5674 19307 5677
rect 5441 5672 13830 5674
rect 5441 5616 5446 5672
rect 5502 5616 13830 5672
rect 5441 5614 13830 5616
rect 5441 5611 5507 5614
rect 13770 5538 13830 5614
rect 13905 5672 19307 5674
rect 13905 5616 13910 5672
rect 13966 5616 19246 5672
rect 19302 5616 19307 5672
rect 13905 5614 19307 5616
rect 13905 5611 13971 5614
rect 19241 5611 19307 5614
rect 24117 5674 24183 5677
rect 32397 5674 32463 5677
rect 24117 5672 32463 5674
rect 24117 5616 24122 5672
rect 24178 5616 32402 5672
rect 32458 5616 32463 5672
rect 24117 5614 32463 5616
rect 24117 5611 24183 5614
rect 32397 5611 32463 5614
rect 14641 5538 14707 5541
rect 13770 5536 14707 5538
rect 13770 5480 14646 5536
rect 14702 5480 14707 5536
rect 13770 5478 14707 5480
rect 14641 5475 14707 5478
rect 7610 5472 7930 5473
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7930 5472
rect 7610 5407 7930 5408
rect 20944 5472 21264 5473
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 5407 21264 5408
rect 34277 5472 34597 5473
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 34277 5407 34597 5408
rect 5073 5266 5139 5269
rect 17401 5266 17467 5269
rect 5073 5264 17467 5266
rect 5073 5208 5078 5264
rect 5134 5208 17406 5264
rect 17462 5208 17467 5264
rect 5073 5206 17467 5208
rect 5073 5203 5139 5206
rect 17401 5203 17467 5206
rect 0 5040 480 5160
rect 24853 5130 24919 5133
rect 614 5128 24919 5130
rect 614 5072 24858 5128
rect 24914 5072 24919 5128
rect 614 5070 24919 5072
rect 614 4858 674 5070
rect 24853 5067 24919 5070
rect 39520 5040 40000 5160
rect 1669 4994 1735 4997
rect 13905 4994 13971 4997
rect 1669 4992 13971 4994
rect 1669 4936 1674 4992
rect 1730 4936 13910 4992
rect 13966 4936 13971 4992
rect 1669 4934 13971 4936
rect 1669 4931 1735 4934
rect 13905 4931 13971 4934
rect 14277 4928 14597 4929
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 4863 14597 4864
rect 27610 4928 27930 4929
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 4863 27930 4864
rect 62 4798 674 4858
rect 62 4208 122 4798
rect 9121 4722 9187 4725
rect 10225 4722 10291 4725
rect 12065 4722 12131 4725
rect 27613 4722 27679 4725
rect 28073 4722 28139 4725
rect 9121 4720 28139 4722
rect 9121 4664 9126 4720
rect 9182 4664 10230 4720
rect 10286 4664 12070 4720
rect 12126 4664 27618 4720
rect 27674 4664 28078 4720
rect 28134 4664 28139 4720
rect 9121 4662 28139 4664
rect 9121 4659 9187 4662
rect 10225 4659 10291 4662
rect 12065 4659 12131 4662
rect 27613 4659 27679 4662
rect 28073 4659 28139 4662
rect 9949 4586 10015 4589
rect 27153 4586 27219 4589
rect 9949 4584 27219 4586
rect 9949 4528 9954 4584
rect 10010 4528 27158 4584
rect 27214 4528 27219 4584
rect 9949 4526 27219 4528
rect 9949 4523 10015 4526
rect 27153 4523 27219 4526
rect 39622 4450 39682 5040
rect 39254 4390 39682 4450
rect 7610 4384 7930 4385
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7930 4384
rect 7610 4319 7930 4320
rect 20944 4384 21264 4385
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 4319 21264 4320
rect 34277 4384 34597 4385
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 34277 4319 34597 4320
rect 0 4088 480 4208
rect 5901 4178 5967 4181
rect 15009 4178 15075 4181
rect 16481 4178 16547 4181
rect 5901 4176 16547 4178
rect 5901 4120 5906 4176
rect 5962 4120 15014 4176
rect 15070 4120 16486 4176
rect 16542 4120 16547 4176
rect 5901 4118 16547 4120
rect 5901 4115 5967 4118
rect 15009 4115 15075 4118
rect 16481 4115 16547 4118
rect 24577 4178 24643 4181
rect 39254 4178 39314 4390
rect 24577 4176 39314 4178
rect 24577 4120 24582 4176
rect 24638 4120 39314 4176
rect 24577 4118 39314 4120
rect 24577 4115 24643 4118
rect 8477 4042 8543 4045
rect 13077 4042 13143 4045
rect 8477 4040 13143 4042
rect 8477 3984 8482 4040
rect 8538 3984 13082 4040
rect 13138 3984 13143 4040
rect 8477 3982 13143 3984
rect 8477 3979 8543 3982
rect 13077 3979 13143 3982
rect 25865 4042 25931 4045
rect 30925 4042 30991 4045
rect 39520 4042 40000 4072
rect 25865 4040 30991 4042
rect 25865 3984 25870 4040
rect 25926 3984 30930 4040
rect 30986 3984 30991 4040
rect 25865 3982 30991 3984
rect 39492 4040 40000 4042
rect 39492 3984 39578 4040
rect 39634 3984 40000 4040
rect 39492 3982 40000 3984
rect 25865 3979 25931 3982
rect 30925 3979 30991 3982
rect 39520 3952 40000 3982
rect 14277 3840 14597 3841
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 3775 14597 3776
rect 27610 3840 27930 3841
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 27610 3775 27930 3776
rect 19517 3498 19583 3501
rect 34145 3498 34211 3501
rect 19517 3496 34211 3498
rect 19517 3440 19522 3496
rect 19578 3440 34150 3496
rect 34206 3440 34211 3496
rect 19517 3438 34211 3440
rect 19517 3435 19583 3438
rect 34145 3435 34211 3438
rect 7610 3296 7930 3297
rect 0 3224 480 3256
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7930 3296
rect 7610 3231 7930 3232
rect 20944 3296 21264 3297
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 3231 21264 3232
rect 34277 3296 34597 3297
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 3231 34597 3232
rect 0 3168 110 3224
rect 166 3168 480 3224
rect 0 3136 480 3168
rect 39520 2818 40000 2848
rect 39492 2816 40000 2818
rect 39492 2760 39578 2816
rect 39634 2760 40000 2816
rect 39492 2758 40000 2760
rect 14277 2752 14597 2753
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2687 14597 2688
rect 27610 2752 27930 2753
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 39520 2728 40000 2758
rect 27610 2687 27930 2688
rect 18413 2410 18479 2413
rect 18413 2408 39682 2410
rect 18413 2352 18418 2408
rect 18474 2352 39682 2408
rect 18413 2350 39682 2352
rect 18413 2347 18479 2350
rect 0 2272 480 2304
rect 0 2216 110 2272
rect 166 2216 480 2272
rect 0 2184 480 2216
rect 7610 2208 7930 2209
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7930 2208
rect 7610 2143 7930 2144
rect 20944 2208 21264 2209
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2143 21264 2144
rect 34277 2208 34597 2209
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 34277 2143 34597 2144
rect 15745 2138 15811 2141
rect 8894 2136 15811 2138
rect 8894 2080 15750 2136
rect 15806 2080 15811 2136
rect 8894 2078 15811 2080
rect 2497 1730 2563 1733
rect 8894 1730 8954 2078
rect 15745 2075 15811 2078
rect 9029 2002 9095 2005
rect 15193 2002 15259 2005
rect 9029 2000 15259 2002
rect 9029 1944 9034 2000
rect 9090 1944 15198 2000
rect 15254 1944 15259 2000
rect 9029 1942 15259 1944
rect 9029 1939 9095 1942
rect 15193 1939 15259 1942
rect 18781 1866 18847 1869
rect 25405 1866 25471 1869
rect 18781 1864 25471 1866
rect 18781 1808 18786 1864
rect 18842 1808 25410 1864
rect 25466 1808 25471 1864
rect 18781 1806 25471 1808
rect 18781 1803 18847 1806
rect 25405 1803 25471 1806
rect 39622 1760 39682 2350
rect 2497 1728 8954 1730
rect 2497 1672 2502 1728
rect 2558 1672 8954 1728
rect 2497 1670 8954 1672
rect 9305 1730 9371 1733
rect 17769 1730 17835 1733
rect 9305 1728 17835 1730
rect 9305 1672 9310 1728
rect 9366 1672 17774 1728
rect 17830 1672 17835 1728
rect 9305 1670 17835 1672
rect 2497 1667 2563 1670
rect 9305 1667 9371 1670
rect 17769 1667 17835 1670
rect 39520 1640 40000 1760
rect 6269 1594 6335 1597
rect 62 1592 6335 1594
rect 62 1536 6274 1592
rect 6330 1536 6335 1592
rect 62 1534 6335 1536
rect 62 1352 122 1534
rect 6269 1531 6335 1534
rect 8477 1594 8543 1597
rect 15101 1594 15167 1597
rect 8477 1592 15167 1594
rect 8477 1536 8482 1592
rect 8538 1536 15106 1592
rect 15162 1536 15167 1592
rect 8477 1534 15167 1536
rect 8477 1531 8543 1534
rect 15101 1531 15167 1534
rect 21817 1458 21883 1461
rect 29637 1458 29703 1461
rect 21817 1456 29703 1458
rect 21817 1400 21822 1456
rect 21878 1400 29642 1456
rect 29698 1400 29703 1456
rect 21817 1398 29703 1400
rect 21817 1395 21883 1398
rect 29637 1395 29703 1398
rect 0 1232 480 1352
rect 9213 1322 9279 1325
rect 16941 1322 17007 1325
rect 9213 1320 17007 1322
rect 9213 1264 9218 1320
rect 9274 1264 16946 1320
rect 17002 1264 17007 1320
rect 9213 1262 17007 1264
rect 9213 1259 9279 1262
rect 16941 1259 17007 1262
rect 27245 1322 27311 1325
rect 38561 1322 38627 1325
rect 27245 1320 38627 1322
rect 27245 1264 27250 1320
rect 27306 1264 38566 1320
rect 38622 1264 38627 1320
rect 27245 1262 38627 1264
rect 27245 1259 27311 1262
rect 38561 1259 38627 1262
rect 6637 1050 6703 1053
rect 62 1048 6703 1050
rect 62 992 6642 1048
rect 6698 992 6703 1048
rect 62 990 6703 992
rect 62 536 122 990
rect 6637 987 6703 990
rect 39520 552 40000 672
rect 0 416 480 536
rect 18321 234 18387 237
rect 39622 234 39682 552
rect 18321 232 39682 234
rect 18321 176 18326 232
rect 18382 176 39682 232
rect 18321 174 39682 176
rect 18321 171 18387 174
<< via3 >>
rect 14285 13628 14349 13632
rect 14285 13572 14289 13628
rect 14289 13572 14345 13628
rect 14345 13572 14349 13628
rect 14285 13568 14349 13572
rect 14365 13628 14429 13632
rect 14365 13572 14369 13628
rect 14369 13572 14425 13628
rect 14425 13572 14429 13628
rect 14365 13568 14429 13572
rect 14445 13628 14509 13632
rect 14445 13572 14449 13628
rect 14449 13572 14505 13628
rect 14505 13572 14509 13628
rect 14445 13568 14509 13572
rect 14525 13628 14589 13632
rect 14525 13572 14529 13628
rect 14529 13572 14585 13628
rect 14585 13572 14589 13628
rect 14525 13568 14589 13572
rect 27618 13628 27682 13632
rect 27618 13572 27622 13628
rect 27622 13572 27678 13628
rect 27678 13572 27682 13628
rect 27618 13568 27682 13572
rect 27698 13628 27762 13632
rect 27698 13572 27702 13628
rect 27702 13572 27758 13628
rect 27758 13572 27762 13628
rect 27698 13568 27762 13572
rect 27778 13628 27842 13632
rect 27778 13572 27782 13628
rect 27782 13572 27838 13628
rect 27838 13572 27842 13628
rect 27778 13568 27842 13572
rect 27858 13628 27922 13632
rect 27858 13572 27862 13628
rect 27862 13572 27918 13628
rect 27918 13572 27922 13628
rect 27858 13568 27922 13572
rect 7618 13084 7682 13088
rect 7618 13028 7622 13084
rect 7622 13028 7678 13084
rect 7678 13028 7682 13084
rect 7618 13024 7682 13028
rect 7698 13084 7762 13088
rect 7698 13028 7702 13084
rect 7702 13028 7758 13084
rect 7758 13028 7762 13084
rect 7698 13024 7762 13028
rect 7778 13084 7842 13088
rect 7778 13028 7782 13084
rect 7782 13028 7838 13084
rect 7838 13028 7842 13084
rect 7778 13024 7842 13028
rect 7858 13084 7922 13088
rect 7858 13028 7862 13084
rect 7862 13028 7918 13084
rect 7918 13028 7922 13084
rect 7858 13024 7922 13028
rect 20952 13084 21016 13088
rect 20952 13028 20956 13084
rect 20956 13028 21012 13084
rect 21012 13028 21016 13084
rect 20952 13024 21016 13028
rect 21032 13084 21096 13088
rect 21032 13028 21036 13084
rect 21036 13028 21092 13084
rect 21092 13028 21096 13084
rect 21032 13024 21096 13028
rect 21112 13084 21176 13088
rect 21112 13028 21116 13084
rect 21116 13028 21172 13084
rect 21172 13028 21176 13084
rect 21112 13024 21176 13028
rect 21192 13084 21256 13088
rect 21192 13028 21196 13084
rect 21196 13028 21252 13084
rect 21252 13028 21256 13084
rect 21192 13024 21256 13028
rect 34285 13084 34349 13088
rect 34285 13028 34289 13084
rect 34289 13028 34345 13084
rect 34345 13028 34349 13084
rect 34285 13024 34349 13028
rect 34365 13084 34429 13088
rect 34365 13028 34369 13084
rect 34369 13028 34425 13084
rect 34425 13028 34429 13084
rect 34365 13024 34429 13028
rect 34445 13084 34509 13088
rect 34445 13028 34449 13084
rect 34449 13028 34505 13084
rect 34505 13028 34509 13084
rect 34445 13024 34509 13028
rect 34525 13084 34589 13088
rect 34525 13028 34529 13084
rect 34529 13028 34585 13084
rect 34585 13028 34589 13084
rect 34525 13024 34589 13028
rect 14285 12540 14349 12544
rect 14285 12484 14289 12540
rect 14289 12484 14345 12540
rect 14345 12484 14349 12540
rect 14285 12480 14349 12484
rect 14365 12540 14429 12544
rect 14365 12484 14369 12540
rect 14369 12484 14425 12540
rect 14425 12484 14429 12540
rect 14365 12480 14429 12484
rect 14445 12540 14509 12544
rect 14445 12484 14449 12540
rect 14449 12484 14505 12540
rect 14505 12484 14509 12540
rect 14445 12480 14509 12484
rect 14525 12540 14589 12544
rect 14525 12484 14529 12540
rect 14529 12484 14585 12540
rect 14585 12484 14589 12540
rect 14525 12480 14589 12484
rect 27618 12540 27682 12544
rect 27618 12484 27622 12540
rect 27622 12484 27678 12540
rect 27678 12484 27682 12540
rect 27618 12480 27682 12484
rect 27698 12540 27762 12544
rect 27698 12484 27702 12540
rect 27702 12484 27758 12540
rect 27758 12484 27762 12540
rect 27698 12480 27762 12484
rect 27778 12540 27842 12544
rect 27778 12484 27782 12540
rect 27782 12484 27838 12540
rect 27838 12484 27842 12540
rect 27778 12480 27842 12484
rect 27858 12540 27922 12544
rect 27858 12484 27862 12540
rect 27862 12484 27918 12540
rect 27918 12484 27922 12540
rect 27858 12480 27922 12484
rect 7618 11996 7682 12000
rect 7618 11940 7622 11996
rect 7622 11940 7678 11996
rect 7678 11940 7682 11996
rect 7618 11936 7682 11940
rect 7698 11996 7762 12000
rect 7698 11940 7702 11996
rect 7702 11940 7758 11996
rect 7758 11940 7762 11996
rect 7698 11936 7762 11940
rect 7778 11996 7842 12000
rect 7778 11940 7782 11996
rect 7782 11940 7838 11996
rect 7838 11940 7842 11996
rect 7778 11936 7842 11940
rect 7858 11996 7922 12000
rect 7858 11940 7862 11996
rect 7862 11940 7918 11996
rect 7918 11940 7922 11996
rect 7858 11936 7922 11940
rect 20952 11996 21016 12000
rect 20952 11940 20956 11996
rect 20956 11940 21012 11996
rect 21012 11940 21016 11996
rect 20952 11936 21016 11940
rect 21032 11996 21096 12000
rect 21032 11940 21036 11996
rect 21036 11940 21092 11996
rect 21092 11940 21096 11996
rect 21032 11936 21096 11940
rect 21112 11996 21176 12000
rect 21112 11940 21116 11996
rect 21116 11940 21172 11996
rect 21172 11940 21176 11996
rect 21112 11936 21176 11940
rect 21192 11996 21256 12000
rect 21192 11940 21196 11996
rect 21196 11940 21252 11996
rect 21252 11940 21256 11996
rect 21192 11936 21256 11940
rect 34285 11996 34349 12000
rect 34285 11940 34289 11996
rect 34289 11940 34345 11996
rect 34345 11940 34349 11996
rect 34285 11936 34349 11940
rect 34365 11996 34429 12000
rect 34365 11940 34369 11996
rect 34369 11940 34425 11996
rect 34425 11940 34429 11996
rect 34365 11936 34429 11940
rect 34445 11996 34509 12000
rect 34445 11940 34449 11996
rect 34449 11940 34505 11996
rect 34505 11940 34509 11996
rect 34445 11936 34509 11940
rect 34525 11996 34589 12000
rect 34525 11940 34529 11996
rect 34529 11940 34585 11996
rect 34585 11940 34589 11996
rect 34525 11936 34589 11940
rect 14285 11452 14349 11456
rect 14285 11396 14289 11452
rect 14289 11396 14345 11452
rect 14345 11396 14349 11452
rect 14285 11392 14349 11396
rect 14365 11452 14429 11456
rect 14365 11396 14369 11452
rect 14369 11396 14425 11452
rect 14425 11396 14429 11452
rect 14365 11392 14429 11396
rect 14445 11452 14509 11456
rect 14445 11396 14449 11452
rect 14449 11396 14505 11452
rect 14505 11396 14509 11452
rect 14445 11392 14509 11396
rect 14525 11452 14589 11456
rect 14525 11396 14529 11452
rect 14529 11396 14585 11452
rect 14585 11396 14589 11452
rect 14525 11392 14589 11396
rect 27618 11452 27682 11456
rect 27618 11396 27622 11452
rect 27622 11396 27678 11452
rect 27678 11396 27682 11452
rect 27618 11392 27682 11396
rect 27698 11452 27762 11456
rect 27698 11396 27702 11452
rect 27702 11396 27758 11452
rect 27758 11396 27762 11452
rect 27698 11392 27762 11396
rect 27778 11452 27842 11456
rect 27778 11396 27782 11452
rect 27782 11396 27838 11452
rect 27838 11396 27842 11452
rect 27778 11392 27842 11396
rect 27858 11452 27922 11456
rect 27858 11396 27862 11452
rect 27862 11396 27918 11452
rect 27918 11396 27922 11452
rect 27858 11392 27922 11396
rect 7618 10908 7682 10912
rect 7618 10852 7622 10908
rect 7622 10852 7678 10908
rect 7678 10852 7682 10908
rect 7618 10848 7682 10852
rect 7698 10908 7762 10912
rect 7698 10852 7702 10908
rect 7702 10852 7758 10908
rect 7758 10852 7762 10908
rect 7698 10848 7762 10852
rect 7778 10908 7842 10912
rect 7778 10852 7782 10908
rect 7782 10852 7838 10908
rect 7838 10852 7842 10908
rect 7778 10848 7842 10852
rect 7858 10908 7922 10912
rect 7858 10852 7862 10908
rect 7862 10852 7918 10908
rect 7918 10852 7922 10908
rect 7858 10848 7922 10852
rect 20952 10908 21016 10912
rect 20952 10852 20956 10908
rect 20956 10852 21012 10908
rect 21012 10852 21016 10908
rect 20952 10848 21016 10852
rect 21032 10908 21096 10912
rect 21032 10852 21036 10908
rect 21036 10852 21092 10908
rect 21092 10852 21096 10908
rect 21032 10848 21096 10852
rect 21112 10908 21176 10912
rect 21112 10852 21116 10908
rect 21116 10852 21172 10908
rect 21172 10852 21176 10908
rect 21112 10848 21176 10852
rect 21192 10908 21256 10912
rect 21192 10852 21196 10908
rect 21196 10852 21252 10908
rect 21252 10852 21256 10908
rect 21192 10848 21256 10852
rect 34285 10908 34349 10912
rect 34285 10852 34289 10908
rect 34289 10852 34345 10908
rect 34345 10852 34349 10908
rect 34285 10848 34349 10852
rect 34365 10908 34429 10912
rect 34365 10852 34369 10908
rect 34369 10852 34425 10908
rect 34425 10852 34429 10908
rect 34365 10848 34429 10852
rect 34445 10908 34509 10912
rect 34445 10852 34449 10908
rect 34449 10852 34505 10908
rect 34505 10852 34509 10908
rect 34445 10848 34509 10852
rect 34525 10908 34589 10912
rect 34525 10852 34529 10908
rect 34529 10852 34585 10908
rect 34585 10852 34589 10908
rect 34525 10848 34589 10852
rect 14285 10364 14349 10368
rect 14285 10308 14289 10364
rect 14289 10308 14345 10364
rect 14345 10308 14349 10364
rect 14285 10304 14349 10308
rect 14365 10364 14429 10368
rect 14365 10308 14369 10364
rect 14369 10308 14425 10364
rect 14425 10308 14429 10364
rect 14365 10304 14429 10308
rect 14445 10364 14509 10368
rect 14445 10308 14449 10364
rect 14449 10308 14505 10364
rect 14505 10308 14509 10364
rect 14445 10304 14509 10308
rect 14525 10364 14589 10368
rect 14525 10308 14529 10364
rect 14529 10308 14585 10364
rect 14585 10308 14589 10364
rect 14525 10304 14589 10308
rect 27618 10364 27682 10368
rect 27618 10308 27622 10364
rect 27622 10308 27678 10364
rect 27678 10308 27682 10364
rect 27618 10304 27682 10308
rect 27698 10364 27762 10368
rect 27698 10308 27702 10364
rect 27702 10308 27758 10364
rect 27758 10308 27762 10364
rect 27698 10304 27762 10308
rect 27778 10364 27842 10368
rect 27778 10308 27782 10364
rect 27782 10308 27838 10364
rect 27838 10308 27842 10364
rect 27778 10304 27842 10308
rect 27858 10364 27922 10368
rect 27858 10308 27862 10364
rect 27862 10308 27918 10364
rect 27918 10308 27922 10364
rect 27858 10304 27922 10308
rect 7618 9820 7682 9824
rect 7618 9764 7622 9820
rect 7622 9764 7678 9820
rect 7678 9764 7682 9820
rect 7618 9760 7682 9764
rect 7698 9820 7762 9824
rect 7698 9764 7702 9820
rect 7702 9764 7758 9820
rect 7758 9764 7762 9820
rect 7698 9760 7762 9764
rect 7778 9820 7842 9824
rect 7778 9764 7782 9820
rect 7782 9764 7838 9820
rect 7838 9764 7842 9820
rect 7778 9760 7842 9764
rect 7858 9820 7922 9824
rect 7858 9764 7862 9820
rect 7862 9764 7918 9820
rect 7918 9764 7922 9820
rect 7858 9760 7922 9764
rect 20952 9820 21016 9824
rect 20952 9764 20956 9820
rect 20956 9764 21012 9820
rect 21012 9764 21016 9820
rect 20952 9760 21016 9764
rect 21032 9820 21096 9824
rect 21032 9764 21036 9820
rect 21036 9764 21092 9820
rect 21092 9764 21096 9820
rect 21032 9760 21096 9764
rect 21112 9820 21176 9824
rect 21112 9764 21116 9820
rect 21116 9764 21172 9820
rect 21172 9764 21176 9820
rect 21112 9760 21176 9764
rect 21192 9820 21256 9824
rect 21192 9764 21196 9820
rect 21196 9764 21252 9820
rect 21252 9764 21256 9820
rect 21192 9760 21256 9764
rect 34285 9820 34349 9824
rect 34285 9764 34289 9820
rect 34289 9764 34345 9820
rect 34345 9764 34349 9820
rect 34285 9760 34349 9764
rect 34365 9820 34429 9824
rect 34365 9764 34369 9820
rect 34369 9764 34425 9820
rect 34425 9764 34429 9820
rect 34365 9760 34429 9764
rect 34445 9820 34509 9824
rect 34445 9764 34449 9820
rect 34449 9764 34505 9820
rect 34505 9764 34509 9820
rect 34445 9760 34509 9764
rect 34525 9820 34589 9824
rect 34525 9764 34529 9820
rect 34529 9764 34585 9820
rect 34585 9764 34589 9820
rect 34525 9760 34589 9764
rect 14285 9276 14349 9280
rect 14285 9220 14289 9276
rect 14289 9220 14345 9276
rect 14345 9220 14349 9276
rect 14285 9216 14349 9220
rect 14365 9276 14429 9280
rect 14365 9220 14369 9276
rect 14369 9220 14425 9276
rect 14425 9220 14429 9276
rect 14365 9216 14429 9220
rect 14445 9276 14509 9280
rect 14445 9220 14449 9276
rect 14449 9220 14505 9276
rect 14505 9220 14509 9276
rect 14445 9216 14509 9220
rect 14525 9276 14589 9280
rect 14525 9220 14529 9276
rect 14529 9220 14585 9276
rect 14585 9220 14589 9276
rect 14525 9216 14589 9220
rect 27618 9276 27682 9280
rect 27618 9220 27622 9276
rect 27622 9220 27678 9276
rect 27678 9220 27682 9276
rect 27618 9216 27682 9220
rect 27698 9276 27762 9280
rect 27698 9220 27702 9276
rect 27702 9220 27758 9276
rect 27758 9220 27762 9276
rect 27698 9216 27762 9220
rect 27778 9276 27842 9280
rect 27778 9220 27782 9276
rect 27782 9220 27838 9276
rect 27838 9220 27842 9276
rect 27778 9216 27842 9220
rect 27858 9276 27922 9280
rect 27858 9220 27862 9276
rect 27862 9220 27918 9276
rect 27918 9220 27922 9276
rect 27858 9216 27922 9220
rect 7618 8732 7682 8736
rect 7618 8676 7622 8732
rect 7622 8676 7678 8732
rect 7678 8676 7682 8732
rect 7618 8672 7682 8676
rect 7698 8732 7762 8736
rect 7698 8676 7702 8732
rect 7702 8676 7758 8732
rect 7758 8676 7762 8732
rect 7698 8672 7762 8676
rect 7778 8732 7842 8736
rect 7778 8676 7782 8732
rect 7782 8676 7838 8732
rect 7838 8676 7842 8732
rect 7778 8672 7842 8676
rect 7858 8732 7922 8736
rect 7858 8676 7862 8732
rect 7862 8676 7918 8732
rect 7918 8676 7922 8732
rect 7858 8672 7922 8676
rect 20952 8732 21016 8736
rect 20952 8676 20956 8732
rect 20956 8676 21012 8732
rect 21012 8676 21016 8732
rect 20952 8672 21016 8676
rect 21032 8732 21096 8736
rect 21032 8676 21036 8732
rect 21036 8676 21092 8732
rect 21092 8676 21096 8732
rect 21032 8672 21096 8676
rect 21112 8732 21176 8736
rect 21112 8676 21116 8732
rect 21116 8676 21172 8732
rect 21172 8676 21176 8732
rect 21112 8672 21176 8676
rect 21192 8732 21256 8736
rect 21192 8676 21196 8732
rect 21196 8676 21252 8732
rect 21252 8676 21256 8732
rect 21192 8672 21256 8676
rect 34285 8732 34349 8736
rect 34285 8676 34289 8732
rect 34289 8676 34345 8732
rect 34345 8676 34349 8732
rect 34285 8672 34349 8676
rect 34365 8732 34429 8736
rect 34365 8676 34369 8732
rect 34369 8676 34425 8732
rect 34425 8676 34429 8732
rect 34365 8672 34429 8676
rect 34445 8732 34509 8736
rect 34445 8676 34449 8732
rect 34449 8676 34505 8732
rect 34505 8676 34509 8732
rect 34445 8672 34509 8676
rect 34525 8732 34589 8736
rect 34525 8676 34529 8732
rect 34529 8676 34585 8732
rect 34585 8676 34589 8732
rect 34525 8672 34589 8676
rect 14285 8188 14349 8192
rect 14285 8132 14289 8188
rect 14289 8132 14345 8188
rect 14345 8132 14349 8188
rect 14285 8128 14349 8132
rect 14365 8188 14429 8192
rect 14365 8132 14369 8188
rect 14369 8132 14425 8188
rect 14425 8132 14429 8188
rect 14365 8128 14429 8132
rect 14445 8188 14509 8192
rect 14445 8132 14449 8188
rect 14449 8132 14505 8188
rect 14505 8132 14509 8188
rect 14445 8128 14509 8132
rect 14525 8188 14589 8192
rect 14525 8132 14529 8188
rect 14529 8132 14585 8188
rect 14585 8132 14589 8188
rect 14525 8128 14589 8132
rect 27618 8188 27682 8192
rect 27618 8132 27622 8188
rect 27622 8132 27678 8188
rect 27678 8132 27682 8188
rect 27618 8128 27682 8132
rect 27698 8188 27762 8192
rect 27698 8132 27702 8188
rect 27702 8132 27758 8188
rect 27758 8132 27762 8188
rect 27698 8128 27762 8132
rect 27778 8188 27842 8192
rect 27778 8132 27782 8188
rect 27782 8132 27838 8188
rect 27838 8132 27842 8188
rect 27778 8128 27842 8132
rect 27858 8188 27922 8192
rect 27858 8132 27862 8188
rect 27862 8132 27918 8188
rect 27918 8132 27922 8188
rect 27858 8128 27922 8132
rect 39620 7652 39684 7716
rect 7618 7644 7682 7648
rect 7618 7588 7622 7644
rect 7622 7588 7678 7644
rect 7678 7588 7682 7644
rect 7618 7584 7682 7588
rect 7698 7644 7762 7648
rect 7698 7588 7702 7644
rect 7702 7588 7758 7644
rect 7758 7588 7762 7644
rect 7698 7584 7762 7588
rect 7778 7644 7842 7648
rect 7778 7588 7782 7644
rect 7782 7588 7838 7644
rect 7838 7588 7842 7644
rect 7778 7584 7842 7588
rect 7858 7644 7922 7648
rect 7858 7588 7862 7644
rect 7862 7588 7918 7644
rect 7918 7588 7922 7644
rect 7858 7584 7922 7588
rect 20952 7644 21016 7648
rect 20952 7588 20956 7644
rect 20956 7588 21012 7644
rect 21012 7588 21016 7644
rect 20952 7584 21016 7588
rect 21032 7644 21096 7648
rect 21032 7588 21036 7644
rect 21036 7588 21092 7644
rect 21092 7588 21096 7644
rect 21032 7584 21096 7588
rect 21112 7644 21176 7648
rect 21112 7588 21116 7644
rect 21116 7588 21172 7644
rect 21172 7588 21176 7644
rect 21112 7584 21176 7588
rect 21192 7644 21256 7648
rect 21192 7588 21196 7644
rect 21196 7588 21252 7644
rect 21252 7588 21256 7644
rect 21192 7584 21256 7588
rect 34285 7644 34349 7648
rect 34285 7588 34289 7644
rect 34289 7588 34345 7644
rect 34345 7588 34349 7644
rect 34285 7584 34349 7588
rect 34365 7644 34429 7648
rect 34365 7588 34369 7644
rect 34369 7588 34425 7644
rect 34425 7588 34429 7644
rect 34365 7584 34429 7588
rect 34445 7644 34509 7648
rect 34445 7588 34449 7644
rect 34449 7588 34505 7644
rect 34505 7588 34509 7644
rect 34445 7584 34509 7588
rect 34525 7644 34589 7648
rect 34525 7588 34529 7644
rect 34529 7588 34585 7644
rect 34585 7588 34589 7644
rect 34525 7584 34589 7588
rect 39620 7380 39684 7444
rect 14285 7100 14349 7104
rect 14285 7044 14289 7100
rect 14289 7044 14345 7100
rect 14345 7044 14349 7100
rect 14285 7040 14349 7044
rect 14365 7100 14429 7104
rect 14365 7044 14369 7100
rect 14369 7044 14425 7100
rect 14425 7044 14429 7100
rect 14365 7040 14429 7044
rect 14445 7100 14509 7104
rect 14445 7044 14449 7100
rect 14449 7044 14505 7100
rect 14505 7044 14509 7100
rect 14445 7040 14509 7044
rect 14525 7100 14589 7104
rect 14525 7044 14529 7100
rect 14529 7044 14585 7100
rect 14585 7044 14589 7100
rect 14525 7040 14589 7044
rect 27618 7100 27682 7104
rect 27618 7044 27622 7100
rect 27622 7044 27678 7100
rect 27678 7044 27682 7100
rect 27618 7040 27682 7044
rect 27698 7100 27762 7104
rect 27698 7044 27702 7100
rect 27702 7044 27758 7100
rect 27758 7044 27762 7100
rect 27698 7040 27762 7044
rect 27778 7100 27842 7104
rect 27778 7044 27782 7100
rect 27782 7044 27838 7100
rect 27838 7044 27842 7100
rect 27778 7040 27842 7044
rect 27858 7100 27922 7104
rect 27858 7044 27862 7100
rect 27862 7044 27918 7100
rect 27918 7044 27922 7100
rect 27858 7040 27922 7044
rect 7618 6556 7682 6560
rect 7618 6500 7622 6556
rect 7622 6500 7678 6556
rect 7678 6500 7682 6556
rect 7618 6496 7682 6500
rect 7698 6556 7762 6560
rect 7698 6500 7702 6556
rect 7702 6500 7758 6556
rect 7758 6500 7762 6556
rect 7698 6496 7762 6500
rect 7778 6556 7842 6560
rect 7778 6500 7782 6556
rect 7782 6500 7838 6556
rect 7838 6500 7842 6556
rect 7778 6496 7842 6500
rect 7858 6556 7922 6560
rect 7858 6500 7862 6556
rect 7862 6500 7918 6556
rect 7918 6500 7922 6556
rect 7858 6496 7922 6500
rect 20952 6556 21016 6560
rect 20952 6500 20956 6556
rect 20956 6500 21012 6556
rect 21012 6500 21016 6556
rect 20952 6496 21016 6500
rect 21032 6556 21096 6560
rect 21032 6500 21036 6556
rect 21036 6500 21092 6556
rect 21092 6500 21096 6556
rect 21032 6496 21096 6500
rect 21112 6556 21176 6560
rect 21112 6500 21116 6556
rect 21116 6500 21172 6556
rect 21172 6500 21176 6556
rect 21112 6496 21176 6500
rect 21192 6556 21256 6560
rect 21192 6500 21196 6556
rect 21196 6500 21252 6556
rect 21252 6500 21256 6556
rect 21192 6496 21256 6500
rect 34285 6556 34349 6560
rect 34285 6500 34289 6556
rect 34289 6500 34345 6556
rect 34345 6500 34349 6556
rect 34285 6496 34349 6500
rect 34365 6556 34429 6560
rect 34365 6500 34369 6556
rect 34369 6500 34425 6556
rect 34425 6500 34429 6556
rect 34365 6496 34429 6500
rect 34445 6556 34509 6560
rect 34445 6500 34449 6556
rect 34449 6500 34505 6556
rect 34505 6500 34509 6556
rect 34445 6496 34509 6500
rect 34525 6556 34589 6560
rect 34525 6500 34529 6556
rect 34529 6500 34585 6556
rect 34585 6500 34589 6556
rect 34525 6496 34589 6500
rect 60 6020 124 6084
rect 14285 6012 14349 6016
rect 14285 5956 14289 6012
rect 14289 5956 14345 6012
rect 14345 5956 14349 6012
rect 14285 5952 14349 5956
rect 14365 6012 14429 6016
rect 14365 5956 14369 6012
rect 14369 5956 14425 6012
rect 14425 5956 14429 6012
rect 14365 5952 14429 5956
rect 14445 6012 14509 6016
rect 14445 5956 14449 6012
rect 14449 5956 14505 6012
rect 14505 5956 14509 6012
rect 14445 5952 14509 5956
rect 14525 6012 14589 6016
rect 14525 5956 14529 6012
rect 14529 5956 14585 6012
rect 14585 5956 14589 6012
rect 14525 5952 14589 5956
rect 27618 6012 27682 6016
rect 27618 5956 27622 6012
rect 27622 5956 27678 6012
rect 27678 5956 27682 6012
rect 27618 5952 27682 5956
rect 27698 6012 27762 6016
rect 27698 5956 27702 6012
rect 27702 5956 27758 6012
rect 27758 5956 27762 6012
rect 27698 5952 27762 5956
rect 27778 6012 27842 6016
rect 27778 5956 27782 6012
rect 27782 5956 27838 6012
rect 27838 5956 27842 6012
rect 27778 5952 27842 5956
rect 27858 6012 27922 6016
rect 27858 5956 27862 6012
rect 27862 5956 27918 6012
rect 27918 5956 27922 6012
rect 27858 5952 27922 5956
rect 60 5748 124 5812
rect 7618 5468 7682 5472
rect 7618 5412 7622 5468
rect 7622 5412 7678 5468
rect 7678 5412 7682 5468
rect 7618 5408 7682 5412
rect 7698 5468 7762 5472
rect 7698 5412 7702 5468
rect 7702 5412 7758 5468
rect 7758 5412 7762 5468
rect 7698 5408 7762 5412
rect 7778 5468 7842 5472
rect 7778 5412 7782 5468
rect 7782 5412 7838 5468
rect 7838 5412 7842 5468
rect 7778 5408 7842 5412
rect 7858 5468 7922 5472
rect 7858 5412 7862 5468
rect 7862 5412 7918 5468
rect 7918 5412 7922 5468
rect 7858 5408 7922 5412
rect 20952 5468 21016 5472
rect 20952 5412 20956 5468
rect 20956 5412 21012 5468
rect 21012 5412 21016 5468
rect 20952 5408 21016 5412
rect 21032 5468 21096 5472
rect 21032 5412 21036 5468
rect 21036 5412 21092 5468
rect 21092 5412 21096 5468
rect 21032 5408 21096 5412
rect 21112 5468 21176 5472
rect 21112 5412 21116 5468
rect 21116 5412 21172 5468
rect 21172 5412 21176 5468
rect 21112 5408 21176 5412
rect 21192 5468 21256 5472
rect 21192 5412 21196 5468
rect 21196 5412 21252 5468
rect 21252 5412 21256 5468
rect 21192 5408 21256 5412
rect 34285 5468 34349 5472
rect 34285 5412 34289 5468
rect 34289 5412 34345 5468
rect 34345 5412 34349 5468
rect 34285 5408 34349 5412
rect 34365 5468 34429 5472
rect 34365 5412 34369 5468
rect 34369 5412 34425 5468
rect 34425 5412 34429 5468
rect 34365 5408 34429 5412
rect 34445 5468 34509 5472
rect 34445 5412 34449 5468
rect 34449 5412 34505 5468
rect 34505 5412 34509 5468
rect 34445 5408 34509 5412
rect 34525 5468 34589 5472
rect 34525 5412 34529 5468
rect 34529 5412 34585 5468
rect 34585 5412 34589 5468
rect 34525 5408 34589 5412
rect 14285 4924 14349 4928
rect 14285 4868 14289 4924
rect 14289 4868 14345 4924
rect 14345 4868 14349 4924
rect 14285 4864 14349 4868
rect 14365 4924 14429 4928
rect 14365 4868 14369 4924
rect 14369 4868 14425 4924
rect 14425 4868 14429 4924
rect 14365 4864 14429 4868
rect 14445 4924 14509 4928
rect 14445 4868 14449 4924
rect 14449 4868 14505 4924
rect 14505 4868 14509 4924
rect 14445 4864 14509 4868
rect 14525 4924 14589 4928
rect 14525 4868 14529 4924
rect 14529 4868 14585 4924
rect 14585 4868 14589 4924
rect 14525 4864 14589 4868
rect 27618 4924 27682 4928
rect 27618 4868 27622 4924
rect 27622 4868 27678 4924
rect 27678 4868 27682 4924
rect 27618 4864 27682 4868
rect 27698 4924 27762 4928
rect 27698 4868 27702 4924
rect 27702 4868 27758 4924
rect 27758 4868 27762 4924
rect 27698 4864 27762 4868
rect 27778 4924 27842 4928
rect 27778 4868 27782 4924
rect 27782 4868 27838 4924
rect 27838 4868 27842 4924
rect 27778 4864 27842 4868
rect 27858 4924 27922 4928
rect 27858 4868 27862 4924
rect 27862 4868 27918 4924
rect 27918 4868 27922 4924
rect 27858 4864 27922 4868
rect 7618 4380 7682 4384
rect 7618 4324 7622 4380
rect 7622 4324 7678 4380
rect 7678 4324 7682 4380
rect 7618 4320 7682 4324
rect 7698 4380 7762 4384
rect 7698 4324 7702 4380
rect 7702 4324 7758 4380
rect 7758 4324 7762 4380
rect 7698 4320 7762 4324
rect 7778 4380 7842 4384
rect 7778 4324 7782 4380
rect 7782 4324 7838 4380
rect 7838 4324 7842 4380
rect 7778 4320 7842 4324
rect 7858 4380 7922 4384
rect 7858 4324 7862 4380
rect 7862 4324 7918 4380
rect 7918 4324 7922 4380
rect 7858 4320 7922 4324
rect 20952 4380 21016 4384
rect 20952 4324 20956 4380
rect 20956 4324 21012 4380
rect 21012 4324 21016 4380
rect 20952 4320 21016 4324
rect 21032 4380 21096 4384
rect 21032 4324 21036 4380
rect 21036 4324 21092 4380
rect 21092 4324 21096 4380
rect 21032 4320 21096 4324
rect 21112 4380 21176 4384
rect 21112 4324 21116 4380
rect 21116 4324 21172 4380
rect 21172 4324 21176 4380
rect 21112 4320 21176 4324
rect 21192 4380 21256 4384
rect 21192 4324 21196 4380
rect 21196 4324 21252 4380
rect 21252 4324 21256 4380
rect 21192 4320 21256 4324
rect 34285 4380 34349 4384
rect 34285 4324 34289 4380
rect 34289 4324 34345 4380
rect 34345 4324 34349 4380
rect 34285 4320 34349 4324
rect 34365 4380 34429 4384
rect 34365 4324 34369 4380
rect 34369 4324 34425 4380
rect 34425 4324 34429 4380
rect 34365 4320 34429 4324
rect 34445 4380 34509 4384
rect 34445 4324 34449 4380
rect 34449 4324 34505 4380
rect 34505 4324 34509 4380
rect 34445 4320 34509 4324
rect 34525 4380 34589 4384
rect 34525 4324 34529 4380
rect 34529 4324 34585 4380
rect 34585 4324 34589 4380
rect 34525 4320 34589 4324
rect 14285 3836 14349 3840
rect 14285 3780 14289 3836
rect 14289 3780 14345 3836
rect 14345 3780 14349 3836
rect 14285 3776 14349 3780
rect 14365 3836 14429 3840
rect 14365 3780 14369 3836
rect 14369 3780 14425 3836
rect 14425 3780 14429 3836
rect 14365 3776 14429 3780
rect 14445 3836 14509 3840
rect 14445 3780 14449 3836
rect 14449 3780 14505 3836
rect 14505 3780 14509 3836
rect 14445 3776 14509 3780
rect 14525 3836 14589 3840
rect 14525 3780 14529 3836
rect 14529 3780 14585 3836
rect 14585 3780 14589 3836
rect 14525 3776 14589 3780
rect 27618 3836 27682 3840
rect 27618 3780 27622 3836
rect 27622 3780 27678 3836
rect 27678 3780 27682 3836
rect 27618 3776 27682 3780
rect 27698 3836 27762 3840
rect 27698 3780 27702 3836
rect 27702 3780 27758 3836
rect 27758 3780 27762 3836
rect 27698 3776 27762 3780
rect 27778 3836 27842 3840
rect 27778 3780 27782 3836
rect 27782 3780 27838 3836
rect 27838 3780 27842 3836
rect 27778 3776 27842 3780
rect 27858 3836 27922 3840
rect 27858 3780 27862 3836
rect 27862 3780 27918 3836
rect 27918 3780 27922 3836
rect 27858 3776 27922 3780
rect 7618 3292 7682 3296
rect 7618 3236 7622 3292
rect 7622 3236 7678 3292
rect 7678 3236 7682 3292
rect 7618 3232 7682 3236
rect 7698 3292 7762 3296
rect 7698 3236 7702 3292
rect 7702 3236 7758 3292
rect 7758 3236 7762 3292
rect 7698 3232 7762 3236
rect 7778 3292 7842 3296
rect 7778 3236 7782 3292
rect 7782 3236 7838 3292
rect 7838 3236 7842 3292
rect 7778 3232 7842 3236
rect 7858 3292 7922 3296
rect 7858 3236 7862 3292
rect 7862 3236 7918 3292
rect 7918 3236 7922 3292
rect 7858 3232 7922 3236
rect 20952 3292 21016 3296
rect 20952 3236 20956 3292
rect 20956 3236 21012 3292
rect 21012 3236 21016 3292
rect 20952 3232 21016 3236
rect 21032 3292 21096 3296
rect 21032 3236 21036 3292
rect 21036 3236 21092 3292
rect 21092 3236 21096 3292
rect 21032 3232 21096 3236
rect 21112 3292 21176 3296
rect 21112 3236 21116 3292
rect 21116 3236 21172 3292
rect 21172 3236 21176 3292
rect 21112 3232 21176 3236
rect 21192 3292 21256 3296
rect 21192 3236 21196 3292
rect 21196 3236 21252 3292
rect 21252 3236 21256 3292
rect 21192 3232 21256 3236
rect 34285 3292 34349 3296
rect 34285 3236 34289 3292
rect 34289 3236 34345 3292
rect 34345 3236 34349 3292
rect 34285 3232 34349 3236
rect 34365 3292 34429 3296
rect 34365 3236 34369 3292
rect 34369 3236 34425 3292
rect 34425 3236 34429 3292
rect 34365 3232 34429 3236
rect 34445 3292 34509 3296
rect 34445 3236 34449 3292
rect 34449 3236 34505 3292
rect 34505 3236 34509 3292
rect 34445 3232 34509 3236
rect 34525 3292 34589 3296
rect 34525 3236 34529 3292
rect 34529 3236 34585 3292
rect 34585 3236 34589 3292
rect 34525 3232 34589 3236
rect 14285 2748 14349 2752
rect 14285 2692 14289 2748
rect 14289 2692 14345 2748
rect 14345 2692 14349 2748
rect 14285 2688 14349 2692
rect 14365 2748 14429 2752
rect 14365 2692 14369 2748
rect 14369 2692 14425 2748
rect 14425 2692 14429 2748
rect 14365 2688 14429 2692
rect 14445 2748 14509 2752
rect 14445 2692 14449 2748
rect 14449 2692 14505 2748
rect 14505 2692 14509 2748
rect 14445 2688 14509 2692
rect 14525 2748 14589 2752
rect 14525 2692 14529 2748
rect 14529 2692 14585 2748
rect 14585 2692 14589 2748
rect 14525 2688 14589 2692
rect 27618 2748 27682 2752
rect 27618 2692 27622 2748
rect 27622 2692 27678 2748
rect 27678 2692 27682 2748
rect 27618 2688 27682 2692
rect 27698 2748 27762 2752
rect 27698 2692 27702 2748
rect 27702 2692 27758 2748
rect 27758 2692 27762 2748
rect 27698 2688 27762 2692
rect 27778 2748 27842 2752
rect 27778 2692 27782 2748
rect 27782 2692 27838 2748
rect 27838 2692 27842 2748
rect 27778 2688 27842 2692
rect 27858 2748 27922 2752
rect 27858 2692 27862 2748
rect 27862 2692 27918 2748
rect 27918 2692 27922 2748
rect 27858 2688 27922 2692
rect 7618 2204 7682 2208
rect 7618 2148 7622 2204
rect 7622 2148 7678 2204
rect 7678 2148 7682 2204
rect 7618 2144 7682 2148
rect 7698 2204 7762 2208
rect 7698 2148 7702 2204
rect 7702 2148 7758 2204
rect 7758 2148 7762 2204
rect 7698 2144 7762 2148
rect 7778 2204 7842 2208
rect 7778 2148 7782 2204
rect 7782 2148 7838 2204
rect 7838 2148 7842 2204
rect 7778 2144 7842 2148
rect 7858 2204 7922 2208
rect 7858 2148 7862 2204
rect 7862 2148 7918 2204
rect 7918 2148 7922 2204
rect 7858 2144 7922 2148
rect 20952 2204 21016 2208
rect 20952 2148 20956 2204
rect 20956 2148 21012 2204
rect 21012 2148 21016 2204
rect 20952 2144 21016 2148
rect 21032 2204 21096 2208
rect 21032 2148 21036 2204
rect 21036 2148 21092 2204
rect 21092 2148 21096 2204
rect 21032 2144 21096 2148
rect 21112 2204 21176 2208
rect 21112 2148 21116 2204
rect 21116 2148 21172 2204
rect 21172 2148 21176 2204
rect 21112 2144 21176 2148
rect 21192 2204 21256 2208
rect 21192 2148 21196 2204
rect 21196 2148 21252 2204
rect 21252 2148 21256 2204
rect 21192 2144 21256 2148
rect 34285 2204 34349 2208
rect 34285 2148 34289 2204
rect 34289 2148 34345 2204
rect 34345 2148 34349 2204
rect 34285 2144 34349 2148
rect 34365 2204 34429 2208
rect 34365 2148 34369 2204
rect 34369 2148 34425 2204
rect 34425 2148 34429 2204
rect 34365 2144 34429 2148
rect 34445 2204 34509 2208
rect 34445 2148 34449 2204
rect 34449 2148 34505 2204
rect 34505 2148 34509 2204
rect 34445 2144 34509 2148
rect 34525 2204 34589 2208
rect 34525 2148 34529 2204
rect 34529 2148 34585 2204
rect 34585 2148 34589 2204
rect 34525 2144 34589 2148
<< metal4 >>
rect 7610 13088 7931 13648
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7931 13088
rect 7610 12000 7931 13024
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7931 12000
rect 7610 10912 7931 11936
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7931 10912
rect 7610 9824 7931 10848
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7931 9824
rect 7610 8736 7931 9760
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7931 8736
rect 7610 7648 7931 8672
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7931 7648
rect 7610 6560 7931 7584
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7931 6560
rect 59 6084 125 6085
rect 59 6020 60 6084
rect 124 6020 125 6084
rect 59 6019 125 6020
rect 62 5813 122 6019
rect 59 5812 125 5813
rect 59 5748 60 5812
rect 124 5748 125 5812
rect 59 5747 125 5748
rect 7610 5472 7931 6496
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7931 5472
rect 7610 4384 7931 5408
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7931 4384
rect 7610 3296 7931 4320
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7931 3296
rect 7610 2208 7931 3232
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7931 2208
rect 7610 2128 7931 2144
rect 14277 13632 14597 13648
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 12544 14597 13568
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 11456 14597 12480
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 10368 14597 11392
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 9280 14597 10304
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 8192 14597 9216
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 7104 14597 8128
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 6016 14597 7040
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 4928 14597 5952
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 3840 14597 4864
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 2752 14597 3776
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2128 14597 2688
rect 20944 13088 21264 13648
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 12000 21264 13024
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 10912 21264 11936
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 9824 21264 10848
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 8736 21264 9760
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 7648 21264 8672
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 6560 21264 7584
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 5472 21264 6496
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 4384 21264 5408
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 3296 21264 4320
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 2208 21264 3232
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2128 21264 2144
rect 27610 13632 27930 13648
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 12544 27930 13568
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 27610 11456 27930 12480
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 27610 10368 27930 11392
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 9280 27930 10304
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 27610 8192 27930 9216
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 7104 27930 8128
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 6016 27930 7040
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 4928 27930 5952
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 3840 27930 4864
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 27610 2752 27930 3776
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 27610 2128 27930 2688
rect 34277 13088 34597 13648
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 34277 12000 34597 13024
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 34277 10912 34597 11936
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 34277 9824 34597 10848
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 34277 8736 34597 9760
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 7648 34597 8672
rect 39619 7716 39685 7717
rect 39619 7652 39620 7716
rect 39684 7652 39685 7716
rect 39619 7651 39685 7652
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 6560 34597 7584
rect 39622 7445 39682 7651
rect 39619 7444 39685 7445
rect 39619 7380 39620 7444
rect 39684 7380 39685 7444
rect 39619 7379 39685 7380
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 34277 5472 34597 6496
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 34277 4384 34597 5408
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 34277 3296 34597 4320
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 2208 34597 3232
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 34277 2128 34597 2144
use scs8hd_decap_4  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use scs8hd_decap_6  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_13 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_12
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2024 0 1 2720
box -38 -48 314 592
use scs8hd_buf_1  _134_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1932 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_17
timestamp 1586364061
transform 1 0 2668 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_16
timestamp 1586364061
transform 1 0 2576 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_1_24
timestamp 1586364061
transform 1 0 3312 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 2852 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 2720
box -38 -48 314 592
use scs8hd_conb_1  _188_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3036 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_30
timestamp 1586364061
transform 1 0 3864 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_42 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4232 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_40
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_36
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_41
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_37
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_inv_8  _123_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 866 592
use scs8hd_inv_8  _071_
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_43
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_55
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__089__C
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 222 592
use scs8hd_or3_4  _089_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7084 0 -1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _088_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6900 0 1 2720
box -38 -48 866 592
use scs8hd_decap_3  FILLER_1_72
timestamp 1586364061
transform 1 0 7728 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_74
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_77
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_78
timestamp 1586364061
transform 1 0 8280 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use scs8hd_buf_1  _069_
timestamp 1586364061
transform 1 0 8556 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_84
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_1  _150_
timestamp 1586364061
transform 1 0 8648 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_88
timestamp 1586364061
transform 1 0 9200 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__C
timestamp 1586364061
transform 1 0 9384 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_44
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_1  _070_
timestamp 1586364061
transform 1 0 9936 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_107
timestamp 1586364061
transform 1 0 10948 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_101
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_103
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_99
timestamp 1586364061
transform 1 0 10212 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 10396 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 10764 0 1 2720
box -38 -48 222 592
use scs8hd_or3_4  _083_
timestamp 1586364061
transform 1 0 9568 0 1 2720
box -38 -48 866 592
use scs8hd_inv_8  _064_
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 866 592
use scs8hd_decap_4  FILLER_1_112
timestamp 1586364061
transform 1 0 11408 0 1 2720
box -38 -48 406 592
use scs8hd_buf_1  _081_
timestamp 1586364061
transform 1 0 11132 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_56
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_45
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_or3_4  _066_
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_132
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_128
timestamp 1586364061
transform 1 0 12880 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__125__D
timestamp 1586364061
transform 1 0 13248 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_1  _077_
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_140
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_136
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__C
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__B
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__C
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use scs8hd_or4_4  _125_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__D
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_157
timestamp 1586364061
transform 1 0 15548 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_153
timestamp 1586364061
transform 1 0 15180 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_160
timestamp 1586364061
transform 1 0 15824 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 15364 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_46
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_8  _092_
timestamp 1586364061
transform 1 0 14352 0 1 2720
box -38 -48 866 592
use scs8hd_nand3_4  _072_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16100 0 -1 2720
box -38 -48 1326 592
use scs8hd_inv_8  _106_
timestamp 1586364061
transform 1 0 16376 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 16192 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__C
timestamp 1586364061
transform 1 0 15916 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_177
timestamp 1586364061
transform 1 0 17388 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_1_161
timestamp 1586364061
transform 1 0 15916 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 17664 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_57
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_182
timestamp 1586364061
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_47
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 18216 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_188
timestamp 1586364061
transform 1 0 18400 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 18584 0 1 2720
box -38 -48 222 592
use scs8hd_or3_4  _149_
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use scs8hd_or3_4  _115_
timestamp 1586364061
transform 1 0 18768 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_205
timestamp 1586364061
transform 1 0 19964 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_201
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_200
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__B
timestamp 1586364061
transform 1 0 19688 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 19780 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_1  _074_
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_207
timestamp 1586364061
transform 1 0 20148 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 20148 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_or3_4  _107_
timestamp 1586364061
transform 1 0 20332 0 1 2720
box -38 -48 866 592
use scs8hd_decap_3  FILLER_1_222
timestamp 1586364061
transform 1 0 21528 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_218
timestamp 1586364061
transform 1 0 21160 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__C
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_48
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_231
timestamp 1586364061
transform 1 0 22356 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_227
timestamp 1586364061
transform 1 0 21988 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__C
timestamp 1586364061
transform 1 0 22172 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 21804 0 1 2720
box -38 -48 222 592
use scs8hd_or3_4  _171_
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 866 592
use scs8hd_inv_8  _154_
timestamp 1586364061
transform 1 0 21988 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_240
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_236
timestamp 1586364061
transform 1 0 22816 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_238
timestamp 1586364061
transform 1 0 23000 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 22540 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22724 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23920 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_58
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_49
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_8  _153_
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_0_258
timestamp 1586364061
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_266
timestamp 1586364061
transform 1 0 25576 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_263
timestamp 1586364061
transform 1 0 25300 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_259
timestamp 1586364061
transform 1 0 24932 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_262
timestamp 1586364061
transform 1 0 25208 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _195_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25576 0 -1 2720
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 24104 0 1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _173_
timestamp 1586364061
transform 1 0 25668 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_276
timestamp 1586364061
transform 1 0 26496 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_274
timestamp 1586364061
transform 1 0 26312 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_270
timestamp 1586364061
transform 1 0 25944 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 26496 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 26128 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_280
timestamp 1586364061
transform 1 0 26864 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_283
timestamp 1586364061
transform 1 0 27140 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_278
timestamp 1586364061
transform 1 0 26680 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 27324 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__B
timestamp 1586364061
transform 1 0 27048 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__B
timestamp 1586364061
transform 1 0 26680 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_50
timestamp 1586364061
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_nor2_4  _174_
timestamp 1586364061
transform 1 0 27232 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_293
timestamp 1586364061
transform 1 0 28060 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_287
timestamp 1586364061
transform 1 0 27508 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__B
timestamp 1586364061
transform 1 0 27692 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_301
timestamp 1586364061
transform 1 0 28796 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_297
timestamp 1586364061
transform 1 0 28428 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_300
timestamp 1586364061
transform 1 0 28704 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28612 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 28888 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__B
timestamp 1586364061
transform 1 0 28980 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28244 0 1 2720
box -38 -48 222 592
use scs8hd_nor2_4  _176_
timestamp 1586364061
transform 1 0 27876 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_0_308
timestamp 1586364061
transform 1 0 29440 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_304
timestamp 1586364061
transform 1 0 29072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 29256 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_59
timestamp 1586364061
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_51
timestamp 1586364061
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_1  _172_
timestamp 1586364061
transform 1 0 29716 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_319
timestamp 1586364061
transform 1 0 30452 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_315
timestamp 1586364061
transform 1 0 30084 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_318
timestamp 1586364061
transform 1 0 30360 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_314
timestamp 1586364061
transform 1 0 29992 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30268 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 30176 0 -1 2720
box -38 -48 222 592
use scs8hd_nor2_4  _177_
timestamp 1586364061
transform 1 0 29256 0 1 2720
box -38 -48 866 592
use scs8hd_conb_1  _180_
timestamp 1586364061
transform 1 0 30820 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30728 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31832 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31188 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_325
timestamp 1586364061
transform 1 0 31004 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_329 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 31372 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_326 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 31096 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_337
timestamp 1586364061
transform 1 0 32108 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_52
timestamp 1586364061
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33120 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32292 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32660 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_342
timestamp 1586364061
transform 1 0 32568 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_354
timestamp 1586364061
transform 1 0 33672 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_341
timestamp 1586364061
transform 1 0 32476 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_345
timestamp 1586364061
transform 1 0 32844 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_350
timestamp 1586364061
transform 1 0 33304 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_53
timestamp 1586364061
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_60
timestamp 1586364061
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_366
timestamp 1586364061
transform 1 0 34776 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_373
timestamp 1586364061
transform 1 0 35420 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_362
timestamp 1586364061
transform 1 0 34408 0 1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_367
timestamp 1586364061
transform 1 0 34868 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_385
timestamp 1586364061
transform 1 0 36524 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_379
timestamp 1586364061
transform 1 0 35972 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_391
timestamp 1586364061
transform 1 0 37076 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 38824 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 38824 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_54
timestamp 1586364061
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_397
timestamp 1586364061
transform 1 0 37628 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_3  FILLER_0_404
timestamp 1586364061
transform 1 0 38272 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_403
timestamp 1586364061
transform 1 0 38180 0 1 2720
box -38 -48 406 592
use scs8hd_nor2_4  _137_
timestamp 1586364061
transform 1 0 2116 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 1564 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1932 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_7
timestamp 1586364061
transform 1 0 1748 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_61
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 4232 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3128 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_20
timestamp 1586364061
transform 1 0 2944 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_24
timestamp 1586364061
transform 1 0 3312 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_30
timestamp 1586364061
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 222 592
use scs8hd_conb_1  _183_
timestamp 1586364061
transform 1 0 5888 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4876 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 4692 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_36
timestamp 1586364061
transform 1 0 4416 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 774 592
use scs8hd_nor2_4  _085_
timestamp 1586364061
transform 1 0 6900 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 6716 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 6348 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_55
timestamp 1586364061
transform 1 0 6164 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_59
timestamp 1586364061
transform 1 0 6532 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_1  _090_
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_72
timestamp 1586364061
transform 1 0 7728 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_6  FILLER_2_83
timestamp 1586364061
transform 1 0 8740 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_89
timestamp 1586364061
transform 1 0 9292 0 -1 3808
box -38 -48 130 592
use scs8hd_inv_8  _065_
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 866 592
use scs8hd_buf_1  _084_
timestamp 1586364061
transform 1 0 9752 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_62
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__080__C
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_97
timestamp 1586364061
transform 1 0 10028 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_101
timestamp 1586364061
transform 1 0 10396 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_104
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 130 592
use scs8hd_or3_4  _086_
timestamp 1586364061
transform 1 0 12328 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__066__C
timestamp 1586364061
transform 1 0 12144 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 11776 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_114
timestamp 1586364061
transform 1 0 11592 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_118
timestamp 1586364061
transform 1 0 11960 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_1  _067_
timestamp 1586364061
transform 1 0 13892 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 13708 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 13340 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_131
timestamp 1586364061
transform 1 0 13156 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_135
timestamp 1586364061
transform 1 0 13524 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_142
timestamp 1586364061
transform 1 0 14168 0 -1 3808
box -38 -48 222 592
use scs8hd_or4_4  _133_
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_63
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__133__C
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_146
timestamp 1586364061
transform 1 0 14536 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_150
timestamp 1586364061
transform 1 0 14904 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__141__C
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__C
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__D
timestamp 1586364061
transform 1 0 17112 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 16744 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_163
timestamp 1586364061
transform 1 0 16100 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_168
timestamp 1586364061
transform 1 0 16560 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_172
timestamp 1586364061
transform 1 0 16928 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_176
timestamp 1586364061
transform 1 0 17296 0 -1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _151_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 17664 0 -1 3808
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_64
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 19412 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 20332 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 19780 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_197
timestamp 1586364061
transform 1 0 19228 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_201
timestamp 1586364061
transform 1 0 19596 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_205
timestamp 1586364061
transform 1 0 19964 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_3  FILLER_2_211
timestamp 1586364061
transform 1 0 20516 0 -1 3808
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_1_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 21804 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21068 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21620 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_219
timestamp 1586364061
transform 1 0 21252 0 -1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23828 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_236
timestamp 1586364061
transform 1 0 22816 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_240
timestamp 1586364061
transform 1 0 23184 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_244
timestamp 1586364061
transform 1 0 23552 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24932 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_256
timestamp 1586364061
transform 1 0 24656 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_261
timestamp 1586364061
transform 1 0 25116 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_267
timestamp 1586364061
transform 1 0 25668 0 -1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _175_
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_65
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__173__B
timestamp 1586364061
transform 1 0 25852 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 26220 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_271
timestamp 1586364061
transform 1 0 26036 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_285
timestamp 1586364061
transform 1 0 27324 0 -1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28060 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27784 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_289
timestamp 1586364061
transform 1 0 27692 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_292
timestamp 1586364061
transform 1 0 27968 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_296
timestamp 1586364061
transform 1 0 28336 0 -1 3808
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29532 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29256 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_304
timestamp 1586364061
transform 1 0 29072 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_308
timestamp 1586364061
transform 1 0 29440 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_318
timestamp 1586364061
transform 1 0 30360 0 -1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32108 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_66
timestamp 1586364061
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__178__B
timestamp 1586364061
transform 1 0 30820 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_322
timestamp 1586364061
transform 1 0 30728 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_325
timestamp 1586364061
transform 1 0 31004 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_2_333
timestamp 1586364061
transform 1 0 31740 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33120 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_340
timestamp 1586364061
transform 1 0 32384 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_12  FILLER_2_351
timestamp 1586364061
transform 1 0 33396 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_363
timestamp 1586364061
transform 1 0 34500 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_375
timestamp 1586364061
transform 1 0 35604 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_387
timestamp 1586364061
transform 1 0 36708 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 38824 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_67
timestamp 1586364061
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_395
timestamp 1586364061
transform 1 0 37444 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_398
timestamp 1586364061
transform 1 0 37720 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_406
timestamp 1586364061
transform 1 0 38456 0 -1 3808
box -38 -48 130 592
use scs8hd_nor2_4  _136_
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_12
timestamp 1586364061
transform 1 0 2208 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_16
timestamp 1586364061
transform 1 0 2576 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2944 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 4048 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2760 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_29
timestamp 1586364061
transform 1 0 3772 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_3_34
timestamp 1586364061
transform 1 0 4232 0 1 3808
box -38 -48 314 592
use scs8hd_nor2_4  _139_
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 5704 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 4508 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_48
timestamp 1586364061
transform 1 0 5520 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_52
timestamp 1586364061
transform 1 0 5888 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_68
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6072 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_56
timestamp 1586364061
transform 1 0 6256 0 1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_3_71
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 406 592
use scs8hd_inv_8  _079_
timestamp 1586364061
transform 1 0 8924 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 8740 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_77
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_81
timestamp 1586364061
transform 1 0 8556 0 1 3808
box -38 -48 222 592
use scs8hd_or3_4  _080_
timestamp 1586364061
transform 1 0 10488 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 10304 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 9936 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_94
timestamp 1586364061
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 222 592
use scs8hd_or3_4  _076_
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_69
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__076__C
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_111
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_115
timestamp 1586364061
transform 1 0 11684 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__C
timestamp 1586364061
transform 1 0 13892 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_136
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_141
timestamp 1586364061
transform 1 0 14076 0 1 3808
box -38 -48 222 592
use scs8hd_or3_4  _093_
timestamp 1586364061
transform 1 0 14812 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 14260 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_145
timestamp 1586364061
transform 1 0 14444 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_158
timestamp 1586364061
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use scs8hd_or4_4  _141_
timestamp 1586364061
transform 1 0 16376 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__C
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_162
timestamp 1586364061
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_175
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _152_
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_70
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__152__D
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 20792 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 19780 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 20148 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_201
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_205
timestamp 1586364061
transform 1 0 19964 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_209
timestamp 1586364061
transform 1 0 20332 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_213
timestamp 1586364061
transform 1 0 20700 0 1 3808
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 20976 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 22172 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_227
timestamp 1586364061
transform 1 0 21988 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_231
timestamp 1586364061
transform 1 0 22356 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_71
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22540 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_235
timestamp 1586364061
transform 1 0 22724 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_240
timestamp 1586364061
transform 1 0 23184 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 25576 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 25392 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24656 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_254
timestamp 1586364061
transform 1 0 24472 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_258
timestamp 1586364061
transform 1 0 24840 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_262
timestamp 1586364061
transform 1 0 25208 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27324 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 26772 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27140 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_277
timestamp 1586364061
transform 1 0 26588 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_281
timestamp 1586364061
transform 1 0 26956 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 28336 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28980 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_294
timestamp 1586364061
transform 1 0 28152 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_298
timestamp 1586364061
transform 1 0 28520 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_302
timestamp 1586364061
transform 1 0 28888 0 1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_72
timestamp 1586364061
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 30268 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 30636 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_315
timestamp 1586364061
transform 1 0 30084 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_319
timestamp 1586364061
transform 1 0 30452 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _178_
timestamp 1586364061
transform 1 0 30820 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32108 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_332
timestamp 1586364061
transform 1 0 31648 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_336
timestamp 1586364061
transform 1 0 32016 0 1 3808
box -38 -48 130 592
use scs8hd_conb_1  _182_
timestamp 1586364061
transform 1 0 32384 0 1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33396 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33856 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32844 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_339
timestamp 1586364061
transform 1 0 32292 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_343
timestamp 1586364061
transform 1 0 32660 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_347
timestamp 1586364061
transform 1 0 33028 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_354
timestamp 1586364061
transform 1 0 33672 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35052 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 34224 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_358
timestamp 1586364061
transform 1 0 34040 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_362
timestamp 1586364061
transform 1 0 34408 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_367
timestamp 1586364061
transform 1 0 34868 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_371
timestamp 1586364061
transform 1 0 35236 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_383
timestamp 1586364061
transform 1 0 36340 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 38824 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_395
timestamp 1586364061
transform 1 0 37444 0 1 3808
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_5_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 1050 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2024 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_7
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 314 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 5612 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__075__B
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_41
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_46
timestamp 1586364061
transform 1 0 5336 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_60
timestamp 1586364061
transform 1 0 6624 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_64
timestamp 1586364061
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 406 592
use scs8hd_nor2_4  _091_
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_72
timestamp 1586364061
transform 1 0 7728 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_88
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 406 592
use scs8hd_buf_1  _087_
timestamp 1586364061
transform 1 0 10028 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_100
timestamp 1586364061
transform 1 0 10304 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_104
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11040 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 12052 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_121
timestamp 1586364061
transform 1 0 12236 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _078_
timestamp 1586364061
transform 1 0 12788 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 13800 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_125
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_136
timestamp 1586364061
transform 1 0 13616 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_140
timestamp 1586364061
transform 1 0 13984 0 -1 4896
box -38 -48 590 592
use scs8hd_or2_4  _124_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 14536 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_148
timestamp 1586364061
transform 1 0 14720 0 -1 4896
box -38 -48 314 592
use scs8hd_or3_4  _155_
timestamp 1586364061
transform 1 0 16652 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__141__D
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_161
timestamp 1586364061
transform 1 0 15916 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_165
timestamp 1586364061
transform 1 0 16284 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_168
timestamp 1586364061
transform 1 0 16560 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 222 592
use scs8hd_or3_4  _163_
timestamp 1586364061
transform 1 0 18768 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__C
timestamp 1586364061
transform 1 0 18400 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 17664 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_182
timestamp 1586364061
transform 1 0 17848 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_186
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 19780 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 20148 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_201
timestamp 1586364061
transform 1 0 19596 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_205
timestamp 1586364061
transform 1 0 19964 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_209
timestamp 1586364061
transform 1 0 20332 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_213
timestamp 1586364061
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_5_.latch
timestamp 1586364061
transform 1 0 21620 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 21436 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23368 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23184 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_234
timestamp 1586364061
transform 1 0 22632 0 -1 4896
box -38 -48 590 592
use scs8hd_inv_1  mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24932 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25668 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_4  FILLER_4_262
timestamp 1586364061
transform 1 0 25208 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_266
timestamp 1586364061
transform 1 0 25576 0 -1 4896
box -38 -48 130 592
use scs8hd_buf_1  _098_
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27232 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_269
timestamp 1586364061
transform 1 0 25852 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_4  FILLER_4_279
timestamp 1586364061
transform 1 0 26772 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_283
timestamp 1586364061
transform 1 0 27140 0 -1 4896
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 27784 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 27600 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_286
timestamp 1586364061
transform 1 0 27416 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_301
timestamp 1586364061
transform 1 0 28796 0 -1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 29532 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29256 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_305
timestamp 1586364061
transform 1 0 29164 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_308
timestamp 1586364061
transform 1 0 29440 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_320
timestamp 1586364061
transform 1 0 30544 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32108 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30728 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_324
timestamp 1586364061
transform 1 0 30912 0 -1 4896
box -38 -48 1142 592
use scs8hd_buf_1  _116_
timestamp 1586364061
transform 1 0 33672 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33120 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_346
timestamp 1586364061
transform 1 0 32936 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_350
timestamp 1586364061
transform 1 0 33304 0 -1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34684 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_357
timestamp 1586364061
transform 1 0 33948 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_12  FILLER_4_368
timestamp 1586364061
transform 1 0 34960 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_380
timestamp 1586364061
transform 1 0 36064 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_4_392
timestamp 1586364061
transform 1 0 37168 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 38824 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_396
timestamp 1586364061
transform 1 0 37536 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_398
timestamp 1586364061
transform 1 0 37720 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_406
timestamp 1586364061
transform 1 0 38456 0 -1 4896
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_4_.latch
timestamp 1586364061
transform 1 0 2392 0 1 4896
box -38 -48 1050 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_6
timestamp 1586364061
transform 1 0 1656 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_10
timestamp 1586364061
transform 1 0 2024 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3956 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_25
timestamp 1586364061
transform 1 0 3404 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_29
timestamp 1586364061
transform 1 0 3772 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _075_
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_36
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_40
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7176 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6992 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6440 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_60
timestamp 1586364061
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8924 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8740 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_77
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_81
timestamp 1586364061
transform 1 0 8556 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_94
timestamp 1586364061
transform 1 0 9752 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_99
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 12604 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 13984 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_138
timestamp 1586364061
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_142
timestamp 1586364061
transform 1 0 14168 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _095_
timestamp 1586364061
transform 1 0 14536 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 15548 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 14352 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_155
timestamp 1586364061
transform 1 0 15364 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 16100 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 15916 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__B
timestamp 1586364061
transform 1 0 17296 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_174
timestamp 1586364061
transform 1 0 17112 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_178
timestamp 1586364061
transform 1 0 17480 0 1 4896
box -38 -48 314 592
use scs8hd_nor2_4  _099_
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_193
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 406 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 19688 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 20700 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_199
timestamp 1586364061
transform 1 0 19412 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_211
timestamp 1586364061
transform 1 0 20516 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_4_.latch
timestamp 1586364061
transform 1 0 21252 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 21068 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_215
timestamp 1586364061
transform 1 0 20884 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_230
timestamp 1586364061
transform 1 0 22264 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_234
timestamp 1586364061
transform 1 0 22632 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_240
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 25668 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 25484 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 25116 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_254
timestamp 1586364061
transform 1 0 24472 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_259
timestamp 1586364061
transform 1 0 24932 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_263
timestamp 1586364061
transform 1 0 25300 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27048 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_278
timestamp 1586364061
transform 1 0 26680 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_284
timestamp 1586364061
transform 1 0 27232 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _169_
timestamp 1586364061
transform 1 0 27600 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 27416 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28980 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28612 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_297
timestamp 1586364061
transform 1 0 28428 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_301
timestamp 1586364061
transform 1 0 28796 0 1 4896
box -38 -48 222 592
use scs8hd_buf_1  _164_
timestamp 1586364061
transform 1 0 29256 0 1 4896
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 30636 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 29716 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 30452 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 30084 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_309
timestamp 1586364061
transform 1 0 29532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_313
timestamp 1586364061
transform 1 0 29900 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_317
timestamp 1586364061
transform 1 0 30268 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32200 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31832 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_332
timestamp 1586364061
transform 1 0 31648 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_336
timestamp 1586364061
transform 1 0 32016 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32384 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33764 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33396 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_349
timestamp 1586364061
transform 1 0 33212 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_353
timestamp 1586364061
transform 1 0 33580 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35420 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34132 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_357
timestamp 1586364061
transform 1 0 33948 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_361
timestamp 1586364061
transform 1 0 34316 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_365
timestamp 1586364061
transform 1 0 34684 0 1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_5_367
timestamp 1586364061
transform 1 0 34868 0 1 4896
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35880 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_376
timestamp 1586364061
transform 1 0 35696 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_380
timestamp 1586364061
transform 1 0 36064 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_392
timestamp 1586364061
transform 1 0 37168 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 38824 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_404
timestamp 1586364061
transform 1 0 38272 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_6
timestamp 1586364061
transform 1 0 1656 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_8
timestamp 1586364061
transform 1 0 1840 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1656 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_10
timestamp 1586364061
transform 1 0 2024 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2024 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_3_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 5984
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_7_23
timestamp 1586364061
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3404 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 3772 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 3956 0 1 5984
box -38 -48 1050 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_41
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_4  FILLER_6_51
timestamp 1586364061
transform 1 0 5796 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_42
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_46
timestamp 1586364061
transform 1 0 5336 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_55
timestamp 1586364061
transform 1 0 6164 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_67
timestamp 1586364061
transform 1 0 7268 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 7084 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6440 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 7268 0 1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8464 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_78
timestamp 1586364061
transform 1 0 8280 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_82
timestamp 1586364061
transform 1 0 8648 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_90
timestamp 1586364061
transform 1 0 9384 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_97
timestamp 1586364061
transform 1 0 10028 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9568 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_105
timestamp 1586364061
transform 1 0 10764 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10948 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9752 0 1 5984
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_7_115
timestamp 1586364061
transform 1 0 11684 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_109
timestamp 1586364061
transform 1 0 11132 0 1 5984
box -38 -48 406 592
use scs8hd_decap_6  FILLER_6_110
timestamp 1586364061
transform 1 0 11224 0 -1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 11500 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_119
timestamp 1586364061
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 11868 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11960 0 -1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _082_
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_132
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_131
timestamp 1586364061
transform 1 0 13156 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_127
timestamp 1586364061
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13340 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_140
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_136
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_135
timestamp 1586364061
transform 1 0 13524 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _097_
timestamp 1586364061
transform 1 0 13616 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 14260 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_160
timestamp 1586364061
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_156
timestamp 1586364061
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15548 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_buf_1  _094_
timestamp 1586364061
transform 1 0 15732 0 -1 5984
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 14444 0 1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 16192 0 1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16744 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_162
timestamp 1586364061
transform 1 0 16008 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_168
timestamp 1586364061
transform 1 0 16560 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_186
timestamp 1586364061
transform 1 0 18216 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_183
timestamp 1586364061
transform 1 0 17940 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_179
timestamp 1586364061
transform 1 0 17572 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 18032 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_193
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_194
timestamp 1586364061
transform 1 0 18952 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18768 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18400 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 19228 0 -1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _145_
timestamp 1586364061
transform 1 0 20148 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 19964 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_206
timestamp 1586364061
transform 1 0 20056 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_4  FILLER_7_197
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_203
timestamp 1586364061
transform 1 0 19780 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 21712 0 1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_3_.latch
timestamp 1586364061
transform 1 0 21436 0 -1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21252 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21252 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_7_216
timestamp 1586364061
transform 1 0 20976 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_221
timestamp 1586364061
transform 1 0 21436 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_239
timestamp 1586364061
transform 1 0 23092 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_235
timestamp 1586364061
transform 1 0 22724 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_236
timestamp 1586364061
transform 1 0 22816 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_232
timestamp 1586364061
transform 1 0 22448 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22632 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 22908 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_249
timestamp 1586364061
transform 1 0 24012 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23184 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_258
timestamp 1586364061
transform 1 0 24840 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_254
timestamp 1586364061
transform 1 0 24472 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_253
timestamp 1586364061
transform 1 0 24380 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24564 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_266
timestamp 1586364061
transform 1 0 25576 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25024 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25208 0 1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _170_
timestamp 1586364061
transform 1 0 24748 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_1  FILLER_7_275
timestamp 1586364061
transform 1 0 26404 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_271
timestamp 1586364061
transform 1 0 26036 0 1 5984
box -38 -48 406 592
use scs8hd_decap_6  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_274
timestamp 1586364061
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26496 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_282
timestamp 1586364061
transform 1 0 27048 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_278
timestamp 1586364061
transform 1 0 26680 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26864 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 27324 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27048 0 -1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 27508 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28704 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28704 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_291
timestamp 1586364061
transform 1 0 27876 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_299
timestamp 1586364061
transform 1 0 28612 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_6_302
timestamp 1586364061
transform 1 0 28888 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_4  FILLER_7_296
timestamp 1586364061
transform 1 0 28336 0 1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_7_302
timestamp 1586364061
transform 1 0 28888 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_309
timestamp 1586364061
transform 1 0 29532 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_308
timestamp 1586364061
transform 1 0 29440 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 29716 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use scs8hd_buf_1  _100_
timestamp 1586364061
transform 1 0 29256 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_7_319
timestamp 1586364061
transform 1 0 30452 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_313
timestamp 1586364061
transform 1 0 29900 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_320
timestamp 1586364061
transform 1 0 30544 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 30268 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30544 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 29532 0 -1 5984
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_7_329
timestamp 1586364061
transform 1 0 31372 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_328
timestamp 1586364061
transform 1 0 31280 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_6_324
timestamp 1586364061
transform 1 0 30912 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31096 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30728 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_333
timestamp 1586364061
transform 1 0 31740 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 31556 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 31924 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32108 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_5_.latch
timestamp 1586364061
transform 1 0 32108 0 1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33764 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33304 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33672 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_346
timestamp 1586364061
transform 1 0 32936 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_354
timestamp 1586364061
transform 1 0 33672 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_348
timestamp 1586364061
transform 1 0 33120 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_352
timestamp 1586364061
transform 1 0 33488 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_356
timestamp 1586364061
transform 1 0 33856 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_362
timestamp 1586364061
transform 1 0 34408 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_364
timestamp 1586364061
transform 1 0 34592 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34224 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_368
timestamp 1586364061
transform 1 0 34960 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35144 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34776 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use scs8hd_conb_1  _186_
timestamp 1586364061
transform 1 0 35328 0 -1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_380
timestamp 1586364061
transform 1 0 36064 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_376
timestamp 1586364061
transform 1 0 35696 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36248 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35880 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_387
timestamp 1586364061
transform 1 0 36708 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_387
timestamp 1586364061
transform 1 0 36708 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36892 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36432 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_391
timestamp 1586364061
transform 1 0 37076 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_375
timestamp 1586364061
transform 1 0 35604 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 38824 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 38824 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_395
timestamp 1586364061
transform 1 0 37444 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_398
timestamp 1586364061
transform 1 0 37720 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_406
timestamp 1586364061
transform 1 0 38456 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_403
timestamp 1586364061
transform 1 0 38180 0 1 5984
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1840 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_6
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_10
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5612 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_8_41
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_58
timestamp 1586364061
transform 1 0 6440 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  FILLER_8_64
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_8_69
timestamp 1586364061
transform 1 0 7452 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_97
timestamp 1586364061
transform 1 0 10028 0 -1 7072
box -38 -48 314 592
use scs8hd_nor2_4  _162_
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_8_109
timestamp 1586364061
transform 1 0 11132 0 -1 7072
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 12880 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13248 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_126
timestamp 1586364061
transform 1 0 12696 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_130
timestamp 1586364061
transform 1 0 13064 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16928 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16284 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_163
timestamp 1586364061
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_167
timestamp 1586364061
transform 1 0 16468 0 -1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_181
timestamp 1586364061
transform 1 0 17756 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_186
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19504 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_198
timestamp 1586364061
transform 1 0 19320 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_6  FILLER_8_208
timestamp 1586364061
transform 1 0 20240 0 -1 7072
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 22264 0 -1 7072
box -38 -48 1050 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21252 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 21712 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 21068 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22080 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_222
timestamp 1586364061
transform 1 0 21528 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_226
timestamp 1586364061
transform 1 0 21896 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24012 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23644 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_241
timestamp 1586364061
transform 1 0 23276 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_247
timestamp 1586364061
transform 1 0 23828 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25208 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25576 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_258
timestamp 1586364061
transform 1 0 24840 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_264
timestamp 1586364061
transform 1 0 25392 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_8_268
timestamp 1586364061
transform 1 0 25760 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_274
timestamp 1586364061
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_285
timestamp 1586364061
transform 1 0 27324 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28704 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 27508 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 28336 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_289
timestamp 1586364061
transform 1 0 27692 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_295
timestamp 1586364061
transform 1 0 28244 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_298
timestamp 1586364061
transform 1 0 28520 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 30268 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30084 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_309
timestamp 1586364061
transform 1 0 29532 0 -1 7072
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_4_.latch
timestamp 1586364061
transform 1 0 32108 0 -1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31740 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_328
timestamp 1586364061
transform 1 0 31280 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_332
timestamp 1586364061
transform 1 0 31648 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_335
timestamp 1586364061
transform 1 0 31924 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_348
timestamp 1586364061
transform 1 0 33120 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_356
timestamp 1586364061
transform 1 0 33856 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34224 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35236 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34040 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_369
timestamp 1586364061
transform 1 0 35052 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_373
timestamp 1586364061
transform 1 0 35420 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35788 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_8_386
timestamp 1586364061
transform 1 0 36616 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 38824 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_394
timestamp 1586364061
transform 1 0 37352 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_398
timestamp 1586364061
transform 1 0 37720 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_406
timestamp 1586364061
transform 1 0 38456 0 -1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2300 0 1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_9
timestamp 1586364061
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_2_.latch
timestamp 1586364061
transform 1 0 3864 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 3680 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 3312 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_22
timestamp 1586364061
transform 1 0 3128 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_26
timestamp 1586364061
transform 1 0 3496 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5428 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5060 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_41
timestamp 1586364061
transform 1 0 4876 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_45
timestamp 1586364061
transform 1 0 5244 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_52
timestamp 1586364061
transform 1 0 5888 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _130_
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6072 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_56
timestamp 1586364061
transform 1 0 6256 0 1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_9_71
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8832 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8648 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_77
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_81
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 130 592
use scs8hd_nor2_4  _160_
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_95
timestamp 1586364061
transform 1 0 9844 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_99
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_112
timestamp 1586364061
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_116
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_120
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13340 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12788 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_129
timestamp 1586364061
transform 1 0 12972 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14536 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14904 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_144
timestamp 1586364061
transform 1 0 14352 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_148
timestamp 1586364061
transform 1 0 14720 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_152
timestamp 1586364061
transform 1 0 15088 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_156
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 16928 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17296 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_170
timestamp 1586364061
transform 1 0 16744 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_174
timestamp 1586364061
transform 1 0 17112 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_178
timestamp 1586364061
transform 1 0 17480 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_193
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 20056 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 19872 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_197
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_201
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_2_.latch
timestamp 1586364061
transform 1 0 21620 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 21436 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_215
timestamp 1586364061
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_219
timestamp 1586364061
transform 1 0 21252 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_234
timestamp 1586364061
transform 1 0 22632 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_238
timestamp 1586364061
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_242
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25208 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_254
timestamp 1586364061
transform 1 0 24472 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_258
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 26496 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 26864 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_271
timestamp 1586364061
transform 1 0 26036 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_275
timestamp 1586364061
transform 1 0 26404 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_278
timestamp 1586364061
transform 1 0 26680 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_282
timestamp 1586364061
transform 1 0 27048 0 1 7072
box -38 -48 406 592
use scs8hd_nor2_4  _118_
timestamp 1586364061
transform 1 0 27600 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 27416 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 28980 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 28612 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_297
timestamp 1586364061
transform 1 0 28428 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_301
timestamp 1586364061
transform 1 0 28796 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 29256 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 30268 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30636 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_315
timestamp 1586364061
transform 1 0 30084 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_319
timestamp 1586364061
transform 1 0 30452 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_3_.latch
timestamp 1586364061
transform 1 0 31740 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 31556 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31188 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_323
timestamp 1586364061
transform 1 0 30820 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_329
timestamp 1586364061
transform 1 0 31372 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33764 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 32936 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33580 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_344
timestamp 1586364061
transform 1 0 32752 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_348
timestamp 1586364061
transform 1 0 33120 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_352
timestamp 1586364061
transform 1 0 33488 0 1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34224 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_358
timestamp 1586364061
transform 1 0 34040 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_362
timestamp 1586364061
transform 1 0 34408 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _197_
timestamp 1586364061
transform 1 0 36432 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 36984 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35880 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36248 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_376
timestamp 1586364061
transform 1 0 35696 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_380
timestamp 1586364061
transform 1 0 36064 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_388
timestamp 1586364061
transform 1 0 36800 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_392
timestamp 1586364061
transform 1 0 37168 0 1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37536 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 38824 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37996 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_399
timestamp 1586364061
transform 1 0 37812 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_403
timestamp 1586364061
transform 1 0 38180 0 1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1656 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_8
timestamp 1586364061
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_2  _198_
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_21
timestamp 1586364061
transform 1 0 3036 0 -1 8160
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5428 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4600 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_36
timestamp 1586364061
transform 1 0 4416 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_40
timestamp 1586364061
transform 1 0 4784 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_46
timestamp 1586364061
transform 1 0 5336 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_58
timestamp 1586364061
transform 1 0 6440 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_10_70
timestamp 1586364061
transform 1 0 7544 0 -1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use scs8hd_fill_1  FILLER_10_74
timestamp 1586364061
transform 1 0 7912 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_102
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_106
timestamp 1586364061
transform 1 0 10856 0 -1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _161_
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_119
timestamp 1586364061
transform 1 0 12052 0 -1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13432 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_125
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_133
timestamp 1586364061
transform 1 0 13340 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_149
timestamp 1586364061
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 16836 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_163
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_10_168
timestamp 1586364061
transform 1 0 16560 0 -1 8160
box -38 -48 314 592
use scs8hd_nor2_4  _114_
timestamp 1586364061
transform 1 0 18952 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18768 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_182
timestamp 1586364061
transform 1 0 17848 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_186
timestamp 1586364061
transform 1 0 18216 0 -1 8160
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19964 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_203
timestamp 1586364061
transform 1 0 19780 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_207
timestamp 1586364061
transform 1 0 20148 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_211
timestamp 1586364061
transform 1 0 20516 0 -1 8160
box -38 -48 130 592
use scs8hd_nor2_4  _146_
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21896 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_224
timestamp 1586364061
transform 1 0 21712 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_228
timestamp 1586364061
transform 1 0 22080 0 -1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 22724 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23920 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22540 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_232
timestamp 1586364061
transform 1 0 22448 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_246
timestamp 1586364061
transform 1 0 23736 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24472 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 25484 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24288 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_250
timestamp 1586364061
transform 1 0 24104 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_263
timestamp 1586364061
transform 1 0 25300 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_267
timestamp 1586364061
transform 1 0 25668 0 -1 8160
box -38 -48 590 592
use scs8hd_nor2_4  _165_
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 26220 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_285
timestamp 1586364061
transform 1 0 27324 0 -1 8160
box -38 -48 314 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 28336 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 27600 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 28152 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_290
timestamp 1586364061
transform 1 0 27784 0 -1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 29900 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 29532 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_305
timestamp 1586364061
transform 1 0 29164 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_311
timestamp 1586364061
transform 1 0 29716 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_2_.latch
timestamp 1586364061
transform 1 0 32108 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31648 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_324
timestamp 1586364061
transform 1 0 30912 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_334
timestamp 1586364061
transform 1 0 31832 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_348
timestamp 1586364061
transform 1 0 33120 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_10_356
timestamp 1586364061
transform 1 0 33856 0 -1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34316 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34132 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35328 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_370
timestamp 1586364061
transform 1 0 35144 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_374
timestamp 1586364061
transform 1 0 35512 0 -1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35880 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_387
timestamp 1586364061
transform 1 0 36708 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 38824 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_395
timestamp 1586364061
transform 1 0 37444 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_398
timestamp 1586364061
transform 1 0 37720 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_406
timestamp 1586364061
transform 1 0 38456 0 -1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_5_.latch
timestamp 1586364061
transform 1 0 2208 0 1 8160
box -38 -48 1050 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 2024 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 1656 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_8
timestamp 1586364061
transform 1 0 1840 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3956 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 3772 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_23
timestamp 1586364061
transform 1 0 3220 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5520 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_40
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_46
timestamp 1586364061
transform 1 0 5336 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7176 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6992 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_55
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_69
timestamp 1586364061
transform 1 0 7452 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_73
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_88
timestamp 1586364061
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10948 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_92
timestamp 1586364061
transform 1 0 9568 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_105
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_109
timestamp 1586364061
transform 1 0 11132 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_134
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_138
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 14352 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_155
timestamp 1586364061
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_159
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_163
timestamp 1586364061
transform 1 0 16100 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_175
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18308 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18768 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_190
timestamp 1586364061
transform 1 0 18584 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_194
timestamp 1586364061
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19320 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 20516 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_209
timestamp 1586364061
transform 1 0 20332 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_213
timestamp 1586364061
transform 1 0 20700 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _148_
timestamp 1586364061
transform 1 0 21068 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 20884 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22080 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_226
timestamp 1586364061
transform 1 0 21896 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_230
timestamp 1586364061
transform 1 0 22264 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23736 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 23092 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22724 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_234
timestamp 1586364061
transform 1 0 22632 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_237
timestamp 1586364061
transform 1 0 22908 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_241
timestamp 1586364061
transform 1 0 23276 0 1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_249
timestamp 1586364061
transform 1 0 24012 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24196 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 24564 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_253
timestamp 1586364061
transform 1 0 24380 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 26496 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 26312 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 25944 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_268
timestamp 1586364061
transform 1 0 25760 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_272
timestamp 1586364061
transform 1 0 26128 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28244 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27692 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28612 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_287
timestamp 1586364061
transform 1 0 27508 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_291
timestamp 1586364061
transform 1 0 27876 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_297
timestamp 1586364061
transform 1 0 28428 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_301
timestamp 1586364061
transform 1 0 28796 0 1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 29532 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_11_306
timestamp 1586364061
transform 1 0 29256 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_320
timestamp 1586364061
transform 1 0 30544 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 31648 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 31464 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30728 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31096 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_324
timestamp 1586364061
transform 1 0 30912 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_328
timestamp 1586364061
transform 1 0 31280 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33764 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 32844 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33212 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33580 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_343
timestamp 1586364061
transform 1 0 32660 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_347
timestamp 1586364061
transform 1 0 33028 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_351
timestamp 1586364061
transform 1 0 33396 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34224 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_358
timestamp 1586364061
transform 1 0 34040 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_362
timestamp 1586364061
transform 1 0 34408 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36432 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36892 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 35880 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_376
timestamp 1586364061
transform 1 0 35696 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_380
timestamp 1586364061
transform 1 0 36064 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_387
timestamp 1586364061
transform 1 0 36708 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_391
timestamp 1586364061
transform 1 0 37076 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37444 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 38824 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37904 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_398
timestamp 1586364061
transform 1 0 37720 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_402
timestamp 1586364061
transform 1 0 38088 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_406
timestamp 1586364061
transform 1 0 38456 0 1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_3_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 1050 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_9
timestamp 1586364061
transform 1 0 1932 0 -1 9248
box -38 -48 130 592
use scs8hd_buf_2  _191_
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4600 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4968 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_36
timestamp 1586364061
transform 1 0 4416 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_40
timestamp 1586364061
transform 1 0 4784 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_2_.latch
timestamp 1586364061
transform 1 0 6900 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6716 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_55
timestamp 1586364061
transform 1 0 6164 0 -1 9248
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8188 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_74
timestamp 1586364061
transform 1 0 7912 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_12_79
timestamp 1586364061
transform 1 0 8372 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_6  FILLER_12_85
timestamp 1586364061
transform 1 0 8924 0 -1 9248
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_91
timestamp 1586364061
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  FILLER_12_114
timestamp 1586364061
transform 1 0 11592 0 -1 9248
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12880 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_126
timestamp 1586364061
transform 1 0 12696 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_130
timestamp 1586364061
transform 1 0 13064 0 -1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_149
timestamp 1586364061
transform 1 0 14812 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _157_
timestamp 1586364061
transform 1 0 16836 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_163
timestamp 1586364061
transform 1 0 16100 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_12_168
timestamp 1586364061
transform 1 0 16560 0 -1 9248
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 19044 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18860 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18400 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_180
timestamp 1586364061
transform 1 0 17664 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_186
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_190
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_206
timestamp 1586364061
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_210
timestamp 1586364061
transform 1 0 20424 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_224
timestamp 1586364061
transform 1 0 21712 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_228
timestamp 1586364061
transform 1 0 22080 0 -1 9248
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_12_236
timestamp 1586364061
transform 1 0 22816 0 -1 9248
box -38 -48 314 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 24840 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 24656 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24288 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_250
timestamp 1586364061
transform 1 0 24104 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_254
timestamp 1586364061
transform 1 0 24472 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_267
timestamp 1586364061
transform 1 0 25668 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25852 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_271
timestamp 1586364061
transform 1 0 26036 0 -1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28244 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_12_287
timestamp 1586364061
transform 1 0 27508 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30452 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29532 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_304
timestamp 1586364061
transform 1 0 29072 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_308
timestamp 1586364061
transform 1 0 29440 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_311
timestamp 1586364061
transform 1 0 29716 0 -1 9248
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 32108 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31832 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_328
timestamp 1586364061
transform 1 0 31280 0 -1 9248
box -38 -48 590 592
use scs8hd_decap_12  FILLER_12_348
timestamp 1586364061
transform 1 0 33120 0 -1 9248
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34316 0 -1 9248
box -38 -48 866 592
use scs8hd_fill_1  FILLER_12_360
timestamp 1586364061
transform 1 0 34224 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_370
timestamp 1586364061
transform 1 0 35144 0 -1 9248
box -38 -48 774 592
use scs8hd_buf_2  _196_
timestamp 1586364061
transform 1 0 35880 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_382
timestamp 1586364061
transform 1 0 36248 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 38824 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_394
timestamp 1586364061
transform 1 0 37352 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_398
timestamp 1586364061
transform 1 0 37720 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_406
timestamp 1586364061
transform 1 0 38456 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_7
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 1564 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_buf_2  _190_
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use scs8hd_decap_3  FILLER_13_11
timestamp 1586364061
transform 1 0 2116 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 1932 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_4_.latch
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 1050 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 2116 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_6  FILLER_14_24
timestamp 1586364061
transform 1 0 3312 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_20
timestamp 1586364061
transform 1 0 2944 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3128 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_30
timestamp 1586364061
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_31
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4140 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4324 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 5612 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 5612 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_44
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_48
timestamp 1586364061
transform 1 0 5520 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_41
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_46
timestamp 1586364061
transform 1 0 5336 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_6  FILLER_14_58
timestamp 1586364061
transform 1 0 6440 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_55
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_70
timestamp 1586364061
transform 1 0 7544 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_66
timestamp 1586364061
transform 1 0 7176 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 -1 10336
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6992 0 1 9248
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8740 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8648 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_75
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_79
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_96
timestamp 1586364061
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_92
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_102
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_107
timestamp 1586364061
transform 1 0 10948 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_103
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10304 0 1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_8  FILLER_14_111
timestamp 1586364061
transform 1 0 11316 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_108
timestamp 1586364061
transform 1 0 11040 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 11132 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11132 0 -1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 12052 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 13432 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13064 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 406 592
use scs8hd_decap_4  FILLER_13_138
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_142
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_128
timestamp 1586364061
transform 1 0 12880 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_132
timestamp 1586364061
transform 1 0 13248 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_149
timestamp 1586364061
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_160
timestamp 1586364061
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_156
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 14444 0 1 9248
box -38 -48 1050 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 16192 0 1 9248
box -38 -48 866 592
use scs8hd_buf_2  _194_
timestamp 1586364061
transform 1 0 16836 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_173
timestamp 1586364061
transform 1 0 17020 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_177
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_163
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_6  FILLER_14_175
timestamp 1586364061
transform 1 0 17204 0 -1 10336
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17848 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_195
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_181
timestamp 1586364061
transform 1 0 17756 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_193
timestamp 1586364061
transform 1 0 18860 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_205
timestamp 1586364061
transform 1 0 19964 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_201
timestamp 1586364061
transform 1 0 19596 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_199
timestamp 1586364061
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 19596 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  _142_
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_213
timestamp 1586364061
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_209
timestamp 1586364061
transform 1 0 20332 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_214
timestamp 1586364061
transform 1 0 20792 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20148 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 19780 0 1 9248
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21528 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20976 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_218
timestamp 1586364061
transform 1 0 21160 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_231
timestamp 1586364061
transform 1 0 22356 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_224
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_13_239
timestamp 1586364061
transform 1 0 23092 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_235
timestamp 1586364061
transform 1 0 22724 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 22908 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 22540 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_248
timestamp 1586364061
transform 1 0 23920 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_245
timestamp 1586364061
transform 1 0 23644 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_241
timestamp 1586364061
transform 1 0 23276 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23736 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _113_
timestamp 1586364061
transform 1 0 22448 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_258
timestamp 1586364061
transform 1 0 24840 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_254
timestamp 1586364061
transform 1 0 24472 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24104 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_265
timestamp 1586364061
transform 1 0 25484 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_261
timestamp 1586364061
transform 1 0 25116 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25024 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 25576 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24288 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25208 0 1 9248
box -38 -48 866 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_274
timestamp 1586364061
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_268
timestamp 1586364061
transform 1 0 25760 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_275
timestamp 1586364061
transform 1 0 26404 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_271
timestamp 1586364061
transform 1 0 26036 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26220 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_284
timestamp 1586364061
transform 1 0 27232 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_280
timestamp 1586364061
transform 1 0 26864 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_279
timestamp 1586364061
transform 1 0 26772 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27048 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 26588 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 26588 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26864 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_293
timestamp 1586364061
transform 1 0 28060 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_289
timestamp 1586364061
transform 1 0 27692 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27876 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_301
timestamp 1586364061
transform 1 0 28796 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_297
timestamp 1586364061
transform 1 0 28428 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_301
timestamp 1586364061
transform 1 0 28796 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_297
timestamp 1586364061
transform 1 0 28428 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28244 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 28612 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 28612 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 28980 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27600 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_312
timestamp 1586364061
transform 1 0 29808 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_306
timestamp 1586364061
transform 1 0 29256 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29532 0 1 9248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_14_314
timestamp 1586364061
transform 1 0 29992 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_316
timestamp 1586364061
transform 1 0 30176 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30544 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30360 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 29992 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30544 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _166_
timestamp 1586364061
transform 1 0 29164 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_6  FILLER_14_325
timestamp 1586364061
transform 1 0 31004 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_329
timestamp 1586364061
transform 1 0 31372 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30728 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_333
timestamp 1586364061
transform 1 0 31740 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_13_333
timestamp 1586364061
transform 1 0 31740 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31556 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32108 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31556 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32108 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_346
timestamp 1586364061
transform 1 0 32936 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_350
timestamp 1586364061
transform 1 0 33304 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_356
timestamp 1586364061
transform 1 0 33856 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_352
timestamp 1586364061
transform 1 0 33488 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_348
timestamp 1586364061
transform 1 0 33120 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33120 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33304 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33672 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32292 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33672 0 -1 10336
box -38 -48 866 592
use scs8hd_buf_2  _192_
timestamp 1586364061
transform 1 0 35420 0 1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35236 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35236 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34040 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_360
timestamp 1586364061
transform 1 0 34224 0 1 9248
box -38 -48 590 592
use scs8hd_decap_4  FILLER_13_367
timestamp 1586364061
transform 1 0 34868 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_363
timestamp 1586364061
transform 1 0 34500 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_374
timestamp 1586364061
transform 1 0 35512 0 -1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 35972 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_377
timestamp 1586364061
transform 1 0 35788 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_381
timestamp 1586364061
transform 1 0 36156 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_386
timestamp 1586364061
transform 1 0 36616 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 38824 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 38824 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_393
timestamp 1586364061
transform 1 0 37260 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_13_405
timestamp 1586364061
transform 1 0 38364 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_394
timestamp 1586364061
transform 1 0 37352 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_398
timestamp 1586364061
transform 1 0 37720 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_406
timestamp 1586364061
transform 1 0 38456 0 -1 10336
box -38 -48 130 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_12
timestamp 1586364061
transform 1 0 2208 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_16
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2944 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_29
timestamp 1586364061
transform 1 0 3772 0 1 10336
box -38 -48 774 592
use scs8hd_nor2_4  _138_
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_37
timestamp 1586364061
transform 1 0 4508 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_40
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_73
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_77
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_90
timestamp 1586364061
transform 1 0 9384 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_95
timestamp 1586364061
transform 1 0 9844 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_101
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_105
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _103_
timestamp 1586364061
transform 1 0 12512 0 1 10336
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11132 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11868 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_112
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_116
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_119
timestamp 1586364061
transform 1 0 12052 0 1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 130 592
use scs8hd_nor2_4  _158_
timestamp 1586364061
transform 1 0 14076 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_133
timestamp 1586364061
transform 1 0 13340 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_137
timestamp 1586364061
transform 1 0 13708 0 1 10336
box -38 -48 222 592
use scs8hd_or3_4  _073_
timestamp 1586364061
transform 1 0 15640 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 15088 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_150
timestamp 1586364061
transform 1 0 14904 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_154
timestamp 1586364061
transform 1 0 15272 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__C
timestamp 1586364061
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17020 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_167
timestamp 1586364061
transform 1 0 16468 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 406 592
use scs8hd_nor2_4  _110_
timestamp 1586364061
transform 1 0 18492 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 18308 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17664 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_15_182
timestamp 1586364061
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20056 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 19504 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 19872 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_198
timestamp 1586364061
transform 1 0 19320 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_202
timestamp 1586364061
transform 1 0 19688 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21068 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_215
timestamp 1586364061
transform 1 0 20884 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_219
timestamp 1586364061
transform 1 0 21252 0 1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_15_231
timestamp 1586364061
transform 1 0 22356 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23736 0 1 10336
box -38 -48 866 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_236
timestamp 1586364061
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_240
timestamp 1586364061
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 130 592
use scs8hd_nor2_4  _167_
timestamp 1586364061
transform 1 0 25576 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_255
timestamp 1586364061
transform 1 0 24564 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_259
timestamp 1586364061
transform 1 0 24932 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_263
timestamp 1586364061
transform 1 0 25300 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26588 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_275
timestamp 1586364061
transform 1 0 26404 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_279
timestamp 1586364061
transform 1 0 26772 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_285
timestamp 1586364061
transform 1 0 27324 0 1 10336
box -38 -48 130 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 27600 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 27416 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 28980 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 28612 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_297
timestamp 1586364061
transform 1 0 28428 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_301
timestamp 1586364061
transform 1 0 28796 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 29256 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_15_315
timestamp 1586364061
transform 1 0 30084 0 1 10336
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 31556 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31004 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31372 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_323
timestamp 1586364061
transform 1 0 30820 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_327
timestamp 1586364061
transform 1 0 31188 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33120 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32568 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33580 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_340
timestamp 1586364061
transform 1 0 32384 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_344
timestamp 1586364061
transform 1 0 32752 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_351
timestamp 1586364061
transform 1 0 33396 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_355
timestamp 1586364061
transform 1 0 33764 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33948 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_359
timestamp 1586364061
transform 1 0 34132 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_365
timestamp 1586364061
transform 1 0 34684 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_367
timestamp 1586364061
transform 1 0 34868 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_379
timestamp 1586364061
transform 1 0 35972 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_391
timestamp 1586364061
transform 1 0 37076 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 38824 0 1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_15_403
timestamp 1586364061
transform 1 0 38180 0 1 10336
box -38 -48 406 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 2116 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_7
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3128 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_20
timestamp 1586364061
transform 1 0 2944 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_24
timestamp 1586364061
transform 1 0 3312 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_30
timestamp 1586364061
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 590 592
use scs8hd_nor2_4  _140_
timestamp 1586364061
transform 1 0 5612 0 -1 11424
box -38 -48 866 592
use scs8hd_inv_1  mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4600 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_41
timestamp 1586364061
transform 1 0 4876 0 -1 11424
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_58
timestamp 1586364061
transform 1 0 6440 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_64
timestamp 1586364061
transform 1 0 6992 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7820 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_72
timestamp 1586364061
transform 1 0 7728 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_82
timestamp 1586364061
transform 1 0 8648 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_86
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_96
timestamp 1586364061
transform 1 0 9936 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_8  FILLER_16_107
timestamp 1586364061
transform 1 0 10948 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11868 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 12512 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_115
timestamp 1586364061
transform 1 0 11684 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_120
timestamp 1586364061
transform 1 0 12144 0 -1 11424
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 12880 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_126
timestamp 1586364061
transform 1 0 12696 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_130
timestamp 1586364061
transform 1 0 13064 0 -1 11424
box -38 -48 1142 592
use scs8hd_buf_1  _156_
timestamp 1586364061
transform 1 0 15548 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_160
timestamp 1586364061
transform 1 0 15824 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16560 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__073__B
timestamp 1586364061
transform 1 0 16008 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_164
timestamp 1586364061
transform 1 0 16192 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_16_171
timestamp 1586364061
transform 1 0 16836 0 -1 11424
box -38 -48 774 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 19136 0 -1 11424
box -38 -48 866 592
use scs8hd_inv_1  mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17664 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 18492 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 18124 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_179
timestamp 1586364061
transform 1 0 17572 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_183
timestamp 1586364061
transform 1 0 17940 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_187
timestamp 1586364061
transform 1 0 18308 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_191
timestamp 1586364061
transform 1 0 18676 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_195
timestamp 1586364061
transform 1 0 19044 0 -1 11424
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_205
timestamp 1586364061
transform 1 0 19964 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_209
timestamp 1586364061
transform 1 0 20332 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_213
timestamp 1586364061
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use scs8hd_conb_1  _189_
timestamp 1586364061
transform 1 0 22080 0 -1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_218
timestamp 1586364061
transform 1 0 21160 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_226
timestamp 1586364061
transform 1 0 21896 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_231
timestamp 1586364061
transform 1 0 22356 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23276 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23736 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_244
timestamp 1586364061
transform 1 0 23552 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_248
timestamp 1586364061
transform 1 0 23920 0 -1 11424
box -38 -48 406 592
use scs8hd_buf_2  _202_
timestamp 1586364061
transform 1 0 24288 0 -1 11424
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_256
timestamp 1586364061
transform 1 0 24656 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_267
timestamp 1586364061
transform 1 0 25668 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 25852 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_271
timestamp 1586364061
transform 1 0 26036 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_16_279
timestamp 1586364061
transform 1 0 26772 0 -1 11424
box -38 -48 774 592
use scs8hd_nor2_4  _168_
timestamp 1586364061
transform 1 0 28152 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 27600 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_287
timestamp 1586364061
transform 1 0 27508 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_290
timestamp 1586364061
transform 1 0 27784 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_3  FILLER_16_303
timestamp 1586364061
transform 1 0 28980 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 29256 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_308
timestamp 1586364061
transform 1 0 29440 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_16_320
timestamp 1586364061
transform 1 0 30544 0 -1 11424
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32108 0 -1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31004 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_324
timestamp 1586364061
transform 1 0 30912 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_328
timestamp 1586364061
transform 1 0 31280 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33304 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_340
timestamp 1586364061
transform 1 0 32384 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_348
timestamp 1586364061
transform 1 0 33120 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_353
timestamp 1586364061
transform 1 0 33580 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_365
timestamp 1586364061
transform 1 0 34684 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_377
timestamp 1586364061
transform 1 0 35788 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_389
timestamp 1586364061
transform 1 0 36892 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 38824 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_398
timestamp 1586364061
transform 1 0 37720 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_406
timestamp 1586364061
transform 1 0 38456 0 -1 11424
box -38 -48 130 592
use scs8hd_buf_2  _199_
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use scs8hd_buf_2  _203_
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_11
timestamp 1586364061
transform 1 0 2116 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 3036 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_19
timestamp 1586364061
transform 1 0 2852 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_23
timestamp 1586364061
transform 1 0 3220 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_35
timestamp 1586364061
transform 1 0 4324 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_47
timestamp 1586364061
transform 1 0 5428 0 1 11424
box -38 -48 774 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_71
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_75
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_82
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9384 0 1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10856 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_93
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_97
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_104
timestamp 1586364061
transform 1 0 10672 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_108
timestamp 1586364061
transform 1 0 11040 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_112
timestamp 1586364061
transform 1 0 11408 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_120
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13800 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_141
timestamp 1586364061
transform 1 0 14076 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _179_
timestamp 1586364061
transform 1 0 14812 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_145
timestamp 1586364061
transform 1 0 14444 0 1 11424
box -38 -48 406 592
use scs8hd_decap_6  FILLER_17_152
timestamp 1586364061
transform 1 0 15088 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_158
timestamp 1586364061
transform 1 0 15640 0 1 11424
box -38 -48 130 592
use scs8hd_conb_1  _184_
timestamp 1586364061
transform 1 0 16560 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17020 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_161
timestamp 1586364061
transform 1 0 15916 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_167
timestamp 1586364061
transform 1 0 16468 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_171
timestamp 1586364061
transform 1 0 16836 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_175
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 590 592
use scs8hd_nor2_4  _109_
timestamp 1586364061
transform 1 0 18124 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_194
timestamp 1586364061
transform 1 0 18952 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19688 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20148 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 20516 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_198
timestamp 1586364061
transform 1 0 19320 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_205
timestamp 1586364061
transform 1 0 19964 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_209
timestamp 1586364061
transform 1 0 20332 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_213
timestamp 1586364061
transform 1 0 20700 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_225
timestamp 1586364061
transform 1 0 21804 0 1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_236
timestamp 1586364061
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_240
timestamp 1586364061
transform 1 0 23184 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_249
timestamp 1586364061
transform 1 0 24012 0 1 11424
box -38 -48 406 592
use scs8hd_buf_1  _068_
timestamp 1586364061
transform 1 0 24380 0 1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 24840 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 25208 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_256
timestamp 1586364061
transform 1 0 24656 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_260
timestamp 1586364061
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_267
timestamp 1586364061
transform 1 0 25668 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _181_
timestamp 1586364061
transform 1 0 27324 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_271
timestamp 1586364061
transform 1 0 26036 0 1 11424
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_17_283
timestamp 1586364061
transform 1 0 27140 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 27784 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_288
timestamp 1586364061
transform 1 0 27600 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_292
timestamp 1586364061
transform 1 0 27968 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_304
timestamp 1586364061
transform 1 0 29072 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_306
timestamp 1586364061
transform 1 0 29256 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_318
timestamp 1586364061
transform 1 0 30360 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_330
timestamp 1586364061
transform 1 0 31464 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_342
timestamp 1586364061
transform 1 0 32568 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_354
timestamp 1586364061
transform 1 0 33672 0 1 11424
box -38 -48 1142 592
use scs8hd_buf_2  _201_
timestamp 1586364061
transform 1 0 35420 0 1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_17_367
timestamp 1586364061
transform 1 0 34868 0 1 11424
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 35972 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_377
timestamp 1586364061
transform 1 0 35788 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_381
timestamp 1586364061
transform 1 0 36156 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 38824 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_393
timestamp 1586364061
transform 1 0 37260 0 1 11424
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_17_405
timestamp 1586364061
transform 1 0 38364 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _187_
timestamp 1586364061
transform 1 0 2668 0 -1 12512
box -38 -48 314 592
use scs8hd_buf_2  _206_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_7
timestamp 1586364061
transform 1 0 1748 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_20
timestamp 1586364061
transform 1 0 2944 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_18_28
timestamp 1586364061
transform 1 0 3680 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7636 0 -1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6624 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_18_63
timestamp 1586364061
transform 1 0 6900 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_18_74
timestamp 1586364061
transform 1 0 7912 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_18_86
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 590 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10672 0 -1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_96
timestamp 1586364061
transform 1 0 9936 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_18_107
timestamp 1586364061
transform 1 0 10948 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_119
timestamp 1586364061
transform 1 0 12052 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_131
timestamp 1586364061
transform 1 0 13156 0 -1 12512
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15732 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_143
timestamp 1586364061
transform 1 0 14260 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_151
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_158
timestamp 1586364061
transform 1 0 15640 0 -1 12512
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16744 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_162
timestamp 1586364061
transform 1 0 16008 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_8  FILLER_18_173
timestamp 1586364061
transform 1 0 17020 0 -1 12512
box -38 -48 774 592
use scs8hd_conb_1  _185_
timestamp 1586364061
transform 1 0 17756 0 -1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18768 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_184
timestamp 1586364061
transform 1 0 18032 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_8  FILLER_18_195
timestamp 1586364061
transform 1 0 19044 0 -1 12512
box -38 -48 774 592
use scs8hd_buf_1  _108_
timestamp 1586364061
transform 1 0 19780 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23460 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_18_246
timestamp 1586364061
transform 1 0 23736 0 -1 12512
box -38 -48 774 592
use scs8hd_buf_1  _104_
timestamp 1586364061
transform 1 0 24472 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_257
timestamp 1586364061
transform 1 0 24748 0 -1 12512
box -38 -48 1142 592
use scs8hd_buf_1  _102_
timestamp 1586364061
transform 1 0 27324 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_18_269
timestamp 1586364061
transform 1 0 25852 0 -1 12512
box -38 -48 590 592
use scs8hd_decap_8  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_284
timestamp 1586364061
transform 1 0 27232 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_288
timestamp 1586364061
transform 1 0 27600 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_300
timestamp 1586364061
transform 1 0 28704 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_312
timestamp 1586364061
transform 1 0 29808 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_324
timestamp 1586364061
transform 1 0 30912 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_337
timestamp 1586364061
transform 1 0 32108 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_349
timestamp 1586364061
transform 1 0 33212 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_361
timestamp 1586364061
transform 1 0 34316 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_373
timestamp 1586364061
transform 1 0 35420 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_385
timestamp 1586364061
transform 1 0 36524 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 38824 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_398
timestamp 1586364061
transform 1 0 37720 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_406
timestamp 1586364061
transform 1 0 38456 0 -1 12512
box -38 -48 130 592
use scs8hd_buf_2  _207_
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 1932 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_11
timestamp 1586364061
transform 1 0 2116 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_23
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_35
timestamp 1586364061
transform 1 0 4324 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_47
timestamp 1586364061
transform 1 0 5428 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_1  _126_
timestamp 1586364061
transform 1 0 7268 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_66
timestamp 1586364061
transform 1 0 7176 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_70
timestamp 1586364061
transform 1 0 7544 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_63
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8280 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 7728 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_81
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_85
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_75
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_87
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_97
timestamp 1586364061
transform 1 0 10028 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_94
timestamp 1586364061
transform 1 0 9752 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_109
timestamp 1586364061
transform 1 0 11132 0 1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_19_121
timestamp 1586364061
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_118
timestamp 1586364061
transform 1 0 11960 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_137
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 15364 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_156
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_171
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_168
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_2  _193_
timestamp 1586364061
transform 1 0 18308 0 1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_191
timestamp 1586364061
transform 1 0 18676 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_195
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_180
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_187
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_207
timestamp 1586364061
transform 1 0 20148 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_199
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_211
timestamp 1586364061
transform 1 0 20516 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_219
timestamp 1586364061
transform 1 0 21252 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_231
timestamp 1586364061
transform 1 0 22356 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_218
timestamp 1586364061
transform 1 0 21160 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_230
timestamp 1586364061
transform 1 0 22264 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 23920 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_243
timestamp 1586364061
transform 1 0 23460 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_242
timestamp 1586364061
transform 1 0 23368 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_249
timestamp 1586364061
transform 1 0 24012 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_261
timestamp 1586364061
transform 1 0 25116 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 26772 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_281
timestamp 1586364061
transform 1 0 26956 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_273
timestamp 1586364061
transform 1 0 26220 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_280
timestamp 1586364061
transform 1 0 26864 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_2  _205_
timestamp 1586364061
transform 1 0 28060 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 28612 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_297
timestamp 1586364061
transform 1 0 28428 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_301
timestamp 1586364061
transform 1 0 28796 0 1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_292
timestamp 1586364061
transform 1 0 27968 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 29624 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_306
timestamp 1586364061
transform 1 0 29256 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_318
timestamp 1586364061
transform 1 0 30360 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_304
timestamp 1586364061
transform 1 0 29072 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_311
timestamp 1586364061
transform 1 0 29716 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_2  _204_
timestamp 1586364061
transform 1 0 31740 0 1 12512
box -38 -48 406 592
use scs8hd_decap_3  FILLER_19_330
timestamp 1586364061
transform 1 0 31464 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_337
timestamp 1586364061
transform 1 0 32108 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_323
timestamp 1586364061
transform 1 0 30820 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_335
timestamp 1586364061
transform 1 0 31924 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 32476 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 32292 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_341
timestamp 1586364061
transform 1 0 32476 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_353
timestamp 1586364061
transform 1 0 33580 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_342
timestamp 1586364061
transform 1 0 32568 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_354
timestamp 1586364061
transform 1 0 33672 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_2  _200_
timestamp 1586364061
transform 1 0 35420 0 1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 35328 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_365
timestamp 1586364061
transform 1 0 34684 0 1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_19_367
timestamp 1586364061
transform 1 0 34868 0 1 12512
box -38 -48 590 592
use scs8hd_decap_6  FILLER_20_366
timestamp 1586364061
transform 1 0 34776 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_373
timestamp 1586364061
transform 1 0 35420 0 -1 13600
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 35972 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_377
timestamp 1586364061
transform 1 0 35788 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_381
timestamp 1586364061
transform 1 0 36156 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_385
timestamp 1586364061
transform 1 0 36524 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 38824 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 38824 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 38180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_393
timestamp 1586364061
transform 1 0 37260 0 1 12512
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_19_405
timestamp 1586364061
transform 1 0 38364 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_397
timestamp 1586364061
transform 1 0 37628 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_3  FILLER_20_404
timestamp 1586364061
transform 1 0 38272 0 -1 13600
box -38 -48 314 592
<< labels >>
rlabel metal3 s 0 416 480 536 6 address[0]
port 0 nsew default input
rlabel metal3 s 0 1232 480 1352 6 address[1]
port 1 nsew default input
rlabel metal2 s 1766 15520 1822 16000 6 address[2]
port 2 nsew default input
rlabel metal3 s 0 2184 480 2304 6 address[3]
port 3 nsew default input
rlabel metal2 s 7102 0 7158 480 6 address[4]
port 4 nsew default input
rlabel metal3 s 39520 552 40000 672 6 address[5]
port 5 nsew default input
rlabel metal3 s 39520 1640 40000 1760 6 address[6]
port 6 nsew default input
rlabel metal3 s 39520 2728 40000 2848 6 bottom_grid_pin_0_
port 7 nsew default tristate
rlabel metal2 s 9034 15520 9090 16000 6 bottom_grid_pin_10_
port 8 nsew default tristate
rlabel metal3 s 0 3136 480 3256 6 bottom_grid_pin_12_
port 9 nsew default tristate
rlabel metal3 s 0 4088 480 4208 6 bottom_grid_pin_14_
port 10 nsew default tristate
rlabel metal2 s 9954 0 10010 480 6 bottom_grid_pin_2_
port 11 nsew default tristate
rlabel metal2 s 12806 0 12862 480 6 bottom_grid_pin_4_
port 12 nsew default tristate
rlabel metal2 s 5354 15520 5410 16000 6 bottom_grid_pin_6_
port 13 nsew default tristate
rlabel metal3 s 39520 3952 40000 4072 6 bottom_grid_pin_8_
port 14 nsew default tristate
rlabel metal3 s 39520 5040 40000 5160 6 chanx_left_in[0]
port 15 nsew default input
rlabel metal2 s 12622 15520 12678 16000 6 chanx_left_in[1]
port 16 nsew default input
rlabel metal3 s 39520 6264 40000 6384 6 chanx_left_in[2]
port 17 nsew default input
rlabel metal2 s 15658 0 15714 480 6 chanx_left_in[3]
port 18 nsew default input
rlabel metal3 s 0 5040 480 5160 6 chanx_left_in[4]
port 19 nsew default input
rlabel metal2 s 18510 0 18566 480 6 chanx_left_in[5]
port 20 nsew default input
rlabel metal2 s 21362 0 21418 480 6 chanx_left_in[6]
port 21 nsew default input
rlabel metal2 s 24214 0 24270 480 6 chanx_left_in[7]
port 22 nsew default input
rlabel metal3 s 0 5992 480 6112 6 chanx_left_in[8]
port 23 nsew default input
rlabel metal3 s 0 6944 480 7064 6 chanx_left_out[0]
port 24 nsew default tristate
rlabel metal3 s 39520 7352 40000 7472 6 chanx_left_out[1]
port 25 nsew default tristate
rlabel metal3 s 39520 8576 40000 8696 6 chanx_left_out[2]
port 26 nsew default tristate
rlabel metal2 s 27066 0 27122 480 6 chanx_left_out[3]
port 27 nsew default tristate
rlabel metal2 s 16302 15520 16358 16000 6 chanx_left_out[4]
port 28 nsew default tristate
rlabel metal2 s 19890 15520 19946 16000 6 chanx_left_out[5]
port 29 nsew default tristate
rlabel metal3 s 39520 9664 40000 9784 6 chanx_left_out[6]
port 30 nsew default tristate
rlabel metal3 s 0 7896 480 8016 6 chanx_left_out[7]
port 31 nsew default tristate
rlabel metal3 s 0 8848 480 8968 6 chanx_left_out[8]
port 32 nsew default tristate
rlabel metal2 s 29918 0 29974 480 6 chanx_right_in[0]
port 33 nsew default input
rlabel metal2 s 32770 0 32826 480 6 chanx_right_in[1]
port 34 nsew default input
rlabel metal2 s 35622 0 35678 480 6 chanx_right_in[2]
port 35 nsew default input
rlabel metal2 s 23570 15520 23626 16000 6 chanx_right_in[3]
port 36 nsew default input
rlabel metal3 s 0 9800 480 9920 6 chanx_right_in[4]
port 37 nsew default input
rlabel metal2 s 27158 15520 27214 16000 6 chanx_right_in[5]
port 38 nsew default input
rlabel metal2 s 30838 15520 30894 16000 6 chanx_right_in[6]
port 39 nsew default input
rlabel metal3 s 39520 10752 40000 10872 6 chanx_right_in[7]
port 40 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_right_in[8]
port 41 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_right_out[0]
port 42 nsew default tristate
rlabel metal3 s 0 12656 480 12776 6 chanx_right_out[1]
port 43 nsew default tristate
rlabel metal3 s 0 13608 480 13728 6 chanx_right_out[2]
port 44 nsew default tristate
rlabel metal2 s 34426 15520 34482 16000 6 chanx_right_out[3]
port 45 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_right_out[4]
port 46 nsew default tristate
rlabel metal3 s 39520 11976 40000 12096 6 chanx_right_out[5]
port 47 nsew default tristate
rlabel metal3 s 39520 13064 40000 13184 6 chanx_right_out[6]
port 48 nsew default tristate
rlabel metal3 s 39520 14288 40000 14408 6 chanx_right_out[7]
port 49 nsew default tristate
rlabel metal3 s 0 15512 480 15632 6 chanx_right_out[8]
port 50 nsew default tristate
rlabel metal2 s 4250 0 4306 480 6 data_in
port 51 nsew default input
rlabel metal2 s 1398 0 1454 480 6 enable
port 52 nsew default input
rlabel metal2 s 38106 15520 38162 16000 6 top_grid_pin_14_
port 53 nsew default tristate
rlabel metal3 s 39520 15376 40000 15496 6 top_grid_pin_2_
port 54 nsew default tristate
rlabel metal2 s 38474 0 38530 480 6 top_grid_pin_6_
port 55 nsew default tristate
rlabel metal4 s 7611 2128 7931 13648 6 vpwr
port 56 nsew default input
rlabel metal4 s 14277 2128 14597 13648 6 vgnd
port 57 nsew default input
<< end >>
