VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_1__0_
  CLASS BLOCK ;
  FOREIGN sb_1__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 140.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 2.400 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 2.400 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 2.400 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 2.400 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 2.400 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 2.400 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 2.400 ;
    END
  END address[6]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 2.400 2.680 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 2.400 7.440 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 2.400 12.880 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 2.400 17.640 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 2.400 23.080 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 2.400 28.520 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 2.400 33.280 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 2.400 38.720 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 2.400 44.160 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 2.400 95.840 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 2.400 100.600 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 2.400 106.040 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 2.400 111.480 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 2.400 116.240 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 2.400 121.680 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 2.400 127.120 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 2.400 131.880 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.720 2.400 137.320 ;
    END
  END chanx_left_out[8]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 6.840 140.000 7.440 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 12.280 140.000 12.880 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 17.040 140.000 17.640 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 22.480 140.000 23.080 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 27.920 140.000 28.520 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 32.680 140.000 33.280 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 38.120 140.000 38.720 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 43.560 140.000 44.160 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 48.320 140.000 48.920 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 95.240 140.000 95.840 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 100.000 140.000 100.600 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 105.440 140.000 106.040 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 110.880 140.000 111.480 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 115.640 140.000 116.240 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 121.080 140.000 121.680 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 126.520 140.000 127.120 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 131.280 140.000 131.880 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 136.720 140.000 137.320 ;
    END
  END chanx_right_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.310 137.600 3.590 140.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.210 137.600 10.490 140.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.110 137.600 17.390 140.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 137.600 24.290 140.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.910 137.600 31.190 140.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.270 137.600 38.550 140.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.170 137.600 45.450 140.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.070 137.600 52.350 140.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.970 137.600 59.250 140.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 80.130 137.600 80.410 140.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.030 137.600 87.310 140.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.930 137.600 94.210 140.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.830 137.600 101.110 140.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.190 137.600 108.470 140.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 115.090 137.600 115.370 140.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.990 137.600 122.270 140.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 128.890 137.600 129.170 140.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 135.790 137.600 136.070 140.000 ;
    END
  END chany_top_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 2.400 ;
    END
  END enable
  PIN left_bottom_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 2.400 80.200 ;
    END
  END left_bottom_grid_pin_11_
  PIN left_bottom_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 2.400 85.640 ;
    END
  END left_bottom_grid_pin_13_
  PIN left_bottom_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 2.400 90.400 ;
    END
  END left_bottom_grid_pin_15_
  PIN left_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 2.400 54.360 ;
    END
  END left_bottom_grid_pin_1_
  PIN left_bottom_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 2.400 59.120 ;
    END
  END left_bottom_grid_pin_3_
  PIN left_bottom_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 2.400 64.560 ;
    END
  END left_bottom_grid_pin_5_
  PIN left_bottom_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 2.400 70.000 ;
    END
  END left_bottom_grid_pin_7_
  PIN left_bottom_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 2.400 74.760 ;
    END
  END left_bottom_grid_pin_9_
  PIN left_top_grid_pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 2.400 48.920 ;
    END
  END left_top_grid_pin_10_
  PIN right_bottom_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 79.600 140.000 80.200 ;
    END
  END right_bottom_grid_pin_11_
  PIN right_bottom_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 85.040 140.000 85.640 ;
    END
  END right_bottom_grid_pin_13_
  PIN right_bottom_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 89.800 140.000 90.400 ;
    END
  END right_bottom_grid_pin_15_
  PIN right_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 53.760 140.000 54.360 ;
    END
  END right_bottom_grid_pin_1_
  PIN right_bottom_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 58.520 140.000 59.120 ;
    END
  END right_bottom_grid_pin_3_
  PIN right_bottom_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 63.960 140.000 64.560 ;
    END
  END right_bottom_grid_pin_5_
  PIN right_bottom_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 69.400 140.000 70.000 ;
    END
  END right_bottom_grid_pin_7_
  PIN right_bottom_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 74.160 140.000 74.760 ;
    END
  END right_bottom_grid_pin_9_
  PIN right_top_grid_pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 2.080 140.000 2.680 ;
    END
  END right_top_grid_pin_10_
  PIN top_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.870 137.600 66.150 140.000 ;
    END
  END top_left_grid_pin_13_
  PIN top_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 73.230 137.600 73.510 140.000 ;
    END
  END top_right_grid_pin_11_
  PIN vpwr
    USE POWER ;
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END vpwr
  PIN vgnd
    USE GROUND ;
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 0.530 0.380 138.850 137.660 ;
      LAYER met2 ;
        RECT 0.550 137.320 3.030 137.770 ;
        RECT 3.870 137.320 9.930 137.770 ;
        RECT 10.770 137.320 16.830 137.770 ;
        RECT 17.670 137.320 23.730 137.770 ;
        RECT 24.570 137.320 30.630 137.770 ;
        RECT 31.470 137.320 37.990 137.770 ;
        RECT 38.830 137.320 44.890 137.770 ;
        RECT 45.730 137.320 51.790 137.770 ;
        RECT 52.630 137.320 58.690 137.770 ;
        RECT 59.530 137.320 65.590 137.770 ;
        RECT 66.430 137.320 72.950 137.770 ;
        RECT 73.790 137.320 79.850 137.770 ;
        RECT 80.690 137.320 86.750 137.770 ;
        RECT 87.590 137.320 93.650 137.770 ;
        RECT 94.490 137.320 100.550 137.770 ;
        RECT 101.390 137.320 107.910 137.770 ;
        RECT 108.750 137.320 114.810 137.770 ;
        RECT 115.650 137.320 121.710 137.770 ;
        RECT 122.550 137.320 128.610 137.770 ;
        RECT 129.450 137.320 135.510 137.770 ;
        RECT 136.350 137.320 138.830 137.770 ;
        RECT 0.550 2.680 138.830 137.320 ;
        RECT 0.550 0.270 7.170 2.680 ;
        RECT 8.010 0.270 22.350 2.680 ;
        RECT 23.190 0.270 37.990 2.680 ;
        RECT 38.830 0.270 53.630 2.680 ;
        RECT 54.470 0.270 69.270 2.680 ;
        RECT 70.110 0.270 84.450 2.680 ;
        RECT 85.290 0.270 100.090 2.680 ;
        RECT 100.930 0.270 115.730 2.680 ;
        RECT 116.570 0.270 131.370 2.680 ;
        RECT 132.210 0.270 138.830 2.680 ;
      LAYER met3 ;
        RECT 2.800 136.320 137.200 136.720 ;
        RECT 0.270 132.280 138.610 136.320 ;
        RECT 2.800 130.880 137.200 132.280 ;
        RECT 0.270 127.520 138.610 130.880 ;
        RECT 2.800 126.120 137.200 127.520 ;
        RECT 0.270 122.080 138.610 126.120 ;
        RECT 2.800 120.680 137.200 122.080 ;
        RECT 0.270 116.640 138.610 120.680 ;
        RECT 2.800 115.240 137.200 116.640 ;
        RECT 0.270 111.880 138.610 115.240 ;
        RECT 2.800 110.480 137.200 111.880 ;
        RECT 0.270 106.440 138.610 110.480 ;
        RECT 2.800 105.040 137.200 106.440 ;
        RECT 0.270 101.000 138.610 105.040 ;
        RECT 2.800 99.600 137.200 101.000 ;
        RECT 0.270 96.240 138.610 99.600 ;
        RECT 2.800 94.840 137.200 96.240 ;
        RECT 0.270 90.800 138.610 94.840 ;
        RECT 2.800 89.400 137.200 90.800 ;
        RECT 0.270 86.040 138.610 89.400 ;
        RECT 2.800 84.640 137.200 86.040 ;
        RECT 0.270 80.600 138.610 84.640 ;
        RECT 2.800 79.200 137.200 80.600 ;
        RECT 0.270 75.160 138.610 79.200 ;
        RECT 2.800 73.760 137.200 75.160 ;
        RECT 0.270 70.400 138.610 73.760 ;
        RECT 2.800 69.000 137.200 70.400 ;
        RECT 0.270 64.960 138.610 69.000 ;
        RECT 2.800 63.560 137.200 64.960 ;
        RECT 0.270 59.520 138.610 63.560 ;
        RECT 2.800 58.120 137.200 59.520 ;
        RECT 0.270 54.760 138.610 58.120 ;
        RECT 2.800 53.360 137.200 54.760 ;
        RECT 0.270 49.320 138.610 53.360 ;
        RECT 2.800 47.920 137.200 49.320 ;
        RECT 0.270 44.560 138.610 47.920 ;
        RECT 2.800 43.160 137.200 44.560 ;
        RECT 0.270 39.120 138.610 43.160 ;
        RECT 2.800 37.720 137.200 39.120 ;
        RECT 0.270 33.680 138.610 37.720 ;
        RECT 2.800 32.280 137.200 33.680 ;
        RECT 0.270 28.920 138.610 32.280 ;
        RECT 2.800 27.520 137.200 28.920 ;
        RECT 0.270 23.480 138.610 27.520 ;
        RECT 2.800 22.080 137.200 23.480 ;
        RECT 0.270 18.040 138.610 22.080 ;
        RECT 2.800 16.640 137.200 18.040 ;
        RECT 0.270 13.280 138.610 16.640 ;
        RECT 2.800 11.880 137.200 13.280 ;
        RECT 0.270 7.840 138.610 11.880 ;
        RECT 2.800 6.440 137.200 7.840 ;
        RECT 0.270 3.080 138.610 6.440 ;
        RECT 2.800 2.680 137.200 3.080 ;
      LAYER met4 ;
        RECT 0.295 10.640 27.655 128.080 ;
        RECT 30.055 10.640 50.985 128.080 ;
        RECT 53.385 10.640 122.985 128.080 ;
  END
END sb_1__0_
END LIBRARY

