VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cby_3__1_
  CLASS BLOCK ;
  FOREIGN cby_3__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 200.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 2.400 6.760 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 2.400 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 2.400 19.000 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.310 197.600 3.590 200.000 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 2.400 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 8.880 80.000 9.480 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 26.560 80.000 27.160 ;
    END
  END address[6]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.750 197.600 10.030 200.000 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 197.600 16.930 200.000 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 2.400 31.240 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 44.920 80.000 45.520 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 2.400 44.160 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 2.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.090 197.600 23.370 200.000 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 2.400 56.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 2.400 68.640 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 29.990 197.600 30.270 200.000 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 36.430 197.600 36.710 200.000 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 43.330 197.600 43.610 200.000 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 63.280 80.000 63.880 ;
    END
  END chany_bottom_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 2.400 81.560 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 2.400 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 2.400 93.800 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 2.400 106.720 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 2.400 118.960 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.770 197.600 50.050 200.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 2.400 131.200 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.670 197.600 56.950 200.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 2.400 144.120 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 80.960 80.000 81.560 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.760 2.400 156.360 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 2.400 168.600 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 2.400 181.520 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 2.400 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 63.110 197.600 63.390 200.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 70.010 197.600 70.290 200.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.450 197.600 76.730 200.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 2.400 ;
    END
  END chany_top_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 2.400 ;
    END
  END enable
  PIN left_grid_pin_1_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 2.400 193.760 ;
    END
  END left_grid_pin_1_
  PIN left_grid_pin_5_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 2.400 ;
    END
  END left_grid_pin_5_
  PIN left_grid_pin_9_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 2.400 ;
    END
  END left_grid_pin_9_
  PIN right_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 99.320 80.000 99.920 ;
    END
  END right_grid_pin_0_
  PIN right_grid_pin_10_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 153.720 80.000 154.320 ;
    END
  END right_grid_pin_10_
  PIN right_grid_pin_12_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 172.080 80.000 172.680 ;
    END
  END right_grid_pin_12_
  PIN right_grid_pin_14_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 190.440 80.000 191.040 ;
    END
  END right_grid_pin_14_
  PIN right_grid_pin_2_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 2.400 ;
    END
  END right_grid_pin_2_
  PIN right_grid_pin_4_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 117.680 80.000 118.280 ;
    END
  END right_grid_pin_4_
  PIN right_grid_pin_6_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 136.040 80.000 136.640 ;
    END
  END right_grid_pin_6_
  PIN right_grid_pin_8_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 2.400 ;
    END
  END right_grid_pin_8_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 18.055 10.640 19.655 187.920 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 31.385 10.640 32.985 187.920 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 74.060 187.765 ;
      LAYER met1 ;
        RECT 0.530 0.380 78.130 198.180 ;
      LAYER met2 ;
        RECT 0.550 197.320 3.030 198.290 ;
        RECT 3.870 197.320 9.470 198.290 ;
        RECT 10.310 197.320 16.370 198.290 ;
        RECT 17.210 197.320 22.810 198.290 ;
        RECT 23.650 197.320 29.710 198.290 ;
        RECT 30.550 197.320 36.150 198.290 ;
        RECT 36.990 197.320 43.050 198.290 ;
        RECT 43.890 197.320 49.490 198.290 ;
        RECT 50.330 197.320 56.390 198.290 ;
        RECT 57.230 197.320 62.830 198.290 ;
        RECT 63.670 197.320 69.730 198.290 ;
        RECT 70.570 197.320 76.170 198.290 ;
        RECT 77.010 197.320 78.100 198.290 ;
        RECT 0.550 2.680 78.100 197.320 ;
        RECT 0.550 0.270 2.110 2.680 ;
        RECT 2.950 0.270 6.710 2.680 ;
        RECT 7.550 0.270 11.310 2.680 ;
        RECT 12.150 0.270 15.910 2.680 ;
        RECT 16.750 0.270 20.510 2.680 ;
        RECT 21.350 0.270 25.570 2.680 ;
        RECT 26.410 0.270 30.170 2.680 ;
        RECT 31.010 0.270 34.770 2.680 ;
        RECT 35.610 0.270 39.370 2.680 ;
        RECT 40.210 0.270 44.430 2.680 ;
        RECT 45.270 0.270 49.030 2.680 ;
        RECT 49.870 0.270 53.630 2.680 ;
        RECT 54.470 0.270 58.230 2.680 ;
        RECT 59.070 0.270 63.290 2.680 ;
        RECT 64.130 0.270 67.890 2.680 ;
        RECT 68.730 0.270 72.490 2.680 ;
        RECT 73.330 0.270 77.090 2.680 ;
        RECT 77.930 0.270 78.100 2.680 ;
      LAYER met3 ;
        RECT 0.270 190.040 77.200 190.905 ;
        RECT 0.270 181.920 77.600 190.040 ;
        RECT 2.800 180.520 77.600 181.920 ;
        RECT 0.270 173.080 77.600 180.520 ;
        RECT 0.270 171.680 77.200 173.080 ;
        RECT 0.270 169.000 77.600 171.680 ;
        RECT 2.800 167.600 77.600 169.000 ;
        RECT 0.270 156.760 77.600 167.600 ;
        RECT 2.800 155.360 77.600 156.760 ;
        RECT 0.270 154.720 77.600 155.360 ;
        RECT 0.270 153.320 77.200 154.720 ;
        RECT 0.270 144.520 77.600 153.320 ;
        RECT 2.800 143.120 77.600 144.520 ;
        RECT 0.270 137.040 77.600 143.120 ;
        RECT 0.270 135.640 77.200 137.040 ;
        RECT 0.270 131.600 77.600 135.640 ;
        RECT 2.800 130.200 77.600 131.600 ;
        RECT 0.270 119.360 77.600 130.200 ;
        RECT 2.800 118.680 77.600 119.360 ;
        RECT 2.800 117.960 77.200 118.680 ;
        RECT 0.270 117.280 77.200 117.960 ;
        RECT 0.270 107.120 77.600 117.280 ;
        RECT 2.800 105.720 77.600 107.120 ;
        RECT 0.270 100.320 77.600 105.720 ;
        RECT 0.270 98.920 77.200 100.320 ;
        RECT 0.270 94.200 77.600 98.920 ;
        RECT 2.800 92.800 77.600 94.200 ;
        RECT 0.270 81.960 77.600 92.800 ;
        RECT 2.800 80.560 77.200 81.960 ;
        RECT 0.270 69.040 77.600 80.560 ;
        RECT 2.800 67.640 77.600 69.040 ;
        RECT 0.270 64.280 77.600 67.640 ;
        RECT 0.270 62.880 77.200 64.280 ;
        RECT 0.270 56.800 77.600 62.880 ;
        RECT 2.800 55.400 77.600 56.800 ;
        RECT 0.270 45.920 77.600 55.400 ;
        RECT 0.270 44.560 77.200 45.920 ;
        RECT 2.800 44.520 77.200 44.560 ;
        RECT 2.800 43.160 77.600 44.520 ;
        RECT 0.270 31.640 77.600 43.160 ;
        RECT 2.800 30.240 77.600 31.640 ;
        RECT 0.270 27.560 77.600 30.240 ;
        RECT 0.270 26.160 77.200 27.560 ;
        RECT 0.270 19.400 77.600 26.160 ;
        RECT 2.800 18.000 77.600 19.400 ;
        RECT 0.270 9.880 77.600 18.000 ;
        RECT 0.270 8.480 77.200 9.880 ;
        RECT 0.270 7.160 77.600 8.480 ;
        RECT 2.800 6.760 77.600 7.160 ;
      LAYER met4 ;
        RECT 0.295 10.240 17.655 187.920 ;
        RECT 20.055 10.240 30.985 187.920 ;
        RECT 33.385 10.240 72.985 187.920 ;
        RECT 0.295 9.015 72.985 10.240 ;
  END
END cby_3__1_
END LIBRARY

