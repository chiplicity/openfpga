* NGSPICE file created from cbx_1__0_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand2_4 abstract view
.subckt scs8hd_nand2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor3_4 abstract view
.subckt scs8hd_nor3_4 A B C Y vgnd vpwr
.ends

.subckt cbx_1__0_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] bottom_grid_pin_0_ bottom_grid_pin_10_ bottom_grid_pin_12_ bottom_grid_pin_14_
+ bottom_grid_pin_2_ bottom_grid_pin_4_ bottom_grid_pin_6_ bottom_grid_pin_8_ chanx_left_in[0]
+ chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_out[0] chanx_left_out[1]
+ chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6]
+ chanx_left_out[7] chanx_left_out[8] chanx_right_in[0] chanx_right_in[1] chanx_right_in[2]
+ chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7]
+ chanx_right_in[8] chanx_right_out[0] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3]
+ chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8]
+ data_in enable top_grid_pin_14_ top_grid_pin_2_ top_grid_pin_6_ vpwr vgnd
XFILLER_10_306 vpwr vgnd scs8hd_fill_2
XFILLER_10_328 vgnd vpwr scs8hd_decap_8
XFILLER_7_7 vgnd vpwr scs8hd_fill_1
XFILLER_18_406 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_7.LATCH_0_.latch/Q mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_12 vpwr vgnd scs8hd_fill_2
XFILLER_5_354 vpwr vgnd scs8hd_fill_2
XFILLER_5_376 vpwr vgnd scs8hd_fill_2
XFILLER_3_89 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_2.LATCH_1_.latch data_in mem_bottom_ipin_2.LATCH_1_.latch/Q _181_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_6_129 vgnd vpwr scs8hd_decap_3
XFILLER_10_103 vpwr vgnd scs8hd_fill_2
XFILLER_10_147 vgnd vpwr scs8hd_decap_4
XFILLER_10_169 vpwr vgnd scs8hd_fill_2
XFILLER_12_10 vpwr vgnd scs8hd_fill_2
XFILLER_2_346 vgnd vpwr scs8hd_decap_8
XFILLER_2_335 vgnd vpwr scs8hd_fill_1
XFILLER_2_313 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_ipin_3.LATCH_3_.latch_SLEEPB _126_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__124__A _070_/X vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_ipin_4.LATCH_3_.latch/Q mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _166_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_200_ chanx_right_in[2] chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_15_228 vpwr vgnd scs8hd_fill_2
XFILLER_15_217 vpwr vgnd scs8hd_fill_2
XFILLER_15_206 vgnd vpwr scs8hd_decap_8
XANTENNA__209__A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
X_131_ _131_/A _131_/X vgnd vpwr scs8hd_buf_1
XFILLER_7_405 vpwr vgnd scs8hd_fill_2
XFILLER_2_154 vpwr vgnd scs8hd_fill_2
XFILLER_0_24 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__119__A _106_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_77 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_242 vgnd vpwr scs8hd_decap_6
X_114_ _114_/A _113_/X _115_/A vgnd vpwr scs8hd_or2_4
Xmem_top_ipin_5.LATCH_0_.latch data_in mem_top_ipin_5.LATCH_0_.latch/Q _146_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_286 vpwr vgnd scs8hd_fill_2
XFILLER_11_297 vpwr vgnd scs8hd_fill_2
XANTENNA__121__B _115_/X vgnd vpwr scs8hd_diode_2
XFILLER_19_342 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _190_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_20_32 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_0_.latch/Q mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_87 vgnd vpwr scs8hd_decap_6
XFILLER_16_389 vgnd vpwr scs8hd_decap_8
Xmem_top_ipin_7.LATCH_3_.latch data_in mem_top_ipin_7.LATCH_3_.latch/Q _159_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_6.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__116__B _115_/X vgnd vpwr scs8hd_diode_2
XANTENNA__132__A _070_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_172 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_ipin_1.LATCH_4_.latch_SLEEPB _103_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _183_/HI mem_bottom_ipin_0.LATCH_5_.latch/Q
+ mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_ipin_4.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_319 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_5.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_186 vpwr vgnd scs8hd_fill_2
XANTENNA__127__A _106_/X vgnd vpwr scs8hd_diode_2
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_385 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_318 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_4.LATCH_1_.latch/Q mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_46 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_5.INVTX1_0_.scs8hd_inv_1 chanx_left_in[3] mux_top_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_369 vgnd vpwr scs8hd_fill_1
XFILLER_18_215 vgnd vpwr scs8hd_decap_12
XANTENNA__124__B _123_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_130 vgnd vpwr scs8hd_decap_3
XFILLER_5_163 vgnd vpwr scs8hd_decap_3
XFILLER_5_174 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_6.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_top_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_380 vpwr vgnd scs8hd_fill_2
XANTENNA__140__A _139_/X vgnd vpwr scs8hd_diode_2
XFILLER_17_281 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_0_ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_130_ _099_/A _175_/B _073_/Y _114_/A _131_/A vgnd vpwr scs8hd_or4_4
XFILLER_2_122 vgnd vpwr scs8hd_fill_1
XFILLER_2_100 vgnd vpwr scs8hd_fill_1
XFILLER_2_188 vpwr vgnd scs8hd_fill_2
XFILLER_2_144 vpwr vgnd scs8hd_fill_2
XFILLER_14_240 vgnd vpwr scs8hd_decap_8
XFILLER_0_58 vpwr vgnd scs8hd_fill_2
XANTENNA__119__B _115_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_23 vpwr vgnd scs8hd_fill_2
XANTENNA__135__A _106_/X vgnd vpwr scs8hd_diode_2
X_113_ _113_/A _113_/X vgnd vpwr scs8hd_buf_1
XFILLER_11_265 vpwr vgnd scs8hd_fill_2
XFILLER_7_258 vpwr vgnd scs8hd_fill_2
XFILLER_19_354 vgnd vpwr scs8hd_decap_12
XFILLER_15_7 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_6.LATCH_0_.latch/Q mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_44 vgnd vpwr scs8hd_decap_12
XFILLER_4_206 vpwr vgnd scs8hd_fill_2
XFILLER_4_228 vgnd vpwr scs8hd_decap_12
XFILLER_6_24 vgnd vpwr scs8hd_decap_6
XANTENNA__132__B _131_/X vgnd vpwr scs8hd_diode_2
XFILLER_19_184 vgnd vpwr scs8hd_decap_12
XFILLER_15_11 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_ipin_3.LATCH_3_.latch/Q mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_16_132 vpwr vgnd scs8hd_fill_2
XFILLER_0_275 vpwr vgnd scs8hd_fill_2
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_154 vgnd vpwr scs8hd_decap_4
XFILLER_12_382 vgnd vpwr scs8hd_decap_12
XANTENNA__127__B _123_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_320 vpwr vgnd scs8hd_fill_2
XANTENNA__143__A _105_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_0.LATCH_4_.latch data_in mem_top_ipin_0.LATCH_4_.latch/Q _081_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_179 vpwr vgnd scs8hd_fill_2
XFILLER_13_157 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_25 vpwr vgnd scs8hd_fill_2
XFILLER_3_58 vgnd vpwr scs8hd_decap_3
XFILLER_3_69 vpwr vgnd scs8hd_fill_2
XANTENNA__138__A _098_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_161 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_ipin_6.LATCH_4_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_109 vpwr vgnd scs8hd_fill_2
XFILLER_12_23 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_2_.latch/Q mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_227 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_ipin_7.LATCH_4_.latch/Q mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_293 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_3.INVTX1_0_.scs8hd_inv_1 chanx_left_in[1] mux_top_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_403 vgnd vpwr scs8hd_decap_4
XFILLER_3_3 vpwr vgnd scs8hd_fill_2
XFILLER_2_167 vgnd vpwr scs8hd_decap_4
XFILLER_14_252 vgnd vpwr scs8hd_fill_1
XFILLER_0_37 vpwr vgnd scs8hd_fill_2
XFILLER_9_35 vpwr vgnd scs8hd_fill_2
X_189_ _189_/HI _189_/LO vgnd vpwr scs8hd_conb_1
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
XANTENNA__135__B _131_/X vgnd vpwr scs8hd_diode_2
XANTENNA__151__A _105_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_211 vgnd vpwr scs8hd_decap_6
Xmux_top_ipin_4.INVTX1_4_.scs8hd_inv_1 chanx_left_in[7] mux_top_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_bottom_ipin_0.LATCH_4_.latch data_in mem_bottom_ipin_0.LATCH_4_.latch/Q _170_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_18_11 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_55 vgnd vpwr scs8hd_decap_12
X_112_ _175_/A address[4] _073_/Y _113_/A vgnd vpwr scs8hd_or3_4
XFILLER_7_204 vpwr vgnd scs8hd_fill_2
XFILLER_11_233 vpwr vgnd scs8hd_fill_2
XFILLER_19_377 vpwr vgnd scs8hd_fill_2
XANTENNA__146__A _110_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _191_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_56 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_ipin_4.LATCH_5_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_3.LATCH_1_.latch/Q mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_47 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_3_295 vpwr vgnd scs8hd_fill_2
XFILLER_19_196 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_1.LATCH_0_.latch data_in mem_top_ipin_1.LATCH_0_.latch/Q _111_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_78 vpwr vgnd scs8hd_fill_2
XFILLER_15_67 vpwr vgnd scs8hd_fill_2
XFILLER_15_45 vgnd vpwr scs8hd_decap_4
XFILLER_15_34 vgnd vpwr scs8hd_fill_1
XFILLER_0_221 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_394 vgnd vpwr scs8hd_decap_3
XFILLER_8_332 vgnd vpwr scs8hd_decap_4
Xmem_top_ipin_3.LATCH_3_.latch data_in mem_top_ipin_3.LATCH_3_.latch/Q _126_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__143__B _146_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_398 vgnd vpwr scs8hd_decap_8
XFILLER_13_136 vpwr vgnd scs8hd_fill_2
XFILLER_13_114 vpwr vgnd scs8hd_fill_2
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_7.LATCH_2_.latch/Q mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_335 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__138__B address[5] vgnd vpwr scs8hd_diode_2
XANTENNA__154__A _110_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_327 vpwr vgnd scs8hd_fill_2
XFILLER_2_305 vpwr vgnd scs8hd_fill_2
XFILLER_5_7 vpwr vgnd scs8hd_fill_2
XFILLER_12_46 vgnd vpwr scs8hd_decap_3
XFILLER_18_239 vgnd vpwr scs8hd_decap_12
XFILLER_1_360 vgnd vpwr scs8hd_decap_4
XFILLER_5_187 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_1.LATCH_0_.latch data_in _166_/A _164_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__149__A _177_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_404 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_5.LATCH_0_.latch/Q mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_188_ _188_/HI _188_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__151__B _150_/B vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_2.LATCH_3_.latch/Q mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
Xmux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_67 vgnd vpwr scs8hd_decap_12
XFILLER_11_212 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_1.INVTX1_0_.scs8hd_inv_1 chanx_left_in[3] mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_7_238 vgnd vpwr scs8hd_decap_4
X_111_ _110_/X _105_/B _111_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_245 vpwr vgnd scs8hd_fill_2
XFILLER_19_367 vgnd vpwr scs8hd_decap_6
XANTENNA__146__B _146_/B vgnd vpwr scs8hd_diode_2
XANTENNA__162__A _174_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_260 vpwr vgnd scs8hd_fill_2
XFILLER_1_81 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_3.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__072__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_16_337 vgnd vpwr scs8hd_decap_12
XFILLER_16_304 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_2.INVTX1_4_.scs8hd_inv_1 chanx_left_in[5] mux_top_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_252 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_7.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_3_274 vpwr vgnd scs8hd_fill_2
XFILLER_15_381 vgnd vpwr scs8hd_decap_12
XANTENNA__157__A _177_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
XANTENNA__067__A address[0] vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_6.LATCH_2_.latch data_in mem_top_ipin_6.LATCH_2_.latch/Q _152_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_ipin_6.LATCH_4_.latch/Q mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_0_299 vgnd vpwr scs8hd_fill_1
XFILLER_0_244 vpwr vgnd scs8hd_fill_2
XFILLER_0_200 vgnd vpwr scs8hd_fill_1
XFILLER_16_145 vgnd vpwr scs8hd_decap_8
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_351 vpwr vgnd scs8hd_fill_2
XFILLER_8_366 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _165_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_358 vpwr vgnd scs8hd_fill_2
XANTENNA__154__B _150_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_152 vgnd vpwr scs8hd_fill_1
XANTENNA__170__A _178_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_3.LATCH_0_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_118 vpwr vgnd scs8hd_fill_2
XANTENNA__080__A _080_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_58 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_ipin_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_SLEEPB _178_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__149__B _150_/B vgnd vpwr scs8hd_diode_2
XANTENNA__165__A _165_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_2.LATCH_1_.latch/Q mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__075__A _075_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_136 vpwr vgnd scs8hd_fill_2
XFILLER_2_125 vpwr vgnd scs8hd_fill_2
XFILLER_2_103 vpwr vgnd scs8hd_fill_2
XFILLER_14_276 vgnd vpwr scs8hd_decap_6
X_187_ _187_/HI _187_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_18_79 vgnd vpwr scs8hd_decap_12
XFILLER_18_35 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_110_ _174_/A _110_/X vgnd vpwr scs8hd_buf_1
XFILLER_7_217 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_5.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA__162__B _156_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_6.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_272 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _183_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _192_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_71 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_ipin_7.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_1.LATCH_1_.latch_SLEEPB _109_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_6.LATCH_2_.latch/Q mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_404 vgnd vpwr scs8hd_decap_3
XFILLER_16_349 vgnd vpwr scs8hd_decap_12
XFILLER_16_316 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_220 vpwr vgnd scs8hd_fill_2
XFILLER_10_91 vgnd vpwr scs8hd_fill_1
XFILLER_19_132 vpwr vgnd scs8hd_fill_2
XFILLER_19_110 vgnd vpwr scs8hd_decap_12
XFILLER_15_393 vgnd vpwr scs8hd_decap_12
XFILLER_15_360 vgnd vpwr scs8hd_fill_1
XANTENNA__157__B _156_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__173__A _108_/A vgnd vpwr scs8hd_diode_2
XANTENNA__083__A _086_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_124 vgnd vpwr scs8hd_decap_8
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_4.LATCH_0_.latch/Q mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_301 vgnd vpwr scs8hd_decap_4
XFILLER_8_389 vgnd vpwr scs8hd_decap_8
Xmux_top_ipin_0.INVTX1_4_.scs8hd_inv_1 chanx_left_in[7] mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__168__A _167_/X vgnd vpwr scs8hd_diode_2
XANTENNA__078__A _070_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_315 vpwr vgnd scs8hd_fill_2
XFILLER_5_326 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_top_ipin_1.LATCH_3_.latch/Q mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XANTENNA__170__B _174_/B vgnd vpwr scs8hd_diode_2
XFILLER_12_182 vpwr vgnd scs8hd_fill_2
XFILLER_8_186 vgnd vpwr scs8hd_decap_3
XFILLER_4_381 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_6.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_top_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_6_ vgnd vpwr scs8hd_inv_1
XFILLER_5_178 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_241 vgnd vpwr scs8hd_decap_3
XANTENNA__181__A _108_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_7.INVTX1_5_.scs8hd_inv_1 chanx_right_in[5] mux_top_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__091__A _094_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_148 vpwr vgnd scs8hd_fill_2
XFILLER_14_222 vpwr vgnd scs8hd_fill_2
XFILLER_9_27 vpwr vgnd scs8hd_fill_2
X_186_ _186_/HI _186_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_170 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_2_.latch/Q mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__176__A _176_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_ipin_5.LATCH_4_.latch/Q mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_18_47 vgnd vpwr scs8hd_decap_4
XANTENNA__086__A _086_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_3 vpwr vgnd scs8hd_fill_2
XFILLER_10_291 vpwr vgnd scs8hd_fill_2
X_169_ _177_/A _174_/B _169_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_328 vgnd vpwr scs8hd_decap_8
XFILLER_3_243 vgnd vpwr scs8hd_fill_1
XANTENNA__173__B _174_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_15_15 vgnd vpwr scs8hd_fill_1
XFILLER_13_309 vpwr vgnd scs8hd_fill_2
XANTENNA__083__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_0_213 vpwr vgnd scs8hd_fill_2
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_169 vpwr vgnd scs8hd_fill_2
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_324 vpwr vgnd scs8hd_fill_2
XFILLER_8_346 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_1.LATCH_1_.latch/Q mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_15_191 vpwr vgnd scs8hd_fill_2
XANTENNA__078__B _094_/A vgnd vpwr scs8hd_diode_2
XANTENNA__094__A _094_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_6.LATCH_1_.latch_SLEEPB _153_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_29 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_2.LATCH_2_.latch data_in mem_top_ipin_2.LATCH_2_.latch/Q _119_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_91 vgnd vpwr scs8hd_fill_1
XANTENNA__179__A _179_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_27 vpwr vgnd scs8hd_fill_2
XANTENNA__089__A address[1] vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_4.LATCH_5_.latch data_in mem_top_ipin_4.LATCH_5_.latch/Q _132_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_146 vpwr vgnd scs8hd_fill_2
XFILLER_5_168 vgnd vpwr scs8hd_decap_3
XANTENNA__181__B _178_/B vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_5.LATCH_2_.latch/Q mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_190 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__091__B _108_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_256 vgnd vpwr scs8hd_decap_8
XFILLER_14_201 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_4.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_top_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_185_ _185_/HI _185_/LO vgnd vpwr scs8hd_conb_1
XFILLER_14_267 vgnd vpwr scs8hd_decap_8
XFILLER_13_92 vgnd vpwr scs8hd_decap_3
XFILLER_9_39 vpwr vgnd scs8hd_fill_2
XFILLER_1_193 vpwr vgnd scs8hd_fill_2
XFILLER_9_260 vpwr vgnd scs8hd_fill_2
XFILLER_9_282 vpwr vgnd scs8hd_fill_2
XFILLER_9_293 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_3.LATCH_0_.latch/Q mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__086__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_2.LATCH_2_.latch data_in mem_bottom_ipin_2.LATCH_2_.latch/Q _180_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_237 vgnd vpwr scs8hd_decap_4
XFILLER_3_403 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_5.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_top_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_4.LATCH_2_.latch_SLEEPB _135_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
X_168_ _167_/X _174_/B vgnd vpwr scs8hd_buf_1
XFILLER_6_241 vgnd vpwr scs8hd_decap_4
XFILLER_6_285 vgnd vpwr scs8hd_decap_8
X_099_ _099_/A address[4] _175_/C _114_/A _099_/X vgnd vpwr scs8hd_or4_4
XFILLER_1_40 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _193_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA__097__A address[6] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_ipin_0.LATCH_3_.latch/Q mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_3_233 vgnd vpwr scs8hd_decap_4
XFILLER_3_255 vpwr vgnd scs8hd_fill_2
XFILLER_3_299 vgnd vpwr scs8hd_decap_4
XFILLER_10_93 vgnd vpwr scs8hd_decap_3
XFILLER_19_123 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_49 vgnd vpwr scs8hd_fill_1
XFILLER_15_27 vgnd vpwr scs8hd_decap_4
XANTENNA__083__C _068_/C vgnd vpwr scs8hd_diode_2
XFILLER_0_269 vgnd vpwr scs8hd_decap_4
XFILLER_0_258 vpwr vgnd scs8hd_fill_2
XFILLER_0_225 vpwr vgnd scs8hd_fill_2
XFILLER_0_203 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_7.LATCH_1_.latch/Q mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_365 vpwr vgnd scs8hd_fill_2
XFILLER_12_321 vgnd vpwr scs8hd_decap_6
XFILLER_12_310 vgnd vpwr scs8hd_decap_8
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_398 vgnd vpwr scs8hd_decap_8
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_15_181 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_5.LATCH_1_.latch data_in mem_top_ipin_5.LATCH_1_.latch/Q _145_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_380 vpwr vgnd scs8hd_fill_2
XANTENNA__094__B _174_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
XFILLER_8_100 vgnd vpwr scs8hd_decap_3
XFILLER_8_166 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_ipin_4.LATCH_4_.latch/Q mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_12_140 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_394 vgnd vpwr scs8hd_decap_3
XANTENNA__179__B _178_/B vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_7.LATCH_4_.latch data_in mem_top_ipin_7.LATCH_4_.latch/Q _158_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__195__A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_2.LATCH_3_.latch_SLEEPB _118_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_309 vgnd vpwr scs8hd_decap_4
XANTENNA__089__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_5_103 vpwr vgnd scs8hd_fill_2
XFILLER_1_353 vgnd vpwr scs8hd_fill_1
XFILLER_5_114 vpwr vgnd scs8hd_fill_2
XFILLER_17_221 vgnd vpwr scs8hd_decap_12
XFILLER_4_84 vpwr vgnd scs8hd_fill_2
XFILLER_4_180 vgnd vpwr scs8hd_decap_4
XFILLER_3_8 vpwr vgnd scs8hd_fill_2
XFILLER_14_213 vgnd vpwr scs8hd_fill_1
X_184_ _184_/HI _184_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_71 vpwr vgnd scs8hd_fill_2
XFILLER_20_249 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_2.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__086__C address[0] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_1_.latch/Q mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_216 vpwr vgnd scs8hd_fill_2
XFILLER_11_249 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
X_167_ _099_/A address[4] _175_/C _175_/D _167_/X vgnd vpwr scs8hd_or4_4
X_098_ _098_/A address[5] _114_/A vgnd vpwr scs8hd_nand2_4
XFILLER_6_264 vgnd vpwr scs8hd_decap_8
XFILLER_10_271 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_96 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_0.LATCH_4_.latch_SLEEPB _081_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_6_ vgnd vpwr scs8hd_inv_1
XFILLER_3_201 vpwr vgnd scs8hd_fill_2
XFILLER_3_289 vgnd vpwr scs8hd_decap_4
XFILLER_10_72 vpwr vgnd scs8hd_fill_2
XFILLER_10_83 vgnd vpwr scs8hd_decap_8
XFILLER_15_363 vgnd vpwr scs8hd_decap_3
XFILLER_15_352 vpwr vgnd scs8hd_fill_2
XFILLER_15_330 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_3.INVTX1_5_.scs8hd_inv_1 chanx_right_in[6] mux_top_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__198__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_18_190 vgnd vpwr scs8hd_decap_12
XFILLER_15_39 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_ipin_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_3.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_355 vgnd vpwr scs8hd_fill_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_4.LATCH_2_.latch/Q mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_ipin_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_7_40 vpwr vgnd scs8hd_fill_2
XFILLER_17_403 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_178 vgnd vpwr scs8hd_decap_6
XFILLER_12_152 vgnd vpwr scs8hd_fill_1
XFILLER_4_340 vpwr vgnd scs8hd_fill_2
XFILLER_4_362 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_2.LATCH_0_.latch/Q mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_SLEEPB _181_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__089__C _068_/C vgnd vpwr scs8hd_diode_2
XFILLER_14_406 vgnd vpwr scs8hd_fill_1
XFILLER_5_126 vpwr vgnd scs8hd_fill_2
XFILLER_1_376 vpwr vgnd scs8hd_fill_2
XFILLER_1_332 vpwr vgnd scs8hd_fill_2
XFILLER_17_233 vgnd vpwr scs8hd_decap_8
XFILLER_1_398 vpwr vgnd scs8hd_fill_2
XFILLER_1_387 vgnd vpwr scs8hd_decap_8
XFILLER_4_41 vpwr vgnd scs8hd_fill_2
XFILLER_4_52 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_7.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_118 vgnd vpwr scs8hd_decap_4
X_183_ _183_/HI _183_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_top_ipin_4.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_0.LATCH_5_.latch data_in mem_top_ipin_0.LATCH_5_.latch/Q _078_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_top_ipin_7.LATCH_3_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_6.LATCH_1_.latch/Q mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_306 vgnd vpwr scs8hd_decap_12
XFILLER_6_210 vpwr vgnd scs8hd_fill_2
X_097_ address[6] _098_/A vgnd vpwr scs8hd_inv_8
X_166_ _166_/A _166_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_20 vpwr vgnd scs8hd_fill_2
XFILLER_1_53 vpwr vgnd scs8hd_fill_2
XFILLER_18_361 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _185_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_SLEEPB _172_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_3.LATCH_4_.latch/Q mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_19_136 vgnd vpwr scs8hd_decap_12
XFILLER_19_60 vgnd vpwr scs8hd_fill_1
XFILLER_15_342 vgnd vpwr scs8hd_decap_6
X_149_ _177_/A _150_/B _149_/Y vgnd vpwr scs8hd_nor2_4
Xmux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_305 vgnd vpwr scs8hd_fill_1
Xmem_bottom_ipin_0.LATCH_5_.latch data_in mem_bottom_ipin_0.LATCH_5_.latch/Q _169_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_150 vgnd vpwr scs8hd_decap_4
XPHY_3 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_7_74 vpwr vgnd scs8hd_fill_2
XFILLER_7_85 vpwr vgnd scs8hd_fill_2
XFILLER_7_393 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_1.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_top_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_319 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_5.LATCH_4_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _193_/HI mem_top_ipin_7.LATCH_5_.latch/Q
+ mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_12_186 vpwr vgnd scs8hd_fill_2
XFILLER_8_146 vgnd vpwr scs8hd_decap_6
XFILLER_8_157 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_12_ vgnd vpwr scs8hd_inv_1
Xmem_top_ipin_1.LATCH_1_.latch data_in mem_top_ipin_1.LATCH_1_.latch/Q _109_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_ipin_7.INVTX1_2_.scs8hd_inv_1 chanx_left_in[1] mux_top_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_245 vgnd vpwr scs8hd_decap_12
XFILLER_17_201 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_3.LATCH_4_.latch data_in mem_top_ipin_3.LATCH_4_.latch/Q _125_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_248 vpwr vgnd scs8hd_fill_2
X_182_ _174_/A _178_/B _182_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_51 vgnd vpwr scs8hd_decap_4
XFILLER_1_174 vgnd vpwr scs8hd_fill_1
XANTENNA__100__A _099_/X vgnd vpwr scs8hd_diode_2
XFILLER_20_218 vgnd vpwr scs8hd_decap_12
XFILLER_13_281 vpwr vgnd scs8hd_fill_2
XFILLER_9_241 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_3.LATCH_2_.latch/Q mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_229 vpwr vgnd scs8hd_fill_2
XFILLER_19_318 vgnd vpwr scs8hd_decap_12
XFILLER_1_7 vpwr vgnd scs8hd_fill_2
X_165_ _165_/A _165_/Y vgnd vpwr scs8hd_inv_8
XFILLER_10_251 vgnd vpwr scs8hd_fill_1
XFILLER_10_295 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_3.LATCH_5_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
X_096_ address[3] _175_/C vgnd vpwr scs8hd_buf_1
XFILLER_18_373 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_1.LATCH_1_.latch data_in _165_/A _163_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_30 vgnd vpwr scs8hd_fill_1
XFILLER_10_41 vgnd vpwr scs8hd_decap_3
XFILLER_19_148 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_1.LATCH_0_.latch/Q mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
X_148_ _147_/X _150_/B vgnd vpwr scs8hd_buf_1
X_079_ address[1] _068_/B address[0] _080_/A vgnd vpwr scs8hd_or3_4
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_107 vgnd vpwr scs8hd_decap_8
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_335 vgnd vpwr scs8hd_fill_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_346 vgnd vpwr scs8hd_decap_3
XFILLER_8_328 vpwr vgnd scs8hd_fill_2
XFILLER_15_173 vgnd vpwr scs8hd_decap_8
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_7_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_165 vpwr vgnd scs8hd_fill_2
XFILLER_8_125 vpwr vgnd scs8hd_fill_2
XFILLER_8_136 vgnd vpwr scs8hd_decap_8
XFILLER_12_110 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_4.LATCH_0_.latch data_in mem_top_ipin_4.LATCH_0_.latch/Q _137_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__103__A _150_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_386 vgnd vpwr scs8hd_decap_8
Xmux_top_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_5.LATCH_1_.latch/Q mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_301 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_356 vpwr vgnd scs8hd_fill_2
XFILLER_17_257 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_6.LATCH_3_.latch data_in mem_top_ipin_6.LATCH_3_.latch/Q _151_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_65 vpwr vgnd scs8hd_fill_2
XFILLER_4_150 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_2.LATCH_4_.latch/Q mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_14_205 vgnd vpwr scs8hd_decap_8
X_181_ _108_/A _178_/B _181_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_197 vpwr vgnd scs8hd_fill_2
XFILLER_1_153 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_5.INVTX1_2_.scs8hd_inv_1 chanx_left_in[7] mux_top_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_220 vpwr vgnd scs8hd_fill_2
XFILLER_9_264 vgnd vpwr scs8hd_decap_4
XFILLER_9_286 vpwr vgnd scs8hd_fill_2
XFILLER_9_297 vpwr vgnd scs8hd_fill_2
XFILLER_18_19 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_3.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__201__A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
X_095_ _175_/A _099_/A vgnd vpwr scs8hd_buf_1
X_164_ _175_/D _113_/X address[0] _164_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_10_230 vgnd vpwr scs8hd_decap_4
XFILLER_18_385 vgnd vpwr scs8hd_decap_12
XFILLER_1_77 vpwr vgnd scs8hd_fill_2
XANTENNA__111__A _110_/X vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _192_/HI mem_top_ipin_6.LATCH_5_.latch/Q
+ mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_3_248 vgnd vpwr scs8hd_decap_4
XFILLER_10_53 vpwr vgnd scs8hd_fill_2
XFILLER_19_62 vgnd vpwr scs8hd_decap_12
XFILLER_19_40 vgnd vpwr scs8hd_fill_1
XFILLER_15_377 vpwr vgnd scs8hd_fill_2
XANTENNA__106__A _106_/A vgnd vpwr scs8hd_diode_2
X_147_ _113_/X _147_/B _147_/X vgnd vpwr scs8hd_or2_4
X_078_ _070_/X _094_/A _078_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_229 vpwr vgnd scs8hd_fill_2
XFILLER_0_207 vgnd vpwr scs8hd_decap_4
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_369 vgnd vpwr scs8hd_decap_4
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_7_21 vpwr vgnd scs8hd_fill_2
XFILLER_7_32 vpwr vgnd scs8hd_fill_2
XFILLER_11_380 vpwr vgnd scs8hd_fill_2
XFILLER_7_65 vpwr vgnd scs8hd_fill_2
XFILLER_7_362 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_2.LATCH_0_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_96 vgnd vpwr scs8hd_decap_8
XFILLER_12_199 vpwr vgnd scs8hd_fill_2
XANTENNA__103__B _105_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_332 vgnd vpwr scs8hd_decap_4
XFILLER_4_398 vgnd vpwr scs8hd_decap_8
Xmux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_2.LATCH_2_.latch/Q mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__204__A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_5_118 vpwr vgnd scs8hd_fill_2
XFILLER_17_269 vgnd vpwr scs8hd_decap_12
XFILLER_4_22 vgnd vpwr scs8hd_decap_3
XFILLER_4_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__114__A _114_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_280 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_0_.latch/Q mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_97 vpwr vgnd scs8hd_fill_2
XFILLER_13_75 vpwr vgnd scs8hd_fill_2
X_180_ _106_/A _178_/B _180_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_5.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_13_294 vpwr vgnd scs8hd_fill_2
XANTENNA__109__A _108_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_254 vgnd vpwr scs8hd_decap_4
X_094_ _094_/A _174_/A _094_/Y vgnd vpwr scs8hd_nor2_4
X_163_ _175_/D _113_/X _068_/C _163_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_6_224 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_4.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_1_.latch_SLEEPB _091_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__111__B _105_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_5.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_3.INVTX1_2_.scs8hd_inv_1 chanx_left_in[5] mux_top_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_ipin_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_216 vpwr vgnd scs8hd_fill_2
XFILLER_10_76 vpwr vgnd scs8hd_fill_2
XFILLER_19_74 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_4.LATCH_1_.latch/Q mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_367 vgnd vpwr scs8hd_decap_4
XFILLER_15_356 vgnd vpwr scs8hd_decap_4
X_146_ _110_/X _146_/B _146_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__122__A _099_/A vgnd vpwr scs8hd_diode_2
X_077_ _077_/A _094_/A vgnd vpwr scs8hd_buf_1
XFILLER_2_271 vpwr vgnd scs8hd_fill_2
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__207__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_308 vgnd vpwr scs8hd_fill_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_6 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_ipin_1.LATCH_4_.latch/Q mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XANTENNA__117__A _150_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_392 vgnd vpwr scs8hd_decap_4
X_129_ _110_/X _123_/X _129_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_8_105 vgnd vpwr scs8hd_decap_3
XFILLER_12_123 vgnd vpwr scs8hd_decap_4
XFILLER_4_344 vpwr vgnd scs8hd_fill_2
XFILLER_4_366 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_160 vpwr vgnd scs8hd_fill_2
XFILLER_1_336 vpwr vgnd scs8hd_fill_2
XANTENNA__114__B _113_/X vgnd vpwr scs8hd_diode_2
XFILLER_0_391 vgnd vpwr scs8hd_decap_12
XFILLER_0_380 vgnd vpwr scs8hd_decap_4
XANTENNA__130__A _099_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_45 vgnd vpwr scs8hd_decap_4
XFILLER_4_163 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _191_/HI mem_top_ipin_5.LATCH_5_.latch/Q
+ mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_16_292 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_7.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_0.LATCH_0_.latch data_in mem_top_ipin_0.LATCH_0_.latch/Q _094_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_229 vgnd vpwr scs8hd_decap_8
XFILLER_14_218 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_7.LATCH_0_.latch_SLEEPB _162_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_406 vgnd vpwr scs8hd_fill_1
XFILLER_1_177 vgnd vpwr scs8hd_decap_4
XFILLER_1_166 vpwr vgnd scs8hd_fill_2
XFILLER_1_100 vpwr vgnd scs8hd_fill_2
XFILLER_8_3 vpwr vgnd scs8hd_fill_2
XANTENNA__109__B _105_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_233 vpwr vgnd scs8hd_fill_2
XANTENNA__125__A _150_/A vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_2.LATCH_3_.latch data_in mem_top_ipin_2.LATCH_3_.latch/Q _118_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_162_ _174_/A _156_/X _162_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_243 vpwr vgnd scs8hd_fill_2
X_093_ _092_/X _174_/A vgnd vpwr scs8hd_buf_1
XFILLER_6_203 vgnd vpwr scs8hd_decap_4
XFILLER_6_247 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_254 vpwr vgnd scs8hd_fill_2
XFILLER_10_287 vpwr vgnd scs8hd_fill_2
XFILLER_1_24 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_398 vgnd vpwr scs8hd_decap_8
XFILLER_1_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_239 vpwr vgnd scs8hd_fill_2
XFILLER_10_22 vpwr vgnd scs8hd_fill_2
XFILLER_10_99 vpwr vgnd scs8hd_fill_2
XFILLER_19_86 vgnd vpwr scs8hd_decap_12
X_145_ _108_/X _146_/B _145_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_1.LATCH_2_.latch/Q mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_076_ _175_/A _175_/B _073_/Y _175_/D _077_/A vgnd vpwr scs8hd_or4_4
XANTENNA__122__B _175_/B vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_0.LATCH_0_.latch data_in mem_bottom_ipin_0.LATCH_0_.latch/Q _174_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_ipin_1.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_top_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_198 vpwr vgnd scs8hd_fill_2
XFILLER_15_187 vpwr vgnd scs8hd_fill_2
XFILLER_15_132 vgnd vpwr scs8hd_decap_4
XPHY_7 vgnd vpwr scs8hd_decap_3
X_128_ _108_/X _123_/X _128_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__117__B _115_/X vgnd vpwr scs8hd_diode_2
XFILLER_7_89 vpwr vgnd scs8hd_fill_2
XANTENNA__133__A _150_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_5.LATCH_1_.latch_SLEEPB _145_/Y vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_2.LATCH_3_.latch data_in mem_bottom_ipin_2.LATCH_3_.latch/Q _179_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__128__A _108_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_315 vpwr vgnd scs8hd_fill_2
XFILLER_17_205 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_142 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__130__B _175_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_186 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_3.LATCH_1_.latch/Q mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_33 vpwr vgnd scs8hd_fill_2
XFILLER_13_88 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_5.LATCH_2_.latch data_in mem_top_ipin_5.LATCH_2_.latch/Q _144_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_13_263 vgnd vpwr scs8hd_fill_1
XANTENNA__125__B _123_/X vgnd vpwr scs8hd_diode_2
XANTENNA__141__A _070_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_3.LATCH_2_.latch_SLEEPB _127_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_7.LATCH_5_.latch data_in mem_top_ipin_7.LATCH_5_.latch/Q _157_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_ipin_0.LATCH_4_.latch/Q mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
X_161_ _108_/A _156_/X _161_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_211 vgnd vpwr scs8hd_fill_1
X_092_ address[1] address[2] address[0] _092_/X vgnd vpwr scs8hd_or3_4
XFILLER_18_300 vgnd vpwr scs8hd_decap_12
XFILLER_1_36 vpwr vgnd scs8hd_fill_2
XANTENNA__136__A _108_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_98 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_7.LATCH_2_.latch/Q mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
X_144_ _106_/X _146_/B _144_/Y vgnd vpwr scs8hd_nor2_4
X_075_ _075_/A _175_/D vgnd vpwr scs8hd_buf_1
XANTENNA__122__C _175_/C vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_0_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_141 vpwr vgnd scs8hd_fill_2
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _190_/HI mem_top_ipin_4.LATCH_5_.latch/Q
+ mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XPHY_8 vgnd vpwr scs8hd_decap_3
X_127_ _106_/X _123_/X _127_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_57 vpwr vgnd scs8hd_fill_2
XANTENNA__133__B _131_/X vgnd vpwr scs8hd_diode_2
XFILLER_7_343 vgnd vpwr scs8hd_decap_4
XFILLER_7_376 vpwr vgnd scs8hd_fill_2
XFILLER_16_3 vgnd vpwr scs8hd_decap_3
XFILLER_12_169 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_1.LATCH_3_.latch_SLEEPB _105_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_180 vgnd vpwr scs8hd_decap_6
XFILLER_4_302 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__128__B _123_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__144__A _106_/X vgnd vpwr scs8hd_diode_2
XFILLER_7_184 vgnd vpwr scs8hd_decap_4
XFILLER_1_349 vgnd vpwr scs8hd_decap_4
XFILLER_9_405 vpwr vgnd scs8hd_fill_2
XFILLER_4_121 vpwr vgnd scs8hd_fill_2
XANTENNA__130__C _073_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_360 vgnd vpwr scs8hd_decap_6
XFILLER_4_69 vpwr vgnd scs8hd_fill_2
XANTENNA__139__A _099_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_13_12 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_2_.latch/Q mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_113 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_9_268 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__141__B _146_/B vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_6.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_top_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_091_ _094_/A _108_/A _091_/Y vgnd vpwr scs8hd_nor2_4
X_160_ _106_/A _156_/X _160_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_201 vpwr vgnd scs8hd_fill_2
XFILLER_10_267 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_312 vgnd vpwr scs8hd_decap_12
XANTENNA__136__B _131_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_260 vgnd vpwr scs8hd_decap_4
XANTENNA__152__A _106_/X vgnd vpwr scs8hd_diode_2
XFILLER_10_46 vgnd vpwr scs8hd_decap_3
XFILLER_10_57 vpwr vgnd scs8hd_fill_2
XFILLER_19_44 vpwr vgnd scs8hd_fill_2
XFILLER_19_22 vgnd vpwr scs8hd_decap_12
XFILLER_19_11 vgnd vpwr scs8hd_decap_4
XFILLER_15_348 vgnd vpwr scs8hd_fill_1
XFILLER_15_304 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_074_ address[6] address[5] _075_/A vgnd vpwr scs8hd_or2_4
X_143_ _105_/A _146_/B _143_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_263 vpwr vgnd scs8hd_fill_2
XANTENNA__122__D _114_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_7 vpwr vgnd scs8hd_fill_2
XANTENNA__147__A _113_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_12_329 vgnd vpwr scs8hd_decap_6
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_20_373 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_ipin_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_ipin_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_156 vpwr vgnd scs8hd_fill_2
XFILLER_7_25 vpwr vgnd scs8hd_fill_2
XFILLER_7_36 vpwr vgnd scs8hd_fill_2
XFILLER_11_362 vpwr vgnd scs8hd_fill_2
X_126_ _105_/A _123_/X _126_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_69 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_2.LATCH_1_.latch/Q mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_SLEEPB _163_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_119 vgnd vpwr scs8hd_decap_4
XFILLER_4_369 vgnd vpwr scs8hd_fill_1
XANTENNA__144__B _146_/B vgnd vpwr scs8hd_diode_2
X_109_ _108_/X _105_/B _109_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__160__A _106_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_380 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_281 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__070__A _177_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__130__D _114_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__155__A _099_/A vgnd vpwr scs8hd_diode_2
XANTENNA__139__B address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_5.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_6.LATCH_2_.latch/Q mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_ipin_6.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XFILLER_13_46 vgnd vpwr scs8hd_decap_3
XFILLER_1_136 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_6.LATCH_3_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
XFILLER_13_243 vgnd vpwr scs8hd_fill_1
XFILLER_13_210 vgnd vpwr scs8hd_decap_4
XFILLER_13_298 vgnd vpwr scs8hd_decap_3
XFILLER_0_180 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _189_/HI mem_top_ipin_3.LATCH_5_.latch/Q
+ mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_090_ _089_/X _108_/A vgnd vpwr scs8hd_buf_1
XFILLER_6_228 vpwr vgnd scs8hd_fill_2
XFILLER_6_3 vgnd vpwr scs8hd_decap_4
XFILLER_18_324 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_1.LATCH_2_.latch data_in mem_top_ipin_1.LATCH_2_.latch/Q _107_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_272 vpwr vgnd scs8hd_fill_2
XANTENNA__152__B _150_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_34 vgnd vpwr scs8hd_decap_6
X_142_ _150_/A _146_/B _142_/Y vgnd vpwr scs8hd_nor2_4
X_211_ chanx_left_in[0] chanx_right_out[0] vgnd vpwr scs8hd_buf_2
X_073_ address[3] _073_/Y vgnd vpwr scs8hd_inv_8
Xmem_top_ipin_3.LATCH_5_.latch data_in mem_top_ipin_3.LATCH_5_.latch/Q _124_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_4.INVTX1_3_.scs8hd_inv_1 chanx_right_in[6] mux_top_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_286 vgnd vpwr scs8hd_decap_6
XFILLER_2_242 vgnd vpwr scs8hd_decap_8
XFILLER_18_154 vgnd vpwr scs8hd_decap_12
XANTENNA__147__B _147_/B vgnd vpwr scs8hd_diode_2
XANTENNA__163__A _175_/D vgnd vpwr scs8hd_diode_2
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_385 vgnd vpwr scs8hd_decap_12
XANTENNA__073__A address[3] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_4_ vgnd vpwr scs8hd_inv_1
X_125_ _150_/A _123_/X _125_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_323 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_ipin_4.LATCH_4_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_190 vgnd vpwr scs8hd_decap_8
XANTENNA__158__A _178_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_68 vgnd vpwr scs8hd_decap_8
XFILLER_16_57 vgnd vpwr scs8hd_decap_8
XFILLER_16_46 vgnd vpwr scs8hd_decap_8
XFILLER_16_35 vpwr vgnd scs8hd_fill_2
XANTENNA__068__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_16_79 vgnd vpwr scs8hd_decap_12
XFILLER_4_348 vgnd vpwr scs8hd_decap_3
X_108_ _108_/A _108_/X vgnd vpwr scs8hd_buf_1
XFILLER_7_153 vgnd vpwr scs8hd_fill_1
XFILLER_7_175 vpwr vgnd scs8hd_fill_2
XANTENNA__160__B _156_/X vgnd vpwr scs8hd_diode_2
XFILLER_3_392 vgnd vpwr scs8hd_decap_4
XFILLER_19_293 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_27 vpwr vgnd scs8hd_fill_2
XFILLER_4_49 vgnd vpwr scs8hd_fill_1
XFILLER_4_167 vpwr vgnd scs8hd_fill_2
XFILLER_16_230 vgnd vpwr scs8hd_decap_12
XANTENNA__139__C _175_/C vgnd vpwr scs8hd_diode_2
XFILLER_16_274 vgnd vpwr scs8hd_fill_1
XANTENNA__155__B _175_/B vgnd vpwr scs8hd_diode_2
XANTENNA__171__A _179_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_406 vgnd vpwr scs8hd_fill_1
XANTENNA__081__A _094_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_7 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_277 vpwr vgnd scs8hd_fill_2
XFILLER_13_266 vgnd vpwr scs8hd_decap_8
XFILLER_13_233 vgnd vpwr scs8hd_decap_4
XFILLER_13_200 vgnd vpwr scs8hd_fill_1
XFILLER_9_237 vgnd vpwr scs8hd_decap_4
XANTENNA__166__A _166_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_2.LATCH_5_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_4.LATCH_1_.latch data_in mem_top_ipin_4.LATCH_1_.latch/Q _136_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__076__A _175_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_207 vgnd vpwr scs8hd_fill_1
XFILLER_10_247 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_1.LATCH_1_.latch/Q mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_240 vpwr vgnd scs8hd_fill_2
XFILLER_5_295 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_391 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_6.LATCH_4_.latch data_in mem_top_ipin_6.LATCH_4_.latch/Q _150_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_26 vpwr vgnd scs8hd_fill_2
XFILLER_15_306 vgnd vpwr scs8hd_decap_12
X_141_ _070_/X _146_/B _141_/Y vgnd vpwr scs8hd_nor2_4
X_210_ chanx_left_in[1] chanx_right_out[1] vgnd vpwr scs8hd_buf_2
X_072_ address[4] _175_/B vgnd vpwr scs8hd_inv_8
XFILLER_18_133 vgnd vpwr scs8hd_decap_8
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_18_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__163__B _113_/X vgnd vpwr scs8hd_diode_2
XFILLER_2_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_342 vgnd vpwr scs8hd_decap_12
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_20_397 vgnd vpwr scs8hd_decap_6
XFILLER_15_169 vpwr vgnd scs8hd_fill_2
XFILLER_15_114 vpwr vgnd scs8hd_fill_2
XFILLER_15_103 vpwr vgnd scs8hd_fill_2
X_124_ _070_/X _123_/X _124_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_302 vgnd vpwr scs8hd_fill_1
XFILLER_7_335 vpwr vgnd scs8hd_fill_2
XFILLER_11_320 vgnd vpwr scs8hd_decap_4
XFILLER_11_342 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_5.LATCH_2_.latch/Q mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_80 vpwr vgnd scs8hd_fill_2
XANTENNA__158__B _156_/X vgnd vpwr scs8hd_diode_2
XANTENNA__174__A _174_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_top_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_0_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__068__B _068_/B vgnd vpwr scs8hd_diode_2
XFILLER_12_106 vpwr vgnd scs8hd_fill_2
XANTENNA__084__A _083_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_316 vgnd vpwr scs8hd_decap_3
X_107_ _106_/X _105_/B _107_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_110 vgnd vpwr scs8hd_fill_1
XFILLER_7_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _188_/HI mem_top_ipin_2.LATCH_5_.latch/Q
+ mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__169__A _177_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_81 vpwr vgnd scs8hd_fill_2
XFILLER_1_319 vpwr vgnd scs8hd_fill_2
XFILLER_17_209 vgnd vpwr scs8hd_decap_12
XANTENNA__079__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_13_404 vgnd vpwr scs8hd_decap_3
XFILLER_4_102 vgnd vpwr scs8hd_decap_3
XFILLER_4_146 vgnd vpwr scs8hd_decap_4
XFILLER_16_242 vgnd vpwr scs8hd_decap_12
XANTENNA__139__D _147_/B vgnd vpwr scs8hd_diode_2
XANTENNA__155__C _175_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__171__B _174_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__081__B _178_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_149 vpwr vgnd scs8hd_fill_2
XFILLER_13_245 vgnd vpwr scs8hd_decap_3
Xmem_top_ipin_7.LATCH_0_.latch data_in mem_top_ipin_7.LATCH_0_.latch/Q _162_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_216 vpwr vgnd scs8hd_fill_2
XANTENNA__182__A _174_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_260 vgnd vpwr scs8hd_decap_8
XFILLER_8_282 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_SLEEPB _179_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_60 vgnd vpwr scs8hd_fill_1
XFILLER_5_82 vpwr vgnd scs8hd_fill_2
XANTENNA__076__B _175_/B vgnd vpwr scs8hd_diode_2
XFILLER_10_215 vpwr vgnd scs8hd_fill_2
XFILLER_10_226 vpwr vgnd scs8hd_fill_2
XANTENNA__092__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_1_29 vpwr vgnd scs8hd_fill_2
XFILLER_18_337 vgnd vpwr scs8hd_decap_12
XANTENNA__177__A _177_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_318 vgnd vpwr scs8hd_decap_12
XANTENNA__087__A _086_/X vgnd vpwr scs8hd_diode_2
X_071_ enable _175_/A vgnd vpwr scs8hd_inv_8
X_140_ _139_/X _146_/B vgnd vpwr scs8hd_buf_1
XFILLER_2_222 vpwr vgnd scs8hd_fill_2
XFILLER_18_145 vgnd vpwr scs8hd_decap_8
XFILLER_18_178 vgnd vpwr scs8hd_decap_12
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__163__C _068_/C vgnd vpwr scs8hd_diode_2
XFILLER_20_354 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_ipin_7.LATCH_5_.latch_SLEEPB _157_/Y vgnd vpwr scs8hd_diode_2
X_123_ _122_/X _123_/X vgnd vpwr scs8hd_buf_1
XFILLER_7_358 vpwr vgnd scs8hd_fill_2
XFILLER_11_376 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_1.LATCH_0_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__174__B _174_/B vgnd vpwr scs8hd_diode_2
XANTENNA__068__C _068_/C vgnd vpwr scs8hd_diode_2
XFILLER_12_129 vpwr vgnd scs8hd_fill_2
XFILLER_4_328 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
X_106_ _106_/A _106_/X vgnd vpwr scs8hd_buf_1
XFILLER_7_188 vgnd vpwr scs8hd_fill_1
XFILLER_11_184 vpwr vgnd scs8hd_fill_2
XFILLER_11_195 vpwr vgnd scs8hd_fill_2
XANTENNA__169__B _174_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_1_.latch/Q mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__079__B _068_/B vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[3] mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__095__A _175_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_4_18 vpwr vgnd scs8hd_fill_2
XFILLER_4_125 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_0_331 vpwr vgnd scs8hd_fill_2
XFILLER_0_320 vgnd vpwr scs8hd_decap_3
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XFILLER_16_254 vgnd vpwr scs8hd_decap_12
XANTENNA__155__D _147_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_16 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_2_ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_6.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_top_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__182__B _178_/B vgnd vpwr scs8hd_diode_2
XANTENNA__092__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__076__C _073_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_205 vgnd vpwr scs8hd_decap_6
XFILLER_18_349 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_4.LATCH_2_.latch/Q mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_7.INVTX1_4_.scs8hd_inv_1 chanx_left_in[5] mux_top_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_ipin_3.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__177__B _178_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_48 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_0.LATCH_1_.latch data_in mem_top_ipin_0.LATCH_1_.latch/Q _091_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_070_ _177_/A _070_/X vgnd vpwr scs8hd_buf_1
XFILLER_2_267 vpwr vgnd scs8hd_fill_2
XFILLER_4_3 vpwr vgnd scs8hd_fill_2
XFILLER_18_113 vgnd vpwr scs8hd_decap_12
XFILLER_18_102 vgnd vpwr scs8hd_decap_8
Xmux_top_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _187_/HI mem_top_ipin_1.LATCH_5_.latch/Q
+ mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_14_396 vgnd vpwr scs8hd_fill_1
XPHY_80 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_199_ chanx_right_in[3] chanx_left_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_84 vpwr vgnd scs8hd_fill_2
XFILLER_20_366 vgnd vpwr scs8hd_decap_6
XFILLER_20_311 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_2.LATCH_4_.latch data_in mem_top_ipin_2.LATCH_4_.latch/Q _117_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__098__A _098_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_138 vgnd vpwr scs8hd_decap_3
XFILLER_7_315 vpwr vgnd scs8hd_fill_2
X_122_ _099_/A _175_/B _175_/C _114_/A _122_/X vgnd vpwr scs8hd_or4_4
XFILLER_11_93 vgnd vpwr scs8hd_decap_4
XFILLER_11_388 vpwr vgnd scs8hd_fill_2
XFILLER_11_399 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_7.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
X_105_ _105_/A _105_/B _105_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_156 vpwr vgnd scs8hd_fill_2
XFILLER_3_351 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_7.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_0.LATCH_1_.latch data_in mem_bottom_ipin_0.LATCH_1_.latch/Q _173_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__079__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_0_387 vpwr vgnd scs8hd_fill_2
XFILLER_0_376 vpwr vgnd scs8hd_fill_2
XFILLER_17_81 vgnd vpwr scs8hd_decap_12
XFILLER_16_266 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_ipin_6.LATCH_0_.latch_SLEEPB _154_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__196__A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_2.LATCH_4_.latch data_in mem_bottom_ipin_2.LATCH_4_.latch/Q _178_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_214 vgnd vpwr scs8hd_fill_1
XFILLER_0_151 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_62 vgnd vpwr scs8hd_decap_3
XFILLER_8_273 vpwr vgnd scs8hd_fill_2
XANTENNA__076__D _175_/D vgnd vpwr scs8hd_diode_2
XANTENNA__092__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_14_93 vgnd vpwr scs8hd_decap_8
XFILLER_5_276 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_3.LATCH_0_.latch data_in mem_top_ipin_3.LATCH_0_.latch/Q _129_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_4.INVTX1_0_.scs8hd_inv_1 chanx_left_in[2] mux_top_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_213 vgnd vpwr scs8hd_fill_1
XFILLER_18_125 vgnd vpwr scs8hd_decap_4
XPHY_70 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_81 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_top_ipin_5.LATCH_3_.latch data_in mem_top_ipin_5.LATCH_3_.latch/Q _143_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_198_ chanx_right_in[4] chanx_left_out[4] vgnd vpwr scs8hd_buf_2
Xmux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_2.LATCH_3_.latch/Q mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_96 vgnd vpwr scs8hd_decap_4
XFILLER_2_41 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_10_ vgnd vpwr scs8hd_inv_1
XFILLER_20_323 vgnd vpwr scs8hd_decap_12
XFILLER_17_191 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_5.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_top_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_4.LATCH_1_.latch_SLEEPB _136_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__098__B address[5] vgnd vpwr scs8hd_diode_2
X_121_ _110_/X _115_/X _121_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_301 vpwr vgnd scs8hd_fill_2
XFILLER_6_371 vpwr vgnd scs8hd_fill_2
XANTENNA__199__A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_16_39 vgnd vpwr scs8hd_decap_4
XFILLER_16_17 vgnd vpwr scs8hd_decap_12
XFILLER_4_308 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_104_ _179_/A _105_/A vgnd vpwr scs8hd_buf_1
XFILLER_7_102 vpwr vgnd scs8hd_fill_2
XFILLER_7_179 vpwr vgnd scs8hd_fill_2
XFILLER_11_164 vpwr vgnd scs8hd_fill_2
XFILLER_11_175 vpwr vgnd scs8hd_fill_2
XFILLER_3_363 vgnd vpwr scs8hd_fill_1
XFILLER_19_220 vgnd vpwr scs8hd_decap_12
XFILLER_8_51 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_3.LATCH_2_.latch/Q mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_366 vgnd vpwr scs8hd_fill_1
XFILLER_17_93 vgnd vpwr scs8hd_decap_6
XFILLER_17_60 vgnd vpwr scs8hd_fill_1
XFILLER_3_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_13_29 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _186_/HI mem_top_ipin_0.LATCH_5_.latch/Q
+ mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_13_259 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_ipin_2.LATCH_2_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_196 vgnd vpwr scs8hd_decap_4
XFILLER_8_241 vpwr vgnd scs8hd_fill_2
XFILLER_2_406 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_299 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_1_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_365 vgnd vpwr scs8hd_decap_8
XFILLER_14_354 vgnd vpwr scs8hd_decap_8
XPHY_60 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_71 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_82 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_14_398 vgnd vpwr scs8hd_decap_8
X_197_ chanx_right_in[5] chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_64 vgnd vpwr scs8hd_decap_4
XFILLER_2_20 vpwr vgnd scs8hd_fill_2
XFILLER_20_335 vgnd vpwr scs8hd_decap_6
XFILLER_9_380 vpwr vgnd scs8hd_fill_2
XFILLER_15_118 vpwr vgnd scs8hd_fill_2
XFILLER_15_107 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_2.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_120_ _108_/X _115_/X _120_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_339 vpwr vgnd scs8hd_fill_2
XFILLER_11_324 vgnd vpwr scs8hd_fill_1
XFILLER_11_346 vgnd vpwr scs8hd_decap_3
XFILLER_11_62 vgnd vpwr scs8hd_decap_3
XFILLER_14_140 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_3_.latch_SLEEPB _085_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_29 vpwr vgnd scs8hd_fill_2
XFILLER_20_187 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_3.INVTX1_4_.scs8hd_inv_1 chanx_left_in[6] mux_top_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_132 vpwr vgnd scs8hd_fill_2
X_103_ _150_/A _105_/B _103_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_114 vpwr vgnd scs8hd_fill_2
XFILLER_7_136 vpwr vgnd scs8hd_fill_2
XFILLER_11_143 vpwr vgnd scs8hd_fill_2
XFILLER_19_232 vgnd vpwr scs8hd_decap_12
XFILLER_8_85 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_8_96 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_0_356 vpwr vgnd scs8hd_fill_2
XFILLER_0_345 vpwr vgnd scs8hd_fill_2
XFILLER_16_202 vgnd vpwr scs8hd_decap_12
XFILLER_3_161 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_SLEEPB _182_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _165_/A mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_0_120 vpwr vgnd scs8hd_fill_2
XFILLER_12_293 vpwr vgnd scs8hd_fill_2
XFILLER_8_286 vpwr vgnd scs8hd_fill_2
XFILLER_5_53 vgnd vpwr scs8hd_fill_1
XFILLER_5_86 vpwr vgnd scs8hd_fill_2
XFILLER_14_84 vgnd vpwr scs8hd_decap_8
XFILLER_5_212 vpwr vgnd scs8hd_fill_2
XFILLER_5_256 vpwr vgnd scs8hd_fill_2
XFILLER_5_267 vgnd vpwr scs8hd_decap_3
XFILLER_5_289 vgnd vpwr scs8hd_decap_4
XFILLER_17_330 vgnd vpwr scs8hd_decap_12
XANTENNA__101__A _070_/X vgnd vpwr scs8hd_diode_2
XFILLER_19_18 vpwr vgnd scs8hd_fill_2
XFILLER_2_259 vpwr vgnd scs8hd_fill_2
XFILLER_2_226 vgnd vpwr scs8hd_decap_3
XFILLER_14_388 vgnd vpwr scs8hd_decap_8
XFILLER_14_377 vgnd vpwr scs8hd_decap_8
XPHY_61 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_ipin_7.LATCH_2_.latch_SLEEPB _160_/Y vgnd vpwr scs8hd_diode_2
XPHY_50 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_72 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_83 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_196_ chanx_right_in[6] chanx_left_out[6] vgnd vpwr scs8hd_buf_2
Xmux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_2.LATCH_2_.latch/Q mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_182 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_11_358 vpwr vgnd scs8hd_fill_2
XFILLER_2_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_SLEEPB _173_/Y vgnd vpwr scs8hd_diode_2
X_179_ _179_/A _178_/B _179_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_384 vpwr vgnd scs8hd_fill_2
XFILLER_10_380 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_1.LATCH_3_.latch data_in mem_top_ipin_1.LATCH_3_.latch/Q _105_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_199 vgnd vpwr scs8hd_decap_12
XFILLER_16_406 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_4.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_3_321 vpwr vgnd scs8hd_fill_2
X_102_ _178_/A _150_/A vgnd vpwr scs8hd_buf_1
XFILLER_11_199 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_0.INVTX1_0_.scs8hd_inv_1 chanx_left_in[2] mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_376 vpwr vgnd scs8hd_fill_2
XFILLER_8_64 vpwr vgnd scs8hd_fill_2
XFILLER_6_181 vpwr vgnd scs8hd_fill_2
XFILLER_4_107 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_335 vpwr vgnd scs8hd_fill_2
XFILLER_0_302 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_40 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_1.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_top_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__104__A _179_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_3.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_5.LATCH_3_.latch_SLEEPB _143_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_4.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_239 vgnd vpwr scs8hd_decap_4
XFILLER_13_217 vgnd vpwr scs8hd_decap_3
XFILLER_5_405 vpwr vgnd scs8hd_fill_2
XFILLER_0_176 vpwr vgnd scs8hd_fill_2
XFILLER_0_165 vpwr vgnd scs8hd_fill_2
XFILLER_8_276 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_7.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_top_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_52 vgnd vpwr scs8hd_decap_8
XFILLER_14_41 vgnd vpwr scs8hd_decap_8
XFILLER_17_342 vgnd vpwr scs8hd_decap_12
XANTENNA__101__B _105_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_205 vpwr vgnd scs8hd_fill_2
XANTENNA__202__A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XPHY_40 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_51 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_73 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_84 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_195_ chanx_right_in[7] chanx_left_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA__112__A _175_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_304 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_393 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_ipin_3.LATCH_4_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_315 vgnd vpwr scs8hd_decap_3
XFILLER_7_319 vgnd vpwr scs8hd_decap_4
XFILLER_11_53 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_4.LATCH_2_.latch data_in mem_top_ipin_4.LATCH_2_.latch/Q _135_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__107__A _106_/X vgnd vpwr scs8hd_diode_2
X_178_ _178_/A _178_/B _178_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_396 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_6.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_20_156 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_0.LATCH_3_.latch/Q mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_top_ipin_6.LATCH_5_.latch data_in mem_top_ipin_6.LATCH_5_.latch/Q _149_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_101_ _070_/X _105_/B _101_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_355 vpwr vgnd scs8hd_fill_2
XFILLER_3_388 vpwr vgnd scs8hd_fill_2
XFILLER_7_149 vgnd vpwr scs8hd_decap_4
XFILLER_19_245 vgnd vpwr scs8hd_decap_12
XFILLER_3_399 vpwr vgnd scs8hd_fill_2
XFILLER_8_32 vpwr vgnd scs8hd_fill_2
XFILLER_0_369 vgnd vpwr scs8hd_decap_3
XFILLER_0_325 vgnd vpwr scs8hd_decap_3
XANTENNA__210__A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_16_215 vgnd vpwr scs8hd_decap_12
XFILLER_3_141 vpwr vgnd scs8hd_fill_2
XFILLER_3_174 vpwr vgnd scs8hd_fill_2
XANTENNA__120__A _108_/X vgnd vpwr scs8hd_diode_2
XFILLER_12_6 vpwr vgnd scs8hd_fill_2
XFILLER_15_292 vpwr vgnd scs8hd_fill_2
XFILLER_15_281 vpwr vgnd scs8hd_fill_2
XFILLER_15_270 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_229 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__205__A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_1.LATCH_2_.latch/Q mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_ipin_1.LATCH_5_.latch_SLEEPB _101_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_200 vgnd vpwr scs8hd_decap_4
XFILLER_8_211 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__115__A _115_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_11 vgnd vpwr scs8hd_decap_4
XFILLER_8_222 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_99 vpwr vgnd scs8hd_fill_2
XFILLER_10_3 vpwr vgnd scs8hd_fill_2
XFILLER_5_225 vpwr vgnd scs8hd_fill_2
XFILLER_5_236 vpwr vgnd scs8hd_fill_2
XFILLER_17_354 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_5.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_top_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_129 vgnd vpwr scs8hd_fill_1
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_52 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_74 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_85 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_194_ chanx_right_in[8] chanx_left_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_1_272 vpwr vgnd scs8hd_fill_2
XANTENNA__112__B address[4] vgnd vpwr scs8hd_diode_2
XFILLER_17_195 vgnd vpwr scs8hd_decap_6
XFILLER_17_184 vgnd vpwr scs8hd_decap_4
XFILLER_17_140 vgnd vpwr scs8hd_fill_1
Xmem_top_ipin_7.LATCH_1_.latch data_in mem_top_ipin_7.LATCH_1_.latch/Q _161_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_1_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_338 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_6.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_top_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_76 vpwr vgnd scs8hd_fill_2
XFILLER_19_405 vpwr vgnd scs8hd_fill_2
XFILLER_14_154 vgnd vpwr scs8hd_decap_6
XFILLER_14_143 vpwr vgnd scs8hd_fill_2
XANTENNA__107__B _105_/B vgnd vpwr scs8hd_diode_2
X_177_ _177_/A _178_/B _177_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__123__A _122_/X vgnd vpwr scs8hd_diode_2
XFILLER_20_168 vgnd vpwr scs8hd_decap_12
XANTENNA__208__A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
X_100_ _099_/X _105_/B vgnd vpwr scs8hd_buf_1
XFILLER_7_106 vpwr vgnd scs8hd_fill_2
XFILLER_11_168 vpwr vgnd scs8hd_fill_2
XFILLER_11_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_334 vgnd vpwr scs8hd_decap_6
XFILLER_19_257 vgnd vpwr scs8hd_decap_12
XANTENNA__118__A _105_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_197 vpwr vgnd scs8hd_fill_2
XANTENNA__120__B _115_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_145 vgnd vpwr scs8hd_decap_4
XFILLER_0_134 vpwr vgnd scs8hd_fill_2
XFILLER_8_245 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_0_.latch/Q mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_34 vpwr vgnd scs8hd_fill_2
XFILLER_5_45 vpwr vgnd scs8hd_fill_2
XFILLER_5_56 vpwr vgnd scs8hd_fill_2
XFILLER_5_67 vpwr vgnd scs8hd_fill_2
XANTENNA__131__A _131_/A vgnd vpwr scs8hd_diode_2
XANTENNA__126__A _105_/A vgnd vpwr scs8hd_diode_2
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_64 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_53 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_42 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_20 vgnd vpwr scs8hd_decap_3
X_193_ _193_/HI _193_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mem_top_ipin_6.LATCH_5_.latch_SLEEPB _149_/Y vgnd vpwr scs8hd_diode_2
XPHY_75 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__112__C _073_/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_240 vpwr vgnd scs8hd_fill_2
XFILLER_2_68 vgnd vpwr scs8hd_fill_1
XFILLER_2_46 vgnd vpwr scs8hd_decap_3
XFILLER_2_24 vgnd vpwr scs8hd_decap_4
XFILLER_17_152 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_380 vgnd vpwr scs8hd_decap_4
XFILLER_9_362 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_0_.latch_SLEEPB _094_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_99 vpwr vgnd scs8hd_fill_2
XFILLER_14_111 vgnd vpwr scs8hd_decap_4
X_176_ _176_/A _178_/B vgnd vpwr scs8hd_buf_1
Xmux_top_ipin_3.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_top_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_398 vgnd vpwr scs8hd_decap_8
XFILLER_20_125 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_1.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_9_170 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_2_.latch/Q mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_11_103 vpwr vgnd scs8hd_fill_2
XFILLER_11_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_5.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_7_118 vpwr vgnd scs8hd_fill_2
XFILLER_11_136 vpwr vgnd scs8hd_fill_2
XFILLER_11_147 vgnd vpwr scs8hd_decap_4
XFILLER_0_3 vpwr vgnd scs8hd_fill_2
XFILLER_19_269 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_0.LATCH_2_.latch data_in mem_top_ipin_0.LATCH_2_.latch/Q _088_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_ipin_4.INVTX1_5_.scs8hd_inv_1 chanx_right_in[7] mux_top_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__118__B _115_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_23 vpwr vgnd scs8hd_fill_2
X_159_ _179_/A _156_/X _159_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_162 vpwr vgnd scs8hd_fill_2
XANTENNA__134__A _105_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_89 vgnd vpwr scs8hd_decap_3
XFILLER_0_349 vgnd vpwr scs8hd_decap_4
XFILLER_17_65 vpwr vgnd scs8hd_fill_2
XFILLER_17_54 vgnd vpwr scs8hd_decap_6
XFILLER_17_21 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_2.LATCH_5_.latch data_in mem_top_ipin_2.LATCH_5_.latch/Q _116_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_7.LATCH_0_.latch/Q mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__129__A _110_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_297 vpwr vgnd scs8hd_fill_2
XFILLER_12_231 vgnd vpwr scs8hd_decap_4
XFILLER_8_268 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_290 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_0.LATCH_2_.latch data_in mem_bottom_ipin_0.LATCH_2_.latch/Q _172_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_367 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_ipin_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__126__B _123_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _150_/A vgnd vpwr scs8hd_diode_2
XPHY_32 vgnd vpwr scs8hd_decap_3
XFILLER_14_337 vgnd vpwr scs8hd_decap_12
XFILLER_14_304 vgnd vpwr scs8hd_decap_12
XPHY_65 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_54 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_43 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_76 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
Xmem_bottom_ipin_2.LATCH_5_.latch data_in mem_bottom_ipin_2.LATCH_5_.latch/Q _177_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_192_ _192_/HI _192_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_285 vpwr vgnd scs8hd_fill_2
XFILLER_17_164 vgnd vpwr scs8hd_decap_12
XFILLER_2_58 vgnd vpwr scs8hd_decap_4
XFILLER_13_392 vpwr vgnd scs8hd_fill_2
XANTENNA__137__A _110_/X vgnd vpwr scs8hd_diode_2
XFILLER_11_12 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_3.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_11_34 vpwr vgnd scs8hd_fill_2
XFILLER_14_101 vgnd vpwr scs8hd_fill_1
X_175_ _175_/A _175_/B _175_/C _175_/D _176_/A vgnd vpwr scs8hd_or4_4
XFILLER_6_388 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_7.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_20_137 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_3.LATCH_1_.latch data_in mem_top_ipin_3.LATCH_1_.latch/Q _128_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ _166_/A mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_ipin_5.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_6.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_ipin_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_8_68 vpwr vgnd scs8hd_fill_2
X_089_ address[1] address[2] _068_/C _089_/X vgnd vpwr scs8hd_or3_4
X_158_ _178_/A _156_/X _158_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_141 vpwr vgnd scs8hd_fill_2
XFILLER_6_185 vgnd vpwr scs8hd_decap_3
XANTENNA__134__B _131_/X vgnd vpwr scs8hd_diode_2
XANTENNA__150__A _150_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_1.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_top_ipin_5.LATCH_4_.latch data_in mem_top_ipin_5.LATCH_4_.latch/Q _142_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_top_ipin_5.LATCH_0_.latch_SLEEPB _146_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_339 vpwr vgnd scs8hd_fill_2
XFILLER_0_306 vpwr vgnd scs8hd_fill_2
XFILLER_17_44 vpwr vgnd scs8hd_fill_2
XFILLER_8_406 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__129__B _123_/X vgnd vpwr scs8hd_diode_2
XANTENNA__145__A _108_/X vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.INVTX1_5_.scs8hd_inv_1 chanx_right_in[5] mux_top_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_103 vpwr vgnd scs8hd_fill_2
XFILLER_0_169 vpwr vgnd scs8hd_fill_2
XFILLER_0_114 vgnd vpwr scs8hd_decap_4
XFILLER_12_276 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_2_ vgnd vpwr scs8hd_inv_1
XFILLER_14_23 vpwr vgnd scs8hd_fill_2
XFILLER_14_12 vpwr vgnd scs8hd_fill_2
XFILLER_17_379 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_2.LATCH_4_.latch/Q mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_250 vpwr vgnd scs8hd_fill_2
XANTENNA__142__B _146_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_209 vpwr vgnd scs8hd_fill_2
XPHY_33 vgnd vpwr scs8hd_decap_3
XFILLER_14_349 vpwr vgnd scs8hd_fill_2
XFILLER_14_316 vgnd vpwr scs8hd_decap_12
XPHY_66 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_55 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_44 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_77 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_191_ _191_/HI _191_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mem_top_ipin_3.LATCH_1_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_297 vpwr vgnd scs8hd_fill_2
XFILLER_1_253 vpwr vgnd scs8hd_fill_2
XFILLER_17_176 vgnd vpwr scs8hd_decap_6
XFILLER_17_132 vgnd vpwr scs8hd_decap_8
XFILLER_17_121 vgnd vpwr scs8hd_fill_1
XANTENNA__137__B _131_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__153__A _108_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_SLEEPB _177_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_57 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_6.LATCH_0_.latch/Q mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_top_ipin_6.LATCH_0_.latch data_in mem_top_ipin_6.LATCH_0_.latch/Q _154_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_352 vgnd vpwr scs8hd_decap_4
X_174_ _174_/A _174_/B _174_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_312 vgnd vpwr scs8hd_decap_4
XFILLER_6_367 vpwr vgnd scs8hd_fill_2
XFILLER_10_363 vpwr vgnd scs8hd_fill_2
XFILLER_10_396 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__148__A _147_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_149 vgnd vpwr scs8hd_decap_6
XFILLER_3_359 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_157_ _177_/A _156_/X _157_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_8_36 vpwr vgnd scs8hd_fill_2
XFILLER_8_47 vpwr vgnd scs8hd_fill_2
XFILLER_10_182 vgnd vpwr scs8hd_decap_4
X_088_ _094_/A _106_/A _088_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__150__B _150_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_34 vgnd vpwr scs8hd_decap_6
XFILLER_3_123 vgnd vpwr scs8hd_decap_3
XFILLER_3_145 vgnd vpwr scs8hd_decap_3
XFILLER_3_178 vgnd vpwr scs8hd_decap_3
XFILLER_15_296 vgnd vpwr scs8hd_decap_8
XFILLER_15_285 vgnd vpwr scs8hd_decap_4
XFILLER_15_274 vpwr vgnd scs8hd_fill_2
X_209_ chanx_left_in[2] chanx_right_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA__145__B _146_/B vgnd vpwr scs8hd_diode_2
XANTENNA__161__A _108_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_1.LATCH_2_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_90 vgnd vpwr scs8hd_decap_6
XANTENNA__071__A enable vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_2_.latch/Q mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_255 vgnd vpwr scs8hd_decap_3
XFILLER_8_204 vgnd vpwr scs8hd_fill_1
XFILLER_10_7 vpwr vgnd scs8hd_fill_2
XANTENNA__156__A _155_/X vgnd vpwr scs8hd_diode_2
XANTENNA__066__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_5_229 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_0.INVTX1_5_.scs8hd_inv_1 chanx_right_in[7] mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_402 vgnd vpwr scs8hd_decap_4
XFILLER_4_240 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_0_.latch/Q mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_12 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XFILLER_14_328 vgnd vpwr scs8hd_decap_8
XPHY_45 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_56 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_67 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_78 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_190_ _190_/HI _190_/LO vgnd vpwr scs8hd_conb_1
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XFILLER_1_210 vgnd vpwr scs8hd_decap_4
XFILLER_2_16 vpwr vgnd scs8hd_fill_2
XFILLER_1_221 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_6.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_top_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__153__B _150_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_332 vgnd vpwr scs8hd_decap_4
XFILLER_9_343 vgnd vpwr scs8hd_decap_4
XFILLER_9_376 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_136 vgnd vpwr scs8hd_decap_4
XFILLER_14_125 vpwr vgnd scs8hd_fill_2
XFILLER_14_169 vgnd vpwr scs8hd_decap_12
XFILLER_14_147 vgnd vpwr scs8hd_decap_6
X_173_ _108_/A _174_/B _173_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_302 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_106 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_2.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__164__A _175_/D vgnd vpwr scs8hd_diode_2
XFILLER_9_140 vpwr vgnd scs8hd_fill_2
XFILLER_9_195 vpwr vgnd scs8hd_fill_2
XANTENNA__074__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_3_316 vgnd vpwr scs8hd_decap_3
X_087_ _086_/X _106_/A vgnd vpwr scs8hd_buf_1
X_156_ _155_/X _156_/X vgnd vpwr scs8hd_buf_1
XFILLER_6_154 vgnd vpwr scs8hd_fill_1
XFILLER_2_382 vgnd vpwr scs8hd_decap_12
XANTENNA__159__A _179_/A vgnd vpwr scs8hd_diode_2
XANTENNA__069__A _069_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _184_/HI _165_/Y mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_157 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_SLEEPB _164_/Y vgnd vpwr scs8hd_diode_2
X_208_ chanx_left_in[3] chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA__161__B _156_/X vgnd vpwr scs8hd_diode_2
X_139_ _099_/A address[4] _175_/C _147_/B _139_/X vgnd vpwr scs8hd_or4_4
XFILLER_0_138 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_1.LATCH_4_.latch data_in mem_top_ipin_1.LATCH_4_.latch/Q _103_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_267 vgnd vpwr scs8hd_decap_8
XFILLER_8_227 vgnd vpwr scs8hd_decap_3
XFILLER_5_49 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _186_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__172__A _106_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_5.LATCH_0_.latch/Q mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_69 vgnd vpwr scs8hd_decap_12
XANTENNA__082__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_5_208 vpwr vgnd scs8hd_fill_2
XFILLER_4_285 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_ipin_6.LATCH_2_.latch_SLEEPB _152_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__167__A _099_/A vgnd vpwr scs8hd_diode_2
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__077__A _077_/A vgnd vpwr scs8hd_diode_2
XPHY_13 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_68 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_79 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_3 vgnd vpwr scs8hd_decap_3
XFILLER_2_28 vgnd vpwr scs8hd_fill_1
XFILLER_13_340 vpwr vgnd scs8hd_fill_2
XFILLER_13_362 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _184_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
X_172_ _106_/A _174_/B _172_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_310 vgnd vpwr scs8hd_decap_8
XFILLER_10_376 vpwr vgnd scs8hd_fill_2
XFILLER_10_398 vgnd vpwr scs8hd_decap_8
XFILLER_20_118 vgnd vpwr scs8hd_decap_6
XFILLER_13_170 vpwr vgnd scs8hd_fill_2
XANTENNA__164__B _113_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_380 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__180__A _106_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_4.INVTX1_2_.scs8hd_inv_1 chanx_left_in[6] mux_top_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_93 vpwr vgnd scs8hd_fill_2
XANTENNA__074__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_11_118 vpwr vgnd scs8hd_fill_2
XFILLER_0_7 vpwr vgnd scs8hd_fill_2
XANTENNA__090__A _089_/X vgnd vpwr scs8hd_diode_2
XFILLER_3_306 vgnd vpwr scs8hd_fill_1
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
X_155_ _099_/A _175_/B _175_/C _147_/B _155_/X vgnd vpwr scs8hd_or4_4
XFILLER_6_177 vpwr vgnd scs8hd_fill_2
XFILLER_6_199 vpwr vgnd scs8hd_fill_2
X_086_ _086_/A address[2] address[0] _086_/X vgnd vpwr scs8hd_or3_4
XFILLER_2_372 vgnd vpwr scs8hd_fill_1
XFILLER_2_394 vgnd vpwr scs8hd_decap_3
XFILLER_18_251 vgnd vpwr scs8hd_decap_12
XANTENNA__159__B _156_/X vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_2.LATCH_0_.latch data_in mem_top_ipin_2.LATCH_0_.latch/Q _121_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__175__A _175_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_4.LATCH_3_.latch_SLEEPB _134_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_69 vgnd vpwr scs8hd_decap_12
XANTENNA__085__A _094_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_114 vpwr vgnd scs8hd_fill_2
XFILLER_15_232 vpwr vgnd scs8hd_fill_2
XFILLER_15_221 vgnd vpwr scs8hd_decap_4
X_207_ chanx_left_in[4] chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_15_265 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_138_ _098_/A address[5] _147_/B vgnd vpwr scs8hd_or2_4
Xmem_top_ipin_4.LATCH_3_.latch data_in mem_top_ipin_4.LATCH_3_.latch/Q _134_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_069_ _069_/A _177_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mem_top_ipin_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_50 vpwr vgnd scs8hd_fill_2
XFILLER_0_72 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_213 vgnd vpwr scs8hd_fill_1
XFILLER_5_28 vgnd vpwr scs8hd_decap_4
XANTENNA__172__B _174_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_294 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_2.LATCH_0_.latch data_in mem_bottom_ipin_2.LATCH_0_.latch/Q _182_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__167__B address[4] vgnd vpwr scs8hd_diode_2
XFILLER_6_82 vpwr vgnd scs8hd_fill_2
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_47 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_69 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_14 vgnd vpwr scs8hd_decap_3
XANTENNA__093__A _092_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_1_245 vgnd vpwr scs8hd_fill_1
XFILLER_17_113 vpwr vgnd scs8hd_fill_2
XFILLER_17_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_2.LATCH_4_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_6.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_289 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _166_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_301 vpwr vgnd scs8hd_fill_2
XFILLER_13_396 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_6.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_7.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__178__A _178_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_0.LATCH_4_.latch/Q mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_16 vpwr vgnd scs8hd_fill_2
XFILLER_11_38 vgnd vpwr scs8hd_decap_4
XANTENNA__088__A _094_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_171_ _179_/A _174_/B _171_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_348 vgnd vpwr scs8hd_decap_6
XFILLER_10_388 vgnd vpwr scs8hd_decap_8
XFILLER_13_193 vgnd vpwr scs8hd_decap_4
XANTENNA__164__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_9_153 vpwr vgnd scs8hd_fill_2
XFILLER_9_175 vpwr vgnd scs8hd_fill_2
XANTENNA__180__B _178_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_208 vgnd vpwr scs8hd_decap_12
XFILLER_6_145 vpwr vgnd scs8hd_fill_2
X_154_ _110_/X _150_/B _154_/Y vgnd vpwr scs8hd_nor2_4
X_085_ _094_/A _179_/A _085_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_12_81 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_4.LATCH_0_.latch/Q mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_263 vgnd vpwr scs8hd_decap_12
XANTENNA__175__B _175_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_48 vgnd vpwr scs8hd_decap_4
Xmem_top_ipin_7.LATCH_2_.latch data_in mem_top_ipin_7.LATCH_2_.latch/Q _160_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_406 vgnd vpwr scs8hd_fill_1
XANTENNA__085__B _179_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_top_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_206_ chanx_left_in[5] chanx_right_out[5] vgnd vpwr scs8hd_buf_2
X_137_ _110_/X _131_/X _137_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_192 vpwr vgnd scs8hd_fill_2
X_068_ address[1] _068_/B _068_/C _069_/A vgnd vpwr scs8hd_or3_4
XANTENNA_mem_top_ipin_0.LATCH_5_.latch_SLEEPB _078_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_3 vpwr vgnd scs8hd_fill_2
XFILLER_0_107 vpwr vgnd scs8hd_fill_2
XFILLER_12_203 vpwr vgnd scs8hd_fill_2
XANTENNA__096__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_20_280 vgnd vpwr scs8hd_decap_12
XFILLER_8_207 vpwr vgnd scs8hd_fill_2
XFILLER_18_91 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_8_ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _187_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_273 vpwr vgnd scs8hd_fill_2
XFILLER_11_280 vgnd vpwr scs8hd_decap_4
XFILLER_14_27 vgnd vpwr scs8hd_decap_4
XFILLER_14_16 vpwr vgnd scs8hd_fill_2
XFILLER_17_306 vgnd vpwr scs8hd_decap_12
XFILLER_4_210 vpwr vgnd scs8hd_fill_2
XFILLER_4_254 vpwr vgnd scs8hd_fill_2
XANTENNA__167__C _175_/C vgnd vpwr scs8hd_diode_2
XFILLER_16_372 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_2_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_59 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_48 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_15 vgnd vpwr scs8hd_decap_3
XFILLER_1_268 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_SLEEPB _180_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_92 vpwr vgnd scs8hd_fill_2
XFILLER_13_353 vpwr vgnd scs8hd_fill_2
XFILLER_13_320 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__178__B _178_/B vgnd vpwr scs8hd_diode_2
XFILLER_16_191 vgnd vpwr scs8hd_decap_8
XANTENNA__194__A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__088__B _106_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_117 vgnd vpwr scs8hd_decap_6
X_170_ _178_/A _174_/B _170_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_316 vgnd vpwr scs8hd_fill_1
XFILLER_9_132 vpwr vgnd scs8hd_fill_2
XFILLER_5_393 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_84 vgnd vpwr scs8hd_decap_3
XANTENNA__099__A _099_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_102 vgnd vpwr scs8hd_decap_4
XFILLER_6_124 vgnd vpwr scs8hd_decap_3
X_153_ _108_/X _150_/B _153_/Y vgnd vpwr scs8hd_nor2_4
X_084_ _083_/X _179_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mem_top_ipin_7.LATCH_4_.latch_SLEEPB _158_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_93 vgnd vpwr scs8hd_decap_4
XFILLER_19_7 vpwr vgnd scs8hd_fill_2
XANTENNA__175__C _175_/C vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_1_.latch/Q mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_245 vgnd vpwr scs8hd_decap_12
X_205_ chanx_left_in[6] chanx_right_out[6] vgnd vpwr scs8hd_buf_2
X_136_ _108_/X _131_/X _136_/Y vgnd vpwr scs8hd_nor2_4
X_067_ address[0] _068_/C vgnd vpwr scs8hd_inv_8
Xmux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_top_ipin_7.LATCH_3_.latch/Q mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_SLEEPB _171_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_30 vgnd vpwr scs8hd_fill_1
XFILLER_0_85 vpwr vgnd scs8hd_fill_2
XFILLER_12_215 vgnd vpwr scs8hd_decap_3
XFILLER_20_292 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.INVTX1_2_.scs8hd_inv_1 chanx_left_in[3] mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_119_ _106_/X _115_/X _119_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_19_381 vgnd vpwr scs8hd_decap_12
XANTENNA__197__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_0.LATCH_3_.latch data_in mem_top_ipin_0.LATCH_3_.latch/Q _085_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_406 vgnd vpwr scs8hd_fill_1
XFILLER_17_318 vgnd vpwr scs8hd_decap_12
XANTENNA__167__D _175_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_5.LATCH_5_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_51 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_16 vgnd vpwr scs8hd_decap_3
XFILLER_1_236 vpwr vgnd scs8hd_fill_2
XFILLER_1_214 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_3.LATCH_0_.latch/Q mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_126 vgnd vpwr scs8hd_decap_4
XFILLER_15_82 vpwr vgnd scs8hd_fill_2
XFILLER_15_71 vgnd vpwr scs8hd_decap_4
XFILLER_13_376 vpwr vgnd scs8hd_fill_2
XFILLER_13_332 vgnd vpwr scs8hd_fill_1
XFILLER_9_336 vgnd vpwr scs8hd_fill_1
XFILLER_9_358 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_0_280 vgnd vpwr scs8hd_decap_4
XFILLER_11_29 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_7.INVTX1_3_.scs8hd_inv_1 chanx_right_in[1] mux_top_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_5.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_3 vgnd vpwr scs8hd_decap_4
XFILLER_6_328 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_140 vpwr vgnd scs8hd_fill_2
XFILLER_9_199 vgnd vpwr scs8hd_decap_4
XFILLER_5_350 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_0.LATCH_3_.latch data_in mem_bottom_ipin_0.LATCH_3_.latch/Q _171_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__099__B address[4] vgnd vpwr scs8hd_diode_2
XFILLER_15_405 vpwr vgnd scs8hd_fill_2
X_083_ _086_/A address[2] _068_/C _083_/X vgnd vpwr scs8hd_or3_4
XFILLER_6_158 vpwr vgnd scs8hd_fill_2
X_152_ _106_/X _150_/B _152_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_165 vpwr vgnd scs8hd_fill_2
XFILLER_2_331 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_7.LATCH_1_.latch/Q mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_276 vgnd vpwr scs8hd_decap_12
XANTENNA__175__D _175_/D vgnd vpwr scs8hd_diode_2
XFILLER_5_191 vgnd vpwr scs8hd_decap_4
XFILLER_17_17 vpwr vgnd scs8hd_fill_2
XFILLER_3_128 vpwr vgnd scs8hd_fill_2
XFILLER_15_202 vpwr vgnd scs8hd_fill_2
XFILLER_15_257 vgnd vpwr scs8hd_decap_8
X_204_ chanx_left_in[7] chanx_right_out[7] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_066_ address[2] _068_/B vgnd vpwr scs8hd_inv_8
X_135_ _106_/X _131_/X _135_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_0_20 vpwr vgnd scs8hd_fill_2
XFILLER_9_73 vpwr vgnd scs8hd_fill_2
XFILLER_12_249 vgnd vpwr scs8hd_decap_4
XFILLER_12_238 vgnd vpwr scs8hd_decap_8
XFILLER_12_227 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_3.LATCH_2_.latch data_in mem_top_ipin_3.LATCH_2_.latch/Q _127_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_18_93 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _188_/HI vgnd vpwr
+ scs8hd_diode_2
X_118_ _105_/A _115_/X _118_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_19_393 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_5.LATCH_5_.latch data_in mem_top_ipin_5.LATCH_5_.latch/Q _141_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_94 vgnd vpwr scs8hd_decap_12
XFILLER_4_267 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_30 vgnd vpwr scs8hd_fill_1
XFILLER_6_63 vgnd vpwr scs8hd_decap_6
XPHY_28 vgnd vpwr scs8hd_decap_3
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_39 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_3.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_13_388 vpwr vgnd scs8hd_fill_2
XFILLER_9_315 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_7.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_8_370 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ _166_/Y mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_14_ vgnd vpwr scs8hd_inv_1
Xmux_top_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_6.LATCH_3_.latch/Q mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_13_174 vgnd vpwr scs8hd_decap_3
XFILLER_5_362 vpwr vgnd scs8hd_fill_2
XFILLER_3_42 vpwr vgnd scs8hd_fill_2
XFILLER_3_53 vgnd vpwr scs8hd_decap_3
XFILLER_3_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_3.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__099__C _175_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_4.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_5.INVTX1_3_.scs8hd_inv_1 chanx_right_in[7] mux_top_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_082_ address[1] _086_/A vgnd vpwr scs8hd_inv_8
X_151_ _105_/A _150_/B _151_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_122 vpwr vgnd scs8hd_fill_2
XFILLER_10_188 vpwr vgnd scs8hd_fill_2
XFILLER_2_365 vgnd vpwr scs8hd_decap_4
XFILLER_2_398 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_ipin_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_4.LATCH_0_.latch_SLEEPB _137_/Y vgnd vpwr scs8hd_diode_2
XFILLER_18_288 vgnd vpwr scs8hd_decap_12
XFILLER_17_29 vgnd vpwr scs8hd_decap_3
XFILLER_3_118 vpwr vgnd scs8hd_fill_2
XFILLER_15_236 vgnd vpwr scs8hd_decap_8
X_203_ chanx_left_in[8] chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_2_140 vpwr vgnd scs8hd_fill_2
X_134_ _105_/A _131_/X _134_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_184 vpwr vgnd scs8hd_fill_2
XFILLER_2_173 vpwr vgnd scs8hd_fill_2
XFILLER_0_32 vgnd vpwr scs8hd_decap_3
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_6.LATCH_1_.latch data_in mem_top_ipin_6.LATCH_1_.latch/Q _153_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_2.LATCH_0_.latch/Q mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_261 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _165_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _185_/HI mem_bottom_ipin_2.LATCH_5_.latch/Q
+ mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_117_ _150_/A _115_/X _117_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_221 vpwr vgnd scs8hd_fill_2
XFILLER_7_254 vpwr vgnd scs8hd_fill_2
XFILLER_11_261 vpwr vgnd scs8hd_fill_2
XFILLER_7_298 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_202 vpwr vgnd scs8hd_fill_2
XFILLER_4_224 vpwr vgnd scs8hd_fill_2
XFILLER_16_364 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_5.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_6_20 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_2.LATCH_1_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_86 vgnd vpwr scs8hd_decap_4
XFILLER_19_180 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XPHY_18 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_6.LATCH_1_.latch/Q mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_249 vpwr vgnd scs8hd_fill_2
XFILLER_9_8 vpwr vgnd scs8hd_fill_2
XFILLER_17_117 vpwr vgnd scs8hd_fill_2
XFILLER_17_106 vpwr vgnd scs8hd_fill_2
XFILLER_15_62 vpwr vgnd scs8hd_fill_2
XFILLER_13_367 vgnd vpwr scs8hd_decap_3
XANTENNA__102__A _178_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_161 vgnd vpwr scs8hd_decap_8
XFILLER_6_308 vpwr vgnd scs8hd_fill_2
XFILLER_10_348 vpwr vgnd scs8hd_fill_2
XFILLER_10_359 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_197 vgnd vpwr scs8hd_fill_1
XFILLER_13_153 vpwr vgnd scs8hd_fill_2
XFILLER_9_157 vpwr vgnd scs8hd_fill_2
XFILLER_5_330 vgnd vpwr scs8hd_decap_3
XFILLER_9_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_65 vpwr vgnd scs8hd_fill_2
XANTENNA__099__D _114_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_150_ _150_/A _150_/B _150_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_081_ _094_/A _178_/A _081_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_149 vpwr vgnd scs8hd_fill_2
XFILLER_12_41 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_182 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_ipin_0.LATCH_2_.latch_SLEEPB _088_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__200__A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
X_133_ _150_/A _131_/X _133_/Y vgnd vpwr scs8hd_nor2_4
X_202_ chanx_right_in[0] chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_2_152 vgnd vpwr scs8hd_fill_1
XFILLER_17_7 vgnd vpwr scs8hd_fill_1
XANTENNA__110__A _174_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_3.INVTX1_3_.scs8hd_inv_1 chanx_right_in[5] mux_top_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_66 vgnd vpwr scs8hd_decap_4
XFILLER_9_53 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_14_ vgnd vpwr scs8hd_inv_1
XFILLER_20_273 vgnd vpwr scs8hd_decap_6
XFILLER_12_207 vgnd vpwr scs8hd_decap_6
XFILLER_4_406 vgnd vpwr scs8hd_fill_1
XFILLER_18_51 vgnd vpwr scs8hd_fill_1
XANTENNA__105__A _105_/A vgnd vpwr scs8hd_diode_2
X_116_ _070_/X _115_/X _116_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_200 vpwr vgnd scs8hd_fill_2
XFILLER_7_277 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _189_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_1_.latch/Q mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_5.LATCH_3_.latch/Q mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_20_63 vgnd vpwr scs8hd_decap_12
XFILLER_16_398 vgnd vpwr scs8hd_decap_8
XFILLER_6_43 vpwr vgnd scs8hd_fill_2
XPHY_19 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_217 vpwr vgnd scs8hd_fill_2
XFILLER_15_96 vgnd vpwr scs8hd_decap_4
XFILLER_13_324 vgnd vpwr scs8hd_decap_8
XFILLER_13_313 vgnd vpwr scs8hd_decap_4
XFILLER_9_339 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_1.LATCH_5_.latch data_in mem_top_ipin_1.LATCH_5_.latch/Q _101_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__203__A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_13_132 vpwr vgnd scs8hd_fill_2
XFILLER_13_110 vpwr vgnd scs8hd_fill_2
XFILLER_9_114 vpwr vgnd scs8hd_fill_2
XFILLER_9_136 vpwr vgnd scs8hd_fill_2
XANTENNA__113__A _113_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_1.LATCH_0_.latch/Q mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_ipin_7.LATCH_1_.latch_SLEEPB _161_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_080_ _080_/A _178_/A vgnd vpwr scs8hd_buf_1
XFILLER_6_106 vgnd vpwr scs8hd_fill_1
XFILLER_10_135 vgnd vpwr scs8hd_decap_12
XFILLER_12_64 vpwr vgnd scs8hd_fill_2
XFILLER_12_75 vgnd vpwr scs8hd_decap_4
XFILLER_12_86 vgnd vpwr scs8hd_decap_6
XFILLER_18_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__108__A _108_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_150 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_SLEEPB _174_/Y vgnd vpwr scs8hd_diode_2
X_132_ _070_/X _131_/X _132_/Y vgnd vpwr scs8hd_nor2_4
X_201_ chanx_right_in[1] chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_14_293 vgnd vpwr scs8hd_decap_8
XFILLER_0_89 vpwr vgnd scs8hd_fill_2
XFILLER_9_43 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_5.LATCH_1_.latch/Q mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_98 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_230 vgnd vpwr scs8hd_decap_12
XANTENNA__211__A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_11_241 vgnd vpwr scs8hd_fill_1
X_115_ _115_/A _115_/X vgnd vpwr scs8hd_buf_1
XANTENNA__105__B _105_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_234 vpwr vgnd scs8hd_fill_2
XANTENNA__121__A _110_/X vgnd vpwr scs8hd_diode_2
XFILLER_19_330 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_ipin_1.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_top_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_top_ipin_2.LATCH_1_.latch data_in mem_top_ipin_2.LATCH_1_.latch/Q _120_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_top_ipin_5.LATCH_2_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__206__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_20_75 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_377 vgnd vpwr scs8hd_decap_12
XANTENNA__116__A _070_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_3_270 vpwr vgnd scs8hd_fill_2
XFILLER_20_3 vgnd vpwr scs8hd_decap_12
XFILLER_19_160 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_4.LATCH_4_.latch data_in mem_top_ipin_4.LATCH_4_.latch/Q _133_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_15_86 vgnd vpwr scs8hd_decap_3
XFILLER_15_53 vpwr vgnd scs8hd_fill_2
XFILLER_15_31 vgnd vpwr scs8hd_fill_1
XFILLER_13_358 vpwr vgnd scs8hd_fill_2
XFILLER_13_347 vgnd vpwr scs8hd_decap_4
XFILLER_13_336 vpwr vgnd scs8hd_fill_2
XFILLER_13_303 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_7.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_top_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_295 vgnd vpwr scs8hd_decap_4
XFILLER_0_262 vpwr vgnd scs8hd_fill_2
XFILLER_0_240 vpwr vgnd scs8hd_fill_2
XFILLER_16_174 vgnd vpwr scs8hd_decap_12
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_351 vgnd vpwr scs8hd_decap_4
.ends

