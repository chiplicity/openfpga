magic
tech EFS8A
magscale 1 2
timestamp 1602523605
<< locali >>
rect 11897 8993 12058 9027
rect 11897 8959 11931 8993
rect 12817 8585 12909 8619
rect 16083 8585 16221 8619
rect 12817 8483 12851 8585
rect 1547 8041 1685 8075
rect 11161 7939 11195 7973
rect 7239 7905 7274 7939
rect 11161 7905 11322 7939
rect 13863 7905 13898 7939
rect 16715 7905 16750 7939
rect 24535 7905 24662 7939
rect 4445 7191 4479 7497
rect 4991 6953 4997 6987
rect 6699 6953 6837 6987
rect 4991 6885 5025 6953
rect 6503 6817 6630 6851
rect 34655 6817 34690 6851
rect 24035 6103 24069 6171
rect 24035 6069 24041 6103
rect 17595 5865 17601 5899
rect 17595 5797 17629 5865
rect 9689 5627 9723 5729
rect 9321 5083 9355 5185
rect 13823 4777 13829 4811
rect 24771 4777 24777 4811
rect 8861 4539 8895 4777
rect 13823 4709 13857 4777
rect 24771 4709 24805 4777
rect 27307 4233 27445 4267
rect 15393 4131 15427 4233
rect 7199 3927 7233 3995
rect 24035 3927 24069 3995
rect 7199 3893 7205 3927
rect 24035 3893 24041 3927
rect 6739 3689 6745 3723
rect 6739 3621 6773 3689
rect 7297 2839 7331 3077
rect 12449 2975 12483 3145
rect 4169 2295 4203 2601
rect 19901 2499 19935 2601
rect 4537 2363 4571 2465
<< viali >>
rect 1593 12937 1627 12971
rect 23857 12937 23891 12971
rect 26433 12937 26467 12971
rect 35633 12937 35667 12971
rect 1409 12733 1443 12767
rect 23673 12733 23707 12767
rect 26249 12733 26283 12767
rect 35449 12733 35483 12767
rect 36001 12733 36035 12767
rect 1961 12597 1995 12631
rect 24317 12597 24351 12631
rect 26801 12597 26835 12631
rect 19349 12257 19383 12291
rect 19533 12053 19567 12087
rect 7021 11849 7055 11883
rect 19441 11849 19475 11883
rect 6837 11645 6871 11679
rect 7389 11509 7423 11543
rect 35633 11305 35667 11339
rect 35449 11169 35483 11203
rect 35449 10625 35483 10659
rect 35633 9129 35667 9163
rect 35449 8993 35483 9027
rect 11897 8925 11931 8959
rect 12127 8789 12161 8823
rect 11161 8585 11195 8619
rect 12909 8585 12943 8619
rect 16221 8585 16255 8619
rect 18613 8585 18647 8619
rect 10517 8517 10551 8551
rect 18199 8517 18233 8551
rect 12817 8449 12851 8483
rect 10333 8381 10367 8415
rect 10793 8381 10827 8415
rect 11380 8381 11414 8415
rect 12495 8381 12529 8415
rect 12587 8381 12621 8415
rect 16012 8381 16046 8415
rect 16405 8381 16439 8415
rect 18128 8381 18162 8415
rect 1685 8245 1719 8279
rect 11483 8245 11517 8279
rect 12081 8245 12115 8279
rect 35449 8245 35483 8279
rect 1685 8041 1719 8075
rect 16819 8041 16853 8075
rect 24041 8041 24075 8075
rect 32321 8041 32355 8075
rect 4721 7973 4755 8007
rect 11161 7973 11195 8007
rect 12173 7973 12207 8007
rect 12357 7973 12391 8007
rect 12449 7973 12483 8007
rect 1476 7905 1510 7939
rect 1869 7905 1903 7939
rect 7205 7905 7239 7939
rect 8585 7905 8619 7939
rect 9689 7905 9723 7939
rect 13829 7905 13863 7939
rect 16681 7905 16715 7939
rect 24501 7905 24535 7939
rect 32137 7905 32171 7939
rect 2789 7837 2823 7871
rect 4629 7837 4663 7871
rect 4905 7837 4939 7871
rect 7757 7837 7791 7871
rect 12817 7837 12851 7871
rect 15301 7837 15335 7871
rect 5641 7769 5675 7803
rect 8769 7769 8803 7803
rect 24731 7769 24765 7803
rect 25421 7769 25455 7803
rect 2513 7701 2547 7735
rect 3249 7701 3283 7735
rect 7343 7701 7377 7735
rect 8125 7701 8159 7735
rect 9873 7701 9907 7735
rect 11391 7701 11425 7735
rect 13277 7701 13311 7735
rect 13967 7701 14001 7735
rect 25053 7701 25087 7735
rect 2789 7497 2823 7531
rect 4445 7497 4479 7531
rect 8585 7497 8619 7531
rect 10701 7497 10735 7531
rect 12265 7497 12299 7531
rect 13461 7497 13495 7531
rect 24685 7497 24719 7531
rect 4261 7429 4295 7463
rect 3065 7361 3099 7395
rect 3341 7361 3375 7395
rect 1409 7293 1443 7327
rect 1961 7293 1995 7327
rect 2513 7225 2547 7259
rect 3157 7225 3191 7259
rect 11805 7429 11839 7463
rect 5549 7361 5583 7395
rect 7665 7361 7699 7395
rect 10885 7361 10919 7395
rect 12541 7361 12575 7395
rect 12817 7361 12851 7395
rect 25053 7361 25087 7395
rect 9848 7293 9882 7327
rect 10333 7293 10367 7327
rect 13921 7293 13955 7327
rect 14080 7293 14114 7327
rect 15612 7293 15646 7327
rect 16037 7293 16071 7327
rect 17024 7293 17058 7327
rect 17877 7293 17911 7327
rect 18153 7293 18187 7327
rect 24016 7293 24050 7327
rect 5273 7225 5307 7259
rect 5365 7225 5399 7259
rect 7757 7225 7791 7259
rect 8309 7225 8343 7259
rect 10977 7225 11011 7259
rect 11529 7225 11563 7259
rect 12633 7225 12667 7259
rect 18061 7225 18095 7259
rect 25145 7225 25179 7259
rect 25697 7225 25731 7259
rect 1593 7157 1627 7191
rect 4445 7157 4479 7191
rect 4629 7157 4663 7191
rect 5089 7157 5123 7191
rect 7297 7157 7331 7191
rect 9597 7157 9631 7191
rect 9919 7157 9953 7191
rect 14151 7157 14185 7191
rect 14565 7157 14599 7191
rect 15715 7157 15749 7191
rect 16681 7157 16715 7191
rect 17095 7157 17129 7191
rect 17509 7157 17543 7191
rect 24087 7157 24121 7191
rect 32229 7157 32263 7191
rect 3801 6953 3835 6987
rect 4997 6953 5031 6987
rect 5549 6953 5583 6987
rect 6837 6953 6871 6987
rect 10885 6953 10919 6987
rect 12173 6953 12207 6987
rect 16497 6953 16531 6987
rect 7481 6885 7515 6919
rect 7757 6885 7791 6919
rect 8309 6885 8343 6919
rect 11574 6885 11608 6919
rect 12541 6885 12575 6919
rect 13185 6885 13219 6919
rect 15393 6885 15427 6919
rect 15485 6885 15519 6919
rect 16037 6885 16071 6919
rect 17601 6885 17635 6919
rect 24961 6885 24995 6919
rect 25053 6885 25087 6919
rect 26709 6885 26743 6919
rect 2605 6817 2639 6851
rect 6469 6817 6503 6851
rect 9781 6817 9815 6851
rect 20913 6817 20947 6851
rect 21373 6817 21407 6851
rect 21925 6817 21959 6851
rect 22109 6817 22143 6851
rect 23800 6817 23834 6851
rect 34621 6817 34655 6851
rect 1593 6749 1627 6783
rect 4629 6749 4663 6783
rect 7665 6749 7699 6783
rect 8585 6749 8619 6783
rect 11253 6749 11287 6783
rect 13093 6749 13127 6783
rect 17509 6749 17543 6783
rect 18981 6749 19015 6783
rect 22385 6749 22419 6783
rect 24225 6749 24259 6783
rect 25605 6749 25639 6783
rect 26617 6749 26651 6783
rect 26893 6749 26927 6783
rect 2789 6681 2823 6715
rect 10241 6681 10275 6715
rect 13645 6681 13679 6715
rect 18061 6681 18095 6715
rect 2329 6613 2363 6647
rect 3065 6613 3099 6647
rect 3525 6613 3559 6647
rect 4353 6613 4387 6647
rect 7113 6613 7147 6647
rect 9965 6613 9999 6647
rect 12817 6613 12851 6647
rect 14381 6613 14415 6647
rect 18429 6613 18463 6647
rect 20177 6613 20211 6647
rect 20637 6613 20671 6647
rect 23903 6613 23937 6647
rect 34759 6613 34793 6647
rect 2053 6409 2087 6443
rect 5457 6409 5491 6443
rect 8125 6409 8159 6443
rect 13369 6409 13403 6443
rect 13645 6409 13679 6443
rect 15393 6409 15427 6443
rect 17509 6409 17543 6443
rect 17877 6409 17911 6443
rect 24593 6409 24627 6443
rect 24961 6409 24995 6443
rect 26617 6409 26651 6443
rect 32045 6409 32079 6443
rect 36093 6409 36127 6443
rect 3617 6341 3651 6375
rect 6653 6341 6687 6375
rect 27629 6341 27663 6375
rect 35633 6341 35667 6375
rect 14381 6273 14415 6307
rect 15025 6273 15059 6307
rect 16497 6273 16531 6307
rect 16865 6273 16899 6307
rect 18153 6273 18187 6307
rect 18521 6273 18555 6307
rect 22293 6273 22327 6307
rect 23673 6273 23707 6307
rect 25513 6273 25547 6307
rect 25789 6273 25823 6307
rect 27077 6273 27111 6307
rect 2513 6205 2547 6239
rect 2697 6205 2731 6239
rect 3065 6205 3099 6239
rect 3433 6205 3467 6239
rect 4537 6205 4571 6239
rect 5733 6205 5767 6239
rect 7205 6205 7239 6239
rect 8769 6205 8803 6239
rect 9873 6205 9907 6239
rect 10149 6205 10183 6239
rect 10425 6205 10459 6239
rect 10793 6205 10827 6239
rect 12449 6205 12483 6239
rect 19993 6205 20027 6239
rect 20177 6205 20211 6239
rect 20637 6205 20671 6239
rect 21189 6205 21223 6239
rect 21373 6205 21407 6239
rect 22661 6205 22695 6239
rect 31560 6205 31594 6239
rect 34713 6205 34747 6239
rect 35449 6205 35483 6239
rect 1777 6137 1811 6171
rect 4445 6137 4479 6171
rect 4899 6137 4933 6171
rect 7526 6137 7560 6171
rect 9505 6137 9539 6171
rect 12173 6137 12207 6171
rect 12770 6137 12804 6171
rect 14473 6137 14507 6171
rect 16313 6137 16347 6171
rect 16589 6137 16623 6171
rect 18245 6137 18279 6171
rect 21649 6137 21683 6171
rect 25329 6137 25363 6171
rect 25605 6137 25639 6171
rect 27169 6137 27203 6171
rect 27997 6137 28031 6171
rect 3985 6069 4019 6103
rect 6101 6069 6135 6103
rect 7021 6069 7055 6103
rect 9045 6069 9079 6103
rect 10977 6069 11011 6103
rect 11345 6069 11379 6103
rect 11713 6069 11747 6103
rect 14197 6069 14231 6103
rect 15669 6069 15703 6103
rect 19717 6069 19751 6103
rect 21925 6069 21959 6103
rect 23029 6069 23063 6103
rect 23397 6069 23431 6103
rect 24041 6069 24075 6103
rect 31631 6069 31665 6103
rect 3157 5865 3191 5899
rect 3525 5865 3559 5899
rect 6745 5865 6779 5899
rect 7205 5865 7239 5899
rect 9137 5865 9171 5899
rect 12265 5865 12299 5899
rect 14381 5865 14415 5899
rect 17601 5865 17635 5899
rect 18153 5865 18187 5899
rect 18429 5865 18463 5899
rect 19993 5865 20027 5899
rect 20637 5865 20671 5899
rect 24133 5865 24167 5899
rect 24777 5865 24811 5899
rect 25099 5865 25133 5899
rect 26341 5865 26375 5899
rect 27629 5865 27663 5899
rect 2599 5797 2633 5831
rect 5549 5797 5583 5831
rect 11529 5797 11563 5831
rect 13782 5797 13816 5831
rect 15117 5797 15151 5831
rect 15761 5797 15795 5831
rect 15853 5797 15887 5831
rect 16405 5797 16439 5831
rect 23534 5797 23568 5831
rect 26709 5797 26743 5831
rect 2237 5729 2271 5763
rect 4261 5729 4295 5763
rect 4537 5729 4571 5763
rect 5089 5729 5123 5763
rect 5273 5729 5307 5763
rect 7205 5729 7239 5763
rect 7389 5729 7423 5763
rect 7941 5729 7975 5763
rect 8125 5729 8159 5763
rect 9413 5729 9447 5763
rect 9689 5729 9723 5763
rect 10333 5729 10367 5763
rect 10609 5729 10643 5763
rect 10885 5729 10919 5763
rect 11253 5729 11287 5763
rect 12392 5729 12426 5763
rect 16773 5729 16807 5763
rect 19809 5729 19843 5763
rect 20913 5729 20947 5763
rect 21373 5729 21407 5763
rect 21925 5729 21959 5763
rect 22109 5729 22143 5763
rect 25028 5729 25062 5763
rect 1777 5661 1811 5695
rect 2053 5661 2087 5695
rect 13461 5661 13495 5695
rect 17233 5661 17267 5695
rect 22385 5661 22419 5695
rect 23213 5661 23247 5695
rect 25421 5661 25455 5695
rect 26617 5661 26651 5695
rect 26893 5661 26927 5695
rect 9689 5593 9723 5627
rect 12495 5593 12529 5627
rect 13185 5593 13219 5627
rect 3893 5525 3927 5559
rect 5825 5525 5859 5559
rect 6469 5525 6503 5559
rect 9965 5525 9999 5559
rect 11897 5525 11931 5559
rect 12817 5525 12851 5559
rect 14657 5525 14691 5559
rect 15485 5525 15519 5559
rect 17141 5525 17175 5559
rect 20269 5525 20303 5559
rect 1593 5321 1627 5355
rect 6193 5321 6227 5355
rect 6561 5321 6595 5355
rect 7113 5321 7147 5355
rect 12265 5321 12299 5355
rect 13645 5321 13679 5355
rect 14197 5321 14231 5355
rect 15209 5321 15243 5355
rect 17417 5321 17451 5355
rect 22201 5321 22235 5355
rect 23213 5321 23247 5355
rect 24041 5321 24075 5355
rect 25145 5321 25179 5355
rect 27353 5321 27387 5355
rect 11345 5253 11379 5287
rect 19901 5253 19935 5287
rect 21833 5253 21867 5287
rect 26985 5253 27019 5287
rect 4077 5185 4111 5219
rect 9321 5185 9355 5219
rect 9413 5185 9447 5219
rect 11069 5185 11103 5219
rect 12725 5185 12759 5219
rect 13185 5185 13219 5219
rect 15761 5185 15795 5219
rect 18061 5185 18095 5219
rect 24225 5185 24259 5219
rect 26065 5185 26099 5219
rect 1409 5117 1443 5151
rect 2881 5117 2915 5151
rect 3065 5117 3099 5151
rect 3433 5117 3467 5151
rect 3801 5117 3835 5151
rect 5089 5117 5123 5151
rect 5641 5117 5675 5151
rect 7481 5117 7515 5151
rect 7665 5117 7699 5151
rect 8769 5117 8803 5151
rect 9873 5117 9907 5151
rect 10057 5117 10091 5151
rect 10425 5117 10459 5151
rect 10793 5117 10827 5151
rect 11713 5117 11747 5151
rect 14289 5117 14323 5151
rect 16221 5117 16255 5151
rect 17141 5117 17175 5151
rect 17877 5117 17911 5151
rect 18153 5117 18187 5151
rect 20085 5117 20119 5151
rect 20637 5117 20671 5151
rect 20913 5117 20947 5151
rect 21465 5117 21499 5151
rect 22569 5117 22603 5151
rect 5917 5049 5951 5083
rect 8309 5049 8343 5083
rect 9321 5049 9355 5083
rect 12817 5049 12851 5083
rect 14610 5049 14644 5083
rect 16037 5049 16071 5083
rect 16542 5049 16576 5083
rect 19165 5049 19199 5083
rect 21557 5049 21591 5083
rect 24546 5049 24580 5083
rect 26157 5049 26191 5083
rect 26709 5049 26743 5083
rect 2053 4981 2087 5015
rect 2421 4981 2455 5015
rect 4353 4981 4387 5015
rect 9045 4981 9079 5015
rect 19533 4981 19567 5015
rect 25513 4981 25547 5015
rect 25789 4981 25823 5015
rect 1685 4777 1719 4811
rect 3433 4777 3467 4811
rect 7205 4777 7239 4811
rect 8861 4777 8895 4811
rect 12265 4777 12299 4811
rect 13277 4777 13311 4811
rect 13829 4777 13863 4811
rect 14381 4777 14415 4811
rect 17049 4777 17083 4811
rect 22661 4777 22695 4811
rect 23213 4777 23247 4811
rect 24225 4777 24259 4811
rect 24777 4777 24811 4811
rect 25329 4777 25363 4811
rect 26065 4777 26099 4811
rect 1961 4641 1995 4675
rect 2973 4641 3007 4675
rect 4629 4641 4663 4675
rect 5089 4641 5123 4675
rect 5641 4641 5675 4675
rect 5825 4641 5859 4675
rect 7481 4641 7515 4675
rect 6101 4573 6135 4607
rect 6377 4573 6411 4607
rect 7849 4573 7883 4607
rect 9045 4709 9079 4743
rect 9413 4709 9447 4743
rect 11161 4709 11195 4743
rect 14657 4709 14691 4743
rect 15393 4709 15427 4743
rect 15485 4709 15519 4743
rect 16037 4709 16071 4743
rect 20085 4709 20119 4743
rect 25605 4709 25639 4743
rect 26709 4709 26743 4743
rect 9965 4641 9999 4675
rect 10149 4641 10183 4675
rect 10701 4641 10735 4675
rect 10885 4641 10919 4675
rect 11989 4641 12023 4675
rect 12173 4641 12207 4675
rect 12817 4641 12851 4675
rect 15025 4641 15059 4675
rect 16497 4641 16531 4675
rect 17233 4641 17267 4675
rect 17417 4641 17451 4675
rect 17785 4641 17819 4675
rect 18153 4641 18187 4675
rect 19324 4641 19358 4675
rect 20545 4641 20579 4675
rect 20913 4641 20947 4675
rect 21373 4641 21407 4675
rect 21925 4641 21959 4675
rect 22109 4641 22143 4675
rect 13461 4573 13495 4607
rect 22385 4573 22419 4607
rect 24409 4573 24443 4607
rect 26617 4573 26651 4607
rect 26893 4573 26927 4607
rect 2697 4505 2731 4539
rect 3157 4505 3191 4539
rect 4261 4505 4295 4539
rect 7941 4505 7975 4539
rect 8861 4505 8895 4539
rect 11529 4505 11563 4539
rect 11805 4505 11839 4539
rect 19717 4505 19751 4539
rect 3801 4437 3835 4471
rect 6837 4437 6871 4471
rect 7619 4437 7653 4471
rect 7757 4437 7791 4471
rect 8769 4437 8803 4471
rect 16773 4437 16807 4471
rect 18705 4437 18739 4471
rect 19165 4437 19199 4471
rect 19395 4437 19429 4471
rect 23673 4437 23707 4471
rect 1869 4233 1903 4267
rect 2605 4233 2639 4267
rect 3709 4233 3743 4267
rect 6653 4233 6687 4267
rect 8861 4233 8895 4267
rect 10793 4233 10827 4267
rect 11529 4233 11563 4267
rect 15393 4233 15427 4267
rect 15485 4233 15519 4267
rect 22569 4233 22603 4267
rect 23489 4233 23523 4267
rect 26341 4233 26375 4267
rect 26709 4233 26743 4267
rect 27445 4233 27479 4267
rect 14105 4165 14139 4199
rect 14473 4165 14507 4199
rect 19901 4165 19935 4199
rect 24869 4165 24903 4199
rect 25237 4165 25271 4199
rect 26985 4165 27019 4199
rect 35081 4165 35115 4199
rect 3065 4097 3099 4131
rect 6009 4097 6043 4131
rect 10517 4097 10551 4131
rect 12817 4097 12851 4131
rect 13185 4097 13219 4131
rect 13829 4097 13863 4131
rect 15393 4097 15427 4131
rect 17141 4097 17175 4131
rect 21925 4097 21959 4131
rect 23673 4097 23707 4131
rect 25421 4097 25455 4131
rect 31401 4097 31435 4131
rect 31677 4097 31711 4131
rect 35541 4097 35575 4131
rect 1685 4029 1719 4063
rect 4261 4029 4295 4063
rect 4813 4029 4847 4063
rect 5089 4029 5123 4063
rect 5641 4029 5675 4063
rect 5733 4029 5767 4063
rect 6837 4029 6871 4063
rect 9045 4029 9079 4063
rect 9781 4029 9815 4063
rect 10057 4029 10091 4063
rect 10241 4029 10275 4063
rect 11345 4029 11379 4063
rect 11805 4029 11839 4063
rect 12173 4029 12207 4063
rect 14289 4029 14323 4063
rect 15945 4029 15979 4063
rect 16129 4029 16163 4063
rect 16497 4029 16531 4063
rect 16865 4029 16899 4063
rect 17417 4029 17451 4063
rect 18245 4029 18279 4063
rect 18521 4029 18555 4063
rect 18889 4029 18923 4063
rect 19257 4029 19291 4063
rect 20729 4029 20763 4063
rect 20913 4029 20947 4063
rect 21465 4029 21499 4063
rect 21649 4029 21683 4063
rect 27236 4029 27270 4063
rect 34897 4029 34931 4063
rect 2789 3961 2823 3995
rect 2881 3961 2915 3995
rect 8493 3961 8527 3995
rect 12909 3961 12943 3995
rect 22201 3961 22235 3995
rect 25742 3961 25776 3995
rect 27721 3961 27755 3995
rect 31493 3961 31527 3995
rect 2145 3893 2179 3927
rect 4077 3893 4111 3927
rect 7205 3893 7239 3927
rect 7757 3893 7791 3927
rect 8125 3893 8159 3927
rect 11253 3893 11287 3927
rect 14933 3893 14967 3927
rect 17785 3893 17819 3927
rect 18153 3893 18187 3927
rect 20361 3893 20395 3927
rect 24041 3893 24075 3927
rect 24593 3893 24627 3927
rect 31217 3893 31251 3927
rect 1961 3689 1995 3723
rect 6745 3689 6779 3723
rect 7665 3689 7699 3723
rect 9413 3689 9447 3723
rect 11069 3689 11103 3723
rect 15025 3689 15059 3723
rect 15485 3689 15519 3723
rect 20177 3689 20211 3723
rect 21741 3689 21775 3723
rect 24685 3689 24719 3723
rect 31401 3689 31435 3723
rect 2237 3621 2271 3655
rect 2605 3621 2639 3655
rect 5825 3621 5859 3655
rect 8033 3621 8067 3655
rect 8677 3621 8711 3655
rect 13737 3621 13771 3655
rect 14289 3621 14323 3655
rect 16313 3621 16347 3655
rect 17141 3621 17175 3655
rect 19717 3621 19751 3655
rect 21373 3621 21407 3655
rect 23851 3621 23885 3655
rect 32321 3621 32355 3655
rect 1476 3553 1510 3587
rect 4077 3553 4111 3587
rect 4813 3553 4847 3587
rect 5089 3553 5123 3587
rect 5457 3553 5491 3587
rect 6377 3553 6411 3587
rect 8125 3553 8159 3587
rect 8309 3553 8343 3587
rect 9137 3553 9171 3587
rect 9781 3553 9815 3587
rect 10425 3553 10459 3587
rect 11529 3553 11563 3587
rect 11897 3553 11931 3587
rect 12081 3553 12115 3587
rect 12449 3553 12483 3587
rect 15301 3553 15335 3587
rect 15853 3553 15887 3587
rect 17049 3553 17083 3587
rect 17877 3553 17911 3587
rect 18245 3553 18279 3587
rect 18429 3553 18463 3587
rect 18797 3553 18831 3587
rect 19165 3553 19199 3587
rect 20980 3553 21014 3587
rect 23489 3553 23523 3587
rect 2513 3485 2547 3519
rect 2789 3485 2823 3519
rect 13001 3485 13035 3519
rect 13645 3485 13679 3519
rect 14657 3485 14691 3519
rect 20453 3485 20487 3519
rect 25237 3485 25271 3519
rect 32229 3485 32263 3519
rect 32505 3485 32539 3519
rect 5457 3417 5491 3451
rect 7297 3417 7331 3451
rect 12633 3417 12667 3451
rect 13369 3417 13403 3451
rect 19349 3417 19383 3451
rect 1547 3349 1581 3383
rect 3433 3349 3467 3383
rect 3893 3349 3927 3383
rect 6193 3349 6227 3383
rect 10793 3349 10827 3383
rect 17417 3349 17451 3383
rect 21051 3349 21085 3383
rect 24409 3349 24443 3383
rect 4353 3145 4387 3179
rect 6101 3145 6135 3179
rect 6469 3145 6503 3179
rect 10241 3145 10275 3179
rect 12265 3145 12299 3179
rect 12449 3145 12483 3179
rect 13645 3145 13679 3179
rect 15301 3145 15335 3179
rect 15669 3145 15703 3179
rect 17417 3145 17451 3179
rect 20177 3145 20211 3179
rect 24225 3145 24259 3179
rect 27077 3145 27111 3179
rect 30849 3145 30883 3179
rect 31309 3145 31343 3179
rect 32735 3145 32769 3179
rect 4721 3077 4755 3111
rect 7297 3077 7331 3111
rect 7803 3077 7837 3111
rect 7941 3077 7975 3111
rect 2145 3009 2179 3043
rect 3065 3009 3099 3043
rect 4813 3009 4847 3043
rect 1501 2941 1535 2975
rect 5733 2941 5767 2975
rect 2973 2873 3007 2907
rect 3427 2873 3461 2907
rect 5175 2873 5209 2907
rect 8033 3009 8067 3043
rect 8677 3009 8711 3043
rect 9321 3009 9355 3043
rect 9965 3009 9999 3043
rect 11161 3009 11195 3043
rect 13185 3077 13219 3111
rect 14749 3077 14783 3111
rect 16313 3077 16347 3111
rect 23949 3077 23983 3111
rect 33149 3077 33183 3111
rect 16497 3009 16531 3043
rect 24961 3009 24995 3043
rect 25145 3009 25179 3043
rect 11897 2941 11931 2975
rect 12449 2941 12483 2975
rect 17877 2941 17911 2975
rect 18337 2941 18371 2975
rect 18521 2941 18555 2975
rect 18889 2941 18923 2975
rect 19257 2941 19291 2975
rect 20453 2941 20487 2975
rect 21960 2941 21994 2975
rect 22385 2941 22419 2975
rect 25789 2941 25823 2975
rect 26684 2941 26718 2975
rect 31125 2941 31159 2975
rect 32137 2941 32171 2975
rect 32664 2941 32698 2975
rect 7665 2873 7699 2907
rect 8401 2873 8435 2907
rect 9045 2873 9079 2907
rect 9413 2873 9447 2907
rect 10885 2873 10919 2907
rect 10977 2873 11011 2907
rect 12633 2873 12667 2907
rect 12725 2873 12759 2907
rect 14197 2873 14231 2907
rect 14289 2873 14323 2907
rect 16589 2873 16623 2907
rect 17141 2873 17175 2907
rect 20361 2873 20395 2907
rect 21741 2873 21775 2907
rect 25237 2873 25271 2907
rect 2421 2805 2455 2839
rect 3985 2805 4019 2839
rect 7205 2805 7239 2839
rect 7297 2805 7331 2839
rect 7481 2805 7515 2839
rect 10701 2805 10735 2839
rect 14013 2805 14047 2839
rect 18153 2805 18187 2839
rect 19809 2805 19843 2839
rect 21465 2805 21499 2839
rect 22063 2805 22097 2839
rect 26755 2805 26789 2839
rect 1593 2601 1627 2635
rect 3893 2601 3927 2635
rect 4169 2601 4203 2635
rect 4445 2601 4479 2635
rect 7113 2601 7147 2635
rect 9965 2601 9999 2635
rect 12449 2601 12483 2635
rect 14197 2601 14231 2635
rect 16313 2601 16347 2635
rect 17417 2601 17451 2635
rect 19901 2601 19935 2635
rect 25145 2601 25179 2635
rect 32229 2601 32263 2635
rect 33241 2601 33275 2635
rect 2421 2533 2455 2567
rect 1409 2465 1443 2499
rect 1869 2465 1903 2499
rect 2237 2465 2271 2499
rect 3065 2465 3099 2499
rect 3525 2329 3559 2363
rect 6377 2533 6411 2567
rect 10609 2533 10643 2567
rect 11155 2533 11189 2567
rect 11989 2533 12023 2567
rect 13001 2533 13035 2567
rect 13369 2533 13403 2567
rect 13921 2533 13955 2567
rect 14933 2533 14967 2567
rect 16818 2533 16852 2567
rect 17693 2533 17727 2567
rect 18153 2533 18187 2567
rect 18521 2533 18555 2567
rect 20637 2533 20671 2567
rect 4261 2465 4295 2499
rect 4537 2465 4571 2499
rect 5181 2465 5215 2499
rect 5365 2465 5399 2499
rect 6745 2465 6779 2499
rect 6929 2465 6963 2499
rect 7481 2465 7515 2499
rect 7941 2465 7975 2499
rect 8088 2465 8122 2499
rect 9781 2465 9815 2499
rect 10241 2465 10275 2499
rect 11713 2465 11747 2499
rect 15552 2465 15586 2499
rect 15945 2465 15979 2499
rect 16497 2465 16531 2499
rect 19073 2465 19107 2499
rect 19901 2465 19935 2499
rect 19993 2465 20027 2499
rect 21189 2465 21223 2499
rect 21281 2465 21315 2499
rect 22201 2465 22235 2499
rect 29745 2465 29779 2499
rect 30297 2465 30331 2499
rect 32597 2465 32631 2499
rect 6009 2397 6043 2431
rect 8309 2397 8343 2431
rect 8677 2397 8711 2431
rect 10793 2397 10827 2431
rect 13277 2397 13311 2431
rect 15301 2397 15335 2431
rect 18429 2397 18463 2431
rect 20913 2397 20947 2431
rect 22753 2397 22787 2431
rect 4537 2329 4571 2363
rect 4813 2329 4847 2363
rect 8217 2329 8251 2363
rect 8953 2329 8987 2363
rect 9321 2329 9355 2363
rect 15623 2329 15657 2363
rect 19349 2329 19383 2363
rect 20177 2329 20211 2363
rect 29929 2329 29963 2363
rect 32781 2329 32815 2363
rect 4169 2261 4203 2295
rect 7849 2261 7883 2295
rect 19717 2261 19751 2295
<< metal1 >>
rect 5626 15512 5632 15564
rect 5684 15552 5690 15564
rect 6638 15552 6644 15564
rect 5684 15524 6644 15552
rect 5684 15512 5690 15524
rect 6638 15512 6644 15524
rect 6696 15512 6702 15564
rect 11054 15512 11060 15564
rect 11112 15552 11118 15564
rect 16482 15552 16488 15564
rect 11112 15524 16488 15552
rect 11112 15512 11118 15524
rect 16482 15512 16488 15524
rect 16540 15512 16546 15564
rect 1104 13626 38824 13648
rect 1104 13574 14315 13626
rect 14367 13574 14379 13626
rect 14431 13574 14443 13626
rect 14495 13574 14507 13626
rect 14559 13574 27648 13626
rect 27700 13574 27712 13626
rect 27764 13574 27776 13626
rect 27828 13574 27840 13626
rect 27892 13574 38824 13626
rect 1104 13552 38824 13574
rect 1104 13082 38824 13104
rect 1104 13030 7648 13082
rect 7700 13030 7712 13082
rect 7764 13030 7776 13082
rect 7828 13030 7840 13082
rect 7892 13030 20982 13082
rect 21034 13030 21046 13082
rect 21098 13030 21110 13082
rect 21162 13030 21174 13082
rect 21226 13030 34315 13082
rect 34367 13030 34379 13082
rect 34431 13030 34443 13082
rect 34495 13030 34507 13082
rect 34559 13030 38824 13082
rect 1104 13008 38824 13030
rect 1578 12968 1584 12980
rect 1539 12940 1584 12968
rect 1578 12928 1584 12940
rect 1636 12928 1642 12980
rect 23845 12971 23903 12977
rect 23845 12937 23857 12971
rect 23891 12968 23903 12971
rect 24118 12968 24124 12980
rect 23891 12940 24124 12968
rect 23891 12937 23903 12940
rect 23845 12931 23903 12937
rect 24118 12928 24124 12940
rect 24176 12928 24182 12980
rect 26421 12971 26479 12977
rect 26421 12937 26433 12971
rect 26467 12968 26479 12971
rect 28534 12968 28540 12980
rect 26467 12940 28540 12968
rect 26467 12937 26479 12940
rect 26421 12931 26479 12937
rect 28534 12928 28540 12940
rect 28592 12928 28598 12980
rect 35618 12968 35624 12980
rect 35579 12940 35624 12968
rect 35618 12928 35624 12940
rect 35676 12928 35682 12980
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12764 1455 12767
rect 23661 12767 23719 12773
rect 1443 12736 1900 12764
rect 1443 12733 1455 12736
rect 1397 12727 1455 12733
rect 1872 12640 1900 12736
rect 23661 12733 23673 12767
rect 23707 12764 23719 12767
rect 24302 12764 24308 12776
rect 23707 12736 24308 12764
rect 23707 12733 23719 12736
rect 23661 12727 23719 12733
rect 24302 12724 24308 12736
rect 24360 12724 24366 12776
rect 26237 12767 26295 12773
rect 26237 12733 26249 12767
rect 26283 12764 26295 12767
rect 26786 12764 26792 12776
rect 26283 12736 26792 12764
rect 26283 12733 26295 12736
rect 26237 12727 26295 12733
rect 26786 12724 26792 12736
rect 26844 12724 26850 12776
rect 35250 12724 35256 12776
rect 35308 12764 35314 12776
rect 35437 12767 35495 12773
rect 35437 12764 35449 12767
rect 35308 12736 35449 12764
rect 35308 12724 35314 12736
rect 35437 12733 35449 12736
rect 35483 12764 35495 12767
rect 35989 12767 36047 12773
rect 35989 12764 36001 12767
rect 35483 12736 36001 12764
rect 35483 12733 35495 12736
rect 35437 12727 35495 12733
rect 35989 12733 36001 12736
rect 36035 12733 36047 12767
rect 35989 12727 36047 12733
rect 16206 12656 16212 12708
rect 16264 12696 16270 12708
rect 39574 12696 39580 12708
rect 16264 12668 39580 12696
rect 16264 12656 16270 12668
rect 39574 12656 39580 12668
rect 39632 12656 39638 12708
rect 1854 12588 1860 12640
rect 1912 12628 1918 12640
rect 1949 12631 2007 12637
rect 1949 12628 1961 12631
rect 1912 12600 1961 12628
rect 1912 12588 1918 12600
rect 1949 12597 1961 12600
rect 1995 12597 2007 12631
rect 24302 12628 24308 12640
rect 24263 12600 24308 12628
rect 1949 12591 2007 12597
rect 24302 12588 24308 12600
rect 24360 12588 24366 12640
rect 26786 12628 26792 12640
rect 26747 12600 26792 12628
rect 26786 12588 26792 12600
rect 26844 12588 26850 12640
rect 1104 12538 38824 12560
rect 1104 12486 14315 12538
rect 14367 12486 14379 12538
rect 14431 12486 14443 12538
rect 14495 12486 14507 12538
rect 14559 12486 27648 12538
rect 27700 12486 27712 12538
rect 27764 12486 27776 12538
rect 27828 12486 27840 12538
rect 27892 12486 38824 12538
rect 1104 12464 38824 12486
rect 19337 12291 19395 12297
rect 19337 12257 19349 12291
rect 19383 12288 19395 12291
rect 19702 12288 19708 12300
rect 19383 12260 19708 12288
rect 19383 12257 19395 12260
rect 19337 12251 19395 12257
rect 19702 12248 19708 12260
rect 19760 12248 19766 12300
rect 19521 12087 19579 12093
rect 19521 12053 19533 12087
rect 19567 12084 19579 12087
rect 39574 12084 39580 12096
rect 19567 12056 39580 12084
rect 19567 12053 19579 12056
rect 19521 12047 19579 12053
rect 39574 12044 39580 12056
rect 39632 12044 39638 12096
rect 1104 11994 38824 12016
rect 1104 11942 7648 11994
rect 7700 11942 7712 11994
rect 7764 11942 7776 11994
rect 7828 11942 7840 11994
rect 7892 11942 20982 11994
rect 21034 11942 21046 11994
rect 21098 11942 21110 11994
rect 21162 11942 21174 11994
rect 21226 11942 34315 11994
rect 34367 11942 34379 11994
rect 34431 11942 34443 11994
rect 34495 11942 34507 11994
rect 34559 11942 38824 11994
rect 1104 11920 38824 11942
rect 7006 11880 7012 11892
rect 6967 11852 7012 11880
rect 7006 11840 7012 11852
rect 7064 11840 7070 11892
rect 19429 11883 19487 11889
rect 19429 11849 19441 11883
rect 19475 11880 19487 11883
rect 19702 11880 19708 11892
rect 19475 11852 19708 11880
rect 19475 11849 19487 11852
rect 19429 11843 19487 11849
rect 19702 11840 19708 11852
rect 19760 11840 19766 11892
rect 6825 11679 6883 11685
rect 6825 11645 6837 11679
rect 6871 11676 6883 11679
rect 6871 11648 7420 11676
rect 6871 11645 6883 11648
rect 6825 11639 6883 11645
rect 7392 11552 7420 11648
rect 7374 11540 7380 11552
rect 7335 11512 7380 11540
rect 7374 11500 7380 11512
rect 7432 11500 7438 11552
rect 1104 11450 38824 11472
rect 1104 11398 14315 11450
rect 14367 11398 14379 11450
rect 14431 11398 14443 11450
rect 14495 11398 14507 11450
rect 14559 11398 27648 11450
rect 27700 11398 27712 11450
rect 27764 11398 27776 11450
rect 27828 11398 27840 11450
rect 27892 11398 38824 11450
rect 1104 11376 38824 11398
rect 35621 11339 35679 11345
rect 35621 11305 35633 11339
rect 35667 11336 35679 11339
rect 39574 11336 39580 11348
rect 35667 11308 39580 11336
rect 35667 11305 35679 11308
rect 35621 11299 35679 11305
rect 39574 11296 39580 11308
rect 39632 11296 39638 11348
rect 35434 11200 35440 11212
rect 35395 11172 35440 11200
rect 35434 11160 35440 11172
rect 35492 11160 35498 11212
rect 1104 10906 38824 10928
rect 1104 10854 7648 10906
rect 7700 10854 7712 10906
rect 7764 10854 7776 10906
rect 7828 10854 7840 10906
rect 7892 10854 20982 10906
rect 21034 10854 21046 10906
rect 21098 10854 21110 10906
rect 21162 10854 21174 10906
rect 21226 10854 34315 10906
rect 34367 10854 34379 10906
rect 34431 10854 34443 10906
rect 34495 10854 34507 10906
rect 34559 10854 38824 10906
rect 1104 10832 38824 10854
rect 35434 10656 35440 10668
rect 35395 10628 35440 10656
rect 35434 10616 35440 10628
rect 35492 10616 35498 10668
rect 1104 10362 38824 10384
rect 1104 10310 14315 10362
rect 14367 10310 14379 10362
rect 14431 10310 14443 10362
rect 14495 10310 14507 10362
rect 14559 10310 27648 10362
rect 27700 10310 27712 10362
rect 27764 10310 27776 10362
rect 27828 10310 27840 10362
rect 27892 10310 38824 10362
rect 1104 10288 38824 10310
rect 1104 9818 38824 9840
rect 1104 9766 7648 9818
rect 7700 9766 7712 9818
rect 7764 9766 7776 9818
rect 7828 9766 7840 9818
rect 7892 9766 20982 9818
rect 21034 9766 21046 9818
rect 21098 9766 21110 9818
rect 21162 9766 21174 9818
rect 21226 9766 34315 9818
rect 34367 9766 34379 9818
rect 34431 9766 34443 9818
rect 34495 9766 34507 9818
rect 34559 9766 38824 9818
rect 1104 9744 38824 9766
rect 1104 9274 38824 9296
rect 1104 9222 14315 9274
rect 14367 9222 14379 9274
rect 14431 9222 14443 9274
rect 14495 9222 14507 9274
rect 14559 9222 27648 9274
rect 27700 9222 27712 9274
rect 27764 9222 27776 9274
rect 27828 9222 27840 9274
rect 27892 9222 38824 9274
rect 1104 9200 38824 9222
rect 35618 9160 35624 9172
rect 35579 9132 35624 9160
rect 35618 9120 35624 9132
rect 35676 9120 35682 9172
rect 35434 9024 35440 9036
rect 35395 8996 35440 9024
rect 35434 8984 35440 8996
rect 35492 8984 35498 9036
rect 11885 8959 11943 8965
rect 11885 8925 11897 8959
rect 11931 8956 11943 8959
rect 12066 8956 12072 8968
rect 11931 8928 12072 8956
rect 11931 8925 11943 8928
rect 11885 8919 11943 8925
rect 12066 8916 12072 8928
rect 12124 8916 12130 8968
rect 12115 8823 12173 8829
rect 12115 8789 12127 8823
rect 12161 8820 12173 8823
rect 13446 8820 13452 8832
rect 12161 8792 13452 8820
rect 12161 8789 12173 8792
rect 12115 8783 12173 8789
rect 13446 8780 13452 8792
rect 13504 8780 13510 8832
rect 1104 8730 38824 8752
rect 1104 8678 7648 8730
rect 7700 8678 7712 8730
rect 7764 8678 7776 8730
rect 7828 8678 7840 8730
rect 7892 8678 20982 8730
rect 21034 8678 21046 8730
rect 21098 8678 21110 8730
rect 21162 8678 21174 8730
rect 21226 8678 34315 8730
rect 34367 8678 34379 8730
rect 34431 8678 34443 8730
rect 34495 8678 34507 8730
rect 34559 8678 38824 8730
rect 1104 8656 38824 8678
rect 11146 8616 11152 8628
rect 11107 8588 11152 8616
rect 11146 8576 11152 8588
rect 11204 8576 11210 8628
rect 12894 8616 12900 8628
rect 12855 8588 12900 8616
rect 12894 8576 12900 8588
rect 12952 8576 12958 8628
rect 16206 8616 16212 8628
rect 16167 8588 16212 8616
rect 16206 8576 16212 8588
rect 16264 8576 16270 8628
rect 18601 8619 18659 8625
rect 18601 8585 18613 8619
rect 18647 8616 18659 8619
rect 19702 8616 19708 8628
rect 18647 8588 19708 8616
rect 18647 8585 18659 8588
rect 18601 8579 18659 8585
rect 10505 8551 10563 8557
rect 10505 8517 10517 8551
rect 10551 8548 10563 8551
rect 12250 8548 12256 8560
rect 10551 8520 12256 8548
rect 10551 8517 10563 8520
rect 10505 8511 10563 8517
rect 12250 8508 12256 8520
rect 12308 8508 12314 8560
rect 12342 8508 12348 8560
rect 12400 8548 12406 8560
rect 18187 8551 18245 8557
rect 18187 8548 18199 8551
rect 12400 8520 18199 8548
rect 12400 8508 12406 8520
rect 18187 8517 18199 8520
rect 18233 8517 18245 8551
rect 18187 8511 18245 8517
rect 12805 8483 12863 8489
rect 12805 8480 12817 8483
rect 12498 8452 12817 8480
rect 9858 8372 9864 8424
rect 9916 8412 9922 8424
rect 10321 8415 10379 8421
rect 10321 8412 10333 8415
rect 9916 8384 10333 8412
rect 9916 8372 9922 8384
rect 10321 8381 10333 8384
rect 10367 8412 10379 8415
rect 10781 8415 10839 8421
rect 10781 8412 10793 8415
rect 10367 8384 10793 8412
rect 10367 8381 10379 8384
rect 10321 8375 10379 8381
rect 10781 8381 10793 8384
rect 10827 8381 10839 8415
rect 10781 8375 10839 8381
rect 11146 8372 11152 8424
rect 11204 8412 11210 8424
rect 12498 8421 12526 8452
rect 12805 8449 12817 8452
rect 12851 8449 12863 8483
rect 12805 8443 12863 8449
rect 11368 8415 11426 8421
rect 11368 8412 11380 8415
rect 11204 8384 11380 8412
rect 11204 8372 11210 8384
rect 11368 8381 11380 8384
rect 11414 8381 11426 8415
rect 11368 8375 11426 8381
rect 12483 8415 12541 8421
rect 12483 8381 12495 8415
rect 12529 8381 12541 8415
rect 12483 8375 12541 8381
rect 12575 8415 12633 8421
rect 12575 8381 12587 8415
rect 12621 8412 12633 8415
rect 12894 8412 12900 8424
rect 12621 8384 12900 8412
rect 12621 8381 12633 8384
rect 12575 8375 12633 8381
rect 11394 8344 11422 8375
rect 12894 8372 12900 8384
rect 12952 8372 12958 8424
rect 16022 8421 16028 8424
rect 16000 8415 16028 8421
rect 16000 8412 16012 8415
rect 15935 8384 16012 8412
rect 16000 8381 16012 8384
rect 16080 8412 16086 8424
rect 16393 8415 16451 8421
rect 16393 8412 16405 8415
rect 16080 8384 16405 8412
rect 16000 8375 16028 8381
rect 16022 8372 16028 8375
rect 16080 8372 16086 8384
rect 16393 8381 16405 8384
rect 16439 8381 16451 8415
rect 16393 8375 16451 8381
rect 18116 8415 18174 8421
rect 18116 8381 18128 8415
rect 18162 8412 18174 8415
rect 18616 8412 18644 8579
rect 19702 8576 19708 8588
rect 19760 8576 19766 8628
rect 18162 8384 18644 8412
rect 18162 8381 18174 8384
rect 18116 8375 18174 8381
rect 15286 8344 15292 8356
rect 11394 8316 15292 8344
rect 15286 8304 15292 8316
rect 15344 8304 15350 8356
rect 1673 8279 1731 8285
rect 1673 8245 1685 8279
rect 1719 8276 1731 8279
rect 2682 8276 2688 8288
rect 1719 8248 2688 8276
rect 1719 8245 1731 8248
rect 1673 8239 1731 8245
rect 2682 8236 2688 8248
rect 2740 8236 2746 8288
rect 11471 8279 11529 8285
rect 11471 8245 11483 8279
rect 11517 8276 11529 8279
rect 11882 8276 11888 8288
rect 11517 8248 11888 8276
rect 11517 8245 11529 8248
rect 11471 8239 11529 8245
rect 11882 8236 11888 8248
rect 11940 8236 11946 8288
rect 12066 8276 12072 8288
rect 11979 8248 12072 8276
rect 12066 8236 12072 8248
rect 12124 8276 12130 8288
rect 12526 8276 12532 8288
rect 12124 8248 12532 8276
rect 12124 8236 12130 8248
rect 12526 8236 12532 8248
rect 12584 8236 12590 8288
rect 35434 8276 35440 8288
rect 35395 8248 35440 8276
rect 35434 8236 35440 8248
rect 35492 8236 35498 8288
rect 1104 8186 38824 8208
rect 1104 8134 14315 8186
rect 14367 8134 14379 8186
rect 14431 8134 14443 8186
rect 14495 8134 14507 8186
rect 14559 8134 27648 8186
rect 27700 8134 27712 8186
rect 27764 8134 27776 8186
rect 27828 8134 27840 8186
rect 27892 8134 38824 8186
rect 1104 8112 38824 8134
rect 1486 8032 1492 8084
rect 1544 8072 1550 8084
rect 1673 8075 1731 8081
rect 1673 8072 1685 8075
rect 1544 8044 1685 8072
rect 1544 8032 1550 8044
rect 1673 8041 1685 8044
rect 1719 8041 1731 8075
rect 1673 8035 1731 8041
rect 16482 8032 16488 8084
rect 16540 8072 16546 8084
rect 16807 8075 16865 8081
rect 16807 8072 16819 8075
rect 16540 8044 16819 8072
rect 16540 8032 16546 8044
rect 16807 8041 16819 8044
rect 16853 8041 16865 8075
rect 16807 8035 16865 8041
rect 24029 8075 24087 8081
rect 24029 8041 24041 8075
rect 24075 8072 24087 8075
rect 24302 8072 24308 8084
rect 24075 8044 24308 8072
rect 24075 8041 24087 8044
rect 24029 8035 24087 8041
rect 24302 8032 24308 8044
rect 24360 8032 24366 8084
rect 32309 8075 32367 8081
rect 32309 8041 32321 8075
rect 32355 8072 32367 8075
rect 33134 8072 33140 8084
rect 32355 8044 33140 8072
rect 32355 8041 32367 8044
rect 32309 8035 32367 8041
rect 33134 8032 33140 8044
rect 33192 8032 33198 8084
rect 4614 7964 4620 8016
rect 4672 8004 4678 8016
rect 4709 8007 4767 8013
rect 4709 8004 4721 8007
rect 4672 7976 4721 8004
rect 4672 7964 4678 7976
rect 4709 7973 4721 7976
rect 4755 7973 4767 8007
rect 4709 7967 4767 7973
rect 5626 7964 5632 8016
rect 5684 8004 5690 8016
rect 5684 7976 8616 8004
rect 5684 7964 5690 7976
rect 8588 7948 8616 7976
rect 11054 7964 11060 8016
rect 11112 8004 11118 8016
rect 11149 8007 11207 8013
rect 11149 8004 11161 8007
rect 11112 7976 11161 8004
rect 11112 7964 11118 7976
rect 11149 7973 11161 7976
rect 11195 7973 11207 8007
rect 11149 7967 11207 7973
rect 12161 8007 12219 8013
rect 12161 7973 12173 8007
rect 12207 8004 12219 8007
rect 12342 8004 12348 8016
rect 12207 7976 12348 8004
rect 12207 7973 12219 7976
rect 12161 7967 12219 7973
rect 12342 7964 12348 7976
rect 12400 7964 12406 8016
rect 12434 7964 12440 8016
rect 12492 8004 12498 8016
rect 12492 7976 12537 8004
rect 12492 7964 12498 7976
rect 1464 7939 1522 7945
rect 1464 7905 1476 7939
rect 1510 7936 1522 7939
rect 1857 7939 1915 7945
rect 1857 7936 1869 7939
rect 1510 7908 1869 7936
rect 1510 7905 1522 7908
rect 1464 7899 1522 7905
rect 1857 7905 1869 7908
rect 1903 7936 1915 7939
rect 3326 7936 3332 7948
rect 1903 7908 3332 7936
rect 1903 7905 1915 7908
rect 1857 7899 1915 7905
rect 3326 7896 3332 7908
rect 3384 7896 3390 7948
rect 7193 7939 7251 7945
rect 7193 7905 7205 7939
rect 7239 7936 7251 7939
rect 7282 7936 7288 7948
rect 7239 7908 7288 7936
rect 7239 7905 7251 7908
rect 7193 7899 7251 7905
rect 7282 7896 7288 7908
rect 7340 7896 7346 7948
rect 8570 7936 8576 7948
rect 8483 7908 8576 7936
rect 8570 7896 8576 7908
rect 8628 7896 8634 7948
rect 9582 7896 9588 7948
rect 9640 7936 9646 7948
rect 9677 7939 9735 7945
rect 9677 7936 9689 7939
rect 9640 7908 9689 7936
rect 9640 7896 9646 7908
rect 9677 7905 9689 7908
rect 9723 7905 9735 7939
rect 9677 7899 9735 7905
rect 13817 7939 13875 7945
rect 13817 7905 13829 7939
rect 13863 7936 13875 7939
rect 13906 7936 13912 7948
rect 13863 7908 13912 7936
rect 13863 7905 13875 7908
rect 13817 7899 13875 7905
rect 13906 7896 13912 7908
rect 13964 7896 13970 7948
rect 16666 7936 16672 7948
rect 16627 7908 16672 7936
rect 16666 7896 16672 7908
rect 16724 7896 16730 7948
rect 24489 7939 24547 7945
rect 24489 7905 24501 7939
rect 24535 7936 24547 7939
rect 24670 7936 24676 7948
rect 24535 7908 24676 7936
rect 24535 7905 24547 7908
rect 24489 7899 24547 7905
rect 24670 7896 24676 7908
rect 24728 7896 24734 7948
rect 32125 7939 32183 7945
rect 32125 7905 32137 7939
rect 32171 7936 32183 7939
rect 32214 7936 32220 7948
rect 32171 7908 32220 7936
rect 32171 7905 32183 7908
rect 32125 7899 32183 7905
rect 32214 7896 32220 7908
rect 32272 7896 32278 7948
rect 2774 7868 2780 7880
rect 2735 7840 2780 7868
rect 2774 7828 2780 7840
rect 2832 7828 2838 7880
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7868 4675 7871
rect 4706 7868 4712 7880
rect 4663 7840 4712 7868
rect 4663 7837 4675 7840
rect 4617 7831 4675 7837
rect 4706 7828 4712 7840
rect 4764 7828 4770 7880
rect 4890 7868 4896 7880
rect 4851 7840 4896 7868
rect 4890 7828 4896 7840
rect 4948 7828 4954 7880
rect 7745 7871 7803 7877
rect 7745 7837 7757 7871
rect 7791 7868 7803 7871
rect 8018 7868 8024 7880
rect 7791 7840 8024 7868
rect 7791 7837 7803 7840
rect 7745 7831 7803 7837
rect 8018 7828 8024 7840
rect 8076 7828 8082 7880
rect 12802 7868 12808 7880
rect 12763 7840 12808 7868
rect 12802 7828 12808 7840
rect 12860 7828 12866 7880
rect 15289 7871 15347 7877
rect 15289 7837 15301 7871
rect 15335 7868 15347 7871
rect 15378 7868 15384 7880
rect 15335 7840 15384 7868
rect 15335 7837 15347 7840
rect 15289 7831 15347 7837
rect 15378 7828 15384 7840
rect 15436 7828 15442 7880
rect 5258 7760 5264 7812
rect 5316 7800 5322 7812
rect 5629 7803 5687 7809
rect 5629 7800 5641 7803
rect 5316 7772 5641 7800
rect 5316 7760 5322 7772
rect 5629 7769 5641 7772
rect 5675 7800 5687 7803
rect 8294 7800 8300 7812
rect 5675 7772 8300 7800
rect 5675 7769 5687 7772
rect 5629 7763 5687 7769
rect 8294 7760 8300 7772
rect 8352 7760 8358 7812
rect 8757 7803 8815 7809
rect 8757 7769 8769 7803
rect 8803 7800 8815 7803
rect 11698 7800 11704 7812
rect 8803 7772 11704 7800
rect 8803 7769 8815 7772
rect 8757 7763 8815 7769
rect 11698 7760 11704 7772
rect 11756 7760 11762 7812
rect 24719 7803 24777 7809
rect 24719 7769 24731 7803
rect 24765 7800 24777 7803
rect 25130 7800 25136 7812
rect 24765 7772 25136 7800
rect 24765 7769 24777 7772
rect 24719 7763 24777 7769
rect 25130 7760 25136 7772
rect 25188 7800 25194 7812
rect 25409 7803 25467 7809
rect 25409 7800 25421 7803
rect 25188 7772 25421 7800
rect 25188 7760 25194 7772
rect 25409 7769 25421 7772
rect 25455 7769 25467 7803
rect 25409 7763 25467 7769
rect 2498 7732 2504 7744
rect 2459 7704 2504 7732
rect 2498 7692 2504 7704
rect 2556 7692 2562 7744
rect 2958 7692 2964 7744
rect 3016 7732 3022 7744
rect 3237 7735 3295 7741
rect 3237 7732 3249 7735
rect 3016 7704 3249 7732
rect 3016 7692 3022 7704
rect 3237 7701 3249 7704
rect 3283 7701 3295 7735
rect 3237 7695 3295 7701
rect 7331 7735 7389 7741
rect 7331 7701 7343 7735
rect 7377 7732 7389 7735
rect 7466 7732 7472 7744
rect 7377 7704 7472 7732
rect 7377 7701 7389 7704
rect 7331 7695 7389 7701
rect 7466 7692 7472 7704
rect 7524 7692 7530 7744
rect 8110 7732 8116 7744
rect 8071 7704 8116 7732
rect 8110 7692 8116 7704
rect 8168 7692 8174 7744
rect 9861 7735 9919 7741
rect 9861 7701 9873 7735
rect 9907 7732 9919 7735
rect 10502 7732 10508 7744
rect 9907 7704 10508 7732
rect 9907 7701 9919 7704
rect 9861 7695 9919 7701
rect 10502 7692 10508 7704
rect 10560 7692 10566 7744
rect 10870 7692 10876 7744
rect 10928 7732 10934 7744
rect 11379 7735 11437 7741
rect 11379 7732 11391 7735
rect 10928 7704 11391 7732
rect 10928 7692 10934 7704
rect 11379 7701 11391 7704
rect 11425 7701 11437 7735
rect 11379 7695 11437 7701
rect 11882 7692 11888 7744
rect 11940 7732 11946 7744
rect 13265 7735 13323 7741
rect 13265 7732 13277 7735
rect 11940 7704 13277 7732
rect 11940 7692 11946 7704
rect 13265 7701 13277 7704
rect 13311 7701 13323 7735
rect 13265 7695 13323 7701
rect 13955 7735 14013 7741
rect 13955 7701 13967 7735
rect 14001 7732 14013 7735
rect 14918 7732 14924 7744
rect 14001 7704 14924 7732
rect 14001 7701 14013 7704
rect 13955 7695 14013 7701
rect 14918 7692 14924 7704
rect 14976 7692 14982 7744
rect 25038 7732 25044 7744
rect 24999 7704 25044 7732
rect 25038 7692 25044 7704
rect 25096 7692 25102 7744
rect 1104 7642 38824 7664
rect 1104 7590 7648 7642
rect 7700 7590 7712 7642
rect 7764 7590 7776 7642
rect 7828 7590 7840 7642
rect 7892 7590 20982 7642
rect 21034 7590 21046 7642
rect 21098 7590 21110 7642
rect 21162 7590 21174 7642
rect 21226 7590 34315 7642
rect 34367 7590 34379 7642
rect 34431 7590 34443 7642
rect 34495 7590 34507 7642
rect 34559 7590 38824 7642
rect 1104 7568 38824 7590
rect 2774 7528 2780 7540
rect 2735 7500 2780 7528
rect 2774 7488 2780 7500
rect 2832 7488 2838 7540
rect 4433 7531 4491 7537
rect 4433 7497 4445 7531
rect 4479 7528 4491 7531
rect 7282 7528 7288 7540
rect 4479 7500 7288 7528
rect 4479 7497 4491 7500
rect 4433 7491 4491 7497
rect 7282 7488 7288 7500
rect 7340 7488 7346 7540
rect 8570 7528 8576 7540
rect 8531 7500 8576 7528
rect 8570 7488 8576 7500
rect 8628 7488 8634 7540
rect 10689 7531 10747 7537
rect 10689 7497 10701 7531
rect 10735 7528 10747 7531
rect 10962 7528 10968 7540
rect 10735 7500 10968 7528
rect 10735 7497 10747 7500
rect 10689 7491 10747 7497
rect 10962 7488 10968 7500
rect 11020 7528 11026 7540
rect 12253 7531 12311 7537
rect 12253 7528 12265 7531
rect 11020 7500 12265 7528
rect 11020 7488 11026 7500
rect 12253 7497 12265 7500
rect 12299 7528 12311 7531
rect 12434 7528 12440 7540
rect 12299 7500 12440 7528
rect 12299 7497 12311 7500
rect 12253 7491 12311 7497
rect 12434 7488 12440 7500
rect 12492 7488 12498 7540
rect 13446 7528 13452 7540
rect 13407 7500 13452 7528
rect 13446 7488 13452 7500
rect 13504 7488 13510 7540
rect 24670 7528 24676 7540
rect 24631 7500 24676 7528
rect 24670 7488 24676 7500
rect 24728 7488 24734 7540
rect 2792 7392 2820 7488
rect 4249 7463 4307 7469
rect 4249 7429 4261 7463
rect 4295 7460 4307 7463
rect 4706 7460 4712 7472
rect 4295 7432 4712 7460
rect 4295 7429 4307 7432
rect 4249 7423 4307 7429
rect 4706 7420 4712 7432
rect 4764 7460 4770 7472
rect 4764 7432 8340 7460
rect 4764 7420 4770 7432
rect 3053 7395 3111 7401
rect 3053 7392 3065 7395
rect 2792 7364 3065 7392
rect 3053 7361 3065 7364
rect 3099 7361 3111 7395
rect 3326 7392 3332 7404
rect 3287 7364 3332 7392
rect 3053 7355 3111 7361
rect 3326 7352 3332 7364
rect 3384 7392 3390 7404
rect 4890 7392 4896 7404
rect 3384 7364 4896 7392
rect 3384 7352 3390 7364
rect 4890 7352 4896 7364
rect 4948 7392 4954 7404
rect 5537 7395 5595 7401
rect 5537 7392 5549 7395
rect 4948 7364 5549 7392
rect 4948 7352 4954 7364
rect 5537 7361 5549 7364
rect 5583 7361 5595 7395
rect 5537 7355 5595 7361
rect 6822 7352 6828 7404
rect 6880 7392 6886 7404
rect 7653 7395 7711 7401
rect 7653 7392 7665 7395
rect 6880 7364 7665 7392
rect 6880 7352 6886 7364
rect 7653 7361 7665 7364
rect 7699 7392 7711 7395
rect 8110 7392 8116 7404
rect 7699 7364 8116 7392
rect 7699 7361 7711 7364
rect 7653 7355 7711 7361
rect 8110 7352 8116 7364
rect 8168 7352 8174 7404
rect 1394 7324 1400 7336
rect 1355 7296 1400 7324
rect 1394 7284 1400 7296
rect 1452 7324 1458 7336
rect 1949 7327 2007 7333
rect 1949 7324 1961 7327
rect 1452 7296 1961 7324
rect 1452 7284 1458 7296
rect 1949 7293 1961 7296
rect 1995 7293 2007 7327
rect 1949 7287 2007 7293
rect 106 7148 112 7200
rect 164 7188 170 7200
rect 1581 7191 1639 7197
rect 1581 7188 1593 7191
rect 164 7160 1593 7188
rect 164 7148 170 7160
rect 1581 7157 1593 7160
rect 1627 7157 1639 7191
rect 1964 7188 1992 7287
rect 2501 7259 2559 7265
rect 2501 7225 2513 7259
rect 2547 7256 2559 7259
rect 3142 7256 3148 7268
rect 2547 7228 3148 7256
rect 2547 7225 2559 7228
rect 2501 7219 2559 7225
rect 3142 7216 3148 7228
rect 3200 7216 3206 7268
rect 5258 7256 5264 7268
rect 5219 7228 5264 7256
rect 5258 7216 5264 7228
rect 5316 7216 5322 7268
rect 5353 7259 5411 7265
rect 5353 7225 5365 7259
rect 5399 7225 5411 7259
rect 5353 7219 5411 7225
rect 7745 7259 7803 7265
rect 7745 7225 7757 7259
rect 7791 7256 7803 7259
rect 8018 7256 8024 7268
rect 7791 7228 8024 7256
rect 7791 7225 7803 7228
rect 7745 7219 7803 7225
rect 4433 7191 4491 7197
rect 4433 7188 4445 7191
rect 1964 7160 4445 7188
rect 1581 7151 1639 7157
rect 4433 7157 4445 7160
rect 4479 7157 4491 7191
rect 4614 7188 4620 7200
rect 4575 7160 4620 7188
rect 4433 7151 4491 7157
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 5077 7191 5135 7197
rect 5077 7157 5089 7191
rect 5123 7188 5135 7191
rect 5368 7188 5396 7219
rect 8018 7216 8024 7228
rect 8076 7216 8082 7268
rect 8312 7265 8340 7432
rect 11054 7420 11060 7472
rect 11112 7460 11118 7472
rect 11793 7463 11851 7469
rect 11793 7460 11805 7463
rect 11112 7432 11805 7460
rect 11112 7420 11118 7432
rect 11793 7429 11805 7432
rect 11839 7460 11851 7463
rect 13998 7460 14004 7472
rect 11839 7432 14004 7460
rect 11839 7429 11851 7432
rect 11793 7423 11851 7429
rect 13998 7420 14004 7432
rect 14056 7420 14062 7472
rect 10870 7392 10876 7404
rect 10831 7364 10876 7392
rect 10870 7352 10876 7364
rect 10928 7352 10934 7404
rect 11882 7352 11888 7404
rect 11940 7392 11946 7404
rect 12529 7395 12587 7401
rect 12529 7392 12541 7395
rect 11940 7364 12541 7392
rect 11940 7352 11946 7364
rect 12529 7361 12541 7364
rect 12575 7361 12587 7395
rect 12802 7392 12808 7404
rect 12763 7364 12808 7392
rect 12529 7355 12587 7361
rect 12802 7352 12808 7364
rect 12860 7352 12866 7404
rect 12986 7352 12992 7404
rect 13044 7392 13050 7404
rect 25041 7395 25099 7401
rect 13044 7364 15643 7392
rect 13044 7352 13050 7364
rect 9836 7327 9894 7333
rect 9836 7293 9848 7327
rect 9882 7324 9894 7327
rect 10321 7327 10379 7333
rect 10321 7324 10333 7327
rect 9882 7296 10333 7324
rect 9882 7293 9894 7296
rect 9836 7287 9894 7293
rect 10321 7293 10333 7296
rect 10367 7324 10379 7327
rect 10594 7324 10600 7336
rect 10367 7296 10600 7324
rect 10367 7293 10379 7296
rect 10321 7287 10379 7293
rect 10594 7284 10600 7296
rect 10652 7284 10658 7336
rect 13906 7324 13912 7336
rect 13867 7296 13912 7324
rect 13906 7284 13912 7296
rect 13964 7284 13970 7336
rect 15615 7333 15643 7364
rect 25041 7361 25053 7395
rect 25087 7392 25099 7395
rect 25130 7392 25136 7404
rect 25087 7364 25136 7392
rect 25087 7361 25099 7364
rect 25041 7355 25099 7361
rect 25130 7352 25136 7364
rect 25188 7352 25194 7404
rect 14068 7327 14126 7333
rect 14068 7293 14080 7327
rect 14114 7324 14126 7327
rect 15600 7327 15658 7333
rect 14114 7296 14596 7324
rect 14114 7293 14126 7296
rect 14068 7287 14126 7293
rect 8297 7259 8355 7265
rect 8297 7225 8309 7259
rect 8343 7256 8355 7259
rect 10962 7256 10968 7268
rect 8343 7228 10364 7256
rect 10923 7228 10968 7256
rect 8343 7225 8355 7228
rect 8297 7219 8355 7225
rect 5534 7188 5540 7200
rect 5123 7160 5540 7188
rect 5123 7157 5135 7160
rect 5077 7151 5135 7157
rect 5534 7148 5540 7160
rect 5592 7148 5598 7200
rect 7282 7188 7288 7200
rect 7243 7160 7288 7188
rect 7282 7148 7288 7160
rect 7340 7148 7346 7200
rect 9582 7188 9588 7200
rect 9543 7160 9588 7188
rect 9582 7148 9588 7160
rect 9640 7148 9646 7200
rect 9674 7148 9680 7200
rect 9732 7188 9738 7200
rect 9907 7191 9965 7197
rect 9907 7188 9919 7191
rect 9732 7160 9919 7188
rect 9732 7148 9738 7160
rect 9907 7157 9919 7160
rect 9953 7157 9965 7191
rect 10336 7188 10364 7228
rect 10962 7216 10968 7228
rect 11020 7216 11026 7268
rect 11517 7259 11575 7265
rect 11517 7225 11529 7259
rect 11563 7256 11575 7259
rect 11606 7256 11612 7268
rect 11563 7228 11612 7256
rect 11563 7225 11575 7228
rect 11517 7219 11575 7225
rect 11532 7188 11560 7219
rect 11606 7216 11612 7228
rect 11664 7216 11670 7268
rect 12618 7216 12624 7268
rect 12676 7256 12682 7268
rect 12676 7228 12721 7256
rect 12676 7216 12682 7228
rect 10336 7160 11560 7188
rect 9907 7151 9965 7157
rect 13906 7148 13912 7200
rect 13964 7188 13970 7200
rect 14568 7197 14596 7296
rect 15600 7293 15612 7327
rect 15646 7324 15658 7327
rect 16025 7327 16083 7333
rect 16025 7324 16037 7327
rect 15646 7296 16037 7324
rect 15646 7293 15658 7296
rect 15600 7287 15658 7293
rect 16025 7293 16037 7296
rect 16071 7293 16083 7327
rect 16025 7287 16083 7293
rect 17012 7327 17070 7333
rect 17012 7293 17024 7327
rect 17058 7324 17070 7327
rect 17865 7327 17923 7333
rect 17058 7296 17540 7324
rect 17058 7293 17070 7296
rect 17012 7287 17070 7293
rect 14139 7191 14197 7197
rect 14139 7188 14151 7191
rect 13964 7160 14151 7188
rect 13964 7148 13970 7160
rect 14139 7157 14151 7160
rect 14185 7157 14197 7191
rect 14139 7151 14197 7157
rect 14553 7191 14611 7197
rect 14553 7157 14565 7191
rect 14599 7188 14611 7191
rect 14734 7188 14740 7200
rect 14599 7160 14740 7188
rect 14599 7157 14611 7160
rect 14553 7151 14611 7157
rect 14734 7148 14740 7160
rect 14792 7148 14798 7200
rect 15562 7148 15568 7200
rect 15620 7188 15626 7200
rect 15703 7191 15761 7197
rect 15703 7188 15715 7191
rect 15620 7160 15715 7188
rect 15620 7148 15626 7160
rect 15703 7157 15715 7160
rect 15749 7157 15761 7191
rect 16666 7188 16672 7200
rect 16627 7160 16672 7188
rect 15703 7151 15761 7157
rect 16666 7148 16672 7160
rect 16724 7148 16730 7200
rect 16758 7148 16764 7200
rect 16816 7188 16822 7200
rect 17512 7197 17540 7296
rect 17865 7293 17877 7327
rect 17911 7324 17923 7327
rect 18141 7327 18199 7333
rect 18141 7324 18153 7327
rect 17911 7296 18153 7324
rect 17911 7293 17923 7296
rect 17865 7287 17923 7293
rect 18141 7293 18153 7296
rect 18187 7324 18199 7327
rect 18230 7324 18236 7336
rect 18187 7296 18236 7324
rect 18187 7293 18199 7296
rect 18141 7287 18199 7293
rect 18230 7284 18236 7296
rect 18288 7284 18294 7336
rect 24004 7327 24062 7333
rect 24004 7293 24016 7327
rect 24050 7324 24062 7327
rect 24302 7324 24308 7336
rect 24050 7296 24308 7324
rect 24050 7293 24062 7296
rect 24004 7287 24062 7293
rect 24302 7284 24308 7296
rect 24360 7284 24366 7336
rect 17586 7216 17592 7268
rect 17644 7256 17650 7268
rect 18049 7259 18107 7265
rect 18049 7256 18061 7259
rect 17644 7228 18061 7256
rect 17644 7216 17650 7228
rect 18049 7225 18061 7228
rect 18095 7225 18107 7259
rect 18049 7219 18107 7225
rect 24394 7216 24400 7268
rect 24452 7256 24458 7268
rect 25038 7256 25044 7268
rect 24452 7228 25044 7256
rect 24452 7216 24458 7228
rect 25038 7216 25044 7228
rect 25096 7256 25102 7268
rect 25133 7259 25191 7265
rect 25133 7256 25145 7259
rect 25096 7228 25145 7256
rect 25096 7216 25102 7228
rect 25133 7225 25145 7228
rect 25179 7225 25191 7259
rect 25133 7219 25191 7225
rect 25685 7259 25743 7265
rect 25685 7225 25697 7259
rect 25731 7256 25743 7259
rect 25774 7256 25780 7268
rect 25731 7228 25780 7256
rect 25731 7225 25743 7228
rect 25685 7219 25743 7225
rect 25774 7216 25780 7228
rect 25832 7216 25838 7268
rect 17083 7191 17141 7197
rect 17083 7188 17095 7191
rect 16816 7160 17095 7188
rect 16816 7148 16822 7160
rect 17083 7157 17095 7160
rect 17129 7157 17141 7191
rect 17083 7151 17141 7157
rect 17497 7191 17555 7197
rect 17497 7157 17509 7191
rect 17543 7188 17555 7191
rect 18322 7188 18328 7200
rect 17543 7160 18328 7188
rect 17543 7157 17555 7160
rect 17497 7151 17555 7157
rect 18322 7148 18328 7160
rect 18380 7148 18386 7200
rect 24075 7191 24133 7197
rect 24075 7157 24087 7191
rect 24121 7188 24133 7191
rect 24486 7188 24492 7200
rect 24121 7160 24492 7188
rect 24121 7157 24133 7160
rect 24075 7151 24133 7157
rect 24486 7148 24492 7160
rect 24544 7148 24550 7200
rect 32214 7188 32220 7200
rect 32175 7160 32220 7188
rect 32214 7148 32220 7160
rect 32272 7148 32278 7200
rect 1104 7098 38824 7120
rect 1104 7046 14315 7098
rect 14367 7046 14379 7098
rect 14431 7046 14443 7098
rect 14495 7046 14507 7098
rect 14559 7046 27648 7098
rect 27700 7046 27712 7098
rect 27764 7046 27776 7098
rect 27828 7046 27840 7098
rect 27892 7046 38824 7098
rect 1104 7024 38824 7046
rect 2498 6944 2504 6996
rect 2556 6984 2562 6996
rect 3789 6987 3847 6993
rect 3789 6984 3801 6987
rect 2556 6956 3801 6984
rect 2556 6944 2562 6956
rect 3789 6953 3801 6956
rect 3835 6953 3847 6987
rect 4982 6984 4988 6996
rect 4943 6956 4988 6984
rect 3789 6947 3847 6953
rect 4982 6944 4988 6956
rect 5040 6944 5046 6996
rect 5534 6984 5540 6996
rect 5495 6956 5540 6984
rect 5534 6944 5540 6956
rect 5592 6944 5598 6996
rect 6822 6984 6828 6996
rect 6783 6956 6828 6984
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 10870 6984 10876 6996
rect 10831 6956 10876 6984
rect 10870 6944 10876 6956
rect 10928 6944 10934 6996
rect 12161 6987 12219 6993
rect 12161 6953 12173 6987
rect 12207 6984 12219 6987
rect 12434 6984 12440 6996
rect 12207 6956 12440 6984
rect 12207 6953 12219 6956
rect 12161 6947 12219 6953
rect 12434 6944 12440 6956
rect 12492 6944 12498 6996
rect 16485 6987 16543 6993
rect 16485 6953 16497 6987
rect 16531 6984 16543 6987
rect 16758 6984 16764 6996
rect 16531 6956 16764 6984
rect 16531 6953 16543 6956
rect 16485 6947 16543 6953
rect 16758 6944 16764 6956
rect 16816 6944 16822 6996
rect 7469 6919 7527 6925
rect 7469 6885 7481 6919
rect 7515 6916 7527 6919
rect 7745 6919 7803 6925
rect 7745 6916 7757 6919
rect 7515 6888 7757 6916
rect 7515 6885 7527 6888
rect 7469 6879 7527 6885
rect 7745 6885 7757 6888
rect 7791 6916 7803 6919
rect 8018 6916 8024 6928
rect 7791 6888 8024 6916
rect 7791 6885 7803 6888
rect 7745 6879 7803 6885
rect 8018 6876 8024 6888
rect 8076 6876 8082 6928
rect 8294 6916 8300 6928
rect 8207 6888 8300 6916
rect 8294 6876 8300 6888
rect 8352 6916 8358 6928
rect 8352 6888 11284 6916
rect 8352 6876 8358 6888
rect 2038 6808 2044 6860
rect 2096 6848 2102 6860
rect 2593 6851 2651 6857
rect 2593 6848 2605 6851
rect 2096 6820 2605 6848
rect 2096 6808 2102 6820
rect 2593 6817 2605 6820
rect 2639 6817 2651 6851
rect 6454 6848 6460 6860
rect 6415 6820 6460 6848
rect 2593 6811 2651 6817
rect 6454 6808 6460 6820
rect 6512 6808 6518 6860
rect 9766 6848 9772 6860
rect 9727 6820 9772 6848
rect 9766 6808 9772 6820
rect 9824 6808 9830 6860
rect 11256 6848 11284 6888
rect 11330 6876 11336 6928
rect 11388 6916 11394 6928
rect 11562 6919 11620 6925
rect 11562 6916 11574 6919
rect 11388 6888 11574 6916
rect 11388 6876 11394 6888
rect 11562 6885 11574 6888
rect 11608 6885 11620 6919
rect 11562 6879 11620 6885
rect 12529 6919 12587 6925
rect 12529 6885 12541 6919
rect 12575 6916 12587 6919
rect 12618 6916 12624 6928
rect 12575 6888 12624 6916
rect 12575 6885 12587 6888
rect 12529 6879 12587 6885
rect 12618 6876 12624 6888
rect 12676 6916 12682 6928
rect 13170 6916 13176 6928
rect 12676 6888 13176 6916
rect 12676 6876 12682 6888
rect 13170 6876 13176 6888
rect 13228 6876 13234 6928
rect 15378 6916 15384 6928
rect 15339 6888 15384 6916
rect 15378 6876 15384 6888
rect 15436 6876 15442 6928
rect 15470 6876 15476 6928
rect 15528 6916 15534 6928
rect 16022 6916 16028 6928
rect 15528 6888 15573 6916
rect 15983 6888 16028 6916
rect 15528 6876 15534 6888
rect 16022 6876 16028 6888
rect 16080 6876 16086 6928
rect 17586 6916 17592 6928
rect 17547 6888 17592 6916
rect 17586 6876 17592 6888
rect 17644 6876 17650 6928
rect 24486 6876 24492 6928
rect 24544 6916 24550 6928
rect 24949 6919 25007 6925
rect 24949 6916 24961 6919
rect 24544 6888 24961 6916
rect 24544 6876 24550 6888
rect 24949 6885 24961 6888
rect 24995 6885 25007 6919
rect 24949 6879 25007 6885
rect 25038 6876 25044 6928
rect 25096 6916 25102 6928
rect 26694 6916 26700 6928
rect 25096 6888 26700 6916
rect 25096 6876 25102 6888
rect 26694 6876 26700 6888
rect 26752 6876 26758 6928
rect 12802 6848 12808 6860
rect 11256 6820 12808 6848
rect 12802 6808 12808 6820
rect 12860 6808 12866 6860
rect 20162 6808 20168 6860
rect 20220 6848 20226 6860
rect 20901 6851 20959 6857
rect 20901 6848 20913 6851
rect 20220 6820 20913 6848
rect 20220 6808 20226 6820
rect 20901 6817 20913 6820
rect 20947 6817 20959 6851
rect 21358 6848 21364 6860
rect 21319 6820 21364 6848
rect 20901 6811 20959 6817
rect 21358 6808 21364 6820
rect 21416 6808 21422 6860
rect 21910 6848 21916 6860
rect 21871 6820 21916 6848
rect 21910 6808 21916 6820
rect 21968 6808 21974 6860
rect 22094 6848 22100 6860
rect 22055 6820 22100 6848
rect 22094 6808 22100 6820
rect 22152 6808 22158 6860
rect 23290 6808 23296 6860
rect 23348 6848 23354 6860
rect 23788 6851 23846 6857
rect 23788 6848 23800 6851
rect 23348 6820 23800 6848
rect 23348 6808 23354 6820
rect 23788 6817 23800 6820
rect 23834 6817 23846 6851
rect 34606 6848 34612 6860
rect 34567 6820 34612 6848
rect 23788 6811 23846 6817
rect 34606 6808 34612 6820
rect 34664 6808 34670 6860
rect 1578 6780 1584 6792
rect 1539 6752 1584 6780
rect 1578 6740 1584 6752
rect 1636 6740 1642 6792
rect 4617 6783 4675 6789
rect 4617 6749 4629 6783
rect 4663 6780 4675 6783
rect 5534 6780 5540 6792
rect 4663 6752 5540 6780
rect 4663 6749 4675 6752
rect 4617 6743 4675 6749
rect 5534 6740 5540 6752
rect 5592 6740 5598 6792
rect 7466 6740 7472 6792
rect 7524 6780 7530 6792
rect 7653 6783 7711 6789
rect 7653 6780 7665 6783
rect 7524 6752 7665 6780
rect 7524 6740 7530 6752
rect 7653 6749 7665 6752
rect 7699 6780 7711 6783
rect 8573 6783 8631 6789
rect 8573 6780 8585 6783
rect 7699 6752 8585 6780
rect 7699 6749 7711 6752
rect 7653 6743 7711 6749
rect 8573 6749 8585 6752
rect 8619 6749 8631 6783
rect 8573 6743 8631 6749
rect 11241 6783 11299 6789
rect 11241 6749 11253 6783
rect 11287 6780 11299 6783
rect 11514 6780 11520 6792
rect 11287 6752 11520 6780
rect 11287 6749 11299 6752
rect 11241 6743 11299 6749
rect 11514 6740 11520 6752
rect 11572 6740 11578 6792
rect 13081 6783 13139 6789
rect 13081 6749 13093 6783
rect 13127 6780 13139 6783
rect 13446 6780 13452 6792
rect 13127 6752 13452 6780
rect 13127 6749 13139 6752
rect 13081 6743 13139 6749
rect 13446 6740 13452 6752
rect 13504 6740 13510 6792
rect 17497 6783 17555 6789
rect 17497 6749 17509 6783
rect 17543 6780 17555 6783
rect 17862 6780 17868 6792
rect 17543 6752 17868 6780
rect 17543 6749 17555 6752
rect 17497 6743 17555 6749
rect 17862 6740 17868 6752
rect 17920 6780 17926 6792
rect 18969 6783 19027 6789
rect 18969 6780 18981 6783
rect 17920 6752 18981 6780
rect 17920 6740 17926 6752
rect 18969 6749 18981 6752
rect 19015 6749 19027 6783
rect 18969 6743 19027 6749
rect 22373 6783 22431 6789
rect 22373 6749 22385 6783
rect 22419 6780 22431 6783
rect 23566 6780 23572 6792
rect 22419 6752 23572 6780
rect 22419 6749 22431 6752
rect 22373 6743 22431 6749
rect 23566 6740 23572 6752
rect 23624 6780 23630 6792
rect 24213 6783 24271 6789
rect 24213 6780 24225 6783
rect 23624 6752 24225 6780
rect 23624 6740 23630 6752
rect 24213 6749 24225 6752
rect 24259 6749 24271 6783
rect 24213 6743 24271 6749
rect 25593 6783 25651 6789
rect 25593 6749 25605 6783
rect 25639 6780 25651 6783
rect 26050 6780 26056 6792
rect 25639 6752 26056 6780
rect 25639 6749 25651 6752
rect 25593 6743 25651 6749
rect 26050 6740 26056 6752
rect 26108 6740 26114 6792
rect 26602 6780 26608 6792
rect 26563 6752 26608 6780
rect 26602 6740 26608 6752
rect 26660 6740 26666 6792
rect 26881 6783 26939 6789
rect 26881 6749 26893 6783
rect 26927 6749 26939 6783
rect 26881 6743 26939 6749
rect 2777 6715 2835 6721
rect 2777 6681 2789 6715
rect 2823 6712 2835 6715
rect 6638 6712 6644 6724
rect 2823 6684 6644 6712
rect 2823 6681 2835 6684
rect 2777 6675 2835 6681
rect 6638 6672 6644 6684
rect 6696 6672 6702 6724
rect 10042 6672 10048 6724
rect 10100 6712 10106 6724
rect 10229 6715 10287 6721
rect 10229 6712 10241 6715
rect 10100 6684 10241 6712
rect 10100 6672 10106 6684
rect 10229 6681 10241 6684
rect 10275 6681 10287 6715
rect 10229 6675 10287 6681
rect 11606 6672 11612 6724
rect 11664 6712 11670 6724
rect 13633 6715 13691 6721
rect 13633 6712 13645 6715
rect 11664 6684 13645 6712
rect 11664 6672 11670 6684
rect 13633 6681 13645 6684
rect 13679 6681 13691 6715
rect 13633 6675 13691 6681
rect 16666 6672 16672 6724
rect 16724 6712 16730 6724
rect 18049 6715 18107 6721
rect 18049 6712 18061 6715
rect 16724 6684 18061 6712
rect 16724 6672 16730 6684
rect 18049 6681 18061 6684
rect 18095 6712 18107 6715
rect 18506 6712 18512 6724
rect 18095 6684 18512 6712
rect 18095 6681 18107 6684
rect 18049 6675 18107 6681
rect 18506 6672 18512 6684
rect 18564 6672 18570 6724
rect 25774 6672 25780 6724
rect 25832 6712 25838 6724
rect 26418 6712 26424 6724
rect 25832 6684 26424 6712
rect 25832 6672 25838 6684
rect 26418 6672 26424 6684
rect 26476 6712 26482 6724
rect 26896 6712 26924 6743
rect 26476 6684 26924 6712
rect 26476 6672 26482 6684
rect 2314 6644 2320 6656
rect 2275 6616 2320 6644
rect 2314 6604 2320 6616
rect 2372 6604 2378 6656
rect 3050 6644 3056 6656
rect 3011 6616 3056 6644
rect 3050 6604 3056 6616
rect 3108 6604 3114 6656
rect 3510 6644 3516 6656
rect 3471 6616 3516 6644
rect 3510 6604 3516 6616
rect 3568 6604 3574 6656
rect 4338 6644 4344 6656
rect 4299 6616 4344 6644
rect 4338 6604 4344 6616
rect 4396 6604 4402 6656
rect 7101 6647 7159 6653
rect 7101 6613 7113 6647
rect 7147 6644 7159 6647
rect 7190 6644 7196 6656
rect 7147 6616 7196 6644
rect 7147 6613 7159 6616
rect 7101 6607 7159 6613
rect 7190 6604 7196 6616
rect 7248 6604 7254 6656
rect 8938 6604 8944 6656
rect 8996 6644 9002 6656
rect 9953 6647 10011 6653
rect 9953 6644 9965 6647
rect 8996 6616 9965 6644
rect 8996 6604 9002 6616
rect 9953 6613 9965 6616
rect 9999 6644 10011 6647
rect 10134 6644 10140 6656
rect 9999 6616 10140 6644
rect 9999 6613 10011 6616
rect 9953 6607 10011 6613
rect 10134 6604 10140 6616
rect 10192 6604 10198 6656
rect 12618 6604 12624 6656
rect 12676 6644 12682 6656
rect 12805 6647 12863 6653
rect 12805 6644 12817 6647
rect 12676 6616 12817 6644
rect 12676 6604 12682 6616
rect 12805 6613 12817 6616
rect 12851 6613 12863 6647
rect 14366 6644 14372 6656
rect 14327 6616 14372 6644
rect 12805 6607 12863 6613
rect 14366 6604 14372 6616
rect 14424 6604 14430 6656
rect 18414 6644 18420 6656
rect 18375 6616 18420 6644
rect 18414 6604 18420 6616
rect 18472 6604 18478 6656
rect 20162 6644 20168 6656
rect 20123 6616 20168 6644
rect 20162 6604 20168 6616
rect 20220 6604 20226 6656
rect 20622 6644 20628 6656
rect 20583 6616 20628 6644
rect 20622 6604 20628 6616
rect 20680 6604 20686 6656
rect 23891 6647 23949 6653
rect 23891 6613 23903 6647
rect 23937 6644 23949 6647
rect 25130 6644 25136 6656
rect 23937 6616 25136 6644
rect 23937 6613 23949 6616
rect 23891 6607 23949 6613
rect 25130 6604 25136 6616
rect 25188 6604 25194 6656
rect 27982 6604 27988 6656
rect 28040 6644 28046 6656
rect 34747 6647 34805 6653
rect 34747 6644 34759 6647
rect 28040 6616 34759 6644
rect 28040 6604 28046 6616
rect 34747 6613 34759 6616
rect 34793 6613 34805 6647
rect 34747 6607 34805 6613
rect 1104 6554 38824 6576
rect 1104 6502 7648 6554
rect 7700 6502 7712 6554
rect 7764 6502 7776 6554
rect 7828 6502 7840 6554
rect 7892 6502 20982 6554
rect 21034 6502 21046 6554
rect 21098 6502 21110 6554
rect 21162 6502 21174 6554
rect 21226 6502 34315 6554
rect 34367 6502 34379 6554
rect 34431 6502 34443 6554
rect 34495 6502 34507 6554
rect 34559 6502 38824 6554
rect 1104 6480 38824 6502
rect 2038 6440 2044 6452
rect 1999 6412 2044 6440
rect 2038 6400 2044 6412
rect 2096 6400 2102 6452
rect 4614 6400 4620 6452
rect 4672 6440 4678 6452
rect 5445 6443 5503 6449
rect 5445 6440 5457 6443
rect 4672 6412 5457 6440
rect 4672 6400 4678 6412
rect 5445 6409 5457 6412
rect 5491 6409 5503 6443
rect 5445 6403 5503 6409
rect 8018 6400 8024 6452
rect 8076 6440 8082 6452
rect 8113 6443 8171 6449
rect 8113 6440 8125 6443
rect 8076 6412 8125 6440
rect 8076 6400 8082 6412
rect 8113 6409 8125 6412
rect 8159 6409 8171 6443
rect 8113 6403 8171 6409
rect 13170 6400 13176 6452
rect 13228 6440 13234 6452
rect 13357 6443 13415 6449
rect 13357 6440 13369 6443
rect 13228 6412 13369 6440
rect 13228 6400 13234 6412
rect 13357 6409 13369 6412
rect 13403 6440 13415 6443
rect 13633 6443 13691 6449
rect 13633 6440 13645 6443
rect 13403 6412 13645 6440
rect 13403 6409 13415 6412
rect 13357 6403 13415 6409
rect 13633 6409 13645 6412
rect 13679 6409 13691 6443
rect 15378 6440 15384 6452
rect 15339 6412 15384 6440
rect 13633 6403 13691 6409
rect 15378 6400 15384 6412
rect 15436 6400 15442 6452
rect 17497 6443 17555 6449
rect 17497 6409 17509 6443
rect 17543 6440 17555 6443
rect 17586 6440 17592 6452
rect 17543 6412 17592 6440
rect 17543 6409 17555 6412
rect 17497 6403 17555 6409
rect 17586 6400 17592 6412
rect 17644 6400 17650 6452
rect 17862 6440 17868 6452
rect 17823 6412 17868 6440
rect 17862 6400 17868 6412
rect 17920 6400 17926 6452
rect 24581 6443 24639 6449
rect 24581 6409 24593 6443
rect 24627 6440 24639 6443
rect 24949 6443 25007 6449
rect 24949 6440 24961 6443
rect 24627 6412 24961 6440
rect 24627 6409 24639 6412
rect 24581 6403 24639 6409
rect 24949 6409 24961 6412
rect 24995 6440 25007 6443
rect 25038 6440 25044 6452
rect 24995 6412 25044 6440
rect 24995 6409 25007 6412
rect 24949 6403 25007 6409
rect 25038 6400 25044 6412
rect 25096 6400 25102 6452
rect 26605 6443 26663 6449
rect 26605 6409 26617 6443
rect 26651 6440 26663 6443
rect 26694 6440 26700 6452
rect 26651 6412 26700 6440
rect 26651 6409 26663 6412
rect 26605 6403 26663 6409
rect 26694 6400 26700 6412
rect 26752 6400 26758 6452
rect 32033 6443 32091 6449
rect 32033 6409 32045 6443
rect 32079 6440 32091 6443
rect 32214 6440 32220 6452
rect 32079 6412 32220 6440
rect 32079 6409 32091 6412
rect 32033 6403 32091 6409
rect 3510 6332 3516 6384
rect 3568 6372 3574 6384
rect 3605 6375 3663 6381
rect 3605 6372 3617 6375
rect 3568 6344 3617 6372
rect 3568 6332 3574 6344
rect 3605 6341 3617 6344
rect 3651 6341 3663 6375
rect 3605 6335 3663 6341
rect 6454 6332 6460 6384
rect 6512 6372 6518 6384
rect 6641 6375 6699 6381
rect 6641 6372 6653 6375
rect 6512 6344 6653 6372
rect 6512 6332 6518 6344
rect 6641 6341 6653 6344
rect 6687 6372 6699 6375
rect 7374 6372 7380 6384
rect 6687 6344 7380 6372
rect 6687 6341 6699 6344
rect 6641 6335 6699 6341
rect 7374 6332 7380 6344
rect 7432 6372 7438 6384
rect 10594 6372 10600 6384
rect 7432 6344 10600 6372
rect 7432 6332 7438 6344
rect 10594 6332 10600 6344
rect 10652 6332 10658 6384
rect 26050 6332 26056 6384
rect 26108 6372 26114 6384
rect 27617 6375 27675 6381
rect 27617 6372 27629 6375
rect 26108 6344 27629 6372
rect 26108 6332 26114 6344
rect 27617 6341 27629 6344
rect 27663 6341 27675 6375
rect 27617 6335 27675 6341
rect 2314 6264 2320 6316
rect 2372 6304 2378 6316
rect 4246 6304 4252 6316
rect 2372 6276 4252 6304
rect 2372 6264 2378 6276
rect 2516 6245 2544 6276
rect 4246 6264 4252 6276
rect 4304 6264 4310 6316
rect 10042 6264 10048 6316
rect 10100 6304 10106 6316
rect 14366 6304 14372 6316
rect 10100 6276 10180 6304
rect 10100 6264 10106 6276
rect 2501 6239 2559 6245
rect 2501 6205 2513 6239
rect 2547 6205 2559 6239
rect 2501 6199 2559 6205
rect 2685 6239 2743 6245
rect 2685 6205 2697 6239
rect 2731 6205 2743 6239
rect 3050 6236 3056 6248
rect 3011 6208 3056 6236
rect 2685 6199 2743 6205
rect 1670 6128 1676 6180
rect 1728 6168 1734 6180
rect 1765 6171 1823 6177
rect 1765 6168 1777 6171
rect 1728 6140 1777 6168
rect 1728 6128 1734 6140
rect 1765 6137 1777 6140
rect 1811 6168 1823 6171
rect 2700 6168 2728 6199
rect 3050 6196 3056 6208
rect 3108 6196 3114 6248
rect 3418 6236 3424 6248
rect 3379 6208 3424 6236
rect 3418 6196 3424 6208
rect 3476 6196 3482 6248
rect 4062 6196 4068 6248
rect 4120 6236 4126 6248
rect 4525 6239 4583 6245
rect 4525 6236 4537 6239
rect 4120 6208 4537 6236
rect 4120 6196 4126 6208
rect 4525 6205 4537 6208
rect 4571 6236 4583 6239
rect 5721 6239 5779 6245
rect 5721 6236 5733 6239
rect 4571 6208 5733 6236
rect 4571 6205 4583 6208
rect 4525 6199 4583 6205
rect 5721 6205 5733 6208
rect 5767 6205 5779 6239
rect 7190 6236 7196 6248
rect 7151 6208 7196 6236
rect 5721 6199 5779 6205
rect 7190 6196 7196 6208
rect 7248 6196 7254 6248
rect 8757 6239 8815 6245
rect 8757 6205 8769 6239
rect 8803 6236 8815 6239
rect 9861 6239 9919 6245
rect 9861 6236 9873 6239
rect 8803 6208 9873 6236
rect 8803 6205 8815 6208
rect 8757 6199 8815 6205
rect 9861 6205 9873 6208
rect 9907 6236 9919 6239
rect 9950 6236 9956 6248
rect 9907 6208 9956 6236
rect 9907 6205 9919 6208
rect 9861 6199 9919 6205
rect 9950 6196 9956 6208
rect 10008 6196 10014 6248
rect 10152 6245 10180 6276
rect 13786 6276 14372 6304
rect 10137 6239 10195 6245
rect 10137 6205 10149 6239
rect 10183 6205 10195 6239
rect 10137 6199 10195 6205
rect 10226 6196 10232 6248
rect 10284 6236 10290 6248
rect 10413 6239 10471 6245
rect 10413 6236 10425 6239
rect 10284 6208 10425 6236
rect 10284 6196 10290 6208
rect 10413 6205 10425 6208
rect 10459 6205 10471 6239
rect 10413 6199 10471 6205
rect 10781 6239 10839 6245
rect 10781 6205 10793 6239
rect 10827 6205 10839 6239
rect 10781 6199 10839 6205
rect 4433 6171 4491 6177
rect 4433 6168 4445 6171
rect 1811 6140 2728 6168
rect 4126 6140 4445 6168
rect 1811 6137 1823 6140
rect 1765 6131 1823 6137
rect 2774 6060 2780 6112
rect 2832 6100 2838 6112
rect 3973 6103 4031 6109
rect 3973 6100 3985 6103
rect 2832 6072 3985 6100
rect 2832 6060 2838 6072
rect 3973 6069 3985 6072
rect 4019 6100 4031 6103
rect 4126 6100 4154 6140
rect 4433 6137 4445 6140
rect 4479 6168 4491 6171
rect 4887 6171 4945 6177
rect 4887 6168 4899 6171
rect 4479 6140 4899 6168
rect 4479 6137 4491 6140
rect 4433 6131 4491 6137
rect 4887 6137 4899 6140
rect 4933 6168 4945 6171
rect 4982 6168 4988 6180
rect 4933 6140 4988 6168
rect 4933 6137 4945 6140
rect 4887 6131 4945 6137
rect 4982 6128 4988 6140
rect 5040 6128 5046 6180
rect 7514 6171 7572 6177
rect 7514 6168 7526 6171
rect 7024 6140 7526 6168
rect 4019 6072 4154 6100
rect 4019 6069 4031 6072
rect 3973 6063 4031 6069
rect 5534 6060 5540 6112
rect 5592 6100 5598 6112
rect 6089 6103 6147 6109
rect 6089 6100 6101 6103
rect 5592 6072 6101 6100
rect 5592 6060 5598 6072
rect 6089 6069 6101 6072
rect 6135 6069 6147 6103
rect 6089 6063 6147 6069
rect 6730 6060 6736 6112
rect 6788 6100 6794 6112
rect 7024 6109 7052 6140
rect 7514 6137 7526 6140
rect 7560 6137 7572 6171
rect 7514 6131 7572 6137
rect 9493 6171 9551 6177
rect 9493 6137 9505 6171
rect 9539 6168 9551 6171
rect 9766 6168 9772 6180
rect 9539 6140 9772 6168
rect 9539 6137 9551 6140
rect 9493 6131 9551 6137
rect 9766 6128 9772 6140
rect 9824 6168 9830 6180
rect 10318 6168 10324 6180
rect 9824 6140 10324 6168
rect 9824 6128 9830 6140
rect 10318 6128 10324 6140
rect 10376 6128 10382 6180
rect 7009 6103 7067 6109
rect 7009 6100 7021 6103
rect 6788 6072 7021 6100
rect 6788 6060 6794 6072
rect 7009 6069 7021 6072
rect 7055 6069 7067 6103
rect 7009 6063 7067 6069
rect 8938 6060 8944 6112
rect 8996 6100 9002 6112
rect 9033 6103 9091 6109
rect 9033 6100 9045 6103
rect 8996 6072 9045 6100
rect 8996 6060 9002 6072
rect 9033 6069 9045 6072
rect 9079 6069 9091 6103
rect 9033 6063 9091 6069
rect 10226 6060 10232 6112
rect 10284 6100 10290 6112
rect 10796 6100 10824 6199
rect 11054 6196 11060 6248
rect 11112 6236 11118 6248
rect 12437 6239 12495 6245
rect 12437 6236 12449 6239
rect 11112 6208 12449 6236
rect 11112 6196 11118 6208
rect 12437 6205 12449 6208
rect 12483 6236 12495 6239
rect 12618 6236 12624 6248
rect 12483 6208 12624 6236
rect 12483 6205 12495 6208
rect 12437 6199 12495 6205
rect 12618 6196 12624 6208
rect 12676 6196 12682 6248
rect 12161 6171 12219 6177
rect 12161 6168 12173 6171
rect 11348 6140 12173 6168
rect 11348 6112 11376 6140
rect 12161 6137 12173 6140
rect 12207 6168 12219 6171
rect 12758 6171 12816 6177
rect 12758 6168 12770 6171
rect 12207 6140 12770 6168
rect 12207 6137 12219 6140
rect 12161 6131 12219 6137
rect 12758 6137 12770 6140
rect 12804 6168 12816 6171
rect 13078 6168 13084 6180
rect 12804 6140 13084 6168
rect 12804 6137 12816 6140
rect 12758 6131 12816 6137
rect 13078 6128 13084 6140
rect 13136 6128 13142 6180
rect 13170 6128 13176 6180
rect 13228 6168 13234 6180
rect 13786 6168 13814 6276
rect 14366 6264 14372 6276
rect 14424 6264 14430 6316
rect 15013 6307 15071 6313
rect 15013 6273 15025 6307
rect 15059 6304 15071 6307
rect 16022 6304 16028 6316
rect 15059 6276 16028 6304
rect 15059 6273 15071 6276
rect 15013 6267 15071 6273
rect 16022 6264 16028 6276
rect 16080 6264 16086 6316
rect 16485 6307 16543 6313
rect 16485 6273 16497 6307
rect 16531 6304 16543 6307
rect 16758 6304 16764 6316
rect 16531 6276 16764 6304
rect 16531 6273 16543 6276
rect 16485 6267 16543 6273
rect 16758 6264 16764 6276
rect 16816 6264 16822 6316
rect 16850 6264 16856 6316
rect 16908 6304 16914 6316
rect 18141 6307 18199 6313
rect 18141 6304 18153 6307
rect 16908 6276 18153 6304
rect 16908 6264 16914 6276
rect 18141 6273 18153 6276
rect 18187 6304 18199 6307
rect 18414 6304 18420 6316
rect 18187 6276 18420 6304
rect 18187 6273 18199 6276
rect 18141 6267 18199 6273
rect 18414 6264 18420 6276
rect 18472 6264 18478 6316
rect 18506 6264 18512 6316
rect 18564 6304 18570 6316
rect 18564 6276 18609 6304
rect 18564 6264 18570 6276
rect 20714 6264 20720 6316
rect 20772 6304 20778 6316
rect 22094 6304 22100 6316
rect 20772 6276 22100 6304
rect 20772 6264 20778 6276
rect 19426 6196 19432 6248
rect 19484 6236 19490 6248
rect 19981 6239 20039 6245
rect 19981 6236 19993 6239
rect 19484 6208 19993 6236
rect 19484 6196 19490 6208
rect 19981 6205 19993 6208
rect 20027 6236 20039 6239
rect 20162 6236 20168 6248
rect 20027 6208 20168 6236
rect 20027 6205 20039 6208
rect 19981 6199 20039 6205
rect 20162 6196 20168 6208
rect 20220 6196 20226 6248
rect 20625 6239 20683 6245
rect 20625 6205 20637 6239
rect 20671 6205 20683 6239
rect 20625 6199 20683 6205
rect 21177 6239 21235 6245
rect 21177 6205 21189 6239
rect 21223 6236 21235 6239
rect 21266 6236 21272 6248
rect 21223 6208 21272 6236
rect 21223 6205 21235 6208
rect 21177 6199 21235 6205
rect 13228 6140 13814 6168
rect 14461 6171 14519 6177
rect 13228 6128 13234 6140
rect 14461 6137 14473 6171
rect 14507 6137 14519 6171
rect 14461 6131 14519 6137
rect 16301 6171 16359 6177
rect 16301 6137 16313 6171
rect 16347 6168 16359 6171
rect 16577 6171 16635 6177
rect 16577 6168 16589 6171
rect 16347 6140 16589 6168
rect 16347 6137 16359 6140
rect 16301 6131 16359 6137
rect 16577 6137 16589 6140
rect 16623 6168 16635 6171
rect 17218 6168 17224 6180
rect 16623 6140 17224 6168
rect 16623 6137 16635 6140
rect 16577 6131 16635 6137
rect 10962 6100 10968 6112
rect 10284 6072 10824 6100
rect 10923 6072 10968 6100
rect 10284 6060 10290 6072
rect 10962 6060 10968 6072
rect 11020 6060 11026 6112
rect 11330 6100 11336 6112
rect 11291 6072 11336 6100
rect 11330 6060 11336 6072
rect 11388 6060 11394 6112
rect 11514 6060 11520 6112
rect 11572 6100 11578 6112
rect 11701 6103 11759 6109
rect 11701 6100 11713 6103
rect 11572 6072 11713 6100
rect 11572 6060 11578 6072
rect 11701 6069 11713 6072
rect 11747 6069 11759 6103
rect 14182 6100 14188 6112
rect 14095 6072 14188 6100
rect 11701 6063 11759 6069
rect 14182 6060 14188 6072
rect 14240 6100 14246 6112
rect 14476 6100 14504 6131
rect 17218 6128 17224 6140
rect 17276 6128 17282 6180
rect 18230 6128 18236 6180
rect 18288 6168 18294 6180
rect 20640 6168 20668 6199
rect 21266 6196 21272 6208
rect 21324 6196 21330 6248
rect 21376 6245 21404 6276
rect 22094 6264 22100 6276
rect 22152 6304 22158 6316
rect 22281 6307 22339 6313
rect 22281 6304 22293 6307
rect 22152 6276 22293 6304
rect 22152 6264 22158 6276
rect 22281 6273 22293 6276
rect 22327 6273 22339 6307
rect 22281 6267 22339 6273
rect 23566 6264 23572 6316
rect 23624 6304 23630 6316
rect 23661 6307 23719 6313
rect 23661 6304 23673 6307
rect 23624 6276 23673 6304
rect 23624 6264 23630 6276
rect 23661 6273 23673 6276
rect 23707 6273 23719 6307
rect 23661 6267 23719 6273
rect 25130 6264 25136 6316
rect 25188 6304 25194 6316
rect 25501 6307 25559 6313
rect 25501 6304 25513 6307
rect 25188 6276 25513 6304
rect 25188 6264 25194 6276
rect 25501 6273 25513 6276
rect 25547 6273 25559 6307
rect 25774 6304 25780 6316
rect 25735 6276 25780 6304
rect 25501 6267 25559 6273
rect 25774 6264 25780 6276
rect 25832 6264 25838 6316
rect 27065 6307 27123 6313
rect 27065 6273 27077 6307
rect 27111 6304 27123 6307
rect 27982 6304 27988 6316
rect 27111 6276 27988 6304
rect 27111 6273 27123 6276
rect 27065 6267 27123 6273
rect 27982 6264 27988 6276
rect 28040 6264 28046 6316
rect 21361 6239 21419 6245
rect 21361 6205 21373 6239
rect 21407 6205 21419 6239
rect 21361 6199 21419 6205
rect 21910 6196 21916 6248
rect 21968 6236 21974 6248
rect 22649 6239 22707 6245
rect 22649 6236 22661 6239
rect 21968 6208 22661 6236
rect 21968 6196 21974 6208
rect 22649 6205 22661 6208
rect 22695 6205 22707 6239
rect 22649 6199 22707 6205
rect 31548 6239 31606 6245
rect 31548 6205 31560 6239
rect 31594 6236 31606 6239
rect 32048 6236 32076 6403
rect 32214 6400 32220 6412
rect 32272 6400 32278 6452
rect 36078 6440 36084 6452
rect 36039 6412 36084 6440
rect 36078 6400 36084 6412
rect 36136 6400 36142 6452
rect 35621 6375 35679 6381
rect 35621 6341 35633 6375
rect 35667 6372 35679 6375
rect 39574 6372 39580 6384
rect 35667 6344 39580 6372
rect 35667 6341 35679 6344
rect 35621 6335 35679 6341
rect 39574 6332 39580 6344
rect 39632 6332 39638 6384
rect 31594 6208 32076 6236
rect 31594 6205 31606 6208
rect 31548 6199 31606 6205
rect 34606 6196 34612 6248
rect 34664 6236 34670 6248
rect 34701 6239 34759 6245
rect 34701 6236 34713 6239
rect 34664 6208 34713 6236
rect 34664 6196 34670 6208
rect 34701 6205 34713 6208
rect 34747 6236 34759 6239
rect 35437 6239 35495 6245
rect 35437 6236 35449 6239
rect 34747 6208 35449 6236
rect 34747 6205 34759 6208
rect 34701 6199 34759 6205
rect 35437 6205 35449 6208
rect 35483 6236 35495 6239
rect 36078 6236 36084 6248
rect 35483 6208 36084 6236
rect 35483 6205 35495 6208
rect 35437 6199 35495 6205
rect 36078 6196 36084 6208
rect 36136 6196 36142 6248
rect 21634 6168 21640 6180
rect 18288 6140 18333 6168
rect 19720 6140 20668 6168
rect 21595 6140 21640 6168
rect 18288 6128 18294 6140
rect 19720 6112 19748 6140
rect 14240 6072 14504 6100
rect 14240 6060 14246 6072
rect 15194 6060 15200 6112
rect 15252 6100 15258 6112
rect 15470 6100 15476 6112
rect 15252 6072 15476 6100
rect 15252 6060 15258 6072
rect 15470 6060 15476 6072
rect 15528 6100 15534 6112
rect 15657 6103 15715 6109
rect 15657 6100 15669 6103
rect 15528 6072 15669 6100
rect 15528 6060 15534 6072
rect 15657 6069 15669 6072
rect 15703 6069 15715 6103
rect 19702 6100 19708 6112
rect 19663 6072 19708 6100
rect 15657 6063 15715 6069
rect 19702 6060 19708 6072
rect 19760 6060 19766 6112
rect 20640 6100 20668 6140
rect 21634 6128 21640 6140
rect 21692 6128 21698 6180
rect 25317 6171 25375 6177
rect 25317 6137 25329 6171
rect 25363 6168 25375 6171
rect 25590 6168 25596 6180
rect 25363 6140 25596 6168
rect 25363 6137 25375 6140
rect 25317 6131 25375 6137
rect 25590 6128 25596 6140
rect 25648 6128 25654 6180
rect 27157 6171 27215 6177
rect 27157 6137 27169 6171
rect 27203 6168 27215 6171
rect 27985 6171 28043 6177
rect 27985 6168 27997 6171
rect 27203 6140 27997 6168
rect 27203 6137 27215 6140
rect 27157 6131 27215 6137
rect 27985 6137 27997 6140
rect 28031 6137 28043 6171
rect 27985 6131 28043 6137
rect 21358 6100 21364 6112
rect 20640 6072 21364 6100
rect 21358 6060 21364 6072
rect 21416 6100 21422 6112
rect 21913 6103 21971 6109
rect 21913 6100 21925 6103
rect 21416 6072 21925 6100
rect 21416 6060 21422 6072
rect 21913 6069 21925 6072
rect 21959 6100 21971 6103
rect 22186 6100 22192 6112
rect 21959 6072 22192 6100
rect 21959 6069 21971 6072
rect 21913 6063 21971 6069
rect 22186 6060 22192 6072
rect 22244 6060 22250 6112
rect 23014 6100 23020 6112
rect 22975 6072 23020 6100
rect 23014 6060 23020 6072
rect 23072 6060 23078 6112
rect 23290 6060 23296 6112
rect 23348 6100 23354 6112
rect 23385 6103 23443 6109
rect 23385 6100 23397 6103
rect 23348 6072 23397 6100
rect 23348 6060 23354 6072
rect 23385 6069 23397 6072
rect 23431 6069 23443 6103
rect 24026 6100 24032 6112
rect 23987 6072 24032 6100
rect 23385 6063 23443 6069
rect 24026 6060 24032 6072
rect 24084 6060 24090 6112
rect 24394 6060 24400 6112
rect 24452 6100 24458 6112
rect 27172 6100 27200 6131
rect 24452 6072 27200 6100
rect 24452 6060 24458 6072
rect 31386 6060 31392 6112
rect 31444 6100 31450 6112
rect 31619 6103 31677 6109
rect 31619 6100 31631 6103
rect 31444 6072 31631 6100
rect 31444 6060 31450 6072
rect 31619 6069 31631 6072
rect 31665 6069 31677 6103
rect 31619 6063 31677 6069
rect 1104 6010 38824 6032
rect 1104 5958 14315 6010
rect 14367 5958 14379 6010
rect 14431 5958 14443 6010
rect 14495 5958 14507 6010
rect 14559 5958 27648 6010
rect 27700 5958 27712 6010
rect 27764 5958 27776 6010
rect 27828 5958 27840 6010
rect 27892 5958 38824 6010
rect 1104 5936 38824 5958
rect 3142 5896 3148 5908
rect 3103 5868 3148 5896
rect 3142 5856 3148 5868
rect 3200 5856 3206 5908
rect 3326 5856 3332 5908
rect 3384 5896 3390 5908
rect 3513 5899 3571 5905
rect 3513 5896 3525 5899
rect 3384 5868 3525 5896
rect 3384 5856 3390 5868
rect 3513 5865 3525 5868
rect 3559 5896 3571 5899
rect 5074 5896 5080 5908
rect 3559 5868 5080 5896
rect 3559 5865 3571 5868
rect 3513 5859 3571 5865
rect 5074 5856 5080 5868
rect 5132 5856 5138 5908
rect 6638 5856 6644 5908
rect 6696 5896 6702 5908
rect 6733 5899 6791 5905
rect 6733 5896 6745 5899
rect 6696 5868 6745 5896
rect 6696 5856 6702 5868
rect 6733 5865 6745 5868
rect 6779 5865 6791 5899
rect 7190 5896 7196 5908
rect 7151 5868 7196 5896
rect 6733 5859 6791 5865
rect 7190 5856 7196 5868
rect 7248 5856 7254 5908
rect 9122 5896 9128 5908
rect 9035 5868 9128 5896
rect 9122 5856 9128 5868
rect 9180 5896 9186 5908
rect 9674 5896 9680 5908
rect 9180 5868 9680 5896
rect 9180 5856 9186 5868
rect 9674 5856 9680 5868
rect 9732 5856 9738 5908
rect 12253 5899 12311 5905
rect 12253 5865 12265 5899
rect 12299 5896 12311 5899
rect 12710 5896 12716 5908
rect 12299 5868 12716 5896
rect 12299 5865 12311 5868
rect 12253 5859 12311 5865
rect 12710 5856 12716 5868
rect 12768 5896 12774 5908
rect 13906 5896 13912 5908
rect 12768 5868 13912 5896
rect 12768 5856 12774 5868
rect 13906 5856 13912 5868
rect 13964 5856 13970 5908
rect 14182 5856 14188 5908
rect 14240 5896 14246 5908
rect 14369 5899 14427 5905
rect 14369 5896 14381 5899
rect 14240 5868 14381 5896
rect 14240 5856 14246 5868
rect 14369 5865 14381 5868
rect 14415 5865 14427 5899
rect 17586 5896 17592 5908
rect 17547 5868 17592 5896
rect 14369 5859 14427 5865
rect 17586 5856 17592 5868
rect 17644 5856 17650 5908
rect 18141 5899 18199 5905
rect 18141 5865 18153 5899
rect 18187 5896 18199 5899
rect 18230 5896 18236 5908
rect 18187 5868 18236 5896
rect 18187 5865 18199 5868
rect 18141 5859 18199 5865
rect 18230 5856 18236 5868
rect 18288 5896 18294 5908
rect 18417 5899 18475 5905
rect 18417 5896 18429 5899
rect 18288 5868 18429 5896
rect 18288 5856 18294 5868
rect 18417 5865 18429 5868
rect 18463 5865 18475 5899
rect 18417 5859 18475 5865
rect 19981 5899 20039 5905
rect 19981 5865 19993 5899
rect 20027 5896 20039 5899
rect 20622 5896 20628 5908
rect 20027 5868 20628 5896
rect 20027 5865 20039 5868
rect 19981 5859 20039 5865
rect 20622 5856 20628 5868
rect 20680 5856 20686 5908
rect 24121 5899 24179 5905
rect 24121 5865 24133 5899
rect 24167 5896 24179 5899
rect 24394 5896 24400 5908
rect 24167 5868 24400 5896
rect 24167 5865 24179 5868
rect 24121 5859 24179 5865
rect 24394 5856 24400 5868
rect 24452 5856 24458 5908
rect 24486 5856 24492 5908
rect 24544 5896 24550 5908
rect 24765 5899 24823 5905
rect 24765 5896 24777 5899
rect 24544 5868 24777 5896
rect 24544 5856 24550 5868
rect 24765 5865 24777 5868
rect 24811 5865 24823 5899
rect 24765 5859 24823 5865
rect 25087 5899 25145 5905
rect 25087 5865 25099 5899
rect 25133 5896 25145 5899
rect 26329 5899 26387 5905
rect 26329 5896 26341 5899
rect 25133 5868 26341 5896
rect 25133 5865 25145 5868
rect 25087 5859 25145 5865
rect 26329 5865 26341 5868
rect 26375 5896 26387 5899
rect 26602 5896 26608 5908
rect 26375 5868 26608 5896
rect 26375 5865 26387 5868
rect 26329 5859 26387 5865
rect 26602 5856 26608 5868
rect 26660 5856 26666 5908
rect 27617 5899 27675 5905
rect 27617 5865 27629 5899
rect 27663 5896 27675 5899
rect 27982 5896 27988 5908
rect 27663 5868 27988 5896
rect 27663 5865 27675 5868
rect 27617 5859 27675 5865
rect 27982 5856 27988 5868
rect 28040 5856 28046 5908
rect 2587 5831 2645 5837
rect 2587 5797 2599 5831
rect 2633 5828 2645 5831
rect 2774 5828 2780 5840
rect 2633 5800 2780 5828
rect 2633 5797 2645 5800
rect 2587 5791 2645 5797
rect 2774 5788 2780 5800
rect 2832 5788 2838 5840
rect 3418 5788 3424 5840
rect 3476 5828 3482 5840
rect 3786 5828 3792 5840
rect 3476 5800 3792 5828
rect 3476 5788 3482 5800
rect 3786 5788 3792 5800
rect 3844 5828 3850 5840
rect 5534 5828 5540 5840
rect 3844 5800 5304 5828
rect 5495 5800 5540 5828
rect 3844 5788 3850 5800
rect 2225 5763 2283 5769
rect 2225 5729 2237 5763
rect 2271 5760 2283 5763
rect 3510 5760 3516 5772
rect 2271 5732 3516 5760
rect 2271 5729 2283 5732
rect 2225 5723 2283 5729
rect 3510 5720 3516 5732
rect 3568 5720 3574 5772
rect 4246 5760 4252 5772
rect 4207 5732 4252 5760
rect 4246 5720 4252 5732
rect 4304 5720 4310 5772
rect 4522 5760 4528 5772
rect 4483 5732 4528 5760
rect 4522 5720 4528 5732
rect 4580 5720 4586 5772
rect 5276 5769 5304 5800
rect 5534 5788 5540 5800
rect 5592 5788 5598 5840
rect 6196 5800 8156 5828
rect 6196 5772 6224 5800
rect 5077 5763 5135 5769
rect 5077 5729 5089 5763
rect 5123 5729 5135 5763
rect 5077 5723 5135 5729
rect 5261 5763 5319 5769
rect 5261 5729 5273 5763
rect 5307 5760 5319 5763
rect 6178 5760 6184 5772
rect 5307 5732 6184 5760
rect 5307 5729 5319 5732
rect 5261 5723 5319 5729
rect 1765 5695 1823 5701
rect 1765 5661 1777 5695
rect 1811 5692 1823 5695
rect 2041 5695 2099 5701
rect 2041 5692 2053 5695
rect 1811 5664 2053 5692
rect 1811 5661 1823 5664
rect 1765 5655 1823 5661
rect 2041 5661 2053 5664
rect 2087 5692 2099 5695
rect 3418 5692 3424 5704
rect 2087 5664 3424 5692
rect 2087 5661 2099 5664
rect 2041 5655 2099 5661
rect 3418 5652 3424 5664
rect 3476 5652 3482 5704
rect 5092 5692 5120 5723
rect 6178 5720 6184 5732
rect 6236 5720 6242 5772
rect 7190 5760 7196 5772
rect 7151 5732 7196 5760
rect 7190 5720 7196 5732
rect 7248 5720 7254 5772
rect 7374 5760 7380 5772
rect 7335 5732 7380 5760
rect 7374 5720 7380 5732
rect 7432 5720 7438 5772
rect 8128 5769 8156 5800
rect 10152 5800 10640 5828
rect 7929 5763 7987 5769
rect 7929 5729 7941 5763
rect 7975 5729 7987 5763
rect 7929 5723 7987 5729
rect 8113 5763 8171 5769
rect 8113 5729 8125 5763
rect 8159 5760 8171 5763
rect 9401 5763 9459 5769
rect 9401 5760 9413 5763
rect 8159 5732 9413 5760
rect 8159 5729 8171 5732
rect 8113 5723 8171 5729
rect 9401 5729 9413 5732
rect 9447 5729 9459 5763
rect 9401 5723 9459 5729
rect 9677 5763 9735 5769
rect 9677 5729 9689 5763
rect 9723 5760 9735 5763
rect 10152 5760 10180 5800
rect 10318 5760 10324 5772
rect 9723 5732 10180 5760
rect 10279 5732 10324 5760
rect 9723 5729 9735 5732
rect 9677 5723 9735 5729
rect 5350 5692 5356 5704
rect 5092 5664 5356 5692
rect 3881 5559 3939 5565
rect 3881 5525 3893 5559
rect 3927 5556 3939 5559
rect 5092 5556 5120 5664
rect 5350 5652 5356 5664
rect 5408 5652 5414 5704
rect 7098 5652 7104 5704
rect 7156 5692 7162 5704
rect 7944 5692 7972 5723
rect 8754 5692 8760 5704
rect 7156 5664 8760 5692
rect 7156 5652 7162 5664
rect 8754 5652 8760 5664
rect 8812 5652 8818 5704
rect 9416 5692 9444 5723
rect 10318 5720 10324 5732
rect 10376 5720 10382 5772
rect 10612 5769 10640 5800
rect 10778 5788 10784 5840
rect 10836 5828 10842 5840
rect 11514 5828 11520 5840
rect 10836 5800 11284 5828
rect 11475 5800 11520 5828
rect 10836 5788 10842 5800
rect 10597 5763 10655 5769
rect 10597 5729 10609 5763
rect 10643 5729 10655 5763
rect 10597 5723 10655 5729
rect 10612 5692 10640 5723
rect 10686 5720 10692 5772
rect 10744 5760 10750 5772
rect 11256 5769 11284 5800
rect 11514 5788 11520 5800
rect 11572 5788 11578 5840
rect 13078 5788 13084 5840
rect 13136 5828 13142 5840
rect 13770 5831 13828 5837
rect 13770 5828 13782 5831
rect 13136 5800 13782 5828
rect 13136 5788 13142 5800
rect 13770 5797 13782 5800
rect 13816 5797 13828 5831
rect 13770 5791 13828 5797
rect 15105 5831 15163 5837
rect 15105 5797 15117 5831
rect 15151 5828 15163 5831
rect 15562 5828 15568 5840
rect 15151 5800 15568 5828
rect 15151 5797 15163 5800
rect 15105 5791 15163 5797
rect 15562 5788 15568 5800
rect 15620 5828 15626 5840
rect 15749 5831 15807 5837
rect 15749 5828 15761 5831
rect 15620 5800 15761 5828
rect 15620 5788 15626 5800
rect 15749 5797 15761 5800
rect 15795 5797 15807 5831
rect 15749 5791 15807 5797
rect 15838 5788 15844 5840
rect 15896 5828 15902 5840
rect 16393 5831 16451 5837
rect 15896 5800 15941 5828
rect 15896 5788 15902 5800
rect 16393 5797 16405 5831
rect 16439 5828 16451 5831
rect 16850 5828 16856 5840
rect 16439 5800 16856 5828
rect 16439 5797 16451 5800
rect 16393 5791 16451 5797
rect 16850 5788 16856 5800
rect 16908 5788 16914 5840
rect 17604 5828 17632 5856
rect 23014 5828 23020 5840
rect 17604 5800 23020 5828
rect 23014 5788 23020 5800
rect 23072 5828 23078 5840
rect 23522 5831 23580 5837
rect 23522 5828 23534 5831
rect 23072 5800 23534 5828
rect 23072 5788 23078 5800
rect 23522 5797 23534 5800
rect 23568 5797 23580 5831
rect 23522 5791 23580 5797
rect 25590 5788 25596 5840
rect 25648 5828 25654 5840
rect 26697 5831 26755 5837
rect 26697 5828 26709 5831
rect 25648 5800 26709 5828
rect 25648 5788 25654 5800
rect 26697 5797 26709 5800
rect 26743 5828 26755 5831
rect 26970 5828 26976 5840
rect 26743 5800 26976 5828
rect 26743 5797 26755 5800
rect 26697 5791 26755 5797
rect 26970 5788 26976 5800
rect 27028 5788 27034 5840
rect 10873 5763 10931 5769
rect 10873 5760 10885 5763
rect 10744 5732 10885 5760
rect 10744 5720 10750 5732
rect 10873 5729 10885 5732
rect 10919 5729 10931 5763
rect 10873 5723 10931 5729
rect 11241 5763 11299 5769
rect 11241 5729 11253 5763
rect 11287 5729 11299 5763
rect 11241 5723 11299 5729
rect 12250 5720 12256 5772
rect 12308 5760 12314 5772
rect 12380 5763 12438 5769
rect 12380 5760 12392 5763
rect 12308 5732 12392 5760
rect 12308 5720 12314 5732
rect 12380 5729 12392 5732
rect 12426 5729 12438 5763
rect 16758 5760 16764 5772
rect 16671 5732 16764 5760
rect 12380 5723 12438 5729
rect 16758 5720 16764 5732
rect 16816 5760 16822 5772
rect 18138 5760 18144 5772
rect 16816 5732 18144 5760
rect 16816 5720 16822 5732
rect 18138 5720 18144 5732
rect 18196 5720 18202 5772
rect 19794 5760 19800 5772
rect 19755 5732 19800 5760
rect 19794 5720 19800 5732
rect 19852 5720 19858 5772
rect 20438 5720 20444 5772
rect 20496 5760 20502 5772
rect 20901 5763 20959 5769
rect 20901 5760 20913 5763
rect 20496 5732 20913 5760
rect 20496 5720 20502 5732
rect 20901 5729 20913 5732
rect 20947 5729 20959 5763
rect 20901 5723 20959 5729
rect 21361 5763 21419 5769
rect 21361 5729 21373 5763
rect 21407 5729 21419 5763
rect 21910 5760 21916 5772
rect 21871 5732 21916 5760
rect 21361 5723 21419 5729
rect 9416 5664 9812 5692
rect 10612 5664 10916 5692
rect 6638 5584 6644 5636
rect 6696 5624 6702 5636
rect 7374 5624 7380 5636
rect 6696 5596 7380 5624
rect 6696 5584 6702 5596
rect 7374 5584 7380 5596
rect 7432 5624 7438 5636
rect 9677 5627 9735 5633
rect 9677 5624 9689 5627
rect 7432 5596 9689 5624
rect 7432 5584 7438 5596
rect 9677 5593 9689 5596
rect 9723 5593 9735 5627
rect 9784 5624 9812 5664
rect 10778 5624 10784 5636
rect 9784 5596 10784 5624
rect 9677 5587 9735 5593
rect 10778 5584 10784 5596
rect 10836 5584 10842 5636
rect 10888 5624 10916 5664
rect 10962 5652 10968 5704
rect 11020 5692 11026 5704
rect 13262 5692 13268 5704
rect 11020 5664 13268 5692
rect 11020 5652 11026 5664
rect 13262 5652 13268 5664
rect 13320 5692 13326 5704
rect 13449 5695 13507 5701
rect 13449 5692 13461 5695
rect 13320 5664 13461 5692
rect 13320 5652 13326 5664
rect 13449 5661 13461 5664
rect 13495 5661 13507 5695
rect 13449 5655 13507 5661
rect 17221 5695 17279 5701
rect 17221 5661 17233 5695
rect 17267 5661 17279 5695
rect 17221 5655 17279 5661
rect 11790 5624 11796 5636
rect 10888 5596 11796 5624
rect 11790 5584 11796 5596
rect 11848 5584 11854 5636
rect 12483 5627 12541 5633
rect 12483 5593 12495 5627
rect 12529 5624 12541 5627
rect 12986 5624 12992 5636
rect 12529 5596 12992 5624
rect 12529 5593 12541 5596
rect 12483 5587 12541 5593
rect 12986 5584 12992 5596
rect 13044 5624 13050 5636
rect 13173 5627 13231 5633
rect 13173 5624 13185 5627
rect 13044 5596 13185 5624
rect 13044 5584 13050 5596
rect 13173 5593 13185 5596
rect 13219 5593 13231 5627
rect 13173 5587 13231 5593
rect 3927 5528 5120 5556
rect 3927 5525 3939 5528
rect 3881 5519 3939 5525
rect 5534 5516 5540 5568
rect 5592 5556 5598 5568
rect 5813 5559 5871 5565
rect 5813 5556 5825 5559
rect 5592 5528 5825 5556
rect 5592 5516 5598 5528
rect 5813 5525 5825 5528
rect 5859 5525 5871 5559
rect 6454 5556 6460 5568
rect 6415 5528 6460 5556
rect 5813 5519 5871 5525
rect 6454 5516 6460 5528
rect 6512 5516 6518 5568
rect 9953 5559 10011 5565
rect 9953 5525 9965 5559
rect 9999 5556 10011 5559
rect 10226 5556 10232 5568
rect 9999 5528 10232 5556
rect 9999 5525 10011 5528
rect 9953 5519 10011 5525
rect 10226 5516 10232 5528
rect 10284 5516 10290 5568
rect 11882 5556 11888 5568
rect 11843 5528 11888 5556
rect 11882 5516 11888 5528
rect 11940 5516 11946 5568
rect 12802 5556 12808 5568
rect 12763 5528 12808 5556
rect 12802 5516 12808 5528
rect 12860 5516 12866 5568
rect 14642 5556 14648 5568
rect 14603 5528 14648 5556
rect 14642 5516 14648 5528
rect 14700 5516 14706 5568
rect 15378 5516 15384 5568
rect 15436 5556 15442 5568
rect 15473 5559 15531 5565
rect 15473 5556 15485 5559
rect 15436 5528 15485 5556
rect 15436 5516 15442 5528
rect 15473 5525 15485 5528
rect 15519 5525 15531 5559
rect 17126 5556 17132 5568
rect 17087 5528 17132 5556
rect 15473 5519 15531 5525
rect 17126 5516 17132 5528
rect 17184 5556 17190 5568
rect 17236 5556 17264 5655
rect 20622 5652 20628 5704
rect 20680 5692 20686 5704
rect 21376 5692 21404 5723
rect 21910 5720 21916 5732
rect 21968 5720 21974 5772
rect 22094 5760 22100 5772
rect 22055 5732 22100 5760
rect 22094 5720 22100 5732
rect 22152 5720 22158 5772
rect 25016 5763 25074 5769
rect 25016 5729 25028 5763
rect 25062 5760 25074 5763
rect 25498 5760 25504 5772
rect 25062 5732 25504 5760
rect 25062 5729 25074 5732
rect 25016 5723 25074 5729
rect 25498 5720 25504 5732
rect 25556 5720 25562 5772
rect 20680 5664 21404 5692
rect 22373 5695 22431 5701
rect 20680 5652 20686 5664
rect 22373 5661 22385 5695
rect 22419 5692 22431 5695
rect 23198 5692 23204 5704
rect 22419 5664 23204 5692
rect 22419 5661 22431 5664
rect 22373 5655 22431 5661
rect 23198 5652 23204 5664
rect 23256 5652 23262 5704
rect 25130 5652 25136 5704
rect 25188 5692 25194 5704
rect 25409 5695 25467 5701
rect 25409 5692 25421 5695
rect 25188 5664 25421 5692
rect 25188 5652 25194 5664
rect 25409 5661 25421 5664
rect 25455 5661 25467 5695
rect 26602 5692 26608 5704
rect 26563 5664 26608 5692
rect 25409 5655 25467 5661
rect 26602 5652 26608 5664
rect 26660 5652 26666 5704
rect 26881 5695 26939 5701
rect 26881 5661 26893 5695
rect 26927 5661 26939 5695
rect 26881 5655 26939 5661
rect 26050 5584 26056 5636
rect 26108 5624 26114 5636
rect 26896 5624 26924 5655
rect 26108 5596 26924 5624
rect 26108 5584 26114 5596
rect 17184 5528 17264 5556
rect 17184 5516 17190 5528
rect 19518 5516 19524 5568
rect 19576 5556 19582 5568
rect 20257 5559 20315 5565
rect 20257 5556 20269 5559
rect 19576 5528 20269 5556
rect 19576 5516 19582 5528
rect 20257 5525 20269 5528
rect 20303 5525 20315 5559
rect 20257 5519 20315 5525
rect 1104 5466 38824 5488
rect 1104 5414 7648 5466
rect 7700 5414 7712 5466
rect 7764 5414 7776 5466
rect 7828 5414 7840 5466
rect 7892 5414 20982 5466
rect 21034 5414 21046 5466
rect 21098 5414 21110 5466
rect 21162 5414 21174 5466
rect 21226 5414 34315 5466
rect 34367 5414 34379 5466
rect 34431 5414 34443 5466
rect 34495 5414 34507 5466
rect 34559 5414 38824 5466
rect 1104 5392 38824 5414
rect 1026 5312 1032 5364
rect 1084 5352 1090 5364
rect 1581 5355 1639 5361
rect 1581 5352 1593 5355
rect 1084 5324 1593 5352
rect 1084 5312 1090 5324
rect 1581 5321 1593 5324
rect 1627 5321 1639 5355
rect 6178 5352 6184 5364
rect 6139 5324 6184 5352
rect 1581 5315 1639 5321
rect 6178 5312 6184 5324
rect 6236 5352 6242 5364
rect 6549 5355 6607 5361
rect 6549 5352 6561 5355
rect 6236 5324 6561 5352
rect 6236 5312 6242 5324
rect 6549 5321 6561 5324
rect 6595 5321 6607 5355
rect 7098 5352 7104 5364
rect 7059 5324 7104 5352
rect 6549 5315 6607 5321
rect 7098 5312 7104 5324
rect 7156 5312 7162 5364
rect 12250 5352 12256 5364
rect 12211 5324 12256 5352
rect 12250 5312 12256 5324
rect 12308 5312 12314 5364
rect 13078 5312 13084 5364
rect 13136 5352 13142 5364
rect 13633 5355 13691 5361
rect 13633 5352 13645 5355
rect 13136 5324 13645 5352
rect 13136 5312 13142 5324
rect 13633 5321 13645 5324
rect 13679 5352 13691 5355
rect 13814 5352 13820 5364
rect 13679 5324 13820 5352
rect 13679 5321 13691 5324
rect 13633 5315 13691 5321
rect 13814 5312 13820 5324
rect 13872 5352 13878 5364
rect 14185 5355 14243 5361
rect 14185 5352 14197 5355
rect 13872 5324 14197 5352
rect 13872 5312 13878 5324
rect 14185 5321 14197 5324
rect 14231 5321 14243 5355
rect 15194 5352 15200 5364
rect 15155 5324 15200 5352
rect 14185 5315 14243 5321
rect 15194 5312 15200 5324
rect 15252 5312 15258 5364
rect 16298 5312 16304 5364
rect 16356 5352 16362 5364
rect 17405 5355 17463 5361
rect 17405 5352 17417 5355
rect 16356 5324 17417 5352
rect 16356 5312 16362 5324
rect 17405 5321 17417 5324
rect 17451 5352 17463 5355
rect 17586 5352 17592 5364
rect 17451 5324 17592 5352
rect 17451 5321 17463 5324
rect 17405 5315 17463 5321
rect 17586 5312 17592 5324
rect 17644 5312 17650 5364
rect 22186 5352 22192 5364
rect 22147 5324 22192 5352
rect 22186 5312 22192 5324
rect 22244 5312 22250 5364
rect 23014 5312 23020 5364
rect 23072 5352 23078 5364
rect 23201 5355 23259 5361
rect 23201 5352 23213 5355
rect 23072 5324 23213 5352
rect 23072 5312 23078 5324
rect 23201 5321 23213 5324
rect 23247 5352 23259 5355
rect 24026 5352 24032 5364
rect 23247 5324 24032 5352
rect 23247 5321 23259 5324
rect 23201 5315 23259 5321
rect 24026 5312 24032 5324
rect 24084 5312 24090 5364
rect 25133 5355 25191 5361
rect 25133 5321 25145 5355
rect 25179 5352 25191 5355
rect 25590 5352 25596 5364
rect 25179 5324 25596 5352
rect 25179 5321 25191 5324
rect 25133 5315 25191 5321
rect 25590 5312 25596 5324
rect 25648 5312 25654 5364
rect 26602 5312 26608 5364
rect 26660 5352 26666 5364
rect 27341 5355 27399 5361
rect 27341 5352 27353 5355
rect 26660 5324 27353 5352
rect 26660 5312 26666 5324
rect 27341 5321 27353 5324
rect 27387 5352 27399 5355
rect 27430 5352 27436 5364
rect 27387 5324 27436 5352
rect 27387 5321 27399 5324
rect 27341 5315 27399 5321
rect 27430 5312 27436 5324
rect 27488 5312 27494 5364
rect 5074 5244 5080 5296
rect 5132 5284 5138 5296
rect 10042 5284 10048 5296
rect 5132 5256 10048 5284
rect 5132 5244 5138 5256
rect 10042 5244 10048 5256
rect 10100 5284 10106 5296
rect 11333 5287 11391 5293
rect 11333 5284 11345 5287
rect 10100 5256 11345 5284
rect 10100 5244 10106 5256
rect 11333 5253 11345 5256
rect 11379 5253 11391 5287
rect 11333 5247 11391 5253
rect 14090 5244 14096 5296
rect 14148 5284 14154 5296
rect 19889 5287 19947 5293
rect 19889 5284 19901 5287
rect 14148 5256 19901 5284
rect 14148 5244 14154 5256
rect 19889 5253 19901 5256
rect 19935 5253 19947 5287
rect 19889 5247 19947 5253
rect 3326 5216 3332 5228
rect 3068 5188 3332 5216
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5148 1455 5151
rect 2038 5148 2044 5160
rect 1443 5120 2044 5148
rect 1443 5117 1455 5120
rect 1397 5111 1455 5117
rect 2038 5108 2044 5120
rect 2096 5108 2102 5160
rect 2866 5148 2872 5160
rect 2827 5120 2872 5148
rect 2866 5108 2872 5120
rect 2924 5108 2930 5160
rect 3068 5157 3096 5188
rect 3326 5176 3332 5188
rect 3384 5176 3390 5228
rect 4062 5216 4068 5228
rect 4023 5188 4068 5216
rect 4062 5176 4068 5188
rect 4120 5176 4126 5228
rect 5000 5188 8800 5216
rect 3053 5151 3111 5157
rect 3053 5117 3065 5151
rect 3099 5117 3111 5151
rect 3053 5111 3111 5117
rect 3142 5108 3148 5160
rect 3200 5148 3206 5160
rect 3421 5151 3479 5157
rect 3421 5148 3433 5151
rect 3200 5120 3433 5148
rect 3200 5108 3206 5120
rect 3421 5117 3433 5120
rect 3467 5117 3479 5151
rect 3786 5148 3792 5160
rect 3747 5120 3792 5148
rect 3421 5111 3479 5117
rect 3786 5108 3792 5120
rect 3844 5108 3850 5160
rect 2884 5080 2912 5108
rect 5000 5080 5028 5188
rect 5077 5151 5135 5157
rect 5077 5117 5089 5151
rect 5123 5148 5135 5151
rect 5626 5148 5632 5160
rect 5123 5120 5632 5148
rect 5123 5117 5135 5120
rect 5077 5111 5135 5117
rect 5626 5108 5632 5120
rect 5684 5148 5690 5160
rect 7466 5148 7472 5160
rect 5684 5120 7328 5148
rect 7379 5120 7472 5148
rect 5684 5108 5690 5120
rect 5902 5080 5908 5092
rect 2884 5052 5028 5080
rect 5863 5052 5908 5080
rect 5902 5040 5908 5052
rect 5960 5040 5966 5092
rect 7300 5080 7328 5120
rect 7466 5108 7472 5120
rect 7524 5148 7530 5160
rect 8772 5157 8800 5188
rect 8938 5176 8944 5228
rect 8996 5216 9002 5228
rect 9309 5219 9367 5225
rect 9309 5216 9321 5219
rect 8996 5188 9321 5216
rect 8996 5176 9002 5188
rect 9309 5185 9321 5188
rect 9355 5216 9367 5219
rect 9401 5219 9459 5225
rect 9401 5216 9413 5219
rect 9355 5188 9413 5216
rect 9355 5185 9367 5188
rect 9309 5179 9367 5185
rect 9401 5185 9413 5188
rect 9447 5185 9459 5219
rect 11054 5216 11060 5228
rect 11015 5188 11060 5216
rect 9401 5179 9459 5185
rect 11054 5176 11060 5188
rect 11112 5176 11118 5228
rect 12710 5216 12716 5228
rect 12671 5188 12716 5216
rect 12710 5176 12716 5188
rect 12768 5176 12774 5228
rect 13170 5216 13176 5228
rect 13131 5188 13176 5216
rect 13170 5176 13176 5188
rect 13228 5176 13234 5228
rect 15749 5219 15807 5225
rect 15749 5185 15761 5219
rect 15795 5216 15807 5219
rect 15838 5216 15844 5228
rect 15795 5188 15844 5216
rect 15795 5185 15807 5188
rect 15749 5179 15807 5185
rect 15838 5176 15844 5188
rect 15896 5216 15902 5228
rect 15896 5188 17172 5216
rect 15896 5176 15902 5188
rect 7653 5151 7711 5157
rect 7653 5148 7665 5151
rect 7524 5120 7665 5148
rect 7524 5108 7530 5120
rect 7653 5117 7665 5120
rect 7699 5117 7711 5151
rect 7653 5111 7711 5117
rect 8757 5151 8815 5157
rect 8757 5117 8769 5151
rect 8803 5148 8815 5151
rect 9858 5148 9864 5160
rect 8803 5120 9864 5148
rect 8803 5117 8815 5120
rect 8757 5111 8815 5117
rect 9858 5108 9864 5120
rect 9916 5108 9922 5160
rect 10042 5148 10048 5160
rect 10003 5120 10048 5148
rect 10042 5108 10048 5120
rect 10100 5108 10106 5160
rect 10134 5108 10140 5160
rect 10192 5148 10198 5160
rect 10413 5151 10471 5157
rect 10413 5148 10425 5151
rect 10192 5120 10425 5148
rect 10192 5108 10198 5120
rect 10413 5117 10425 5120
rect 10459 5117 10471 5151
rect 10778 5148 10784 5160
rect 10739 5120 10784 5148
rect 10413 5111 10471 5117
rect 10778 5108 10784 5120
rect 10836 5148 10842 5160
rect 11701 5151 11759 5157
rect 11701 5148 11713 5151
rect 10836 5120 11713 5148
rect 10836 5108 10842 5120
rect 11701 5117 11713 5120
rect 11747 5117 11759 5151
rect 11701 5111 11759 5117
rect 13722 5108 13728 5160
rect 13780 5148 13786 5160
rect 14277 5151 14335 5157
rect 14277 5148 14289 5151
rect 13780 5120 14289 5148
rect 13780 5108 13786 5120
rect 14277 5117 14289 5120
rect 14323 5117 14335 5151
rect 14277 5111 14335 5117
rect 16209 5151 16267 5157
rect 16209 5117 16221 5151
rect 16255 5148 16267 5151
rect 16758 5148 16764 5160
rect 16255 5120 16764 5148
rect 16255 5117 16267 5120
rect 16209 5111 16267 5117
rect 16758 5108 16764 5120
rect 16816 5108 16822 5160
rect 17144 5157 17172 5188
rect 17218 5176 17224 5228
rect 17276 5216 17282 5228
rect 18049 5219 18107 5225
rect 18049 5216 18061 5219
rect 17276 5188 18061 5216
rect 17276 5176 17282 5188
rect 18049 5185 18061 5188
rect 18095 5185 18107 5219
rect 18049 5179 18107 5185
rect 17129 5151 17187 5157
rect 17129 5117 17141 5151
rect 17175 5148 17187 5151
rect 17865 5151 17923 5157
rect 17865 5148 17877 5151
rect 17175 5120 17877 5148
rect 17175 5117 17187 5120
rect 17129 5111 17187 5117
rect 17865 5117 17877 5120
rect 17911 5148 17923 5151
rect 18141 5151 18199 5157
rect 18141 5148 18153 5151
rect 17911 5120 18153 5148
rect 17911 5117 17923 5120
rect 17865 5111 17923 5117
rect 18141 5117 18153 5120
rect 18187 5117 18199 5151
rect 19904 5148 19932 5247
rect 20438 5244 20444 5296
rect 20496 5284 20502 5296
rect 21821 5287 21879 5293
rect 21821 5284 21833 5287
rect 20496 5256 21833 5284
rect 20496 5244 20502 5256
rect 21821 5253 21833 5256
rect 21867 5253 21879 5287
rect 26970 5284 26976 5296
rect 26931 5256 26976 5284
rect 21821 5247 21879 5253
rect 26970 5244 26976 5256
rect 27028 5244 27034 5296
rect 21634 5176 21640 5228
rect 21692 5216 21698 5228
rect 24210 5216 24216 5228
rect 21692 5188 24216 5216
rect 21692 5176 21698 5188
rect 24210 5176 24216 5188
rect 24268 5176 24274 5228
rect 26050 5216 26056 5228
rect 26011 5188 26056 5216
rect 26050 5176 26056 5188
rect 26108 5176 26114 5228
rect 20073 5151 20131 5157
rect 20073 5148 20085 5151
rect 19904 5120 20085 5148
rect 18141 5111 18199 5117
rect 20073 5117 20085 5120
rect 20119 5148 20131 5151
rect 20438 5148 20444 5160
rect 20119 5120 20444 5148
rect 20119 5117 20131 5120
rect 20073 5111 20131 5117
rect 20438 5108 20444 5120
rect 20496 5108 20502 5160
rect 20622 5148 20628 5160
rect 20583 5120 20628 5148
rect 20622 5108 20628 5120
rect 20680 5108 20686 5160
rect 20901 5151 20959 5157
rect 20901 5117 20913 5151
rect 20947 5117 20959 5151
rect 20901 5111 20959 5117
rect 21453 5151 21511 5157
rect 21453 5117 21465 5151
rect 21499 5148 21511 5151
rect 22094 5148 22100 5160
rect 21499 5120 22100 5148
rect 21499 5117 21511 5120
rect 21453 5111 21511 5117
rect 8110 5080 8116 5092
rect 7300 5052 8116 5080
rect 8110 5040 8116 5052
rect 8168 5040 8174 5092
rect 8294 5080 8300 5092
rect 8255 5052 8300 5080
rect 8294 5040 8300 5052
rect 8352 5040 8358 5092
rect 9309 5083 9367 5089
rect 9309 5049 9321 5083
rect 9355 5080 9367 5083
rect 10686 5080 10692 5092
rect 9355 5052 10692 5080
rect 9355 5049 9367 5052
rect 9309 5043 9367 5049
rect 10686 5040 10692 5052
rect 10744 5040 10750 5092
rect 12802 5040 12808 5092
rect 12860 5080 12866 5092
rect 12860 5052 12905 5080
rect 12860 5040 12866 5052
rect 13814 5040 13820 5092
rect 13872 5080 13878 5092
rect 14598 5083 14656 5089
rect 14598 5080 14610 5083
rect 13872 5052 14610 5080
rect 13872 5040 13878 5052
rect 14598 5049 14610 5052
rect 14644 5080 14656 5083
rect 16025 5083 16083 5089
rect 16025 5080 16037 5083
rect 14644 5052 16037 5080
rect 14644 5049 14656 5052
rect 14598 5043 14656 5049
rect 16025 5049 16037 5052
rect 16071 5080 16083 5083
rect 16298 5080 16304 5092
rect 16071 5052 16304 5080
rect 16071 5049 16083 5052
rect 16025 5043 16083 5049
rect 16298 5040 16304 5052
rect 16356 5080 16362 5092
rect 16530 5083 16588 5089
rect 16530 5080 16542 5083
rect 16356 5052 16542 5080
rect 16356 5040 16362 5052
rect 16530 5049 16542 5052
rect 16576 5049 16588 5083
rect 16530 5043 16588 5049
rect 16850 5040 16856 5092
rect 16908 5080 16914 5092
rect 19153 5083 19211 5089
rect 19153 5080 19165 5083
rect 16908 5052 19165 5080
rect 16908 5040 16914 5052
rect 19153 5049 19165 5052
rect 19199 5080 19211 5083
rect 19794 5080 19800 5092
rect 19199 5052 19800 5080
rect 19199 5049 19211 5052
rect 19153 5043 19211 5049
rect 19794 5040 19800 5052
rect 19852 5040 19858 5092
rect 2038 5012 2044 5024
rect 1999 4984 2044 5012
rect 2038 4972 2044 4984
rect 2096 4972 2102 5024
rect 2409 5015 2467 5021
rect 2409 4981 2421 5015
rect 2455 5012 2467 5015
rect 2774 5012 2780 5024
rect 2455 4984 2780 5012
rect 2455 4981 2467 4984
rect 2409 4975 2467 4981
rect 2774 4972 2780 4984
rect 2832 4972 2838 5024
rect 4246 4972 4252 5024
rect 4304 5012 4310 5024
rect 4341 5015 4399 5021
rect 4341 5012 4353 5015
rect 4304 4984 4353 5012
rect 4304 4972 4310 4984
rect 4341 4981 4353 4984
rect 4387 4981 4399 5015
rect 4341 4975 4399 4981
rect 8754 4972 8760 5024
rect 8812 5012 8818 5024
rect 9033 5015 9091 5021
rect 9033 5012 9045 5015
rect 8812 4984 9045 5012
rect 8812 4972 8818 4984
rect 9033 4981 9045 4984
rect 9079 4981 9091 5015
rect 19518 5012 19524 5024
rect 19479 4984 19524 5012
rect 9033 4975 9091 4981
rect 19518 4972 19524 4984
rect 19576 5012 19582 5024
rect 20916 5012 20944 5111
rect 22094 5108 22100 5120
rect 22152 5148 22158 5160
rect 22557 5151 22615 5157
rect 22557 5148 22569 5151
rect 22152 5120 22569 5148
rect 22152 5108 22158 5120
rect 22557 5117 22569 5120
rect 22603 5117 22615 5151
rect 22557 5111 22615 5117
rect 24026 5108 24032 5160
rect 24084 5148 24090 5160
rect 24084 5120 24577 5148
rect 24084 5108 24090 5120
rect 21545 5083 21603 5089
rect 21545 5049 21557 5083
rect 21591 5080 21603 5083
rect 24394 5080 24400 5092
rect 21591 5052 24400 5080
rect 21591 5049 21603 5052
rect 21545 5043 21603 5049
rect 24394 5040 24400 5052
rect 24452 5040 24458 5092
rect 24549 5089 24577 5120
rect 24534 5083 24592 5089
rect 24534 5049 24546 5083
rect 24580 5080 24592 5083
rect 24762 5080 24768 5092
rect 24580 5052 24768 5080
rect 24580 5049 24592 5052
rect 24534 5043 24592 5049
rect 24762 5040 24768 5052
rect 24820 5040 24826 5092
rect 26145 5083 26203 5089
rect 26145 5049 26157 5083
rect 26191 5049 26203 5083
rect 26145 5043 26203 5049
rect 26697 5083 26755 5089
rect 26697 5049 26709 5083
rect 26743 5080 26755 5083
rect 26878 5080 26884 5092
rect 26743 5052 26884 5080
rect 26743 5049 26755 5052
rect 26697 5043 26755 5049
rect 21266 5012 21272 5024
rect 19576 4984 21272 5012
rect 19576 4972 19582 4984
rect 21266 4972 21272 4984
rect 21324 4972 21330 5024
rect 25498 5012 25504 5024
rect 25459 4984 25504 5012
rect 25498 4972 25504 4984
rect 25556 4972 25562 5024
rect 25774 5012 25780 5024
rect 25735 4984 25780 5012
rect 25774 4972 25780 4984
rect 25832 5012 25838 5024
rect 26160 5012 26188 5043
rect 26878 5040 26884 5052
rect 26936 5040 26942 5092
rect 25832 4984 26188 5012
rect 25832 4972 25838 4984
rect 1104 4922 38824 4944
rect 1104 4870 14315 4922
rect 14367 4870 14379 4922
rect 14431 4870 14443 4922
rect 14495 4870 14507 4922
rect 14559 4870 27648 4922
rect 27700 4870 27712 4922
rect 27764 4870 27776 4922
rect 27828 4870 27840 4922
rect 27892 4870 38824 4922
rect 1104 4848 38824 4870
rect 1670 4808 1676 4820
rect 1631 4780 1676 4808
rect 1670 4768 1676 4780
rect 1728 4768 1734 4820
rect 2866 4768 2872 4820
rect 2924 4808 2930 4820
rect 3421 4811 3479 4817
rect 3421 4808 3433 4811
rect 2924 4780 3433 4808
rect 2924 4768 2930 4780
rect 3421 4777 3433 4780
rect 3467 4808 3479 4811
rect 3510 4808 3516 4820
rect 3467 4780 3516 4808
rect 3467 4777 3479 4780
rect 3421 4771 3479 4777
rect 3510 4768 3516 4780
rect 3568 4768 3574 4820
rect 7190 4808 7196 4820
rect 7151 4780 7196 4808
rect 7190 4768 7196 4780
rect 7248 4808 7254 4820
rect 8849 4811 8907 4817
rect 8849 4808 8861 4811
rect 7248 4780 8861 4808
rect 7248 4768 7254 4780
rect 8849 4777 8861 4780
rect 8895 4777 8907 4811
rect 8849 4771 8907 4777
rect 9582 4768 9588 4820
rect 9640 4808 9646 4820
rect 12253 4811 12311 4817
rect 12253 4808 12265 4811
rect 9640 4780 12265 4808
rect 9640 4768 9646 4780
rect 12253 4777 12265 4780
rect 12299 4777 12311 4811
rect 13262 4808 13268 4820
rect 13223 4780 13268 4808
rect 12253 4771 12311 4777
rect 13262 4768 13268 4780
rect 13320 4768 13326 4820
rect 13814 4808 13820 4820
rect 13775 4780 13820 4808
rect 13814 4768 13820 4780
rect 13872 4768 13878 4820
rect 14369 4811 14427 4817
rect 14369 4777 14381 4811
rect 14415 4808 14427 4811
rect 15010 4808 15016 4820
rect 14415 4780 15016 4808
rect 14415 4777 14427 4780
rect 14369 4771 14427 4777
rect 15010 4768 15016 4780
rect 15068 4808 15074 4820
rect 17034 4808 17040 4820
rect 15068 4780 15516 4808
rect 16995 4780 17040 4808
rect 15068 4768 15074 4780
rect 7098 4740 7104 4752
rect 1964 4712 3004 4740
rect 1964 4684 1992 4712
rect 1946 4672 1952 4684
rect 1907 4644 1952 4672
rect 1946 4632 1952 4644
rect 2004 4632 2010 4684
rect 2498 4632 2504 4684
rect 2556 4672 2562 4684
rect 2866 4672 2872 4684
rect 2556 4644 2872 4672
rect 2556 4632 2562 4644
rect 2866 4632 2872 4644
rect 2924 4632 2930 4684
rect 2976 4681 3004 4712
rect 5644 4712 7104 4740
rect 2961 4675 3019 4681
rect 2961 4641 2973 4675
rect 3007 4672 3019 4675
rect 3694 4672 3700 4684
rect 3007 4644 3700 4672
rect 3007 4641 3019 4644
rect 2961 4635 3019 4641
rect 3694 4632 3700 4644
rect 3752 4632 3758 4684
rect 4617 4675 4675 4681
rect 4617 4672 4629 4675
rect 4264 4644 4629 4672
rect 4264 4548 4292 4644
rect 4617 4641 4629 4644
rect 4663 4641 4675 4675
rect 5074 4672 5080 4684
rect 5035 4644 5080 4672
rect 4617 4635 4675 4641
rect 5074 4632 5080 4644
rect 5132 4632 5138 4684
rect 5350 4632 5356 4684
rect 5408 4672 5414 4684
rect 5644 4681 5672 4712
rect 7098 4700 7104 4712
rect 7156 4700 7162 4752
rect 9033 4743 9091 4749
rect 9033 4740 9045 4743
rect 7392 4712 9045 4740
rect 5629 4675 5687 4681
rect 5629 4672 5641 4675
rect 5408 4644 5641 4672
rect 5408 4632 5414 4644
rect 5629 4641 5641 4644
rect 5675 4641 5687 4675
rect 5629 4635 5687 4641
rect 5718 4632 5724 4684
rect 5776 4672 5782 4684
rect 5813 4675 5871 4681
rect 5813 4672 5825 4675
rect 5776 4644 5825 4672
rect 5776 4632 5782 4644
rect 5813 4641 5825 4644
rect 5859 4672 5871 4675
rect 7006 4672 7012 4684
rect 5859 4644 7012 4672
rect 5859 4641 5871 4644
rect 5813 4635 5871 4641
rect 7006 4632 7012 4644
rect 7064 4672 7070 4684
rect 7392 4672 7420 4712
rect 9033 4709 9045 4712
rect 9079 4740 9091 4743
rect 9401 4743 9459 4749
rect 9401 4740 9413 4743
rect 9079 4712 9413 4740
rect 9079 4709 9091 4712
rect 9033 4703 9091 4709
rect 9401 4709 9413 4712
rect 9447 4740 9459 4743
rect 10226 4740 10232 4752
rect 9447 4712 10232 4740
rect 9447 4709 9459 4712
rect 9401 4703 9459 4709
rect 10226 4700 10232 4712
rect 10284 4740 10290 4752
rect 11149 4743 11207 4749
rect 10284 4712 10916 4740
rect 10284 4700 10290 4712
rect 7064 4644 7420 4672
rect 7469 4675 7527 4681
rect 7064 4632 7070 4644
rect 7469 4641 7481 4675
rect 7515 4672 7527 4675
rect 8018 4672 8024 4684
rect 7515 4644 8024 4672
rect 7515 4641 7527 4644
rect 7469 4635 7527 4641
rect 8018 4632 8024 4644
rect 8076 4632 8082 4684
rect 9950 4672 9956 4684
rect 9911 4644 9956 4672
rect 9950 4632 9956 4644
rect 10008 4632 10014 4684
rect 10042 4632 10048 4684
rect 10100 4672 10106 4684
rect 10137 4675 10195 4681
rect 10137 4672 10149 4675
rect 10100 4644 10149 4672
rect 10100 4632 10106 4644
rect 10137 4641 10149 4644
rect 10183 4641 10195 4675
rect 10686 4672 10692 4684
rect 10647 4644 10692 4672
rect 10137 4635 10195 4641
rect 10686 4632 10692 4644
rect 10744 4632 10750 4684
rect 10888 4681 10916 4712
rect 11149 4709 11161 4743
rect 11195 4740 11207 4743
rect 13722 4740 13728 4752
rect 11195 4712 13728 4740
rect 11195 4709 11207 4712
rect 11149 4703 11207 4709
rect 13722 4700 13728 4712
rect 13780 4740 13786 4752
rect 14645 4743 14703 4749
rect 14645 4740 14657 4743
rect 13780 4712 14657 4740
rect 13780 4700 13786 4712
rect 14645 4709 14657 4712
rect 14691 4709 14703 4743
rect 15378 4740 15384 4752
rect 15339 4712 15384 4740
rect 14645 4703 14703 4709
rect 15378 4700 15384 4712
rect 15436 4700 15442 4752
rect 15488 4749 15516 4780
rect 17034 4768 17040 4780
rect 17092 4768 17098 4820
rect 21910 4768 21916 4820
rect 21968 4808 21974 4820
rect 22554 4808 22560 4820
rect 21968 4780 22560 4808
rect 21968 4768 21974 4780
rect 22554 4768 22560 4780
rect 22612 4808 22618 4820
rect 22649 4811 22707 4817
rect 22649 4808 22661 4811
rect 22612 4780 22661 4808
rect 22612 4768 22618 4780
rect 22649 4777 22661 4780
rect 22695 4777 22707 4811
rect 23198 4808 23204 4820
rect 23159 4780 23204 4808
rect 22649 4771 22707 4777
rect 23198 4768 23204 4780
rect 23256 4768 23262 4820
rect 24210 4808 24216 4820
rect 24171 4780 24216 4808
rect 24210 4768 24216 4780
rect 24268 4768 24274 4820
rect 24762 4808 24768 4820
rect 24723 4780 24768 4808
rect 24762 4768 24768 4780
rect 24820 4768 24826 4820
rect 25317 4811 25375 4817
rect 25317 4777 25329 4811
rect 25363 4808 25375 4811
rect 25774 4808 25780 4820
rect 25363 4780 25780 4808
rect 25363 4777 25375 4780
rect 25317 4771 25375 4777
rect 25774 4768 25780 4780
rect 25832 4768 25838 4820
rect 26050 4808 26056 4820
rect 26011 4780 26056 4808
rect 26050 4768 26056 4780
rect 26108 4768 26114 4820
rect 15473 4743 15531 4749
rect 15473 4709 15485 4743
rect 15519 4709 15531 4743
rect 16022 4740 16028 4752
rect 15983 4712 16028 4740
rect 15473 4703 15531 4709
rect 16022 4700 16028 4712
rect 16080 4700 16086 4752
rect 16574 4700 16580 4752
rect 16632 4740 16638 4752
rect 19702 4740 19708 4752
rect 16632 4712 19708 4740
rect 16632 4700 16638 4712
rect 19702 4700 19708 4712
rect 19760 4740 19766 4752
rect 20073 4743 20131 4749
rect 20073 4740 20085 4743
rect 19760 4712 20085 4740
rect 19760 4700 19766 4712
rect 20073 4709 20085 4712
rect 20119 4740 20131 4743
rect 20622 4740 20628 4752
rect 20119 4712 20628 4740
rect 20119 4709 20131 4712
rect 20073 4703 20131 4709
rect 20622 4700 20628 4712
rect 20680 4700 20686 4752
rect 10873 4675 10931 4681
rect 10873 4641 10885 4675
rect 10919 4641 10931 4675
rect 11974 4672 11980 4684
rect 11935 4644 11980 4672
rect 10873 4635 10931 4641
rect 11974 4632 11980 4644
rect 12032 4632 12038 4684
rect 12161 4675 12219 4681
rect 12161 4641 12173 4675
rect 12207 4672 12219 4675
rect 12805 4675 12863 4681
rect 12805 4672 12817 4675
rect 12207 4644 12817 4672
rect 12207 4641 12219 4644
rect 12161 4635 12219 4641
rect 12805 4641 12817 4644
rect 12851 4641 12863 4675
rect 12805 4635 12863 4641
rect 6089 4607 6147 4613
rect 6089 4573 6101 4607
rect 6135 4604 6147 4607
rect 6362 4604 6368 4616
rect 6135 4576 6368 4604
rect 6135 4573 6147 4576
rect 6089 4567 6147 4573
rect 6362 4564 6368 4576
rect 6420 4564 6426 4616
rect 6638 4564 6644 4616
rect 6696 4604 6702 4616
rect 7282 4604 7288 4616
rect 6696 4576 7288 4604
rect 6696 4564 6702 4576
rect 7282 4564 7288 4576
rect 7340 4604 7346 4616
rect 7837 4607 7895 4613
rect 7837 4604 7849 4607
rect 7340 4576 7849 4604
rect 7340 4564 7346 4576
rect 7837 4573 7849 4576
rect 7883 4573 7895 4607
rect 7837 4567 7895 4573
rect 8294 4564 8300 4616
rect 8352 4604 8358 4616
rect 12176 4604 12204 4635
rect 14918 4632 14924 4684
rect 14976 4672 14982 4684
rect 15013 4675 15071 4681
rect 15013 4672 15025 4675
rect 14976 4644 15025 4672
rect 14976 4632 14982 4644
rect 15013 4641 15025 4644
rect 15059 4641 15071 4675
rect 15013 4635 15071 4641
rect 16485 4675 16543 4681
rect 16485 4641 16497 4675
rect 16531 4672 16543 4675
rect 17218 4672 17224 4684
rect 16531 4644 17224 4672
rect 16531 4641 16543 4644
rect 16485 4635 16543 4641
rect 17218 4632 17224 4644
rect 17276 4632 17282 4684
rect 17310 4632 17316 4684
rect 17368 4672 17374 4684
rect 17405 4675 17463 4681
rect 17405 4672 17417 4675
rect 17368 4644 17417 4672
rect 17368 4632 17374 4644
rect 17405 4641 17417 4644
rect 17451 4641 17463 4675
rect 17770 4672 17776 4684
rect 17731 4644 17776 4672
rect 17405 4635 17463 4641
rect 17770 4632 17776 4644
rect 17828 4632 17834 4684
rect 18141 4675 18199 4681
rect 18141 4641 18153 4675
rect 18187 4641 18199 4675
rect 18141 4635 18199 4641
rect 8352 4576 12204 4604
rect 8352 4564 8358 4576
rect 12618 4564 12624 4616
rect 12676 4604 12682 4616
rect 13449 4607 13507 4613
rect 13449 4604 13461 4607
rect 12676 4576 13461 4604
rect 12676 4564 12682 4576
rect 13449 4573 13461 4576
rect 13495 4573 13507 4607
rect 13449 4567 13507 4573
rect 17494 4564 17500 4616
rect 17552 4604 17558 4616
rect 18156 4604 18184 4635
rect 18322 4632 18328 4684
rect 18380 4672 18386 4684
rect 19312 4675 19370 4681
rect 19312 4672 19324 4675
rect 18380 4644 19324 4672
rect 18380 4632 18386 4644
rect 19312 4641 19324 4644
rect 19358 4672 19370 4675
rect 19886 4672 19892 4684
rect 19358 4644 19892 4672
rect 19358 4641 19370 4644
rect 19312 4635 19370 4641
rect 19886 4632 19892 4644
rect 19944 4632 19950 4684
rect 20533 4675 20591 4681
rect 20533 4641 20545 4675
rect 20579 4672 20591 4675
rect 20714 4672 20720 4684
rect 20579 4644 20720 4672
rect 20579 4641 20591 4644
rect 20533 4635 20591 4641
rect 20714 4632 20720 4644
rect 20772 4672 20778 4684
rect 20901 4675 20959 4681
rect 20901 4672 20913 4675
rect 20772 4644 20913 4672
rect 20772 4632 20778 4644
rect 20901 4641 20913 4644
rect 20947 4641 20959 4675
rect 21358 4672 21364 4684
rect 21319 4644 21364 4672
rect 20901 4635 20959 4641
rect 21358 4632 21364 4644
rect 21416 4632 21422 4684
rect 21726 4632 21732 4684
rect 21784 4672 21790 4684
rect 21928 4681 21956 4768
rect 24394 4700 24400 4752
rect 24452 4740 24458 4752
rect 25406 4740 25412 4752
rect 24452 4712 25412 4740
rect 24452 4700 24458 4712
rect 25406 4700 25412 4712
rect 25464 4740 25470 4752
rect 25593 4743 25651 4749
rect 25593 4740 25605 4743
rect 25464 4712 25605 4740
rect 25464 4700 25470 4712
rect 25593 4709 25605 4712
rect 25639 4709 25651 4743
rect 26694 4740 26700 4752
rect 26655 4712 26700 4740
rect 25593 4703 25651 4709
rect 26694 4700 26700 4712
rect 26752 4700 26758 4752
rect 21913 4675 21971 4681
rect 21913 4672 21925 4675
rect 21784 4644 21925 4672
rect 21784 4632 21790 4644
rect 21913 4641 21925 4644
rect 21959 4641 21971 4675
rect 22094 4672 22100 4684
rect 22055 4644 22100 4672
rect 21913 4635 21971 4641
rect 22094 4632 22100 4644
rect 22152 4632 22158 4684
rect 19518 4604 19524 4616
rect 17552 4576 19524 4604
rect 17552 4564 17558 4576
rect 19518 4564 19524 4576
rect 19576 4564 19582 4616
rect 21634 4564 21640 4616
rect 21692 4604 21698 4616
rect 22112 4604 22140 4632
rect 21692 4576 22140 4604
rect 22373 4607 22431 4613
rect 21692 4564 21698 4576
rect 22373 4573 22385 4607
rect 22419 4604 22431 4607
rect 24397 4607 24455 4613
rect 24397 4604 24409 4607
rect 22419 4576 24409 4604
rect 22419 4573 22431 4576
rect 22373 4567 22431 4573
rect 24397 4573 24409 4576
rect 24443 4604 24455 4607
rect 24670 4604 24676 4616
rect 24443 4576 24676 4604
rect 24443 4573 24455 4576
rect 24397 4567 24455 4573
rect 24670 4564 24676 4576
rect 24728 4564 24734 4616
rect 26418 4564 26424 4616
rect 26476 4604 26482 4616
rect 26605 4607 26663 4613
rect 26605 4604 26617 4607
rect 26476 4576 26617 4604
rect 26476 4564 26482 4576
rect 26605 4573 26617 4576
rect 26651 4573 26663 4607
rect 26878 4604 26884 4616
rect 26839 4576 26884 4604
rect 26605 4567 26663 4573
rect 26878 4564 26884 4576
rect 26936 4564 26942 4616
rect 2685 4539 2743 4545
rect 2685 4505 2697 4539
rect 2731 4536 2743 4539
rect 3050 4536 3056 4548
rect 2731 4508 3056 4536
rect 2731 4505 2743 4508
rect 2685 4499 2743 4505
rect 3050 4496 3056 4508
rect 3108 4496 3114 4548
rect 3145 4539 3203 4545
rect 3145 4505 3157 4539
rect 3191 4536 3203 4539
rect 3326 4536 3332 4548
rect 3191 4508 3332 4536
rect 3191 4505 3203 4508
rect 3145 4499 3203 4505
rect 3326 4496 3332 4508
rect 3384 4496 3390 4548
rect 4246 4536 4252 4548
rect 4207 4508 4252 4536
rect 4246 4496 4252 4508
rect 4304 4496 4310 4548
rect 6914 4496 6920 4548
rect 6972 4536 6978 4548
rect 7929 4539 7987 4545
rect 7929 4536 7941 4539
rect 6972 4508 7941 4536
rect 6972 4496 6978 4508
rect 7929 4505 7941 4508
rect 7975 4505 7987 4539
rect 7929 4499 7987 4505
rect 8849 4539 8907 4545
rect 8849 4505 8861 4539
rect 8895 4536 8907 4539
rect 10318 4536 10324 4548
rect 8895 4508 10324 4536
rect 8895 4505 8907 4508
rect 8849 4499 8907 4505
rect 10318 4496 10324 4508
rect 10376 4536 10382 4548
rect 11514 4536 11520 4548
rect 10376 4508 11520 4536
rect 10376 4496 10382 4508
rect 11514 4496 11520 4508
rect 11572 4496 11578 4548
rect 11790 4536 11796 4548
rect 11751 4508 11796 4536
rect 11790 4496 11796 4508
rect 11848 4496 11854 4548
rect 16482 4496 16488 4548
rect 16540 4536 16546 4548
rect 19705 4539 19763 4545
rect 19705 4536 19717 4539
rect 16540 4508 19717 4536
rect 16540 4496 16546 4508
rect 19705 4505 19717 4508
rect 19751 4505 19763 4539
rect 19705 4499 19763 4505
rect 1670 4428 1676 4480
rect 1728 4468 1734 4480
rect 3789 4471 3847 4477
rect 3789 4468 3801 4471
rect 1728 4440 3801 4468
rect 1728 4428 1734 4440
rect 3789 4437 3801 4440
rect 3835 4468 3847 4471
rect 4522 4468 4528 4480
rect 3835 4440 4528 4468
rect 3835 4437 3847 4440
rect 3789 4431 3847 4437
rect 4522 4428 4528 4440
rect 4580 4428 4586 4480
rect 6730 4428 6736 4480
rect 6788 4468 6794 4480
rect 6825 4471 6883 4477
rect 6825 4468 6837 4471
rect 6788 4440 6837 4468
rect 6788 4428 6794 4440
rect 6825 4437 6837 4440
rect 6871 4437 6883 4471
rect 6825 4431 6883 4437
rect 7466 4428 7472 4480
rect 7524 4468 7530 4480
rect 7607 4471 7665 4477
rect 7607 4468 7619 4471
rect 7524 4440 7619 4468
rect 7524 4428 7530 4440
rect 7607 4437 7619 4440
rect 7653 4437 7665 4471
rect 7607 4431 7665 4437
rect 7745 4471 7803 4477
rect 7745 4437 7757 4471
rect 7791 4468 7803 4471
rect 8110 4468 8116 4480
rect 7791 4440 8116 4468
rect 7791 4437 7803 4440
rect 7745 4431 7803 4437
rect 8110 4428 8116 4440
rect 8168 4428 8174 4480
rect 8754 4468 8760 4480
rect 8715 4440 8760 4468
rect 8754 4428 8760 4440
rect 8812 4428 8818 4480
rect 14182 4428 14188 4480
rect 14240 4468 14246 4480
rect 16761 4471 16819 4477
rect 16761 4468 16773 4471
rect 14240 4440 16773 4468
rect 14240 4428 14246 4440
rect 16761 4437 16773 4440
rect 16807 4468 16819 4471
rect 17770 4468 17776 4480
rect 16807 4440 17776 4468
rect 16807 4437 16819 4440
rect 16761 4431 16819 4437
rect 17770 4428 17776 4440
rect 17828 4428 17834 4480
rect 18414 4428 18420 4480
rect 18472 4468 18478 4480
rect 18693 4471 18751 4477
rect 18693 4468 18705 4471
rect 18472 4440 18705 4468
rect 18472 4428 18478 4440
rect 18693 4437 18705 4440
rect 18739 4437 18751 4471
rect 19150 4468 19156 4480
rect 19111 4440 19156 4468
rect 18693 4431 18751 4437
rect 19150 4428 19156 4440
rect 19208 4428 19214 4480
rect 19242 4428 19248 4480
rect 19300 4468 19306 4480
rect 19383 4471 19441 4477
rect 19383 4468 19395 4471
rect 19300 4440 19395 4468
rect 19300 4428 19306 4440
rect 19383 4437 19395 4440
rect 19429 4437 19441 4471
rect 23658 4468 23664 4480
rect 23619 4440 23664 4468
rect 19383 4431 19441 4437
rect 23658 4428 23664 4440
rect 23716 4428 23722 4480
rect 1104 4378 38824 4400
rect 1104 4326 7648 4378
rect 7700 4326 7712 4378
rect 7764 4326 7776 4378
rect 7828 4326 7840 4378
rect 7892 4326 20982 4378
rect 21034 4326 21046 4378
rect 21098 4326 21110 4378
rect 21162 4326 21174 4378
rect 21226 4326 34315 4378
rect 34367 4326 34379 4378
rect 34431 4326 34443 4378
rect 34495 4326 34507 4378
rect 34559 4326 38824 4378
rect 1104 4304 38824 4326
rect 1854 4264 1860 4276
rect 1815 4236 1860 4264
rect 1854 4224 1860 4236
rect 1912 4224 1918 4276
rect 2593 4267 2651 4273
rect 2593 4233 2605 4267
rect 2639 4264 2651 4267
rect 3326 4264 3332 4276
rect 2639 4236 3332 4264
rect 2639 4233 2651 4236
rect 2593 4227 2651 4233
rect 3326 4224 3332 4236
rect 3384 4224 3390 4276
rect 3694 4264 3700 4276
rect 3655 4236 3700 4264
rect 3694 4224 3700 4236
rect 3752 4224 3758 4276
rect 6638 4264 6644 4276
rect 6599 4236 6644 4264
rect 6638 4224 6644 4236
rect 6696 4224 6702 4276
rect 8849 4267 8907 4273
rect 8849 4264 8861 4267
rect 8312 4236 8861 4264
rect 2682 4156 2688 4208
rect 2740 4196 2746 4208
rect 2740 4168 3096 4196
rect 2740 4156 2746 4168
rect 3068 4137 3096 4168
rect 4246 4156 4252 4208
rect 4304 4196 4310 4208
rect 8312 4196 8340 4236
rect 8849 4233 8861 4236
rect 8895 4264 8907 4267
rect 9030 4264 9036 4276
rect 8895 4236 9036 4264
rect 8895 4233 8907 4236
rect 8849 4227 8907 4233
rect 9030 4224 9036 4236
rect 9088 4224 9094 4276
rect 9950 4224 9956 4276
rect 10008 4264 10014 4276
rect 10781 4267 10839 4273
rect 10781 4264 10793 4267
rect 10008 4236 10793 4264
rect 10008 4224 10014 4236
rect 10781 4233 10793 4236
rect 10827 4233 10839 4267
rect 10781 4227 10839 4233
rect 11517 4267 11575 4273
rect 11517 4233 11529 4267
rect 11563 4264 11575 4267
rect 15381 4267 15439 4273
rect 15381 4264 15393 4267
rect 11563 4236 15393 4264
rect 11563 4233 11575 4236
rect 11517 4227 11575 4233
rect 15381 4233 15393 4236
rect 15427 4264 15439 4267
rect 15473 4267 15531 4273
rect 15473 4264 15485 4267
rect 15427 4236 15485 4264
rect 15427 4233 15439 4236
rect 15381 4227 15439 4233
rect 15473 4233 15485 4236
rect 15519 4233 15531 4267
rect 15473 4227 15531 4233
rect 15562 4224 15568 4276
rect 15620 4264 15626 4276
rect 19426 4264 19432 4276
rect 15620 4236 19432 4264
rect 15620 4224 15626 4236
rect 19426 4224 19432 4236
rect 19484 4224 19490 4276
rect 22554 4264 22560 4276
rect 22515 4236 22560 4264
rect 22554 4224 22560 4236
rect 22612 4224 22618 4276
rect 23477 4267 23535 4273
rect 23477 4233 23489 4267
rect 23523 4264 23535 4267
rect 24026 4264 24032 4276
rect 23523 4236 24032 4264
rect 23523 4233 23535 4236
rect 23477 4227 23535 4233
rect 24026 4224 24032 4236
rect 24084 4224 24090 4276
rect 26329 4267 26387 4273
rect 24631 4236 25820 4264
rect 4304 4168 8340 4196
rect 4304 4156 4310 4168
rect 8754 4156 8760 4208
rect 8812 4196 8818 4208
rect 8812 4168 10088 4196
rect 8812 4156 8818 4168
rect 3053 4131 3111 4137
rect 3053 4128 3065 4131
rect 3031 4100 3065 4128
rect 3053 4097 3065 4100
rect 3099 4097 3111 4131
rect 3053 4091 3111 4097
rect 3142 4088 3148 4140
rect 3200 4128 3206 4140
rect 5997 4131 6055 4137
rect 5997 4128 6009 4131
rect 3200 4100 6009 4128
rect 3200 4088 3206 4100
rect 1673 4063 1731 4069
rect 1673 4029 1685 4063
rect 1719 4029 1731 4063
rect 4246 4060 4252 4072
rect 1673 4023 1731 4029
rect 4080 4032 4252 4060
rect 1394 3884 1400 3936
rect 1452 3924 1458 3936
rect 1688 3924 1716 4023
rect 2777 3995 2835 4001
rect 2777 3961 2789 3995
rect 2823 3961 2835 3995
rect 2777 3955 2835 3961
rect 2133 3927 2191 3933
rect 2133 3924 2145 3927
rect 1452 3896 2145 3924
rect 1452 3884 1458 3896
rect 2133 3893 2145 3896
rect 2179 3893 2191 3927
rect 2792 3924 2820 3955
rect 2866 3952 2872 4004
rect 2924 3992 2930 4004
rect 3050 3992 3056 4004
rect 2924 3964 3056 3992
rect 2924 3952 2930 3964
rect 3050 3952 3056 3964
rect 3108 3952 3114 4004
rect 2958 3924 2964 3936
rect 2792 3896 2964 3924
rect 2133 3887 2191 3893
rect 2958 3884 2964 3896
rect 3016 3884 3022 3936
rect 3694 3884 3700 3936
rect 3752 3924 3758 3936
rect 4080 3933 4108 4032
rect 4246 4020 4252 4032
rect 4304 4020 4310 4072
rect 4798 4060 4804 4072
rect 4759 4032 4804 4060
rect 4798 4020 4804 4032
rect 4856 4020 4862 4072
rect 5092 4069 5120 4100
rect 5997 4097 6009 4100
rect 6043 4128 6055 4131
rect 8938 4128 8944 4140
rect 6043 4100 8944 4128
rect 6043 4097 6055 4100
rect 5997 4091 6055 4097
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 9950 4128 9956 4140
rect 9646 4100 9956 4128
rect 5077 4063 5135 4069
rect 5077 4029 5089 4063
rect 5123 4029 5135 4063
rect 5626 4060 5632 4072
rect 5587 4032 5632 4060
rect 5077 4023 5135 4029
rect 5626 4020 5632 4032
rect 5684 4020 5690 4072
rect 5721 4063 5779 4069
rect 5721 4029 5733 4063
rect 5767 4060 5779 4063
rect 6454 4060 6460 4072
rect 5767 4032 6460 4060
rect 5767 4029 5779 4032
rect 5721 4023 5779 4029
rect 6454 4020 6460 4032
rect 6512 4060 6518 4072
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6512 4032 6837 4060
rect 6512 4020 6518 4032
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 9030 4060 9036 4072
rect 8991 4032 9036 4060
rect 6825 4023 6883 4029
rect 9030 4020 9036 4032
rect 9088 4060 9094 4072
rect 9646 4060 9674 4100
rect 9950 4088 9956 4100
rect 10008 4088 10014 4140
rect 10060 4128 10088 4168
rect 10318 4156 10324 4208
rect 10376 4196 10382 4208
rect 10594 4196 10600 4208
rect 10376 4168 10600 4196
rect 10376 4156 10382 4168
rect 10594 4156 10600 4168
rect 10652 4156 10658 4208
rect 14093 4199 14151 4205
rect 14093 4196 14105 4199
rect 12636 4168 14105 4196
rect 12636 4140 12664 4168
rect 14093 4165 14105 4168
rect 14139 4165 14151 4199
rect 14093 4159 14151 4165
rect 14461 4199 14519 4205
rect 14461 4165 14473 4199
rect 14507 4196 14519 4199
rect 17494 4196 17500 4208
rect 14507 4168 17500 4196
rect 14507 4165 14519 4168
rect 14461 4159 14519 4165
rect 17494 4156 17500 4168
rect 17552 4156 17558 4208
rect 18874 4156 18880 4208
rect 18932 4196 18938 4208
rect 19886 4196 19892 4208
rect 18932 4168 19288 4196
rect 19799 4168 19892 4196
rect 18932 4156 18938 4168
rect 10134 4128 10140 4140
rect 10060 4100 10140 4128
rect 10060 4069 10088 4100
rect 10134 4088 10140 4100
rect 10192 4088 10198 4140
rect 10505 4131 10563 4137
rect 10505 4097 10517 4131
rect 10551 4128 10563 4131
rect 12618 4128 12624 4140
rect 10551 4100 12624 4128
rect 10551 4097 10563 4100
rect 10505 4091 10563 4097
rect 12618 4088 12624 4100
rect 12676 4088 12682 4140
rect 12805 4131 12863 4137
rect 12805 4097 12817 4131
rect 12851 4128 12863 4131
rect 12894 4128 12900 4140
rect 12851 4100 12900 4128
rect 12851 4097 12863 4100
rect 12805 4091 12863 4097
rect 12894 4088 12900 4100
rect 12952 4088 12958 4140
rect 13170 4128 13176 4140
rect 13131 4100 13176 4128
rect 13170 4088 13176 4100
rect 13228 4088 13234 4140
rect 13814 4128 13820 4140
rect 13775 4100 13820 4128
rect 13814 4088 13820 4100
rect 13872 4088 13878 4140
rect 15381 4131 15439 4137
rect 15381 4097 15393 4131
rect 15427 4128 15439 4131
rect 17126 4128 17132 4140
rect 15427 4100 16896 4128
rect 17087 4100 17132 4128
rect 15427 4097 15439 4100
rect 15381 4091 15439 4097
rect 9088 4032 9674 4060
rect 9769 4063 9827 4069
rect 9088 4020 9094 4032
rect 9769 4029 9781 4063
rect 9815 4029 9827 4063
rect 9769 4023 9827 4029
rect 10045 4063 10103 4069
rect 10045 4029 10057 4063
rect 10091 4029 10103 4063
rect 10226 4060 10232 4072
rect 10187 4032 10232 4060
rect 10045 4023 10103 4029
rect 4816 3992 4844 4020
rect 5258 3992 5264 4004
rect 4816 3964 5264 3992
rect 5258 3952 5264 3964
rect 5316 3952 5322 4004
rect 8018 3952 8024 4004
rect 8076 3992 8082 4004
rect 8478 3992 8484 4004
rect 8076 3964 8484 3992
rect 8076 3952 8082 3964
rect 8478 3952 8484 3964
rect 8536 3952 8542 4004
rect 9784 3992 9812 4023
rect 10226 4020 10232 4032
rect 10284 4020 10290 4072
rect 10410 4020 10416 4072
rect 10468 4060 10474 4072
rect 11333 4063 11391 4069
rect 11333 4060 11345 4063
rect 10468 4032 11345 4060
rect 10468 4020 10474 4032
rect 11333 4029 11345 4032
rect 11379 4060 11391 4063
rect 11793 4063 11851 4069
rect 11793 4060 11805 4063
rect 11379 4032 11805 4060
rect 11379 4029 11391 4032
rect 11333 4023 11391 4029
rect 11793 4029 11805 4032
rect 11839 4029 11851 4063
rect 11793 4023 11851 4029
rect 11974 4020 11980 4072
rect 12032 4060 12038 4072
rect 12161 4063 12219 4069
rect 12161 4060 12173 4063
rect 12032 4032 12173 4060
rect 12032 4020 12038 4032
rect 12161 4029 12173 4032
rect 12207 4029 12219 4063
rect 12161 4023 12219 4029
rect 13998 4020 14004 4072
rect 14056 4060 14062 4072
rect 14277 4063 14335 4069
rect 14277 4060 14289 4063
rect 14056 4032 14289 4060
rect 14056 4020 14062 4032
rect 14277 4029 14289 4032
rect 14323 4060 14335 4063
rect 15930 4060 15936 4072
rect 14323 4032 14964 4060
rect 15891 4032 15936 4060
rect 14323 4029 14335 4032
rect 14277 4023 14335 4029
rect 12894 3992 12900 4004
rect 9784 3964 11284 3992
rect 12855 3964 12900 3992
rect 11256 3936 11284 3964
rect 12894 3952 12900 3964
rect 12952 3952 12958 4004
rect 4065 3927 4123 3933
rect 4065 3924 4077 3927
rect 3752 3896 4077 3924
rect 3752 3884 3758 3896
rect 4065 3893 4077 3896
rect 4111 3893 4123 3927
rect 7190 3924 7196 3936
rect 7151 3896 7196 3924
rect 4065 3887 4123 3893
rect 7190 3884 7196 3896
rect 7248 3884 7254 3936
rect 7742 3924 7748 3936
rect 7703 3896 7748 3924
rect 7742 3884 7748 3896
rect 7800 3884 7806 3936
rect 8113 3927 8171 3933
rect 8113 3893 8125 3927
rect 8159 3924 8171 3927
rect 8202 3924 8208 3936
rect 8159 3896 8208 3924
rect 8159 3893 8171 3896
rect 8113 3887 8171 3893
rect 8202 3884 8208 3896
rect 8260 3884 8266 3936
rect 11238 3924 11244 3936
rect 11199 3896 11244 3924
rect 11238 3884 11244 3896
rect 11296 3884 11302 3936
rect 12342 3884 12348 3936
rect 12400 3924 12406 3936
rect 14826 3924 14832 3936
rect 12400 3896 14832 3924
rect 12400 3884 12406 3896
rect 14826 3884 14832 3896
rect 14884 3884 14890 3936
rect 14936 3933 14964 4032
rect 15930 4020 15936 4032
rect 15988 4020 15994 4072
rect 16868 4069 16896 4100
rect 17126 4088 17132 4100
rect 17184 4088 17190 4140
rect 17218 4088 17224 4140
rect 17276 4128 17282 4140
rect 19150 4128 19156 4140
rect 17276 4100 19156 4128
rect 17276 4088 17282 4100
rect 18248 4072 18276 4100
rect 19150 4088 19156 4100
rect 19208 4088 19214 4140
rect 16117 4063 16175 4069
rect 16117 4029 16129 4063
rect 16163 4029 16175 4063
rect 16117 4023 16175 4029
rect 16485 4063 16543 4069
rect 16485 4029 16497 4063
rect 16531 4029 16543 4063
rect 16485 4023 16543 4029
rect 16853 4063 16911 4069
rect 16853 4029 16865 4063
rect 16899 4060 16911 4063
rect 17402 4060 17408 4072
rect 16899 4032 17408 4060
rect 16899 4029 16911 4032
rect 16853 4023 16911 4029
rect 15838 3952 15844 4004
rect 15896 3992 15902 4004
rect 16132 3992 16160 4023
rect 15896 3964 16160 3992
rect 16500 3992 16528 4023
rect 17402 4020 17408 4032
rect 17460 4020 17466 4072
rect 18230 4060 18236 4072
rect 18191 4032 18236 4060
rect 18230 4020 18236 4032
rect 18288 4020 18294 4072
rect 18414 4020 18420 4072
rect 18472 4060 18478 4072
rect 18509 4063 18567 4069
rect 18509 4060 18521 4063
rect 18472 4032 18521 4060
rect 18472 4020 18478 4032
rect 18509 4029 18521 4032
rect 18555 4029 18567 4063
rect 18509 4023 18567 4029
rect 18877 4063 18935 4069
rect 18877 4029 18889 4063
rect 18923 4060 18935 4063
rect 19058 4060 19064 4072
rect 18923 4032 19064 4060
rect 18923 4029 18935 4032
rect 18877 4023 18935 4029
rect 18892 3992 18920 4023
rect 19058 4020 19064 4032
rect 19116 4020 19122 4072
rect 19260 4069 19288 4168
rect 19886 4156 19892 4168
rect 19944 4196 19950 4208
rect 24631 4196 24659 4236
rect 19944 4168 24659 4196
rect 19944 4156 19950 4168
rect 24762 4156 24768 4208
rect 24820 4196 24826 4208
rect 24857 4199 24915 4205
rect 24857 4196 24869 4199
rect 24820 4168 24869 4196
rect 24820 4156 24826 4168
rect 24857 4165 24869 4168
rect 24903 4196 24915 4199
rect 25225 4199 25283 4205
rect 25225 4196 25237 4199
rect 24903 4168 25237 4196
rect 24903 4165 24915 4168
rect 24857 4159 24915 4165
rect 25225 4165 25237 4168
rect 25271 4165 25283 4199
rect 25225 4159 25283 4165
rect 21913 4131 21971 4137
rect 21913 4097 21925 4131
rect 21959 4128 21971 4131
rect 23658 4128 23664 4140
rect 21959 4100 23664 4128
rect 21959 4097 21971 4100
rect 21913 4091 21971 4097
rect 23658 4088 23664 4100
rect 23716 4088 23722 4140
rect 19245 4063 19303 4069
rect 19245 4029 19257 4063
rect 19291 4029 19303 4063
rect 19245 4023 19303 4029
rect 19426 4020 19432 4072
rect 19484 4060 19490 4072
rect 20714 4060 20720 4072
rect 19484 4032 20720 4060
rect 19484 4020 19490 4032
rect 20714 4020 20720 4032
rect 20772 4020 20778 4072
rect 20901 4063 20959 4069
rect 20901 4029 20913 4063
rect 20947 4029 20959 4063
rect 20901 4023 20959 4029
rect 20916 3992 20944 4023
rect 21266 4020 21272 4072
rect 21324 4060 21330 4072
rect 21453 4063 21511 4069
rect 21453 4060 21465 4063
rect 21324 4032 21465 4060
rect 21324 4020 21330 4032
rect 21453 4029 21465 4032
rect 21499 4029 21511 4063
rect 21634 4060 21640 4072
rect 21595 4032 21640 4060
rect 21453 4023 21511 4029
rect 21358 3992 21364 4004
rect 16500 3964 18920 3992
rect 20456 3964 21364 3992
rect 15896 3952 15902 3964
rect 14921 3927 14979 3933
rect 14921 3893 14933 3927
rect 14967 3924 14979 3927
rect 15194 3924 15200 3936
rect 14967 3896 15200 3924
rect 14967 3893 14979 3896
rect 14921 3887 14979 3893
rect 15194 3884 15200 3896
rect 15252 3884 15258 3936
rect 15654 3884 15660 3936
rect 15712 3924 15718 3936
rect 16500 3924 16528 3964
rect 20456 3936 20484 3964
rect 21358 3952 21364 3964
rect 21416 3952 21422 4004
rect 21468 3992 21496 4023
rect 21634 4020 21640 4032
rect 21692 4020 21698 4072
rect 22189 3995 22247 4001
rect 22189 3992 22201 3995
rect 21468 3964 22201 3992
rect 22189 3961 22201 3964
rect 22235 3961 22247 3995
rect 25240 3992 25268 4159
rect 25406 4128 25412 4140
rect 25367 4100 25412 4128
rect 25406 4088 25412 4100
rect 25464 4088 25470 4140
rect 25792 4128 25820 4236
rect 26329 4233 26341 4267
rect 26375 4264 26387 4267
rect 26694 4264 26700 4276
rect 26375 4236 26700 4264
rect 26375 4233 26387 4236
rect 26329 4227 26387 4233
rect 26694 4224 26700 4236
rect 26752 4224 26758 4276
rect 27430 4264 27436 4276
rect 27391 4236 27436 4264
rect 27430 4224 27436 4236
rect 27488 4224 27494 4276
rect 26418 4156 26424 4208
rect 26476 4196 26482 4208
rect 26973 4199 27031 4205
rect 26973 4196 26985 4199
rect 26476 4168 26985 4196
rect 26476 4156 26482 4168
rect 26973 4165 26985 4168
rect 27019 4165 27031 4199
rect 35069 4199 35127 4205
rect 26973 4159 27031 4165
rect 28966 4168 34928 4196
rect 26786 4128 26792 4140
rect 25792 4100 26792 4128
rect 26786 4088 26792 4100
rect 26844 4088 26850 4140
rect 27224 4063 27282 4069
rect 27224 4029 27236 4063
rect 27270 4060 27282 4063
rect 27270 4032 27752 4060
rect 27270 4029 27282 4032
rect 27224 4023 27282 4029
rect 27724 4001 27752 4032
rect 25730 3995 25788 4001
rect 25730 3992 25742 3995
rect 25240 3964 25742 3992
rect 22189 3955 22247 3961
rect 25730 3961 25742 3964
rect 25776 3961 25788 3995
rect 25730 3955 25788 3961
rect 27709 3995 27767 4001
rect 27709 3961 27721 3995
rect 27755 3992 27767 3995
rect 28966 3992 28994 4168
rect 31386 4128 31392 4140
rect 31347 4100 31392 4128
rect 31386 4088 31392 4100
rect 31444 4088 31450 4140
rect 31662 4128 31668 4140
rect 31623 4100 31668 4128
rect 31662 4088 31668 4100
rect 31720 4088 31726 4140
rect 34900 4128 34928 4168
rect 35069 4165 35081 4199
rect 35115 4196 35127 4199
rect 36078 4196 36084 4208
rect 35115 4168 36084 4196
rect 35115 4165 35127 4168
rect 35069 4159 35127 4165
rect 36078 4156 36084 4168
rect 36136 4156 36142 4208
rect 35526 4128 35532 4140
rect 34900 4100 35532 4128
rect 34900 4069 34928 4100
rect 35526 4088 35532 4100
rect 35584 4088 35590 4140
rect 34885 4063 34943 4069
rect 34885 4029 34897 4063
rect 34931 4029 34943 4063
rect 34885 4023 34943 4029
rect 27755 3964 28994 3992
rect 27755 3961 27767 3964
rect 27709 3955 27767 3961
rect 31478 3952 31484 4004
rect 31536 3992 31542 4004
rect 31536 3964 31581 3992
rect 31536 3952 31542 3964
rect 15712 3896 16528 3924
rect 15712 3884 15718 3896
rect 17126 3884 17132 3936
rect 17184 3924 17190 3936
rect 17310 3924 17316 3936
rect 17184 3896 17316 3924
rect 17184 3884 17190 3896
rect 17310 3884 17316 3896
rect 17368 3884 17374 3936
rect 17678 3884 17684 3936
rect 17736 3924 17742 3936
rect 17773 3927 17831 3933
rect 17773 3924 17785 3927
rect 17736 3896 17785 3924
rect 17736 3884 17742 3896
rect 17773 3893 17785 3896
rect 17819 3893 17831 3927
rect 18138 3924 18144 3936
rect 18099 3896 18144 3924
rect 17773 3887 17831 3893
rect 18138 3884 18144 3896
rect 18196 3884 18202 3936
rect 20349 3927 20407 3933
rect 20349 3893 20361 3927
rect 20395 3924 20407 3927
rect 20438 3924 20444 3936
rect 20395 3896 20444 3924
rect 20395 3893 20407 3896
rect 20349 3887 20407 3893
rect 20438 3884 20444 3896
rect 20496 3884 20502 3936
rect 24026 3924 24032 3936
rect 23987 3896 24032 3924
rect 24026 3884 24032 3896
rect 24084 3884 24090 3936
rect 24578 3924 24584 3936
rect 24539 3896 24584 3924
rect 24578 3884 24584 3896
rect 24636 3884 24642 3936
rect 31205 3927 31263 3933
rect 31205 3893 31217 3927
rect 31251 3924 31263 3927
rect 31294 3924 31300 3936
rect 31251 3896 31300 3924
rect 31251 3893 31263 3896
rect 31205 3887 31263 3893
rect 31294 3884 31300 3896
rect 31352 3884 31358 3936
rect 1104 3834 38824 3856
rect 1104 3782 14315 3834
rect 14367 3782 14379 3834
rect 14431 3782 14443 3834
rect 14495 3782 14507 3834
rect 14559 3782 27648 3834
rect 27700 3782 27712 3834
rect 27764 3782 27776 3834
rect 27828 3782 27840 3834
rect 27892 3782 38824 3834
rect 1104 3760 38824 3782
rect 1946 3720 1952 3732
rect 1907 3692 1952 3720
rect 1946 3680 1952 3692
rect 2004 3680 2010 3732
rect 6730 3720 6736 3732
rect 6691 3692 6736 3720
rect 6730 3680 6736 3692
rect 6788 3680 6794 3732
rect 7653 3723 7711 3729
rect 7653 3689 7665 3723
rect 7699 3720 7711 3723
rect 8110 3720 8116 3732
rect 7699 3692 8116 3720
rect 7699 3689 7711 3692
rect 7653 3683 7711 3689
rect 8110 3680 8116 3692
rect 8168 3680 8174 3732
rect 8938 3680 8944 3732
rect 8996 3720 9002 3732
rect 9401 3723 9459 3729
rect 9401 3720 9413 3723
rect 8996 3692 9413 3720
rect 8996 3680 9002 3692
rect 9401 3689 9413 3692
rect 9447 3689 9459 3723
rect 9401 3683 9459 3689
rect 10502 3680 10508 3732
rect 10560 3720 10566 3732
rect 11057 3723 11115 3729
rect 11057 3720 11069 3723
rect 10560 3692 11069 3720
rect 10560 3680 10566 3692
rect 11057 3689 11069 3692
rect 11103 3720 11115 3723
rect 12066 3720 12072 3732
rect 11103 3692 12072 3720
rect 11103 3689 11115 3692
rect 11057 3683 11115 3689
rect 12066 3680 12072 3692
rect 12124 3720 12130 3732
rect 14182 3720 14188 3732
rect 12124 3692 14188 3720
rect 12124 3680 12130 3692
rect 14182 3680 14188 3692
rect 14240 3680 14246 3732
rect 15010 3720 15016 3732
rect 14971 3692 15016 3720
rect 15010 3680 15016 3692
rect 15068 3680 15074 3732
rect 15473 3723 15531 3729
rect 15473 3689 15485 3723
rect 15519 3720 15531 3723
rect 19978 3720 19984 3732
rect 15519 3692 19984 3720
rect 15519 3689 15531 3692
rect 15473 3683 15531 3689
rect 19978 3680 19984 3692
rect 20036 3680 20042 3732
rect 20165 3723 20223 3729
rect 20165 3689 20177 3723
rect 20211 3720 20223 3723
rect 21634 3720 21640 3732
rect 20211 3692 21640 3720
rect 20211 3689 20223 3692
rect 20165 3683 20223 3689
rect 21634 3680 21640 3692
rect 21692 3720 21698 3732
rect 21729 3723 21787 3729
rect 21729 3720 21741 3723
rect 21692 3692 21741 3720
rect 21692 3680 21698 3692
rect 21729 3689 21741 3692
rect 21775 3689 21787 3723
rect 24670 3720 24676 3732
rect 24631 3692 24676 3720
rect 21729 3683 21787 3689
rect 24670 3680 24676 3692
rect 24728 3680 24734 3732
rect 31386 3720 31392 3732
rect 31347 3692 31392 3720
rect 31386 3680 31392 3692
rect 31444 3680 31450 3732
rect 1578 3612 1584 3664
rect 1636 3652 1642 3664
rect 2225 3655 2283 3661
rect 2225 3652 2237 3655
rect 1636 3624 2237 3652
rect 1636 3612 1642 3624
rect 2225 3621 2237 3624
rect 2271 3621 2283 3655
rect 2225 3615 2283 3621
rect 1464 3587 1522 3593
rect 1464 3553 1476 3587
rect 1510 3553 1522 3587
rect 1464 3547 1522 3553
rect 1479 3448 1507 3547
rect 2240 3516 2268 3615
rect 2498 3612 2504 3664
rect 2556 3652 2562 3664
rect 2593 3655 2651 3661
rect 2593 3652 2605 3655
rect 2556 3624 2605 3652
rect 2556 3612 2562 3624
rect 2593 3621 2605 3624
rect 2639 3621 2651 3655
rect 5813 3655 5871 3661
rect 5813 3652 5825 3655
rect 2593 3615 2651 3621
rect 5368 3624 5825 3652
rect 5368 3596 5396 3624
rect 5813 3621 5825 3624
rect 5859 3621 5871 3655
rect 8018 3652 8024 3664
rect 7979 3624 8024 3652
rect 5813 3615 5871 3621
rect 8018 3612 8024 3624
rect 8076 3652 8082 3664
rect 8665 3655 8723 3661
rect 8076 3624 8156 3652
rect 8076 3612 8082 3624
rect 3510 3584 3516 3596
rect 3423 3556 3516 3584
rect 2501 3519 2559 3525
rect 2501 3516 2513 3519
rect 2240 3488 2513 3516
rect 2501 3485 2513 3488
rect 2547 3485 2559 3519
rect 2501 3479 2559 3485
rect 2777 3519 2835 3525
rect 2777 3485 2789 3519
rect 2823 3485 2835 3519
rect 2777 3479 2835 3485
rect 2682 3448 2688 3460
rect 1479 3420 2688 3448
rect 2682 3408 2688 3420
rect 2740 3448 2746 3460
rect 2792 3448 2820 3479
rect 2740 3420 2820 3448
rect 2740 3408 2746 3420
rect 106 3340 112 3392
rect 164 3380 170 3392
rect 1535 3383 1593 3389
rect 1535 3380 1547 3383
rect 164 3352 1547 3380
rect 164 3340 170 3352
rect 1535 3349 1547 3352
rect 1581 3349 1593 3383
rect 1535 3343 1593 3349
rect 2130 3340 2136 3392
rect 2188 3380 2194 3392
rect 3436 3389 3464 3556
rect 3510 3544 3516 3556
rect 3568 3584 3574 3596
rect 4065 3587 4123 3593
rect 4065 3584 4077 3587
rect 3568 3556 4077 3584
rect 3568 3544 3574 3556
rect 4065 3553 4077 3556
rect 4111 3553 4123 3587
rect 4798 3584 4804 3596
rect 4711 3556 4804 3584
rect 4065 3547 4123 3553
rect 4798 3544 4804 3556
rect 4856 3544 4862 3596
rect 5077 3587 5135 3593
rect 5077 3553 5089 3587
rect 5123 3584 5135 3587
rect 5350 3584 5356 3596
rect 5123 3556 5356 3584
rect 5123 3553 5135 3556
rect 5077 3547 5135 3553
rect 5350 3544 5356 3556
rect 5408 3544 5414 3596
rect 5445 3587 5503 3593
rect 5445 3553 5457 3587
rect 5491 3584 5503 3587
rect 5626 3584 5632 3596
rect 5491 3556 5632 3584
rect 5491 3553 5503 3556
rect 5445 3547 5503 3553
rect 5626 3544 5632 3556
rect 5684 3544 5690 3596
rect 6362 3584 6368 3596
rect 6323 3556 6368 3584
rect 6362 3544 6368 3556
rect 6420 3544 6426 3596
rect 8128 3593 8156 3624
rect 8665 3621 8677 3655
rect 8711 3652 8723 3655
rect 12618 3652 12624 3664
rect 8711 3624 12624 3652
rect 8711 3621 8723 3624
rect 8665 3615 8723 3621
rect 12618 3612 12624 3624
rect 12676 3612 12682 3664
rect 13630 3652 13636 3664
rect 13004 3624 13636 3652
rect 8113 3587 8171 3593
rect 8113 3553 8125 3587
rect 8159 3553 8171 3587
rect 8113 3547 8171 3553
rect 8202 3544 8208 3596
rect 8260 3584 8266 3596
rect 8297 3587 8355 3593
rect 8297 3584 8309 3587
rect 8260 3556 8309 3584
rect 8260 3544 8266 3556
rect 8297 3553 8309 3556
rect 8343 3553 8355 3587
rect 8297 3547 8355 3553
rect 9125 3587 9183 3593
rect 9125 3553 9137 3587
rect 9171 3584 9183 3587
rect 9214 3584 9220 3596
rect 9171 3556 9220 3584
rect 9171 3553 9183 3556
rect 9125 3547 9183 3553
rect 9214 3544 9220 3556
rect 9272 3544 9278 3596
rect 9766 3584 9772 3596
rect 9727 3556 9772 3584
rect 9766 3544 9772 3556
rect 9824 3544 9830 3596
rect 10410 3584 10416 3596
rect 10371 3556 10416 3584
rect 10410 3544 10416 3556
rect 10468 3544 10474 3596
rect 11514 3584 11520 3596
rect 11475 3556 11520 3584
rect 11514 3544 11520 3556
rect 11572 3544 11578 3596
rect 11882 3584 11888 3596
rect 11843 3556 11888 3584
rect 11882 3544 11888 3556
rect 11940 3544 11946 3596
rect 12066 3584 12072 3596
rect 12027 3556 12072 3584
rect 12066 3544 12072 3556
rect 12124 3544 12130 3596
rect 12250 3544 12256 3596
rect 12308 3584 12314 3596
rect 12437 3587 12495 3593
rect 12437 3584 12449 3587
rect 12308 3556 12449 3584
rect 12308 3544 12314 3556
rect 12437 3553 12449 3556
rect 12483 3553 12495 3587
rect 12437 3547 12495 3553
rect 4816 3516 4844 3544
rect 12894 3516 12900 3528
rect 4816 3488 6132 3516
rect 4798 3408 4804 3460
rect 4856 3448 4862 3460
rect 5445 3451 5503 3457
rect 5445 3448 5457 3451
rect 4856 3420 5457 3448
rect 4856 3408 4862 3420
rect 5445 3417 5457 3420
rect 5491 3448 5503 3451
rect 5534 3448 5540 3460
rect 5491 3420 5540 3448
rect 5491 3417 5503 3420
rect 5445 3411 5503 3417
rect 5534 3408 5540 3420
rect 5592 3408 5598 3460
rect 6104 3392 6132 3488
rect 11117 3488 12900 3516
rect 7285 3451 7343 3457
rect 7285 3417 7297 3451
rect 7331 3448 7343 3451
rect 11117 3448 11145 3488
rect 12894 3476 12900 3488
rect 12952 3516 12958 3528
rect 13004 3525 13032 3624
rect 13630 3612 13636 3624
rect 13688 3652 13694 3664
rect 13725 3655 13783 3661
rect 13725 3652 13737 3655
rect 13688 3624 13737 3652
rect 13688 3612 13694 3624
rect 13725 3621 13737 3624
rect 13771 3621 13783 3655
rect 13725 3615 13783 3621
rect 14277 3655 14335 3661
rect 14277 3621 14289 3655
rect 14323 3652 14335 3655
rect 14734 3652 14740 3664
rect 14323 3624 14740 3652
rect 14323 3621 14335 3624
rect 14277 3615 14335 3621
rect 14734 3612 14740 3624
rect 14792 3652 14798 3664
rect 15378 3652 15384 3664
rect 14792 3624 15384 3652
rect 14792 3612 14798 3624
rect 15378 3612 15384 3624
rect 15436 3612 15442 3664
rect 15930 3612 15936 3664
rect 15988 3652 15994 3664
rect 16301 3655 16359 3661
rect 16301 3652 16313 3655
rect 15988 3624 16313 3652
rect 15988 3612 15994 3624
rect 16301 3621 16313 3624
rect 16347 3652 16359 3655
rect 17129 3655 17187 3661
rect 17129 3652 17141 3655
rect 16347 3624 17141 3652
rect 16347 3621 16359 3624
rect 16301 3615 16359 3621
rect 17129 3621 17141 3624
rect 17175 3652 17187 3655
rect 17218 3652 17224 3664
rect 17175 3624 17224 3652
rect 17175 3621 17187 3624
rect 17129 3615 17187 3621
rect 17218 3612 17224 3624
rect 17276 3612 17282 3664
rect 17770 3612 17776 3664
rect 17828 3652 17834 3664
rect 17828 3624 18828 3652
rect 17828 3612 17834 3624
rect 15286 3584 15292 3596
rect 15247 3556 15292 3584
rect 15286 3544 15292 3556
rect 15344 3544 15350 3596
rect 15838 3584 15844 3596
rect 15799 3556 15844 3584
rect 15838 3544 15844 3556
rect 15896 3544 15902 3596
rect 17037 3587 17095 3593
rect 17037 3553 17049 3587
rect 17083 3584 17095 3587
rect 17310 3584 17316 3596
rect 17083 3556 17316 3584
rect 17083 3553 17095 3556
rect 17037 3547 17095 3553
rect 17310 3544 17316 3556
rect 17368 3544 17374 3596
rect 17678 3544 17684 3596
rect 17736 3584 17742 3596
rect 17865 3587 17923 3593
rect 17865 3584 17877 3587
rect 17736 3556 17877 3584
rect 17736 3544 17742 3556
rect 17865 3553 17877 3556
rect 17911 3553 17923 3587
rect 18230 3584 18236 3596
rect 18191 3556 18236 3584
rect 17865 3547 17923 3553
rect 18230 3544 18236 3556
rect 18288 3544 18294 3596
rect 18414 3584 18420 3596
rect 18375 3556 18420 3584
rect 18414 3544 18420 3556
rect 18472 3544 18478 3596
rect 18800 3593 18828 3624
rect 19058 3612 19064 3664
rect 19116 3652 19122 3664
rect 19705 3655 19763 3661
rect 19705 3652 19717 3655
rect 19116 3624 19717 3652
rect 19116 3612 19122 3624
rect 19705 3621 19717 3624
rect 19751 3621 19763 3655
rect 19705 3615 19763 3621
rect 20714 3612 20720 3664
rect 20772 3652 20778 3664
rect 21361 3655 21419 3661
rect 21361 3652 21373 3655
rect 20772 3624 21373 3652
rect 20772 3612 20778 3624
rect 21361 3621 21373 3624
rect 21407 3621 21419 3655
rect 21361 3615 21419 3621
rect 23839 3655 23897 3661
rect 23839 3621 23851 3655
rect 23885 3652 23897 3655
rect 24026 3652 24032 3664
rect 23885 3624 24032 3652
rect 23885 3621 23897 3624
rect 23839 3615 23897 3621
rect 24026 3612 24032 3624
rect 24084 3612 24090 3664
rect 32306 3652 32312 3664
rect 32267 3624 32312 3652
rect 32306 3612 32312 3624
rect 32364 3612 32370 3664
rect 18785 3587 18843 3593
rect 18785 3553 18797 3587
rect 18831 3584 18843 3587
rect 18874 3584 18880 3596
rect 18831 3556 18880 3584
rect 18831 3553 18843 3556
rect 18785 3547 18843 3553
rect 18874 3544 18880 3556
rect 18932 3544 18938 3596
rect 18966 3544 18972 3596
rect 19024 3584 19030 3596
rect 19153 3587 19211 3593
rect 19153 3584 19165 3587
rect 19024 3556 19165 3584
rect 19024 3544 19030 3556
rect 19153 3553 19165 3556
rect 19199 3553 19211 3587
rect 19153 3547 19211 3553
rect 19334 3544 19340 3596
rect 19392 3584 19398 3596
rect 20968 3587 21026 3593
rect 19392 3556 20852 3584
rect 19392 3544 19398 3556
rect 12989 3519 13047 3525
rect 12989 3516 13001 3519
rect 12952 3488 13001 3516
rect 12952 3476 12958 3488
rect 12989 3485 13001 3488
rect 13035 3485 13047 3519
rect 12989 3479 13047 3485
rect 13633 3519 13691 3525
rect 13633 3485 13645 3519
rect 13679 3516 13691 3519
rect 14645 3519 14703 3525
rect 14645 3516 14657 3519
rect 13679 3488 14657 3516
rect 13679 3485 13691 3488
rect 13633 3479 13691 3485
rect 14645 3485 14657 3488
rect 14691 3516 14703 3519
rect 19242 3516 19248 3528
rect 14691 3488 19248 3516
rect 14691 3485 14703 3488
rect 14645 3479 14703 3485
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 20438 3516 20444 3528
rect 20399 3488 20444 3516
rect 20438 3476 20444 3488
rect 20496 3476 20502 3528
rect 20824 3516 20852 3556
rect 20968 3553 20980 3587
rect 21014 3584 21026 3587
rect 21450 3584 21456 3596
rect 21014 3556 21456 3584
rect 21014 3553 21026 3556
rect 20968 3547 21026 3553
rect 21450 3544 21456 3556
rect 21508 3544 21514 3596
rect 23474 3544 23480 3596
rect 23532 3584 23538 3596
rect 25498 3584 25504 3596
rect 23532 3556 23577 3584
rect 25056 3556 25504 3584
rect 23532 3544 23538 3556
rect 25056 3516 25084 3556
rect 25498 3544 25504 3556
rect 25556 3544 25562 3596
rect 25222 3516 25228 3528
rect 20824 3488 25084 3516
rect 25183 3488 25228 3516
rect 25222 3476 25228 3488
rect 25280 3476 25286 3528
rect 32214 3516 32220 3528
rect 32175 3488 32220 3516
rect 32214 3476 32220 3488
rect 32272 3476 32278 3528
rect 32493 3519 32551 3525
rect 32493 3485 32505 3519
rect 32539 3485 32551 3519
rect 32493 3479 32551 3485
rect 7331 3420 11145 3448
rect 7331 3417 7343 3420
rect 7285 3411 7343 3417
rect 11238 3408 11244 3460
rect 11296 3448 11302 3460
rect 11296 3420 11836 3448
rect 11296 3408 11302 3420
rect 3421 3383 3479 3389
rect 3421 3380 3433 3383
rect 2188 3352 3433 3380
rect 2188 3340 2194 3352
rect 3421 3349 3433 3352
rect 3467 3349 3479 3383
rect 3878 3380 3884 3392
rect 3839 3352 3884 3380
rect 3421 3343 3479 3349
rect 3878 3340 3884 3352
rect 3936 3340 3942 3392
rect 6086 3340 6092 3392
rect 6144 3380 6150 3392
rect 6181 3383 6239 3389
rect 6181 3380 6193 3383
rect 6144 3352 6193 3380
rect 6144 3340 6150 3352
rect 6181 3349 6193 3352
rect 6227 3349 6239 3383
rect 6181 3343 6239 3349
rect 9398 3340 9404 3392
rect 9456 3380 9462 3392
rect 10781 3383 10839 3389
rect 10781 3380 10793 3383
rect 9456 3352 10793 3380
rect 9456 3340 9462 3352
rect 10781 3349 10793 3352
rect 10827 3380 10839 3383
rect 11698 3380 11704 3392
rect 10827 3352 11704 3380
rect 10827 3349 10839 3352
rect 10781 3343 10839 3349
rect 11698 3340 11704 3352
rect 11756 3340 11762 3392
rect 11808 3380 11836 3420
rect 12434 3408 12440 3460
rect 12492 3448 12498 3460
rect 12621 3451 12679 3457
rect 12621 3448 12633 3451
rect 12492 3420 12633 3448
rect 12492 3408 12498 3420
rect 12621 3417 12633 3420
rect 12667 3417 12679 3451
rect 12621 3411 12679 3417
rect 12710 3408 12716 3460
rect 12768 3448 12774 3460
rect 13357 3451 13415 3457
rect 13357 3448 13369 3451
rect 12768 3420 13369 3448
rect 12768 3408 12774 3420
rect 13357 3417 13369 3420
rect 13403 3417 13415 3451
rect 13357 3411 13415 3417
rect 14182 3408 14188 3460
rect 14240 3448 14246 3460
rect 19337 3451 19395 3457
rect 14240 3420 18552 3448
rect 14240 3408 14246 3420
rect 14660 3392 14688 3420
rect 14550 3380 14556 3392
rect 11808 3352 14556 3380
rect 14550 3340 14556 3352
rect 14608 3340 14614 3392
rect 14642 3340 14648 3392
rect 14700 3340 14706 3392
rect 15838 3340 15844 3392
rect 15896 3380 15902 3392
rect 17126 3380 17132 3392
rect 15896 3352 17132 3380
rect 15896 3340 15902 3352
rect 17126 3340 17132 3352
rect 17184 3380 17190 3392
rect 17405 3383 17463 3389
rect 17405 3380 17417 3383
rect 17184 3352 17417 3380
rect 17184 3340 17190 3352
rect 17405 3349 17417 3352
rect 17451 3380 17463 3383
rect 18414 3380 18420 3392
rect 17451 3352 18420 3380
rect 17451 3349 17463 3352
rect 17405 3343 17463 3349
rect 18414 3340 18420 3352
rect 18472 3340 18478 3392
rect 18524 3380 18552 3420
rect 19337 3417 19349 3451
rect 19383 3448 19395 3451
rect 20898 3448 20904 3460
rect 19383 3420 20904 3448
rect 19383 3417 19395 3420
rect 19337 3411 19395 3417
rect 20898 3408 20904 3420
rect 20956 3408 20962 3460
rect 31662 3408 31668 3460
rect 31720 3448 31726 3460
rect 32508 3448 32536 3479
rect 31720 3420 32536 3448
rect 31720 3408 31726 3420
rect 21039 3383 21097 3389
rect 21039 3380 21051 3383
rect 18524 3352 21051 3380
rect 21039 3349 21051 3352
rect 21085 3349 21097 3383
rect 21039 3343 21097 3349
rect 24397 3383 24455 3389
rect 24397 3349 24409 3383
rect 24443 3380 24455 3383
rect 30834 3380 30840 3392
rect 24443 3352 30840 3380
rect 24443 3349 24455 3352
rect 24397 3343 24455 3349
rect 30834 3340 30840 3352
rect 30892 3340 30898 3392
rect 1104 3290 38824 3312
rect 1104 3238 7648 3290
rect 7700 3238 7712 3290
rect 7764 3238 7776 3290
rect 7828 3238 7840 3290
rect 7892 3238 20982 3290
rect 21034 3238 21046 3290
rect 21098 3238 21110 3290
rect 21162 3238 21174 3290
rect 21226 3238 34315 3290
rect 34367 3238 34379 3290
rect 34431 3238 34443 3290
rect 34495 3238 34507 3290
rect 34559 3238 38824 3290
rect 1104 3216 38824 3238
rect 3878 3136 3884 3188
rect 3936 3176 3942 3188
rect 4341 3179 4399 3185
rect 4341 3176 4353 3179
rect 3936 3148 4353 3176
rect 3936 3136 3942 3148
rect 4341 3145 4353 3148
rect 4387 3176 4399 3179
rect 5626 3176 5632 3188
rect 4387 3148 5632 3176
rect 4387 3145 4399 3148
rect 4341 3139 4399 3145
rect 5626 3136 5632 3148
rect 5684 3136 5690 3188
rect 6086 3176 6092 3188
rect 6047 3148 6092 3176
rect 6086 3136 6092 3148
rect 6144 3136 6150 3188
rect 6457 3179 6515 3185
rect 6457 3145 6469 3179
rect 6503 3176 6515 3179
rect 6730 3176 6736 3188
rect 6503 3148 6736 3176
rect 6503 3145 6515 3148
rect 6457 3139 6515 3145
rect 4709 3111 4767 3117
rect 4709 3077 4721 3111
rect 4755 3108 4767 3111
rect 6472 3108 6500 3139
rect 6730 3136 6736 3148
rect 6788 3136 6794 3188
rect 9766 3176 9772 3188
rect 7161 3148 9772 3176
rect 4755 3080 6500 3108
rect 4755 3077 4767 3080
rect 4709 3071 4767 3077
rect 2130 3040 2136 3052
rect 2091 3012 2136 3040
rect 2130 3000 2136 3012
rect 2188 3000 2194 3052
rect 3053 3043 3111 3049
rect 3053 3009 3065 3043
rect 3099 3040 3111 3043
rect 4338 3040 4344 3052
rect 3099 3012 4344 3040
rect 3099 3009 3111 3012
rect 3053 3003 3111 3009
rect 4338 3000 4344 3012
rect 4396 3000 4402 3052
rect 4798 3040 4804 3052
rect 4759 3012 4804 3040
rect 4798 3000 4804 3012
rect 4856 3000 4862 3052
rect 1394 2932 1400 2984
rect 1452 2972 1458 2984
rect 1489 2975 1547 2981
rect 1489 2972 1501 2975
rect 1452 2944 1501 2972
rect 1452 2932 1458 2944
rect 1489 2941 1501 2944
rect 1535 2941 1547 2975
rect 1489 2935 1547 2941
rect 2774 2864 2780 2916
rect 2832 2904 2838 2916
rect 2961 2907 3019 2913
rect 2961 2904 2973 2907
rect 2832 2876 2973 2904
rect 2832 2864 2838 2876
rect 2961 2873 2973 2876
rect 3007 2904 3019 2907
rect 3415 2907 3473 2913
rect 3415 2904 3427 2907
rect 3007 2876 3427 2904
rect 3007 2873 3019 2876
rect 2961 2867 3019 2873
rect 3415 2873 3427 2876
rect 3461 2904 3473 2907
rect 3510 2904 3516 2916
rect 3461 2876 3516 2904
rect 3461 2873 3473 2876
rect 3415 2867 3473 2873
rect 3510 2864 3516 2876
rect 3568 2904 3574 2916
rect 5178 2913 5206 3080
rect 5626 3000 5632 3052
rect 5684 3040 5690 3052
rect 7161 3040 7189 3148
rect 9766 3136 9772 3148
rect 9824 3176 9830 3188
rect 10229 3179 10287 3185
rect 10229 3176 10241 3179
rect 9824 3148 10241 3176
rect 9824 3136 9830 3148
rect 10229 3145 10241 3148
rect 10275 3145 10287 3179
rect 12250 3176 12256 3188
rect 12211 3148 12256 3176
rect 10229 3139 10287 3145
rect 12250 3136 12256 3148
rect 12308 3136 12314 3188
rect 12437 3179 12495 3185
rect 12437 3145 12449 3179
rect 12483 3176 12495 3179
rect 13630 3176 13636 3188
rect 12483 3148 13308 3176
rect 13591 3148 13636 3176
rect 12483 3145 12495 3148
rect 12437 3139 12495 3145
rect 7282 3068 7288 3120
rect 7340 3108 7346 3120
rect 7791 3111 7849 3117
rect 7791 3108 7803 3111
rect 7340 3080 7803 3108
rect 7340 3068 7346 3080
rect 7791 3077 7803 3080
rect 7837 3077 7849 3111
rect 7926 3108 7932 3120
rect 7887 3080 7932 3108
rect 7791 3071 7849 3077
rect 7926 3068 7932 3080
rect 7984 3068 7990 3120
rect 12710 3108 12716 3120
rect 9048 3080 12716 3108
rect 5684 3012 7189 3040
rect 5684 3000 5690 3012
rect 7466 3000 7472 3052
rect 7524 3040 7530 3052
rect 8021 3043 8079 3049
rect 8021 3040 8033 3043
rect 7524 3012 8033 3040
rect 7524 3000 7530 3012
rect 8021 3009 8033 3012
rect 8067 3040 8079 3043
rect 8202 3040 8208 3052
rect 8067 3012 8208 3040
rect 8067 3009 8079 3012
rect 8021 3003 8079 3009
rect 8202 3000 8208 3012
rect 8260 3040 8266 3052
rect 8665 3043 8723 3049
rect 8665 3040 8677 3043
rect 8260 3012 8677 3040
rect 8260 3000 8266 3012
rect 8665 3009 8677 3012
rect 8711 3009 8723 3043
rect 8665 3003 8723 3009
rect 5721 2975 5779 2981
rect 5721 2941 5733 2975
rect 5767 2972 5779 2975
rect 9048 2972 9076 3080
rect 12710 3068 12716 3080
rect 12768 3068 12774 3120
rect 13170 3108 13176 3120
rect 13131 3080 13176 3108
rect 13170 3068 13176 3080
rect 13228 3068 13234 3120
rect 13280 3108 13308 3148
rect 13630 3136 13636 3148
rect 13688 3136 13694 3188
rect 15286 3176 15292 3188
rect 13786 3148 14964 3176
rect 15247 3148 15292 3176
rect 13786 3108 13814 3148
rect 14734 3108 14740 3120
rect 13280 3080 13814 3108
rect 14695 3080 14740 3108
rect 14734 3068 14740 3080
rect 14792 3068 14798 3120
rect 14936 3108 14964 3148
rect 15286 3136 15292 3148
rect 15344 3136 15350 3188
rect 15654 3176 15660 3188
rect 15615 3148 15660 3176
rect 15654 3136 15660 3148
rect 15712 3136 15718 3188
rect 17402 3176 17408 3188
rect 17363 3148 17408 3176
rect 17402 3136 17408 3148
rect 17460 3136 17466 3188
rect 18874 3136 18880 3188
rect 18932 3176 18938 3188
rect 20165 3179 20223 3185
rect 20165 3176 20177 3179
rect 18932 3148 20177 3176
rect 18932 3136 18938 3148
rect 20165 3145 20177 3148
rect 20211 3145 20223 3179
rect 20165 3139 20223 3145
rect 23474 3136 23480 3188
rect 23532 3176 23538 3188
rect 24213 3179 24271 3185
rect 24213 3176 24225 3179
rect 23532 3148 24225 3176
rect 23532 3136 23538 3148
rect 24213 3145 24225 3148
rect 24259 3145 24271 3179
rect 24213 3139 24271 3145
rect 26878 3136 26884 3188
rect 26936 3176 26942 3188
rect 27065 3179 27123 3185
rect 27065 3176 27077 3179
rect 26936 3148 27077 3176
rect 26936 3136 26942 3148
rect 27065 3145 27077 3148
rect 27111 3145 27123 3179
rect 30834 3176 30840 3188
rect 30795 3148 30840 3176
rect 27065 3139 27123 3145
rect 30834 3136 30840 3148
rect 30892 3136 30898 3188
rect 31294 3176 31300 3188
rect 31255 3148 31300 3176
rect 31294 3136 31300 3148
rect 31352 3136 31358 3188
rect 32214 3136 32220 3188
rect 32272 3176 32278 3188
rect 32723 3179 32781 3185
rect 32723 3176 32735 3179
rect 32272 3148 32735 3176
rect 32272 3136 32278 3148
rect 32723 3145 32735 3148
rect 32769 3145 32781 3179
rect 32723 3139 32781 3145
rect 16301 3111 16359 3117
rect 16301 3108 16313 3111
rect 14936 3080 16313 3108
rect 16301 3077 16313 3080
rect 16347 3108 16359 3111
rect 17310 3108 17316 3120
rect 16347 3080 17316 3108
rect 16347 3077 16359 3080
rect 16301 3071 16359 3077
rect 17310 3068 17316 3080
rect 17368 3068 17374 3120
rect 17420 3108 17448 3136
rect 19242 3108 19248 3120
rect 17420 3080 19248 3108
rect 19242 3068 19248 3080
rect 19300 3068 19306 3120
rect 23937 3111 23995 3117
rect 23937 3077 23949 3111
rect 23983 3108 23995 3111
rect 24026 3108 24032 3120
rect 23983 3080 24032 3108
rect 23983 3077 23995 3080
rect 23937 3071 23995 3077
rect 24026 3068 24032 3080
rect 24084 3068 24090 3120
rect 33137 3111 33195 3117
rect 33137 3077 33149 3111
rect 33183 3108 33195 3111
rect 33226 3108 33232 3120
rect 33183 3080 33232 3108
rect 33183 3077 33195 3080
rect 33137 3071 33195 3077
rect 9122 3000 9128 3052
rect 9180 3040 9186 3052
rect 9309 3043 9367 3049
rect 9309 3040 9321 3043
rect 9180 3012 9321 3040
rect 9180 3000 9186 3012
rect 9309 3009 9321 3012
rect 9355 3009 9367 3043
rect 9309 3003 9367 3009
rect 9953 3043 10011 3049
rect 9953 3009 9965 3043
rect 9999 3040 10011 3043
rect 11149 3043 11207 3049
rect 11149 3040 11161 3043
rect 9999 3012 11161 3040
rect 9999 3009 10011 3012
rect 9953 3003 10011 3009
rect 11149 3009 11161 3012
rect 11195 3040 11207 3043
rect 16482 3040 16488 3052
rect 11195 3012 16488 3040
rect 11195 3009 11207 3012
rect 11149 3003 11207 3009
rect 16482 3000 16488 3012
rect 16540 3000 16546 3052
rect 24949 3043 25007 3049
rect 19076 3012 20576 3040
rect 5767 2944 9076 2972
rect 5767 2941 5779 2944
rect 5721 2935 5779 2941
rect 11514 2932 11520 2984
rect 11572 2972 11578 2984
rect 11885 2975 11943 2981
rect 11885 2972 11897 2975
rect 11572 2944 11897 2972
rect 11572 2932 11578 2944
rect 11885 2941 11897 2944
rect 11931 2972 11943 2975
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 11931 2944 12449 2972
rect 11931 2941 11943 2944
rect 11885 2935 11943 2941
rect 12437 2941 12449 2944
rect 12483 2941 12495 2975
rect 12437 2935 12495 2941
rect 17310 2932 17316 2984
rect 17368 2972 17374 2984
rect 17865 2975 17923 2981
rect 17865 2972 17877 2975
rect 17368 2944 17877 2972
rect 17368 2932 17374 2944
rect 17865 2941 17877 2944
rect 17911 2972 17923 2975
rect 18322 2972 18328 2984
rect 17911 2944 18328 2972
rect 17911 2941 17923 2944
rect 17865 2935 17923 2941
rect 18322 2932 18328 2944
rect 18380 2932 18386 2984
rect 18414 2932 18420 2984
rect 18472 2972 18478 2984
rect 18509 2975 18567 2981
rect 18509 2972 18521 2975
rect 18472 2944 18521 2972
rect 18472 2932 18478 2944
rect 18509 2941 18521 2944
rect 18555 2941 18567 2975
rect 18874 2972 18880 2984
rect 18835 2944 18880 2972
rect 18509 2935 18567 2941
rect 18874 2932 18880 2944
rect 18932 2932 18938 2984
rect 19076 2916 19104 3012
rect 19242 2972 19248 2984
rect 19203 2944 19248 2972
rect 19242 2932 19248 2944
rect 19300 2932 19306 2984
rect 19334 2932 19340 2984
rect 19392 2972 19398 2984
rect 20441 2975 20499 2981
rect 20441 2972 20453 2975
rect 19392 2944 20453 2972
rect 19392 2932 19398 2944
rect 20441 2941 20453 2944
rect 20487 2941 20499 2975
rect 20548 2972 20576 3012
rect 24949 3009 24961 3043
rect 24995 3040 25007 3043
rect 25133 3043 25191 3049
rect 25133 3040 25145 3043
rect 24995 3012 25145 3040
rect 24995 3009 25007 3012
rect 24949 3003 25007 3009
rect 25133 3009 25145 3012
rect 25179 3040 25191 3043
rect 25222 3040 25228 3052
rect 25179 3012 25228 3040
rect 25179 3009 25191 3012
rect 25133 3003 25191 3009
rect 25222 3000 25228 3012
rect 25280 3000 25286 3052
rect 21948 2975 22006 2981
rect 21948 2972 21960 2975
rect 20548 2944 21960 2972
rect 20441 2935 20499 2941
rect 21948 2941 21960 2944
rect 21994 2972 22006 2975
rect 22373 2975 22431 2981
rect 22373 2972 22385 2975
rect 21994 2944 22385 2972
rect 21994 2941 22006 2944
rect 21948 2935 22006 2941
rect 22373 2941 22385 2944
rect 22419 2941 22431 2975
rect 22373 2935 22431 2941
rect 25777 2975 25835 2981
rect 25777 2941 25789 2975
rect 25823 2972 25835 2975
rect 26672 2975 26730 2981
rect 26672 2972 26684 2975
rect 25823 2944 26684 2972
rect 25823 2941 25835 2944
rect 25777 2935 25835 2941
rect 26672 2941 26684 2944
rect 26718 2972 26730 2975
rect 26878 2972 26884 2984
rect 26718 2944 26884 2972
rect 26718 2941 26730 2944
rect 26672 2935 26730 2941
rect 5163 2907 5221 2913
rect 5163 2904 5175 2907
rect 3568 2876 5175 2904
rect 3568 2864 3574 2876
rect 5163 2873 5175 2876
rect 5209 2873 5221 2907
rect 5163 2867 5221 2873
rect 5902 2864 5908 2916
rect 5960 2904 5966 2916
rect 7653 2907 7711 2913
rect 7653 2904 7665 2907
rect 5960 2876 7665 2904
rect 5960 2864 5966 2876
rect 7653 2873 7665 2876
rect 7699 2904 7711 2907
rect 8202 2904 8208 2916
rect 7699 2876 8208 2904
rect 7699 2873 7711 2876
rect 7653 2867 7711 2873
rect 8202 2864 8208 2876
rect 8260 2864 8266 2916
rect 8386 2904 8392 2916
rect 8347 2876 8392 2904
rect 8386 2864 8392 2876
rect 8444 2864 8450 2916
rect 9030 2904 9036 2916
rect 8991 2876 9036 2904
rect 9030 2864 9036 2876
rect 9088 2864 9094 2916
rect 9398 2904 9404 2916
rect 9359 2876 9404 2904
rect 9398 2864 9404 2876
rect 9456 2864 9462 2916
rect 10870 2904 10876 2916
rect 10831 2876 10876 2904
rect 10870 2864 10876 2876
rect 10928 2864 10934 2916
rect 10962 2864 10968 2916
rect 11020 2904 11026 2916
rect 12621 2907 12679 2913
rect 11020 2876 11065 2904
rect 11020 2864 11026 2876
rect 12621 2873 12633 2907
rect 12667 2873 12679 2907
rect 12621 2867 12679 2873
rect 2406 2836 2412 2848
rect 2367 2808 2412 2836
rect 2406 2796 2412 2808
rect 2464 2796 2470 2848
rect 3050 2796 3056 2848
rect 3108 2836 3114 2848
rect 3973 2839 4031 2845
rect 3973 2836 3985 2839
rect 3108 2808 3985 2836
rect 3108 2796 3114 2808
rect 3973 2805 3985 2808
rect 4019 2805 4031 2839
rect 7190 2836 7196 2848
rect 7151 2808 7196 2836
rect 3973 2799 4031 2805
rect 7190 2796 7196 2808
rect 7248 2836 7254 2848
rect 7285 2839 7343 2845
rect 7285 2836 7297 2839
rect 7248 2808 7297 2836
rect 7248 2796 7254 2808
rect 7285 2805 7297 2808
rect 7331 2805 7343 2839
rect 7466 2836 7472 2848
rect 7427 2808 7472 2836
rect 7285 2799 7343 2805
rect 7466 2796 7472 2808
rect 7524 2796 7530 2848
rect 10689 2839 10747 2845
rect 10689 2805 10701 2839
rect 10735 2836 10747 2839
rect 10980 2836 11008 2864
rect 10735 2808 11008 2836
rect 12636 2836 12664 2867
rect 12710 2864 12716 2916
rect 12768 2904 12774 2916
rect 14182 2904 14188 2916
rect 12768 2876 13814 2904
rect 14143 2876 14188 2904
rect 12768 2864 12774 2876
rect 12802 2836 12808 2848
rect 12636 2808 12808 2836
rect 10735 2805 10747 2808
rect 10689 2799 10747 2805
rect 12802 2796 12808 2808
rect 12860 2796 12866 2848
rect 13786 2836 13814 2876
rect 14182 2864 14188 2876
rect 14240 2864 14246 2916
rect 14277 2907 14335 2913
rect 14277 2873 14289 2907
rect 14323 2873 14335 2907
rect 14277 2867 14335 2873
rect 16577 2907 16635 2913
rect 16577 2873 16589 2907
rect 16623 2904 16635 2907
rect 16942 2904 16948 2916
rect 16623 2876 16948 2904
rect 16623 2873 16635 2876
rect 16577 2867 16635 2873
rect 14001 2839 14059 2845
rect 14001 2836 14013 2839
rect 13786 2808 14013 2836
rect 14001 2805 14013 2808
rect 14047 2836 14059 2839
rect 14292 2836 14320 2867
rect 16942 2864 16948 2876
rect 17000 2864 17006 2916
rect 17129 2907 17187 2913
rect 17129 2873 17141 2907
rect 17175 2904 17187 2907
rect 19058 2904 19064 2916
rect 17175 2876 19064 2904
rect 17175 2873 17187 2876
rect 17129 2867 17187 2873
rect 19058 2864 19064 2876
rect 19116 2864 19122 2916
rect 20346 2904 20352 2916
rect 20307 2876 20352 2904
rect 20346 2864 20352 2876
rect 20404 2864 20410 2916
rect 20456 2904 20484 2935
rect 26878 2932 26884 2944
rect 26936 2932 26942 2984
rect 30834 2932 30840 2984
rect 30892 2972 30898 2984
rect 31113 2975 31171 2981
rect 31113 2972 31125 2975
rect 30892 2944 31125 2972
rect 30892 2932 30898 2944
rect 31113 2941 31125 2944
rect 31159 2972 31171 2975
rect 32125 2975 32183 2981
rect 32125 2972 32137 2975
rect 31159 2944 32137 2972
rect 31159 2941 31171 2944
rect 31113 2935 31171 2941
rect 32125 2941 32137 2944
rect 32171 2972 32183 2975
rect 32306 2972 32312 2984
rect 32171 2944 32312 2972
rect 32171 2941 32183 2944
rect 32125 2935 32183 2941
rect 32306 2932 32312 2944
rect 32364 2932 32370 2984
rect 32652 2975 32710 2981
rect 32652 2941 32664 2975
rect 32698 2972 32710 2975
rect 33152 2972 33180 3071
rect 33226 3068 33232 3080
rect 33284 3108 33290 3120
rect 34698 3108 34704 3120
rect 33284 3080 34704 3108
rect 33284 3068 33290 3080
rect 34698 3068 34704 3080
rect 34756 3068 34762 3120
rect 32698 2944 33180 2972
rect 32698 2941 32710 2944
rect 32652 2935 32710 2941
rect 21729 2907 21787 2913
rect 21729 2904 21741 2907
rect 20456 2876 21741 2904
rect 21729 2873 21741 2876
rect 21775 2873 21787 2907
rect 21729 2867 21787 2873
rect 24578 2864 24584 2916
rect 24636 2904 24642 2916
rect 25130 2904 25136 2916
rect 24636 2876 25136 2904
rect 24636 2864 24642 2876
rect 25130 2864 25136 2876
rect 25188 2904 25194 2916
rect 25225 2907 25283 2913
rect 25225 2904 25237 2907
rect 25188 2876 25237 2904
rect 25188 2864 25194 2876
rect 25225 2873 25237 2876
rect 25271 2873 25283 2907
rect 25225 2867 25283 2873
rect 14047 2808 14320 2836
rect 14047 2805 14059 2808
rect 14001 2799 14059 2805
rect 17862 2796 17868 2848
rect 17920 2836 17926 2848
rect 18141 2839 18199 2845
rect 18141 2836 18153 2839
rect 17920 2808 18153 2836
rect 17920 2796 17926 2808
rect 18141 2805 18153 2808
rect 18187 2805 18199 2839
rect 18141 2799 18199 2805
rect 18414 2796 18420 2848
rect 18472 2836 18478 2848
rect 19797 2839 19855 2845
rect 19797 2836 19809 2839
rect 18472 2808 19809 2836
rect 18472 2796 18478 2808
rect 19797 2805 19809 2808
rect 19843 2805 19855 2839
rect 21450 2836 21456 2848
rect 21411 2808 21456 2836
rect 19797 2799 19855 2805
rect 21450 2796 21456 2808
rect 21508 2796 21514 2848
rect 22051 2839 22109 2845
rect 22051 2805 22063 2839
rect 22097 2836 22109 2839
rect 22278 2836 22284 2848
rect 22097 2808 22284 2836
rect 22097 2805 22109 2808
rect 22051 2799 22109 2805
rect 22278 2796 22284 2808
rect 22336 2796 22342 2848
rect 26743 2839 26801 2845
rect 26743 2805 26755 2839
rect 26789 2836 26801 2839
rect 29914 2836 29920 2848
rect 26789 2808 29920 2836
rect 26789 2805 26801 2808
rect 26743 2799 26801 2805
rect 29914 2796 29920 2808
rect 29972 2796 29978 2848
rect 1104 2746 38824 2768
rect 1104 2694 14315 2746
rect 14367 2694 14379 2746
rect 14431 2694 14443 2746
rect 14495 2694 14507 2746
rect 14559 2694 27648 2746
rect 27700 2694 27712 2746
rect 27764 2694 27776 2746
rect 27828 2694 27840 2746
rect 27892 2694 38824 2746
rect 1104 2672 38824 2694
rect 1581 2635 1639 2641
rect 1581 2601 1593 2635
rect 1627 2632 1639 2635
rect 3694 2632 3700 2644
rect 1627 2604 3700 2632
rect 1627 2601 1639 2604
rect 1581 2595 1639 2601
rect 3694 2592 3700 2604
rect 3752 2592 3758 2644
rect 3878 2632 3884 2644
rect 3839 2604 3884 2632
rect 3878 2592 3884 2604
rect 3936 2592 3942 2644
rect 4157 2635 4215 2641
rect 4157 2601 4169 2635
rect 4203 2632 4215 2635
rect 4433 2635 4491 2641
rect 4433 2632 4445 2635
rect 4203 2604 4445 2632
rect 4203 2601 4215 2604
rect 4157 2595 4215 2601
rect 4433 2601 4445 2604
rect 4479 2632 4491 2635
rect 5350 2632 5356 2644
rect 4479 2604 5356 2632
rect 4479 2601 4491 2604
rect 4433 2595 4491 2601
rect 5350 2592 5356 2604
rect 5408 2592 5414 2644
rect 7098 2632 7104 2644
rect 7059 2604 7104 2632
rect 7098 2592 7104 2604
rect 7156 2592 7162 2644
rect 9953 2635 10011 2641
rect 9953 2601 9965 2635
rect 9999 2632 10011 2635
rect 10686 2632 10692 2644
rect 9999 2604 10692 2632
rect 9999 2601 10011 2604
rect 9953 2595 10011 2601
rect 10686 2592 10692 2604
rect 10744 2592 10750 2644
rect 10888 2604 11192 2632
rect 2406 2564 2412 2576
rect 2367 2536 2412 2564
rect 2406 2524 2412 2536
rect 2464 2524 2470 2576
rect 6365 2567 6423 2573
rect 6365 2533 6377 2567
rect 6411 2564 6423 2567
rect 8294 2564 8300 2576
rect 6411 2536 8300 2564
rect 6411 2533 6423 2536
rect 6365 2527 6423 2533
rect 1394 2496 1400 2508
rect 1355 2468 1400 2496
rect 1394 2456 1400 2468
rect 1452 2496 1458 2508
rect 1857 2499 1915 2505
rect 1857 2496 1869 2499
rect 1452 2468 1869 2496
rect 1452 2456 1458 2468
rect 1857 2465 1869 2468
rect 1903 2496 1915 2499
rect 2225 2499 2283 2505
rect 2225 2496 2237 2499
rect 1903 2468 2237 2496
rect 1903 2465 1915 2468
rect 1857 2459 1915 2465
rect 2225 2465 2237 2468
rect 2271 2465 2283 2499
rect 3050 2496 3056 2508
rect 3011 2468 3056 2496
rect 2225 2459 2283 2465
rect 3050 2456 3056 2468
rect 3108 2456 3114 2508
rect 4249 2499 4307 2505
rect 4249 2465 4261 2499
rect 4295 2496 4307 2499
rect 4525 2499 4583 2505
rect 4525 2496 4537 2499
rect 4295 2468 4537 2496
rect 4295 2465 4307 2468
rect 4249 2459 4307 2465
rect 4525 2465 4537 2468
rect 4571 2465 4583 2499
rect 4525 2459 4583 2465
rect 5169 2499 5227 2505
rect 5169 2465 5181 2499
rect 5215 2496 5227 2499
rect 5353 2499 5411 2505
rect 5353 2496 5365 2499
rect 5215 2468 5365 2496
rect 5215 2465 5227 2468
rect 5169 2459 5227 2465
rect 5353 2465 5365 2468
rect 5399 2465 5411 2499
rect 5353 2459 5411 2465
rect 6733 2499 6791 2505
rect 6733 2465 6745 2499
rect 6779 2496 6791 2499
rect 6914 2496 6920 2508
rect 6779 2468 6920 2496
rect 6779 2465 6791 2468
rect 6733 2459 6791 2465
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 5184 2428 5212 2459
rect 6914 2456 6920 2468
rect 6972 2456 6978 2508
rect 7469 2499 7527 2505
rect 7469 2465 7481 2499
rect 7515 2496 7527 2499
rect 7926 2496 7932 2508
rect 7515 2468 7932 2496
rect 7515 2465 7527 2468
rect 7469 2459 7527 2465
rect 1360 2400 5212 2428
rect 5997 2431 6055 2437
rect 1360 2388 1366 2400
rect 5997 2397 6009 2431
rect 6043 2428 6055 2431
rect 7484 2428 7512 2459
rect 7926 2456 7932 2468
rect 7984 2456 7990 2508
rect 8091 2505 8119 2536
rect 8294 2524 8300 2536
rect 8352 2524 8358 2576
rect 10594 2564 10600 2576
rect 10555 2536 10600 2564
rect 10594 2524 10600 2536
rect 10652 2524 10658 2576
rect 8076 2499 8134 2505
rect 8076 2465 8088 2499
rect 8122 2465 8134 2499
rect 8076 2459 8134 2465
rect 8386 2456 8392 2508
rect 8444 2496 8450 2508
rect 9769 2499 9827 2505
rect 9769 2496 9781 2499
rect 8444 2468 9781 2496
rect 8444 2456 8450 2468
rect 9769 2465 9781 2468
rect 9815 2496 9827 2499
rect 10229 2499 10287 2505
rect 10229 2496 10241 2499
rect 9815 2468 10241 2496
rect 9815 2465 9827 2468
rect 9769 2459 9827 2465
rect 10229 2465 10241 2468
rect 10275 2465 10287 2499
rect 10612 2496 10640 2524
rect 10888 2496 10916 2604
rect 11164 2573 11192 2604
rect 11238 2592 11244 2644
rect 11296 2632 11302 2644
rect 12434 2632 12440 2644
rect 11296 2604 12440 2632
rect 11296 2592 11302 2604
rect 12434 2592 12440 2604
rect 12492 2592 12498 2644
rect 12802 2592 12808 2644
rect 12860 2632 12866 2644
rect 14185 2635 14243 2641
rect 14185 2632 14197 2635
rect 12860 2604 14197 2632
rect 12860 2592 12866 2604
rect 14185 2601 14197 2604
rect 14231 2601 14243 2635
rect 16298 2632 16304 2644
rect 16259 2604 16304 2632
rect 14185 2595 14243 2601
rect 16298 2592 16304 2604
rect 16356 2632 16362 2644
rect 16356 2604 16849 2632
rect 16356 2592 16362 2604
rect 11143 2567 11201 2573
rect 11143 2533 11155 2567
rect 11189 2533 11201 2567
rect 11143 2527 11201 2533
rect 11882 2524 11888 2576
rect 11940 2564 11946 2576
rect 11977 2567 12035 2573
rect 11977 2564 11989 2567
rect 11940 2536 11989 2564
rect 11940 2524 11946 2536
rect 11977 2533 11989 2536
rect 12023 2533 12035 2567
rect 12986 2564 12992 2576
rect 12947 2536 12992 2564
rect 11977 2527 12035 2533
rect 12986 2524 12992 2536
rect 13044 2564 13050 2576
rect 13357 2567 13415 2573
rect 13357 2564 13369 2567
rect 13044 2536 13369 2564
rect 13044 2524 13050 2536
rect 13357 2533 13369 2536
rect 13403 2533 13415 2567
rect 13357 2527 13415 2533
rect 13909 2567 13967 2573
rect 13909 2533 13921 2567
rect 13955 2564 13967 2567
rect 14734 2564 14740 2576
rect 13955 2536 14740 2564
rect 13955 2533 13967 2536
rect 13909 2527 13967 2533
rect 14734 2524 14740 2536
rect 14792 2524 14798 2576
rect 16821 2573 16849 2604
rect 16942 2592 16948 2644
rect 17000 2632 17006 2644
rect 17405 2635 17463 2641
rect 17405 2632 17417 2635
rect 17000 2604 17417 2632
rect 17000 2592 17006 2604
rect 17405 2601 17417 2604
rect 17451 2632 17463 2635
rect 19334 2632 19340 2644
rect 17451 2604 19340 2632
rect 17451 2601 17463 2604
rect 17405 2595 17463 2601
rect 19334 2592 19340 2604
rect 19392 2592 19398 2644
rect 19889 2635 19947 2641
rect 19889 2601 19901 2635
rect 19935 2632 19947 2635
rect 25130 2632 25136 2644
rect 19935 2604 20668 2632
rect 25091 2604 25136 2632
rect 19935 2601 19947 2604
rect 19889 2595 19947 2601
rect 14921 2567 14979 2573
rect 14921 2533 14933 2567
rect 14967 2564 14979 2567
rect 16806 2567 16864 2573
rect 14967 2536 16528 2564
rect 14967 2533 14979 2536
rect 14921 2527 14979 2533
rect 11698 2496 11704 2508
rect 10612 2468 10916 2496
rect 11659 2468 11704 2496
rect 10229 2459 10287 2465
rect 11698 2456 11704 2468
rect 11756 2456 11762 2508
rect 15194 2456 15200 2508
rect 15252 2496 15258 2508
rect 16500 2505 16528 2536
rect 16806 2533 16818 2567
rect 16852 2533 16864 2567
rect 16806 2527 16864 2533
rect 17126 2524 17132 2576
rect 17184 2564 17190 2576
rect 17681 2567 17739 2573
rect 17681 2564 17693 2567
rect 17184 2536 17693 2564
rect 17184 2524 17190 2536
rect 17681 2533 17693 2536
rect 17727 2533 17739 2567
rect 17681 2527 17739 2533
rect 18141 2567 18199 2573
rect 18141 2533 18153 2567
rect 18187 2564 18199 2567
rect 18509 2567 18567 2573
rect 18509 2564 18521 2567
rect 18187 2536 18521 2564
rect 18187 2533 18199 2536
rect 18141 2527 18199 2533
rect 18509 2533 18521 2536
rect 18555 2564 18567 2567
rect 20346 2564 20352 2576
rect 18555 2536 20352 2564
rect 18555 2533 18567 2536
rect 18509 2527 18567 2533
rect 20346 2524 20352 2536
rect 20404 2524 20410 2576
rect 20640 2573 20668 2604
rect 25130 2592 25136 2604
rect 25188 2592 25194 2644
rect 32214 2632 32220 2644
rect 32175 2604 32220 2632
rect 32214 2592 32220 2604
rect 32272 2592 32278 2644
rect 33226 2632 33232 2644
rect 33187 2604 33232 2632
rect 33226 2592 33232 2604
rect 33284 2592 33290 2644
rect 20625 2567 20683 2573
rect 20625 2533 20637 2567
rect 20671 2564 20683 2567
rect 21450 2564 21456 2576
rect 20671 2536 21456 2564
rect 20671 2533 20683 2536
rect 20625 2527 20683 2533
rect 21450 2524 21456 2536
rect 21508 2524 21514 2576
rect 15540 2499 15598 2505
rect 15540 2496 15552 2499
rect 15252 2468 15552 2496
rect 15252 2456 15258 2468
rect 15540 2465 15552 2468
rect 15586 2496 15598 2499
rect 15933 2499 15991 2505
rect 15933 2496 15945 2499
rect 15586 2468 15945 2496
rect 15586 2465 15598 2468
rect 15540 2459 15598 2465
rect 15933 2465 15945 2468
rect 15979 2465 15991 2499
rect 15933 2459 15991 2465
rect 16485 2499 16543 2505
rect 16485 2465 16497 2499
rect 16531 2496 16543 2499
rect 17862 2496 17868 2508
rect 16531 2468 17868 2496
rect 16531 2465 16543 2468
rect 16485 2459 16543 2465
rect 17862 2456 17868 2468
rect 17920 2456 17926 2508
rect 19058 2456 19064 2508
rect 19116 2496 19122 2508
rect 19889 2499 19947 2505
rect 19116 2468 19161 2496
rect 19116 2456 19122 2468
rect 19889 2465 19901 2499
rect 19935 2496 19947 2499
rect 19981 2499 20039 2505
rect 19981 2496 19993 2499
rect 19935 2468 19993 2496
rect 19935 2465 19947 2468
rect 19889 2459 19947 2465
rect 19981 2465 19993 2468
rect 20027 2465 20039 2499
rect 19981 2459 20039 2465
rect 20070 2456 20076 2508
rect 20128 2496 20134 2508
rect 21177 2499 21235 2505
rect 21177 2496 21189 2499
rect 20128 2468 21189 2496
rect 20128 2456 20134 2468
rect 21177 2465 21189 2468
rect 21223 2465 21235 2499
rect 21177 2459 21235 2465
rect 21266 2456 21272 2508
rect 21324 2496 21330 2508
rect 22189 2499 22247 2505
rect 22189 2496 22201 2499
rect 21324 2468 22201 2496
rect 21324 2456 21330 2468
rect 22189 2465 22201 2468
rect 22235 2465 22247 2499
rect 22189 2459 22247 2465
rect 25498 2456 25504 2508
rect 25556 2496 25562 2508
rect 29733 2499 29791 2505
rect 29733 2496 29745 2499
rect 25556 2468 29745 2496
rect 25556 2456 25562 2468
rect 29733 2465 29745 2468
rect 29779 2496 29791 2499
rect 30285 2499 30343 2505
rect 30285 2496 30297 2499
rect 29779 2468 30297 2496
rect 29779 2465 29791 2468
rect 29733 2459 29791 2465
rect 30285 2465 30297 2468
rect 30331 2465 30343 2499
rect 30285 2459 30343 2465
rect 32585 2499 32643 2505
rect 32585 2465 32597 2499
rect 32631 2496 32643 2499
rect 33244 2496 33272 2592
rect 32631 2468 33272 2496
rect 32631 2465 32643 2468
rect 32585 2459 32643 2465
rect 8297 2431 8355 2437
rect 8297 2428 8309 2431
rect 6043 2400 7512 2428
rect 8036 2400 8309 2428
rect 6043 2397 6055 2400
rect 5997 2391 6055 2397
rect 3513 2363 3571 2369
rect 3513 2329 3525 2363
rect 3559 2360 3571 2363
rect 4525 2363 4583 2369
rect 3559 2332 3924 2360
rect 3559 2329 3571 2332
rect 3513 2323 3571 2329
rect 3896 2292 3924 2332
rect 4525 2329 4537 2363
rect 4571 2360 4583 2363
rect 4801 2363 4859 2369
rect 4801 2360 4813 2363
rect 4571 2332 4813 2360
rect 4571 2329 4583 2332
rect 4525 2323 4583 2329
rect 4801 2329 4813 2332
rect 4847 2360 4859 2363
rect 5626 2360 5632 2372
rect 4847 2332 5632 2360
rect 4847 2329 4859 2332
rect 4801 2323 4859 2329
rect 5626 2320 5632 2332
rect 5684 2320 5690 2372
rect 4157 2295 4215 2301
rect 4157 2292 4169 2295
rect 3896 2264 4169 2292
rect 4157 2261 4169 2264
rect 4203 2261 4215 2295
rect 4157 2255 4215 2261
rect 7190 2252 7196 2304
rect 7248 2292 7254 2304
rect 7837 2295 7895 2301
rect 7837 2292 7849 2295
rect 7248 2264 7849 2292
rect 7248 2252 7254 2264
rect 7837 2261 7849 2264
rect 7883 2292 7895 2295
rect 8036 2292 8064 2400
rect 8297 2397 8309 2400
rect 8343 2397 8355 2431
rect 8662 2428 8668 2440
rect 8623 2400 8668 2428
rect 8297 2391 8355 2397
rect 8662 2388 8668 2400
rect 8720 2388 8726 2440
rect 10781 2431 10839 2437
rect 10781 2397 10793 2431
rect 10827 2428 10839 2431
rect 11054 2428 11060 2440
rect 10827 2400 11060 2428
rect 10827 2397 10839 2400
rect 10781 2391 10839 2397
rect 11054 2388 11060 2400
rect 11112 2388 11118 2440
rect 13265 2431 13323 2437
rect 13265 2397 13277 2431
rect 13311 2428 13323 2431
rect 14918 2428 14924 2440
rect 13311 2400 14924 2428
rect 13311 2397 13323 2400
rect 13265 2391 13323 2397
rect 14918 2388 14924 2400
rect 14976 2388 14982 2440
rect 15289 2431 15347 2437
rect 15289 2397 15301 2431
rect 15335 2428 15347 2431
rect 16942 2428 16948 2440
rect 15335 2400 16948 2428
rect 15335 2397 15347 2400
rect 15289 2391 15347 2397
rect 16942 2388 16948 2400
rect 17000 2388 17006 2440
rect 18417 2431 18475 2437
rect 18417 2397 18429 2431
rect 18463 2428 18475 2431
rect 20901 2431 20959 2437
rect 20901 2428 20913 2431
rect 18463 2400 20913 2428
rect 18463 2397 18475 2400
rect 18417 2391 18475 2397
rect 20901 2397 20913 2400
rect 20947 2428 20959 2431
rect 22741 2431 22799 2437
rect 22741 2428 22753 2431
rect 20947 2400 22753 2428
rect 20947 2397 20959 2400
rect 20901 2391 20959 2397
rect 22741 2397 22753 2400
rect 22787 2397 22799 2431
rect 22741 2391 22799 2397
rect 8202 2360 8208 2372
rect 8163 2332 8208 2360
rect 8202 2320 8208 2332
rect 8260 2360 8266 2372
rect 8941 2363 8999 2369
rect 8941 2360 8953 2363
rect 8260 2332 8953 2360
rect 8260 2320 8266 2332
rect 8941 2329 8953 2332
rect 8987 2360 8999 2363
rect 9309 2363 9367 2369
rect 9309 2360 9321 2363
rect 8987 2332 9321 2360
rect 8987 2329 8999 2332
rect 8941 2323 8999 2329
rect 9309 2329 9321 2332
rect 9355 2329 9367 2363
rect 9309 2323 9367 2329
rect 10870 2320 10876 2372
rect 10928 2360 10934 2372
rect 11974 2360 11980 2372
rect 10928 2332 11980 2360
rect 10928 2320 10934 2332
rect 11974 2320 11980 2332
rect 12032 2360 12038 2372
rect 15611 2363 15669 2369
rect 15611 2360 15623 2363
rect 12032 2332 15623 2360
rect 12032 2320 12038 2332
rect 15611 2329 15623 2332
rect 15657 2329 15669 2363
rect 15611 2323 15669 2329
rect 18874 2320 18880 2372
rect 18932 2360 18938 2372
rect 19337 2363 19395 2369
rect 19337 2360 19349 2363
rect 18932 2332 19349 2360
rect 18932 2320 18938 2332
rect 19337 2329 19349 2332
rect 19383 2329 19395 2363
rect 19337 2323 19395 2329
rect 20165 2363 20223 2369
rect 20165 2329 20177 2363
rect 20211 2360 20223 2363
rect 22370 2360 22376 2372
rect 20211 2332 22376 2360
rect 20211 2329 20223 2332
rect 20165 2323 20223 2329
rect 22370 2320 22376 2332
rect 22428 2320 22434 2372
rect 29917 2363 29975 2369
rect 29917 2329 29929 2363
rect 29963 2360 29975 2363
rect 31754 2360 31760 2372
rect 29963 2332 31760 2360
rect 29963 2329 29975 2332
rect 29917 2323 29975 2329
rect 31754 2320 31760 2332
rect 31812 2320 31818 2372
rect 32769 2363 32827 2369
rect 32769 2329 32781 2363
rect 32815 2360 32827 2363
rect 34146 2360 34152 2372
rect 32815 2332 34152 2360
rect 32815 2329 32827 2332
rect 32769 2323 32827 2329
rect 34146 2320 34152 2332
rect 34204 2320 34210 2372
rect 11514 2292 11520 2304
rect 7883 2264 11520 2292
rect 7883 2261 7895 2264
rect 7837 2255 7895 2261
rect 11514 2252 11520 2264
rect 11572 2252 11578 2304
rect 18230 2252 18236 2304
rect 18288 2292 18294 2304
rect 19705 2295 19763 2301
rect 19705 2292 19717 2295
rect 18288 2264 19717 2292
rect 18288 2252 18294 2264
rect 19705 2261 19717 2264
rect 19751 2261 19763 2295
rect 19705 2255 19763 2261
rect 1104 2202 38824 2224
rect 1104 2150 7648 2202
rect 7700 2150 7712 2202
rect 7764 2150 7776 2202
rect 7828 2150 7840 2202
rect 7892 2150 20982 2202
rect 21034 2150 21046 2202
rect 21098 2150 21110 2202
rect 21162 2150 21174 2202
rect 21226 2150 34315 2202
rect 34367 2150 34379 2202
rect 34431 2150 34443 2202
rect 34495 2150 34507 2202
rect 34559 2150 38824 2202
rect 1104 2128 38824 2150
rect 8110 76 8116 128
rect 8168 116 8174 128
rect 12158 116 12164 128
rect 8168 88 12164 116
rect 8168 76 8174 88
rect 12158 76 12164 88
rect 12216 76 12222 128
<< via1 >>
rect 5632 15512 5684 15564
rect 6644 15512 6696 15564
rect 11060 15512 11112 15564
rect 16488 15512 16540 15564
rect 14315 13574 14367 13626
rect 14379 13574 14431 13626
rect 14443 13574 14495 13626
rect 14507 13574 14559 13626
rect 27648 13574 27700 13626
rect 27712 13574 27764 13626
rect 27776 13574 27828 13626
rect 27840 13574 27892 13626
rect 7648 13030 7700 13082
rect 7712 13030 7764 13082
rect 7776 13030 7828 13082
rect 7840 13030 7892 13082
rect 20982 13030 21034 13082
rect 21046 13030 21098 13082
rect 21110 13030 21162 13082
rect 21174 13030 21226 13082
rect 34315 13030 34367 13082
rect 34379 13030 34431 13082
rect 34443 13030 34495 13082
rect 34507 13030 34559 13082
rect 1584 12971 1636 12980
rect 1584 12937 1593 12971
rect 1593 12937 1627 12971
rect 1627 12937 1636 12971
rect 1584 12928 1636 12937
rect 24124 12928 24176 12980
rect 28540 12928 28592 12980
rect 35624 12971 35676 12980
rect 35624 12937 35633 12971
rect 35633 12937 35667 12971
rect 35667 12937 35676 12971
rect 35624 12928 35676 12937
rect 24308 12724 24360 12776
rect 26792 12724 26844 12776
rect 35256 12724 35308 12776
rect 16212 12656 16264 12708
rect 39580 12656 39632 12708
rect 1860 12588 1912 12640
rect 24308 12631 24360 12640
rect 24308 12597 24317 12631
rect 24317 12597 24351 12631
rect 24351 12597 24360 12631
rect 24308 12588 24360 12597
rect 26792 12631 26844 12640
rect 26792 12597 26801 12631
rect 26801 12597 26835 12631
rect 26835 12597 26844 12631
rect 26792 12588 26844 12597
rect 14315 12486 14367 12538
rect 14379 12486 14431 12538
rect 14443 12486 14495 12538
rect 14507 12486 14559 12538
rect 27648 12486 27700 12538
rect 27712 12486 27764 12538
rect 27776 12486 27828 12538
rect 27840 12486 27892 12538
rect 19708 12248 19760 12300
rect 39580 12044 39632 12096
rect 7648 11942 7700 11994
rect 7712 11942 7764 11994
rect 7776 11942 7828 11994
rect 7840 11942 7892 11994
rect 20982 11942 21034 11994
rect 21046 11942 21098 11994
rect 21110 11942 21162 11994
rect 21174 11942 21226 11994
rect 34315 11942 34367 11994
rect 34379 11942 34431 11994
rect 34443 11942 34495 11994
rect 34507 11942 34559 11994
rect 7012 11883 7064 11892
rect 7012 11849 7021 11883
rect 7021 11849 7055 11883
rect 7055 11849 7064 11883
rect 7012 11840 7064 11849
rect 19708 11840 19760 11892
rect 7380 11543 7432 11552
rect 7380 11509 7389 11543
rect 7389 11509 7423 11543
rect 7423 11509 7432 11543
rect 7380 11500 7432 11509
rect 14315 11398 14367 11450
rect 14379 11398 14431 11450
rect 14443 11398 14495 11450
rect 14507 11398 14559 11450
rect 27648 11398 27700 11450
rect 27712 11398 27764 11450
rect 27776 11398 27828 11450
rect 27840 11398 27892 11450
rect 39580 11296 39632 11348
rect 35440 11203 35492 11212
rect 35440 11169 35449 11203
rect 35449 11169 35483 11203
rect 35483 11169 35492 11203
rect 35440 11160 35492 11169
rect 7648 10854 7700 10906
rect 7712 10854 7764 10906
rect 7776 10854 7828 10906
rect 7840 10854 7892 10906
rect 20982 10854 21034 10906
rect 21046 10854 21098 10906
rect 21110 10854 21162 10906
rect 21174 10854 21226 10906
rect 34315 10854 34367 10906
rect 34379 10854 34431 10906
rect 34443 10854 34495 10906
rect 34507 10854 34559 10906
rect 35440 10659 35492 10668
rect 35440 10625 35449 10659
rect 35449 10625 35483 10659
rect 35483 10625 35492 10659
rect 35440 10616 35492 10625
rect 14315 10310 14367 10362
rect 14379 10310 14431 10362
rect 14443 10310 14495 10362
rect 14507 10310 14559 10362
rect 27648 10310 27700 10362
rect 27712 10310 27764 10362
rect 27776 10310 27828 10362
rect 27840 10310 27892 10362
rect 7648 9766 7700 9818
rect 7712 9766 7764 9818
rect 7776 9766 7828 9818
rect 7840 9766 7892 9818
rect 20982 9766 21034 9818
rect 21046 9766 21098 9818
rect 21110 9766 21162 9818
rect 21174 9766 21226 9818
rect 34315 9766 34367 9818
rect 34379 9766 34431 9818
rect 34443 9766 34495 9818
rect 34507 9766 34559 9818
rect 14315 9222 14367 9274
rect 14379 9222 14431 9274
rect 14443 9222 14495 9274
rect 14507 9222 14559 9274
rect 27648 9222 27700 9274
rect 27712 9222 27764 9274
rect 27776 9222 27828 9274
rect 27840 9222 27892 9274
rect 35624 9163 35676 9172
rect 35624 9129 35633 9163
rect 35633 9129 35667 9163
rect 35667 9129 35676 9163
rect 35624 9120 35676 9129
rect 35440 9027 35492 9036
rect 35440 8993 35449 9027
rect 35449 8993 35483 9027
rect 35483 8993 35492 9027
rect 35440 8984 35492 8993
rect 12072 8916 12124 8968
rect 13452 8780 13504 8832
rect 7648 8678 7700 8730
rect 7712 8678 7764 8730
rect 7776 8678 7828 8730
rect 7840 8678 7892 8730
rect 20982 8678 21034 8730
rect 21046 8678 21098 8730
rect 21110 8678 21162 8730
rect 21174 8678 21226 8730
rect 34315 8678 34367 8730
rect 34379 8678 34431 8730
rect 34443 8678 34495 8730
rect 34507 8678 34559 8730
rect 11152 8619 11204 8628
rect 11152 8585 11161 8619
rect 11161 8585 11195 8619
rect 11195 8585 11204 8619
rect 11152 8576 11204 8585
rect 12900 8619 12952 8628
rect 12900 8585 12909 8619
rect 12909 8585 12943 8619
rect 12943 8585 12952 8619
rect 12900 8576 12952 8585
rect 16212 8619 16264 8628
rect 16212 8585 16221 8619
rect 16221 8585 16255 8619
rect 16255 8585 16264 8619
rect 16212 8576 16264 8585
rect 12256 8508 12308 8560
rect 12348 8508 12400 8560
rect 9864 8372 9916 8424
rect 11152 8372 11204 8424
rect 12900 8372 12952 8424
rect 16028 8415 16080 8424
rect 16028 8381 16046 8415
rect 16046 8381 16080 8415
rect 16028 8372 16080 8381
rect 19708 8576 19760 8628
rect 15292 8304 15344 8356
rect 2688 8236 2740 8288
rect 11888 8236 11940 8288
rect 12072 8279 12124 8288
rect 12072 8245 12081 8279
rect 12081 8245 12115 8279
rect 12115 8245 12124 8279
rect 12072 8236 12124 8245
rect 12532 8236 12584 8288
rect 35440 8279 35492 8288
rect 35440 8245 35449 8279
rect 35449 8245 35483 8279
rect 35483 8245 35492 8279
rect 35440 8236 35492 8245
rect 14315 8134 14367 8186
rect 14379 8134 14431 8186
rect 14443 8134 14495 8186
rect 14507 8134 14559 8186
rect 27648 8134 27700 8186
rect 27712 8134 27764 8186
rect 27776 8134 27828 8186
rect 27840 8134 27892 8186
rect 1492 8032 1544 8084
rect 16488 8032 16540 8084
rect 24308 8032 24360 8084
rect 33140 8032 33192 8084
rect 4620 7964 4672 8016
rect 5632 7964 5684 8016
rect 11060 7964 11112 8016
rect 12348 8007 12400 8016
rect 12348 7973 12357 8007
rect 12357 7973 12391 8007
rect 12391 7973 12400 8007
rect 12348 7964 12400 7973
rect 12440 8007 12492 8016
rect 12440 7973 12449 8007
rect 12449 7973 12483 8007
rect 12483 7973 12492 8007
rect 12440 7964 12492 7973
rect 3332 7896 3384 7948
rect 7288 7896 7340 7948
rect 8576 7939 8628 7948
rect 8576 7905 8585 7939
rect 8585 7905 8619 7939
rect 8619 7905 8628 7939
rect 8576 7896 8628 7905
rect 9588 7896 9640 7948
rect 13912 7896 13964 7948
rect 16672 7939 16724 7948
rect 16672 7905 16681 7939
rect 16681 7905 16715 7939
rect 16715 7905 16724 7939
rect 16672 7896 16724 7905
rect 24676 7896 24728 7948
rect 32220 7896 32272 7948
rect 2780 7871 2832 7880
rect 2780 7837 2789 7871
rect 2789 7837 2823 7871
rect 2823 7837 2832 7871
rect 2780 7828 2832 7837
rect 4712 7828 4764 7880
rect 4896 7871 4948 7880
rect 4896 7837 4905 7871
rect 4905 7837 4939 7871
rect 4939 7837 4948 7871
rect 4896 7828 4948 7837
rect 8024 7828 8076 7880
rect 12808 7871 12860 7880
rect 12808 7837 12817 7871
rect 12817 7837 12851 7871
rect 12851 7837 12860 7871
rect 12808 7828 12860 7837
rect 15384 7828 15436 7880
rect 5264 7760 5316 7812
rect 8300 7760 8352 7812
rect 11704 7760 11756 7812
rect 25136 7760 25188 7812
rect 2504 7735 2556 7744
rect 2504 7701 2513 7735
rect 2513 7701 2547 7735
rect 2547 7701 2556 7735
rect 2504 7692 2556 7701
rect 2964 7692 3016 7744
rect 7472 7692 7524 7744
rect 8116 7735 8168 7744
rect 8116 7701 8125 7735
rect 8125 7701 8159 7735
rect 8159 7701 8168 7735
rect 8116 7692 8168 7701
rect 10508 7692 10560 7744
rect 10876 7692 10928 7744
rect 11888 7692 11940 7744
rect 14924 7692 14976 7744
rect 25044 7735 25096 7744
rect 25044 7701 25053 7735
rect 25053 7701 25087 7735
rect 25087 7701 25096 7735
rect 25044 7692 25096 7701
rect 7648 7590 7700 7642
rect 7712 7590 7764 7642
rect 7776 7590 7828 7642
rect 7840 7590 7892 7642
rect 20982 7590 21034 7642
rect 21046 7590 21098 7642
rect 21110 7590 21162 7642
rect 21174 7590 21226 7642
rect 34315 7590 34367 7642
rect 34379 7590 34431 7642
rect 34443 7590 34495 7642
rect 34507 7590 34559 7642
rect 2780 7531 2832 7540
rect 2780 7497 2789 7531
rect 2789 7497 2823 7531
rect 2823 7497 2832 7531
rect 2780 7488 2832 7497
rect 7288 7488 7340 7540
rect 8576 7531 8628 7540
rect 8576 7497 8585 7531
rect 8585 7497 8619 7531
rect 8619 7497 8628 7531
rect 8576 7488 8628 7497
rect 10968 7488 11020 7540
rect 12440 7488 12492 7540
rect 13452 7531 13504 7540
rect 13452 7497 13461 7531
rect 13461 7497 13495 7531
rect 13495 7497 13504 7531
rect 13452 7488 13504 7497
rect 24676 7531 24728 7540
rect 24676 7497 24685 7531
rect 24685 7497 24719 7531
rect 24719 7497 24728 7531
rect 24676 7488 24728 7497
rect 4712 7420 4764 7472
rect 3332 7395 3384 7404
rect 3332 7361 3341 7395
rect 3341 7361 3375 7395
rect 3375 7361 3384 7395
rect 3332 7352 3384 7361
rect 4896 7352 4948 7404
rect 6828 7352 6880 7404
rect 8116 7352 8168 7404
rect 1400 7327 1452 7336
rect 1400 7293 1409 7327
rect 1409 7293 1443 7327
rect 1443 7293 1452 7327
rect 1400 7284 1452 7293
rect 112 7148 164 7200
rect 3148 7259 3200 7268
rect 3148 7225 3157 7259
rect 3157 7225 3191 7259
rect 3191 7225 3200 7259
rect 3148 7216 3200 7225
rect 5264 7259 5316 7268
rect 5264 7225 5273 7259
rect 5273 7225 5307 7259
rect 5307 7225 5316 7259
rect 5264 7216 5316 7225
rect 4620 7191 4672 7200
rect 4620 7157 4629 7191
rect 4629 7157 4663 7191
rect 4663 7157 4672 7191
rect 4620 7148 4672 7157
rect 8024 7216 8076 7268
rect 11060 7420 11112 7472
rect 14004 7420 14056 7472
rect 10876 7395 10928 7404
rect 10876 7361 10885 7395
rect 10885 7361 10919 7395
rect 10919 7361 10928 7395
rect 10876 7352 10928 7361
rect 11888 7352 11940 7404
rect 12808 7395 12860 7404
rect 12808 7361 12817 7395
rect 12817 7361 12851 7395
rect 12851 7361 12860 7395
rect 12808 7352 12860 7361
rect 12992 7352 13044 7404
rect 10600 7284 10652 7336
rect 13912 7327 13964 7336
rect 13912 7293 13921 7327
rect 13921 7293 13955 7327
rect 13955 7293 13964 7327
rect 13912 7284 13964 7293
rect 25136 7352 25188 7404
rect 10968 7259 11020 7268
rect 5540 7148 5592 7200
rect 7288 7191 7340 7200
rect 7288 7157 7297 7191
rect 7297 7157 7331 7191
rect 7331 7157 7340 7191
rect 7288 7148 7340 7157
rect 9588 7191 9640 7200
rect 9588 7157 9597 7191
rect 9597 7157 9631 7191
rect 9631 7157 9640 7191
rect 9588 7148 9640 7157
rect 9680 7148 9732 7200
rect 10968 7225 10977 7259
rect 10977 7225 11011 7259
rect 11011 7225 11020 7259
rect 10968 7216 11020 7225
rect 11612 7216 11664 7268
rect 12624 7259 12676 7268
rect 12624 7225 12633 7259
rect 12633 7225 12667 7259
rect 12667 7225 12676 7259
rect 12624 7216 12676 7225
rect 13912 7148 13964 7200
rect 14740 7148 14792 7200
rect 15568 7148 15620 7200
rect 16672 7191 16724 7200
rect 16672 7157 16681 7191
rect 16681 7157 16715 7191
rect 16715 7157 16724 7191
rect 16672 7148 16724 7157
rect 16764 7148 16816 7200
rect 18236 7284 18288 7336
rect 24308 7284 24360 7336
rect 17592 7216 17644 7268
rect 24400 7216 24452 7268
rect 25044 7216 25096 7268
rect 25780 7216 25832 7268
rect 18328 7148 18380 7200
rect 24492 7148 24544 7200
rect 32220 7191 32272 7200
rect 32220 7157 32229 7191
rect 32229 7157 32263 7191
rect 32263 7157 32272 7191
rect 32220 7148 32272 7157
rect 14315 7046 14367 7098
rect 14379 7046 14431 7098
rect 14443 7046 14495 7098
rect 14507 7046 14559 7098
rect 27648 7046 27700 7098
rect 27712 7046 27764 7098
rect 27776 7046 27828 7098
rect 27840 7046 27892 7098
rect 2504 6944 2556 6996
rect 4988 6987 5040 6996
rect 4988 6953 4997 6987
rect 4997 6953 5031 6987
rect 5031 6953 5040 6987
rect 4988 6944 5040 6953
rect 5540 6987 5592 6996
rect 5540 6953 5549 6987
rect 5549 6953 5583 6987
rect 5583 6953 5592 6987
rect 5540 6944 5592 6953
rect 6828 6987 6880 6996
rect 6828 6953 6837 6987
rect 6837 6953 6871 6987
rect 6871 6953 6880 6987
rect 6828 6944 6880 6953
rect 10876 6987 10928 6996
rect 10876 6953 10885 6987
rect 10885 6953 10919 6987
rect 10919 6953 10928 6987
rect 10876 6944 10928 6953
rect 12440 6944 12492 6996
rect 16764 6944 16816 6996
rect 8024 6876 8076 6928
rect 8300 6919 8352 6928
rect 8300 6885 8309 6919
rect 8309 6885 8343 6919
rect 8343 6885 8352 6919
rect 8300 6876 8352 6885
rect 2044 6808 2096 6860
rect 6460 6851 6512 6860
rect 6460 6817 6469 6851
rect 6469 6817 6503 6851
rect 6503 6817 6512 6851
rect 6460 6808 6512 6817
rect 9772 6851 9824 6860
rect 9772 6817 9781 6851
rect 9781 6817 9815 6851
rect 9815 6817 9824 6851
rect 9772 6808 9824 6817
rect 11336 6876 11388 6928
rect 12624 6876 12676 6928
rect 13176 6919 13228 6928
rect 13176 6885 13185 6919
rect 13185 6885 13219 6919
rect 13219 6885 13228 6919
rect 13176 6876 13228 6885
rect 15384 6919 15436 6928
rect 15384 6885 15393 6919
rect 15393 6885 15427 6919
rect 15427 6885 15436 6919
rect 15384 6876 15436 6885
rect 15476 6919 15528 6928
rect 15476 6885 15485 6919
rect 15485 6885 15519 6919
rect 15519 6885 15528 6919
rect 16028 6919 16080 6928
rect 15476 6876 15528 6885
rect 16028 6885 16037 6919
rect 16037 6885 16071 6919
rect 16071 6885 16080 6919
rect 16028 6876 16080 6885
rect 17592 6919 17644 6928
rect 17592 6885 17601 6919
rect 17601 6885 17635 6919
rect 17635 6885 17644 6919
rect 17592 6876 17644 6885
rect 24492 6876 24544 6928
rect 25044 6919 25096 6928
rect 25044 6885 25053 6919
rect 25053 6885 25087 6919
rect 25087 6885 25096 6919
rect 26700 6919 26752 6928
rect 25044 6876 25096 6885
rect 26700 6885 26709 6919
rect 26709 6885 26743 6919
rect 26743 6885 26752 6919
rect 26700 6876 26752 6885
rect 12808 6808 12860 6860
rect 20168 6808 20220 6860
rect 21364 6851 21416 6860
rect 21364 6817 21373 6851
rect 21373 6817 21407 6851
rect 21407 6817 21416 6851
rect 21364 6808 21416 6817
rect 21916 6851 21968 6860
rect 21916 6817 21925 6851
rect 21925 6817 21959 6851
rect 21959 6817 21968 6851
rect 21916 6808 21968 6817
rect 22100 6851 22152 6860
rect 22100 6817 22109 6851
rect 22109 6817 22143 6851
rect 22143 6817 22152 6851
rect 22100 6808 22152 6817
rect 23296 6808 23348 6860
rect 34612 6851 34664 6860
rect 34612 6817 34621 6851
rect 34621 6817 34655 6851
rect 34655 6817 34664 6851
rect 34612 6808 34664 6817
rect 1584 6783 1636 6792
rect 1584 6749 1593 6783
rect 1593 6749 1627 6783
rect 1627 6749 1636 6783
rect 1584 6740 1636 6749
rect 5540 6740 5592 6792
rect 7472 6740 7524 6792
rect 11520 6740 11572 6792
rect 13452 6740 13504 6792
rect 17868 6740 17920 6792
rect 23572 6740 23624 6792
rect 26056 6740 26108 6792
rect 26608 6783 26660 6792
rect 26608 6749 26617 6783
rect 26617 6749 26651 6783
rect 26651 6749 26660 6783
rect 26608 6740 26660 6749
rect 6644 6672 6696 6724
rect 10048 6672 10100 6724
rect 11612 6672 11664 6724
rect 16672 6672 16724 6724
rect 18512 6672 18564 6724
rect 25780 6672 25832 6724
rect 26424 6672 26476 6724
rect 2320 6647 2372 6656
rect 2320 6613 2329 6647
rect 2329 6613 2363 6647
rect 2363 6613 2372 6647
rect 2320 6604 2372 6613
rect 3056 6647 3108 6656
rect 3056 6613 3065 6647
rect 3065 6613 3099 6647
rect 3099 6613 3108 6647
rect 3056 6604 3108 6613
rect 3516 6647 3568 6656
rect 3516 6613 3525 6647
rect 3525 6613 3559 6647
rect 3559 6613 3568 6647
rect 3516 6604 3568 6613
rect 4344 6647 4396 6656
rect 4344 6613 4353 6647
rect 4353 6613 4387 6647
rect 4387 6613 4396 6647
rect 4344 6604 4396 6613
rect 7196 6604 7248 6656
rect 8944 6604 8996 6656
rect 10140 6604 10192 6656
rect 12624 6604 12676 6656
rect 14372 6647 14424 6656
rect 14372 6613 14381 6647
rect 14381 6613 14415 6647
rect 14415 6613 14424 6647
rect 14372 6604 14424 6613
rect 18420 6647 18472 6656
rect 18420 6613 18429 6647
rect 18429 6613 18463 6647
rect 18463 6613 18472 6647
rect 18420 6604 18472 6613
rect 20168 6647 20220 6656
rect 20168 6613 20177 6647
rect 20177 6613 20211 6647
rect 20211 6613 20220 6647
rect 20168 6604 20220 6613
rect 20628 6647 20680 6656
rect 20628 6613 20637 6647
rect 20637 6613 20671 6647
rect 20671 6613 20680 6647
rect 20628 6604 20680 6613
rect 25136 6604 25188 6656
rect 27988 6604 28040 6656
rect 7648 6502 7700 6554
rect 7712 6502 7764 6554
rect 7776 6502 7828 6554
rect 7840 6502 7892 6554
rect 20982 6502 21034 6554
rect 21046 6502 21098 6554
rect 21110 6502 21162 6554
rect 21174 6502 21226 6554
rect 34315 6502 34367 6554
rect 34379 6502 34431 6554
rect 34443 6502 34495 6554
rect 34507 6502 34559 6554
rect 2044 6443 2096 6452
rect 2044 6409 2053 6443
rect 2053 6409 2087 6443
rect 2087 6409 2096 6443
rect 2044 6400 2096 6409
rect 4620 6400 4672 6452
rect 8024 6400 8076 6452
rect 13176 6400 13228 6452
rect 15384 6443 15436 6452
rect 15384 6409 15393 6443
rect 15393 6409 15427 6443
rect 15427 6409 15436 6443
rect 15384 6400 15436 6409
rect 17592 6400 17644 6452
rect 17868 6443 17920 6452
rect 17868 6409 17877 6443
rect 17877 6409 17911 6443
rect 17911 6409 17920 6443
rect 17868 6400 17920 6409
rect 25044 6400 25096 6452
rect 26700 6400 26752 6452
rect 3516 6332 3568 6384
rect 6460 6332 6512 6384
rect 7380 6332 7432 6384
rect 10600 6332 10652 6384
rect 26056 6332 26108 6384
rect 2320 6264 2372 6316
rect 4252 6264 4304 6316
rect 10048 6264 10100 6316
rect 14372 6307 14424 6316
rect 3056 6239 3108 6248
rect 1676 6128 1728 6180
rect 3056 6205 3065 6239
rect 3065 6205 3099 6239
rect 3099 6205 3108 6239
rect 3056 6196 3108 6205
rect 3424 6239 3476 6248
rect 3424 6205 3433 6239
rect 3433 6205 3467 6239
rect 3467 6205 3476 6239
rect 3424 6196 3476 6205
rect 4068 6196 4120 6248
rect 7196 6239 7248 6248
rect 7196 6205 7205 6239
rect 7205 6205 7239 6239
rect 7239 6205 7248 6239
rect 7196 6196 7248 6205
rect 9956 6196 10008 6248
rect 10232 6196 10284 6248
rect 2780 6060 2832 6112
rect 4988 6128 5040 6180
rect 5540 6060 5592 6112
rect 6736 6060 6788 6112
rect 9772 6128 9824 6180
rect 10324 6128 10376 6180
rect 8944 6060 8996 6112
rect 10232 6060 10284 6112
rect 11060 6196 11112 6248
rect 12624 6196 12676 6248
rect 13084 6128 13136 6180
rect 13176 6128 13228 6180
rect 14372 6273 14381 6307
rect 14381 6273 14415 6307
rect 14415 6273 14424 6307
rect 14372 6264 14424 6273
rect 16028 6264 16080 6316
rect 16764 6264 16816 6316
rect 16856 6307 16908 6316
rect 16856 6273 16865 6307
rect 16865 6273 16899 6307
rect 16899 6273 16908 6307
rect 16856 6264 16908 6273
rect 18420 6264 18472 6316
rect 18512 6307 18564 6316
rect 18512 6273 18521 6307
rect 18521 6273 18555 6307
rect 18555 6273 18564 6307
rect 18512 6264 18564 6273
rect 20720 6264 20772 6316
rect 19432 6196 19484 6248
rect 20168 6239 20220 6248
rect 20168 6205 20177 6239
rect 20177 6205 20211 6239
rect 20211 6205 20220 6239
rect 20168 6196 20220 6205
rect 10968 6103 11020 6112
rect 10968 6069 10977 6103
rect 10977 6069 11011 6103
rect 11011 6069 11020 6103
rect 10968 6060 11020 6069
rect 11336 6103 11388 6112
rect 11336 6069 11345 6103
rect 11345 6069 11379 6103
rect 11379 6069 11388 6103
rect 11336 6060 11388 6069
rect 11520 6060 11572 6112
rect 14188 6103 14240 6112
rect 14188 6069 14197 6103
rect 14197 6069 14231 6103
rect 14231 6069 14240 6103
rect 17224 6128 17276 6180
rect 18236 6171 18288 6180
rect 18236 6137 18245 6171
rect 18245 6137 18279 6171
rect 18279 6137 18288 6171
rect 21272 6196 21324 6248
rect 22100 6264 22152 6316
rect 23572 6264 23624 6316
rect 25136 6264 25188 6316
rect 25780 6307 25832 6316
rect 25780 6273 25789 6307
rect 25789 6273 25823 6307
rect 25823 6273 25832 6307
rect 25780 6264 25832 6273
rect 27988 6264 28040 6316
rect 21916 6196 21968 6248
rect 32220 6400 32272 6452
rect 36084 6443 36136 6452
rect 36084 6409 36093 6443
rect 36093 6409 36127 6443
rect 36127 6409 36136 6443
rect 36084 6400 36136 6409
rect 39580 6332 39632 6384
rect 34612 6196 34664 6248
rect 36084 6196 36136 6248
rect 21640 6171 21692 6180
rect 18236 6128 18288 6137
rect 14188 6060 14240 6069
rect 15200 6060 15252 6112
rect 15476 6060 15528 6112
rect 19708 6103 19760 6112
rect 19708 6069 19717 6103
rect 19717 6069 19751 6103
rect 19751 6069 19760 6103
rect 19708 6060 19760 6069
rect 21640 6137 21649 6171
rect 21649 6137 21683 6171
rect 21683 6137 21692 6171
rect 21640 6128 21692 6137
rect 25596 6171 25648 6180
rect 25596 6137 25605 6171
rect 25605 6137 25639 6171
rect 25639 6137 25648 6171
rect 25596 6128 25648 6137
rect 21364 6060 21416 6112
rect 22192 6060 22244 6112
rect 23020 6103 23072 6112
rect 23020 6069 23029 6103
rect 23029 6069 23063 6103
rect 23063 6069 23072 6103
rect 23020 6060 23072 6069
rect 23296 6060 23348 6112
rect 24032 6103 24084 6112
rect 24032 6069 24041 6103
rect 24041 6069 24075 6103
rect 24075 6069 24084 6103
rect 24032 6060 24084 6069
rect 24400 6060 24452 6112
rect 31392 6060 31444 6112
rect 14315 5958 14367 6010
rect 14379 5958 14431 6010
rect 14443 5958 14495 6010
rect 14507 5958 14559 6010
rect 27648 5958 27700 6010
rect 27712 5958 27764 6010
rect 27776 5958 27828 6010
rect 27840 5958 27892 6010
rect 3148 5899 3200 5908
rect 3148 5865 3157 5899
rect 3157 5865 3191 5899
rect 3191 5865 3200 5899
rect 3148 5856 3200 5865
rect 3332 5856 3384 5908
rect 5080 5856 5132 5908
rect 6644 5856 6696 5908
rect 7196 5899 7248 5908
rect 7196 5865 7205 5899
rect 7205 5865 7239 5899
rect 7239 5865 7248 5899
rect 7196 5856 7248 5865
rect 9128 5899 9180 5908
rect 9128 5865 9137 5899
rect 9137 5865 9171 5899
rect 9171 5865 9180 5899
rect 9128 5856 9180 5865
rect 9680 5856 9732 5908
rect 12716 5856 12768 5908
rect 13912 5856 13964 5908
rect 14188 5856 14240 5908
rect 17592 5899 17644 5908
rect 17592 5865 17601 5899
rect 17601 5865 17635 5899
rect 17635 5865 17644 5899
rect 17592 5856 17644 5865
rect 18236 5856 18288 5908
rect 20628 5899 20680 5908
rect 20628 5865 20637 5899
rect 20637 5865 20671 5899
rect 20671 5865 20680 5899
rect 20628 5856 20680 5865
rect 24400 5856 24452 5908
rect 24492 5856 24544 5908
rect 26608 5856 26660 5908
rect 27988 5856 28040 5908
rect 2780 5788 2832 5840
rect 3424 5788 3476 5840
rect 3792 5788 3844 5840
rect 5540 5831 5592 5840
rect 3516 5720 3568 5772
rect 4252 5763 4304 5772
rect 4252 5729 4261 5763
rect 4261 5729 4295 5763
rect 4295 5729 4304 5763
rect 4252 5720 4304 5729
rect 4528 5763 4580 5772
rect 4528 5729 4537 5763
rect 4537 5729 4571 5763
rect 4571 5729 4580 5763
rect 4528 5720 4580 5729
rect 5540 5797 5549 5831
rect 5549 5797 5583 5831
rect 5583 5797 5592 5831
rect 5540 5788 5592 5797
rect 3424 5652 3476 5704
rect 6184 5720 6236 5772
rect 7196 5763 7248 5772
rect 7196 5729 7205 5763
rect 7205 5729 7239 5763
rect 7239 5729 7248 5763
rect 7196 5720 7248 5729
rect 7380 5763 7432 5772
rect 7380 5729 7389 5763
rect 7389 5729 7423 5763
rect 7423 5729 7432 5763
rect 7380 5720 7432 5729
rect 10324 5763 10376 5772
rect 5356 5652 5408 5704
rect 7104 5652 7156 5704
rect 8760 5652 8812 5704
rect 10324 5729 10333 5763
rect 10333 5729 10367 5763
rect 10367 5729 10376 5763
rect 10324 5720 10376 5729
rect 10784 5788 10836 5840
rect 11520 5831 11572 5840
rect 10692 5720 10744 5772
rect 11520 5797 11529 5831
rect 11529 5797 11563 5831
rect 11563 5797 11572 5831
rect 11520 5788 11572 5797
rect 13084 5788 13136 5840
rect 15568 5788 15620 5840
rect 15844 5831 15896 5840
rect 15844 5797 15853 5831
rect 15853 5797 15887 5831
rect 15887 5797 15896 5831
rect 15844 5788 15896 5797
rect 16856 5788 16908 5840
rect 23020 5788 23072 5840
rect 25596 5788 25648 5840
rect 26976 5788 27028 5840
rect 12256 5720 12308 5772
rect 16764 5763 16816 5772
rect 16764 5729 16773 5763
rect 16773 5729 16807 5763
rect 16807 5729 16816 5763
rect 16764 5720 16816 5729
rect 18144 5720 18196 5772
rect 19800 5763 19852 5772
rect 19800 5729 19809 5763
rect 19809 5729 19843 5763
rect 19843 5729 19852 5763
rect 19800 5720 19852 5729
rect 20444 5720 20496 5772
rect 21916 5763 21968 5772
rect 6644 5584 6696 5636
rect 7380 5584 7432 5636
rect 10784 5584 10836 5636
rect 10968 5652 11020 5704
rect 13268 5652 13320 5704
rect 11796 5584 11848 5636
rect 12992 5584 13044 5636
rect 5540 5516 5592 5568
rect 6460 5559 6512 5568
rect 6460 5525 6469 5559
rect 6469 5525 6503 5559
rect 6503 5525 6512 5559
rect 6460 5516 6512 5525
rect 10232 5516 10284 5568
rect 11888 5559 11940 5568
rect 11888 5525 11897 5559
rect 11897 5525 11931 5559
rect 11931 5525 11940 5559
rect 11888 5516 11940 5525
rect 12808 5559 12860 5568
rect 12808 5525 12817 5559
rect 12817 5525 12851 5559
rect 12851 5525 12860 5559
rect 12808 5516 12860 5525
rect 14648 5559 14700 5568
rect 14648 5525 14657 5559
rect 14657 5525 14691 5559
rect 14691 5525 14700 5559
rect 14648 5516 14700 5525
rect 15384 5516 15436 5568
rect 17132 5559 17184 5568
rect 17132 5525 17141 5559
rect 17141 5525 17175 5559
rect 17175 5525 17184 5559
rect 20628 5652 20680 5704
rect 21916 5729 21925 5763
rect 21925 5729 21959 5763
rect 21959 5729 21968 5763
rect 21916 5720 21968 5729
rect 22100 5763 22152 5772
rect 22100 5729 22109 5763
rect 22109 5729 22143 5763
rect 22143 5729 22152 5763
rect 22100 5720 22152 5729
rect 25504 5720 25556 5772
rect 23204 5695 23256 5704
rect 23204 5661 23213 5695
rect 23213 5661 23247 5695
rect 23247 5661 23256 5695
rect 23204 5652 23256 5661
rect 25136 5652 25188 5704
rect 26608 5695 26660 5704
rect 26608 5661 26617 5695
rect 26617 5661 26651 5695
rect 26651 5661 26660 5695
rect 26608 5652 26660 5661
rect 26056 5584 26108 5636
rect 17132 5516 17184 5525
rect 19524 5516 19576 5568
rect 7648 5414 7700 5466
rect 7712 5414 7764 5466
rect 7776 5414 7828 5466
rect 7840 5414 7892 5466
rect 20982 5414 21034 5466
rect 21046 5414 21098 5466
rect 21110 5414 21162 5466
rect 21174 5414 21226 5466
rect 34315 5414 34367 5466
rect 34379 5414 34431 5466
rect 34443 5414 34495 5466
rect 34507 5414 34559 5466
rect 1032 5312 1084 5364
rect 6184 5355 6236 5364
rect 6184 5321 6193 5355
rect 6193 5321 6227 5355
rect 6227 5321 6236 5355
rect 6184 5312 6236 5321
rect 7104 5355 7156 5364
rect 7104 5321 7113 5355
rect 7113 5321 7147 5355
rect 7147 5321 7156 5355
rect 7104 5312 7156 5321
rect 12256 5355 12308 5364
rect 12256 5321 12265 5355
rect 12265 5321 12299 5355
rect 12299 5321 12308 5355
rect 12256 5312 12308 5321
rect 13084 5312 13136 5364
rect 13820 5312 13872 5364
rect 15200 5355 15252 5364
rect 15200 5321 15209 5355
rect 15209 5321 15243 5355
rect 15243 5321 15252 5355
rect 15200 5312 15252 5321
rect 16304 5312 16356 5364
rect 17592 5312 17644 5364
rect 22192 5355 22244 5364
rect 22192 5321 22201 5355
rect 22201 5321 22235 5355
rect 22235 5321 22244 5355
rect 22192 5312 22244 5321
rect 23020 5312 23072 5364
rect 24032 5355 24084 5364
rect 24032 5321 24041 5355
rect 24041 5321 24075 5355
rect 24075 5321 24084 5355
rect 24032 5312 24084 5321
rect 25596 5312 25648 5364
rect 26608 5312 26660 5364
rect 27436 5312 27488 5364
rect 5080 5244 5132 5296
rect 10048 5244 10100 5296
rect 14096 5244 14148 5296
rect 2044 5108 2096 5160
rect 2872 5151 2924 5160
rect 2872 5117 2881 5151
rect 2881 5117 2915 5151
rect 2915 5117 2924 5151
rect 2872 5108 2924 5117
rect 3332 5176 3384 5228
rect 4068 5219 4120 5228
rect 4068 5185 4077 5219
rect 4077 5185 4111 5219
rect 4111 5185 4120 5219
rect 4068 5176 4120 5185
rect 3148 5108 3200 5160
rect 3792 5151 3844 5160
rect 3792 5117 3801 5151
rect 3801 5117 3835 5151
rect 3835 5117 3844 5151
rect 3792 5108 3844 5117
rect 5632 5151 5684 5160
rect 5632 5117 5641 5151
rect 5641 5117 5675 5151
rect 5675 5117 5684 5151
rect 7472 5151 7524 5160
rect 5632 5108 5684 5117
rect 5908 5083 5960 5092
rect 5908 5049 5917 5083
rect 5917 5049 5951 5083
rect 5951 5049 5960 5083
rect 5908 5040 5960 5049
rect 7472 5117 7481 5151
rect 7481 5117 7515 5151
rect 7515 5117 7524 5151
rect 8944 5176 8996 5228
rect 11060 5219 11112 5228
rect 11060 5185 11069 5219
rect 11069 5185 11103 5219
rect 11103 5185 11112 5219
rect 11060 5176 11112 5185
rect 12716 5219 12768 5228
rect 12716 5185 12725 5219
rect 12725 5185 12759 5219
rect 12759 5185 12768 5219
rect 12716 5176 12768 5185
rect 13176 5219 13228 5228
rect 13176 5185 13185 5219
rect 13185 5185 13219 5219
rect 13219 5185 13228 5219
rect 13176 5176 13228 5185
rect 15844 5176 15896 5228
rect 7472 5108 7524 5117
rect 9864 5151 9916 5160
rect 9864 5117 9873 5151
rect 9873 5117 9907 5151
rect 9907 5117 9916 5151
rect 9864 5108 9916 5117
rect 10048 5151 10100 5160
rect 10048 5117 10057 5151
rect 10057 5117 10091 5151
rect 10091 5117 10100 5151
rect 10048 5108 10100 5117
rect 10140 5108 10192 5160
rect 10784 5151 10836 5160
rect 10784 5117 10793 5151
rect 10793 5117 10827 5151
rect 10827 5117 10836 5151
rect 10784 5108 10836 5117
rect 13728 5108 13780 5160
rect 16764 5108 16816 5160
rect 17224 5176 17276 5228
rect 20444 5244 20496 5296
rect 26976 5287 27028 5296
rect 26976 5253 26985 5287
rect 26985 5253 27019 5287
rect 27019 5253 27028 5287
rect 26976 5244 27028 5253
rect 21640 5176 21692 5228
rect 24216 5219 24268 5228
rect 24216 5185 24225 5219
rect 24225 5185 24259 5219
rect 24259 5185 24268 5219
rect 24216 5176 24268 5185
rect 26056 5219 26108 5228
rect 26056 5185 26065 5219
rect 26065 5185 26099 5219
rect 26099 5185 26108 5219
rect 26056 5176 26108 5185
rect 20444 5108 20496 5160
rect 20628 5151 20680 5160
rect 20628 5117 20637 5151
rect 20637 5117 20671 5151
rect 20671 5117 20680 5151
rect 20628 5108 20680 5117
rect 8116 5040 8168 5092
rect 8300 5083 8352 5092
rect 8300 5049 8309 5083
rect 8309 5049 8343 5083
rect 8343 5049 8352 5083
rect 8300 5040 8352 5049
rect 10692 5040 10744 5092
rect 12808 5083 12860 5092
rect 12808 5049 12817 5083
rect 12817 5049 12851 5083
rect 12851 5049 12860 5083
rect 12808 5040 12860 5049
rect 13820 5040 13872 5092
rect 16304 5040 16356 5092
rect 16856 5040 16908 5092
rect 19800 5040 19852 5092
rect 2044 5015 2096 5024
rect 2044 4981 2053 5015
rect 2053 4981 2087 5015
rect 2087 4981 2096 5015
rect 2044 4972 2096 4981
rect 2780 4972 2832 5024
rect 4252 4972 4304 5024
rect 8760 4972 8812 5024
rect 19524 5015 19576 5024
rect 19524 4981 19533 5015
rect 19533 4981 19567 5015
rect 19567 4981 19576 5015
rect 22100 5108 22152 5160
rect 24032 5108 24084 5160
rect 24400 5040 24452 5092
rect 24768 5040 24820 5092
rect 19524 4972 19576 4981
rect 21272 4972 21324 5024
rect 25504 5015 25556 5024
rect 25504 4981 25513 5015
rect 25513 4981 25547 5015
rect 25547 4981 25556 5015
rect 25504 4972 25556 4981
rect 25780 5015 25832 5024
rect 25780 4981 25789 5015
rect 25789 4981 25823 5015
rect 25823 4981 25832 5015
rect 26884 5040 26936 5092
rect 25780 4972 25832 4981
rect 14315 4870 14367 4922
rect 14379 4870 14431 4922
rect 14443 4870 14495 4922
rect 14507 4870 14559 4922
rect 27648 4870 27700 4922
rect 27712 4870 27764 4922
rect 27776 4870 27828 4922
rect 27840 4870 27892 4922
rect 1676 4811 1728 4820
rect 1676 4777 1685 4811
rect 1685 4777 1719 4811
rect 1719 4777 1728 4811
rect 1676 4768 1728 4777
rect 2872 4768 2924 4820
rect 3516 4768 3568 4820
rect 7196 4811 7248 4820
rect 7196 4777 7205 4811
rect 7205 4777 7239 4811
rect 7239 4777 7248 4811
rect 7196 4768 7248 4777
rect 9588 4768 9640 4820
rect 13268 4811 13320 4820
rect 13268 4777 13277 4811
rect 13277 4777 13311 4811
rect 13311 4777 13320 4811
rect 13268 4768 13320 4777
rect 13820 4811 13872 4820
rect 13820 4777 13829 4811
rect 13829 4777 13863 4811
rect 13863 4777 13872 4811
rect 13820 4768 13872 4777
rect 15016 4768 15068 4820
rect 17040 4811 17092 4820
rect 1952 4675 2004 4684
rect 1952 4641 1961 4675
rect 1961 4641 1995 4675
rect 1995 4641 2004 4675
rect 1952 4632 2004 4641
rect 2504 4632 2556 4684
rect 2872 4632 2924 4684
rect 3700 4632 3752 4684
rect 5080 4675 5132 4684
rect 5080 4641 5089 4675
rect 5089 4641 5123 4675
rect 5123 4641 5132 4675
rect 5080 4632 5132 4641
rect 5356 4632 5408 4684
rect 7104 4700 7156 4752
rect 5724 4632 5776 4684
rect 7012 4632 7064 4684
rect 10232 4700 10284 4752
rect 8024 4632 8076 4684
rect 9956 4675 10008 4684
rect 9956 4641 9965 4675
rect 9965 4641 9999 4675
rect 9999 4641 10008 4675
rect 9956 4632 10008 4641
rect 10048 4632 10100 4684
rect 10692 4675 10744 4684
rect 10692 4641 10701 4675
rect 10701 4641 10735 4675
rect 10735 4641 10744 4675
rect 10692 4632 10744 4641
rect 13728 4700 13780 4752
rect 15384 4743 15436 4752
rect 15384 4709 15393 4743
rect 15393 4709 15427 4743
rect 15427 4709 15436 4743
rect 15384 4700 15436 4709
rect 17040 4777 17049 4811
rect 17049 4777 17083 4811
rect 17083 4777 17092 4811
rect 17040 4768 17092 4777
rect 21916 4768 21968 4820
rect 22560 4768 22612 4820
rect 23204 4811 23256 4820
rect 23204 4777 23213 4811
rect 23213 4777 23247 4811
rect 23247 4777 23256 4811
rect 23204 4768 23256 4777
rect 24216 4811 24268 4820
rect 24216 4777 24225 4811
rect 24225 4777 24259 4811
rect 24259 4777 24268 4811
rect 24216 4768 24268 4777
rect 24768 4811 24820 4820
rect 24768 4777 24777 4811
rect 24777 4777 24811 4811
rect 24811 4777 24820 4811
rect 24768 4768 24820 4777
rect 25780 4768 25832 4820
rect 26056 4811 26108 4820
rect 26056 4777 26065 4811
rect 26065 4777 26099 4811
rect 26099 4777 26108 4811
rect 26056 4768 26108 4777
rect 16028 4743 16080 4752
rect 16028 4709 16037 4743
rect 16037 4709 16071 4743
rect 16071 4709 16080 4743
rect 16028 4700 16080 4709
rect 16580 4700 16632 4752
rect 19708 4700 19760 4752
rect 20628 4700 20680 4752
rect 11980 4675 12032 4684
rect 11980 4641 11989 4675
rect 11989 4641 12023 4675
rect 12023 4641 12032 4675
rect 11980 4632 12032 4641
rect 6368 4607 6420 4616
rect 6368 4573 6377 4607
rect 6377 4573 6411 4607
rect 6411 4573 6420 4607
rect 6368 4564 6420 4573
rect 6644 4564 6696 4616
rect 7288 4564 7340 4616
rect 8300 4564 8352 4616
rect 14924 4632 14976 4684
rect 17224 4675 17276 4684
rect 17224 4641 17233 4675
rect 17233 4641 17267 4675
rect 17267 4641 17276 4675
rect 17224 4632 17276 4641
rect 17316 4632 17368 4684
rect 17776 4675 17828 4684
rect 17776 4641 17785 4675
rect 17785 4641 17819 4675
rect 17819 4641 17828 4675
rect 17776 4632 17828 4641
rect 12624 4564 12676 4616
rect 17500 4564 17552 4616
rect 18328 4632 18380 4684
rect 19892 4632 19944 4684
rect 20720 4632 20772 4684
rect 21364 4675 21416 4684
rect 21364 4641 21373 4675
rect 21373 4641 21407 4675
rect 21407 4641 21416 4675
rect 21364 4632 21416 4641
rect 21732 4632 21784 4684
rect 24400 4700 24452 4752
rect 25412 4700 25464 4752
rect 26700 4743 26752 4752
rect 26700 4709 26709 4743
rect 26709 4709 26743 4743
rect 26743 4709 26752 4743
rect 26700 4700 26752 4709
rect 22100 4675 22152 4684
rect 22100 4641 22109 4675
rect 22109 4641 22143 4675
rect 22143 4641 22152 4675
rect 22100 4632 22152 4641
rect 19524 4564 19576 4616
rect 21640 4564 21692 4616
rect 24676 4564 24728 4616
rect 26424 4564 26476 4616
rect 26884 4607 26936 4616
rect 26884 4573 26893 4607
rect 26893 4573 26927 4607
rect 26927 4573 26936 4607
rect 26884 4564 26936 4573
rect 3056 4496 3108 4548
rect 3332 4496 3384 4548
rect 4252 4539 4304 4548
rect 4252 4505 4261 4539
rect 4261 4505 4295 4539
rect 4295 4505 4304 4539
rect 4252 4496 4304 4505
rect 6920 4496 6972 4548
rect 10324 4496 10376 4548
rect 11520 4539 11572 4548
rect 11520 4505 11529 4539
rect 11529 4505 11563 4539
rect 11563 4505 11572 4539
rect 11520 4496 11572 4505
rect 11796 4539 11848 4548
rect 11796 4505 11805 4539
rect 11805 4505 11839 4539
rect 11839 4505 11848 4539
rect 11796 4496 11848 4505
rect 16488 4496 16540 4548
rect 1676 4428 1728 4480
rect 4528 4428 4580 4480
rect 6736 4428 6788 4480
rect 7472 4428 7524 4480
rect 8116 4428 8168 4480
rect 8760 4471 8812 4480
rect 8760 4437 8769 4471
rect 8769 4437 8803 4471
rect 8803 4437 8812 4471
rect 8760 4428 8812 4437
rect 14188 4428 14240 4480
rect 17776 4428 17828 4480
rect 18420 4428 18472 4480
rect 19156 4471 19208 4480
rect 19156 4437 19165 4471
rect 19165 4437 19199 4471
rect 19199 4437 19208 4471
rect 19156 4428 19208 4437
rect 19248 4428 19300 4480
rect 23664 4471 23716 4480
rect 23664 4437 23673 4471
rect 23673 4437 23707 4471
rect 23707 4437 23716 4471
rect 23664 4428 23716 4437
rect 7648 4326 7700 4378
rect 7712 4326 7764 4378
rect 7776 4326 7828 4378
rect 7840 4326 7892 4378
rect 20982 4326 21034 4378
rect 21046 4326 21098 4378
rect 21110 4326 21162 4378
rect 21174 4326 21226 4378
rect 34315 4326 34367 4378
rect 34379 4326 34431 4378
rect 34443 4326 34495 4378
rect 34507 4326 34559 4378
rect 1860 4267 1912 4276
rect 1860 4233 1869 4267
rect 1869 4233 1903 4267
rect 1903 4233 1912 4267
rect 1860 4224 1912 4233
rect 3332 4224 3384 4276
rect 3700 4267 3752 4276
rect 3700 4233 3709 4267
rect 3709 4233 3743 4267
rect 3743 4233 3752 4267
rect 3700 4224 3752 4233
rect 6644 4267 6696 4276
rect 6644 4233 6653 4267
rect 6653 4233 6687 4267
rect 6687 4233 6696 4267
rect 6644 4224 6696 4233
rect 2688 4156 2740 4208
rect 4252 4156 4304 4208
rect 9036 4224 9088 4276
rect 9956 4224 10008 4276
rect 15568 4224 15620 4276
rect 19432 4224 19484 4276
rect 22560 4267 22612 4276
rect 22560 4233 22569 4267
rect 22569 4233 22603 4267
rect 22603 4233 22612 4267
rect 22560 4224 22612 4233
rect 24032 4224 24084 4276
rect 8760 4156 8812 4208
rect 3148 4088 3200 4140
rect 4252 4063 4304 4072
rect 1400 3884 1452 3936
rect 2872 3995 2924 4004
rect 2872 3961 2881 3995
rect 2881 3961 2915 3995
rect 2915 3961 2924 3995
rect 2872 3952 2924 3961
rect 3056 3952 3108 4004
rect 2964 3884 3016 3936
rect 3700 3884 3752 3936
rect 4252 4029 4261 4063
rect 4261 4029 4295 4063
rect 4295 4029 4304 4063
rect 4252 4020 4304 4029
rect 4804 4063 4856 4072
rect 4804 4029 4813 4063
rect 4813 4029 4847 4063
rect 4847 4029 4856 4063
rect 4804 4020 4856 4029
rect 8944 4088 8996 4140
rect 5632 4063 5684 4072
rect 5632 4029 5641 4063
rect 5641 4029 5675 4063
rect 5675 4029 5684 4063
rect 5632 4020 5684 4029
rect 6460 4020 6512 4072
rect 9036 4063 9088 4072
rect 9036 4029 9045 4063
rect 9045 4029 9079 4063
rect 9079 4029 9088 4063
rect 9956 4088 10008 4140
rect 10324 4156 10376 4208
rect 10600 4156 10652 4208
rect 17500 4156 17552 4208
rect 18880 4156 18932 4208
rect 19892 4199 19944 4208
rect 10140 4088 10192 4140
rect 12624 4088 12676 4140
rect 12900 4088 12952 4140
rect 13176 4131 13228 4140
rect 13176 4097 13185 4131
rect 13185 4097 13219 4131
rect 13219 4097 13228 4131
rect 13176 4088 13228 4097
rect 13820 4131 13872 4140
rect 13820 4097 13829 4131
rect 13829 4097 13863 4131
rect 13863 4097 13872 4131
rect 13820 4088 13872 4097
rect 17132 4131 17184 4140
rect 9036 4020 9088 4029
rect 10232 4063 10284 4072
rect 5264 3952 5316 4004
rect 8024 3952 8076 4004
rect 8484 3995 8536 4004
rect 8484 3961 8493 3995
rect 8493 3961 8527 3995
rect 8527 3961 8536 3995
rect 8484 3952 8536 3961
rect 10232 4029 10241 4063
rect 10241 4029 10275 4063
rect 10275 4029 10284 4063
rect 10232 4020 10284 4029
rect 10416 4020 10468 4072
rect 11980 4020 12032 4072
rect 14004 4020 14056 4072
rect 15936 4063 15988 4072
rect 12900 3995 12952 4004
rect 12900 3961 12909 3995
rect 12909 3961 12943 3995
rect 12943 3961 12952 3995
rect 12900 3952 12952 3961
rect 7196 3927 7248 3936
rect 7196 3893 7205 3927
rect 7205 3893 7239 3927
rect 7239 3893 7248 3927
rect 7196 3884 7248 3893
rect 7748 3927 7800 3936
rect 7748 3893 7757 3927
rect 7757 3893 7791 3927
rect 7791 3893 7800 3927
rect 7748 3884 7800 3893
rect 8208 3884 8260 3936
rect 11244 3927 11296 3936
rect 11244 3893 11253 3927
rect 11253 3893 11287 3927
rect 11287 3893 11296 3927
rect 11244 3884 11296 3893
rect 12348 3884 12400 3936
rect 14832 3884 14884 3936
rect 15936 4029 15945 4063
rect 15945 4029 15979 4063
rect 15979 4029 15988 4063
rect 15936 4020 15988 4029
rect 17132 4097 17141 4131
rect 17141 4097 17175 4131
rect 17175 4097 17184 4131
rect 17132 4088 17184 4097
rect 17224 4088 17276 4140
rect 19156 4088 19208 4140
rect 17408 4063 17460 4072
rect 15844 3952 15896 4004
rect 17408 4029 17417 4063
rect 17417 4029 17451 4063
rect 17451 4029 17460 4063
rect 17408 4020 17460 4029
rect 18236 4063 18288 4072
rect 18236 4029 18245 4063
rect 18245 4029 18279 4063
rect 18279 4029 18288 4063
rect 18236 4020 18288 4029
rect 18420 4020 18472 4072
rect 19064 4020 19116 4072
rect 19892 4165 19901 4199
rect 19901 4165 19935 4199
rect 19935 4165 19944 4199
rect 19892 4156 19944 4165
rect 24768 4156 24820 4208
rect 23664 4131 23716 4140
rect 23664 4097 23673 4131
rect 23673 4097 23707 4131
rect 23707 4097 23716 4131
rect 23664 4088 23716 4097
rect 19432 4020 19484 4072
rect 20720 4063 20772 4072
rect 20720 4029 20729 4063
rect 20729 4029 20763 4063
rect 20763 4029 20772 4063
rect 20720 4020 20772 4029
rect 21272 4020 21324 4072
rect 21640 4063 21692 4072
rect 15200 3884 15252 3936
rect 15660 3884 15712 3936
rect 21364 3952 21416 4004
rect 21640 4029 21649 4063
rect 21649 4029 21683 4063
rect 21683 4029 21692 4063
rect 21640 4020 21692 4029
rect 25412 4131 25464 4140
rect 25412 4097 25421 4131
rect 25421 4097 25455 4131
rect 25455 4097 25464 4131
rect 25412 4088 25464 4097
rect 26700 4267 26752 4276
rect 26700 4233 26709 4267
rect 26709 4233 26743 4267
rect 26743 4233 26752 4267
rect 26700 4224 26752 4233
rect 27436 4267 27488 4276
rect 27436 4233 27445 4267
rect 27445 4233 27479 4267
rect 27479 4233 27488 4267
rect 27436 4224 27488 4233
rect 26424 4156 26476 4208
rect 26792 4088 26844 4140
rect 31392 4131 31444 4140
rect 31392 4097 31401 4131
rect 31401 4097 31435 4131
rect 31435 4097 31444 4131
rect 31392 4088 31444 4097
rect 31668 4131 31720 4140
rect 31668 4097 31677 4131
rect 31677 4097 31711 4131
rect 31711 4097 31720 4131
rect 31668 4088 31720 4097
rect 36084 4156 36136 4208
rect 35532 4131 35584 4140
rect 35532 4097 35541 4131
rect 35541 4097 35575 4131
rect 35575 4097 35584 4131
rect 35532 4088 35584 4097
rect 31484 3995 31536 4004
rect 31484 3961 31493 3995
rect 31493 3961 31527 3995
rect 31527 3961 31536 3995
rect 31484 3952 31536 3961
rect 17132 3884 17184 3936
rect 17316 3884 17368 3936
rect 17684 3884 17736 3936
rect 18144 3927 18196 3936
rect 18144 3893 18153 3927
rect 18153 3893 18187 3927
rect 18187 3893 18196 3927
rect 18144 3884 18196 3893
rect 20444 3884 20496 3936
rect 24032 3927 24084 3936
rect 24032 3893 24041 3927
rect 24041 3893 24075 3927
rect 24075 3893 24084 3927
rect 24032 3884 24084 3893
rect 24584 3927 24636 3936
rect 24584 3893 24593 3927
rect 24593 3893 24627 3927
rect 24627 3893 24636 3927
rect 24584 3884 24636 3893
rect 31300 3884 31352 3936
rect 14315 3782 14367 3834
rect 14379 3782 14431 3834
rect 14443 3782 14495 3834
rect 14507 3782 14559 3834
rect 27648 3782 27700 3834
rect 27712 3782 27764 3834
rect 27776 3782 27828 3834
rect 27840 3782 27892 3834
rect 1952 3723 2004 3732
rect 1952 3689 1961 3723
rect 1961 3689 1995 3723
rect 1995 3689 2004 3723
rect 1952 3680 2004 3689
rect 6736 3723 6788 3732
rect 6736 3689 6745 3723
rect 6745 3689 6779 3723
rect 6779 3689 6788 3723
rect 6736 3680 6788 3689
rect 8116 3680 8168 3732
rect 8944 3680 8996 3732
rect 10508 3680 10560 3732
rect 12072 3680 12124 3732
rect 14188 3680 14240 3732
rect 15016 3723 15068 3732
rect 15016 3689 15025 3723
rect 15025 3689 15059 3723
rect 15059 3689 15068 3723
rect 15016 3680 15068 3689
rect 19984 3680 20036 3732
rect 21640 3680 21692 3732
rect 24676 3723 24728 3732
rect 24676 3689 24685 3723
rect 24685 3689 24719 3723
rect 24719 3689 24728 3723
rect 24676 3680 24728 3689
rect 31392 3723 31444 3732
rect 31392 3689 31401 3723
rect 31401 3689 31435 3723
rect 31435 3689 31444 3723
rect 31392 3680 31444 3689
rect 1584 3612 1636 3664
rect 2504 3612 2556 3664
rect 8024 3655 8076 3664
rect 8024 3621 8033 3655
rect 8033 3621 8067 3655
rect 8067 3621 8076 3655
rect 8024 3612 8076 3621
rect 2688 3408 2740 3460
rect 112 3340 164 3392
rect 2136 3340 2188 3392
rect 3516 3544 3568 3596
rect 4804 3587 4856 3596
rect 4804 3553 4813 3587
rect 4813 3553 4847 3587
rect 4847 3553 4856 3587
rect 4804 3544 4856 3553
rect 5356 3544 5408 3596
rect 5632 3544 5684 3596
rect 6368 3587 6420 3596
rect 6368 3553 6377 3587
rect 6377 3553 6411 3587
rect 6411 3553 6420 3587
rect 6368 3544 6420 3553
rect 12624 3612 12676 3664
rect 8208 3544 8260 3596
rect 9220 3544 9272 3596
rect 9772 3587 9824 3596
rect 9772 3553 9781 3587
rect 9781 3553 9815 3587
rect 9815 3553 9824 3587
rect 9772 3544 9824 3553
rect 10416 3587 10468 3596
rect 10416 3553 10425 3587
rect 10425 3553 10459 3587
rect 10459 3553 10468 3587
rect 10416 3544 10468 3553
rect 11520 3587 11572 3596
rect 11520 3553 11529 3587
rect 11529 3553 11563 3587
rect 11563 3553 11572 3587
rect 11520 3544 11572 3553
rect 11888 3587 11940 3596
rect 11888 3553 11897 3587
rect 11897 3553 11931 3587
rect 11931 3553 11940 3587
rect 11888 3544 11940 3553
rect 12072 3587 12124 3596
rect 12072 3553 12081 3587
rect 12081 3553 12115 3587
rect 12115 3553 12124 3587
rect 12072 3544 12124 3553
rect 12256 3544 12308 3596
rect 4804 3408 4856 3460
rect 5540 3408 5592 3460
rect 12900 3476 12952 3528
rect 13636 3612 13688 3664
rect 14740 3612 14792 3664
rect 15384 3612 15436 3664
rect 15936 3612 15988 3664
rect 17224 3612 17276 3664
rect 17776 3612 17828 3664
rect 15292 3587 15344 3596
rect 15292 3553 15301 3587
rect 15301 3553 15335 3587
rect 15335 3553 15344 3587
rect 15292 3544 15344 3553
rect 15844 3587 15896 3596
rect 15844 3553 15853 3587
rect 15853 3553 15887 3587
rect 15887 3553 15896 3587
rect 15844 3544 15896 3553
rect 17316 3544 17368 3596
rect 17684 3544 17736 3596
rect 18236 3587 18288 3596
rect 18236 3553 18245 3587
rect 18245 3553 18279 3587
rect 18279 3553 18288 3587
rect 18236 3544 18288 3553
rect 18420 3587 18472 3596
rect 18420 3553 18429 3587
rect 18429 3553 18463 3587
rect 18463 3553 18472 3587
rect 18420 3544 18472 3553
rect 19064 3612 19116 3664
rect 20720 3612 20772 3664
rect 24032 3612 24084 3664
rect 32312 3655 32364 3664
rect 32312 3621 32321 3655
rect 32321 3621 32355 3655
rect 32355 3621 32364 3655
rect 32312 3612 32364 3621
rect 18880 3544 18932 3596
rect 18972 3544 19024 3596
rect 19340 3544 19392 3596
rect 19248 3476 19300 3528
rect 20444 3519 20496 3528
rect 20444 3485 20453 3519
rect 20453 3485 20487 3519
rect 20487 3485 20496 3519
rect 20444 3476 20496 3485
rect 21456 3544 21508 3596
rect 23480 3587 23532 3596
rect 23480 3553 23489 3587
rect 23489 3553 23523 3587
rect 23523 3553 23532 3587
rect 23480 3544 23532 3553
rect 25504 3544 25556 3596
rect 25228 3519 25280 3528
rect 25228 3485 25237 3519
rect 25237 3485 25271 3519
rect 25271 3485 25280 3519
rect 25228 3476 25280 3485
rect 32220 3519 32272 3528
rect 32220 3485 32229 3519
rect 32229 3485 32263 3519
rect 32263 3485 32272 3519
rect 32220 3476 32272 3485
rect 11244 3408 11296 3460
rect 3884 3383 3936 3392
rect 3884 3349 3893 3383
rect 3893 3349 3927 3383
rect 3927 3349 3936 3383
rect 3884 3340 3936 3349
rect 6092 3340 6144 3392
rect 9404 3340 9456 3392
rect 11704 3340 11756 3392
rect 12440 3408 12492 3460
rect 12716 3408 12768 3460
rect 14188 3408 14240 3460
rect 14556 3340 14608 3392
rect 14648 3340 14700 3392
rect 15844 3340 15896 3392
rect 17132 3340 17184 3392
rect 18420 3340 18472 3392
rect 20904 3408 20956 3460
rect 31668 3408 31720 3460
rect 30840 3340 30892 3392
rect 7648 3238 7700 3290
rect 7712 3238 7764 3290
rect 7776 3238 7828 3290
rect 7840 3238 7892 3290
rect 20982 3238 21034 3290
rect 21046 3238 21098 3290
rect 21110 3238 21162 3290
rect 21174 3238 21226 3290
rect 34315 3238 34367 3290
rect 34379 3238 34431 3290
rect 34443 3238 34495 3290
rect 34507 3238 34559 3290
rect 3884 3136 3936 3188
rect 5632 3136 5684 3188
rect 6092 3179 6144 3188
rect 6092 3145 6101 3179
rect 6101 3145 6135 3179
rect 6135 3145 6144 3179
rect 6092 3136 6144 3145
rect 6736 3136 6788 3188
rect 2136 3043 2188 3052
rect 2136 3009 2145 3043
rect 2145 3009 2179 3043
rect 2179 3009 2188 3043
rect 2136 3000 2188 3009
rect 4344 3000 4396 3052
rect 4804 3043 4856 3052
rect 4804 3009 4813 3043
rect 4813 3009 4847 3043
rect 4847 3009 4856 3043
rect 4804 3000 4856 3009
rect 1400 2932 1452 2984
rect 2780 2864 2832 2916
rect 3516 2864 3568 2916
rect 5632 3000 5684 3052
rect 9772 3136 9824 3188
rect 12256 3179 12308 3188
rect 12256 3145 12265 3179
rect 12265 3145 12299 3179
rect 12299 3145 12308 3179
rect 12256 3136 12308 3145
rect 13636 3179 13688 3188
rect 7288 3111 7340 3120
rect 7288 3077 7297 3111
rect 7297 3077 7331 3111
rect 7331 3077 7340 3111
rect 7288 3068 7340 3077
rect 7932 3111 7984 3120
rect 7932 3077 7941 3111
rect 7941 3077 7975 3111
rect 7975 3077 7984 3111
rect 7932 3068 7984 3077
rect 7472 3000 7524 3052
rect 8208 3000 8260 3052
rect 12716 3068 12768 3120
rect 13176 3111 13228 3120
rect 13176 3077 13185 3111
rect 13185 3077 13219 3111
rect 13219 3077 13228 3111
rect 13176 3068 13228 3077
rect 13636 3145 13645 3179
rect 13645 3145 13679 3179
rect 13679 3145 13688 3179
rect 13636 3136 13688 3145
rect 15292 3179 15344 3188
rect 14740 3111 14792 3120
rect 14740 3077 14749 3111
rect 14749 3077 14783 3111
rect 14783 3077 14792 3111
rect 14740 3068 14792 3077
rect 15292 3145 15301 3179
rect 15301 3145 15335 3179
rect 15335 3145 15344 3179
rect 15292 3136 15344 3145
rect 15660 3179 15712 3188
rect 15660 3145 15669 3179
rect 15669 3145 15703 3179
rect 15703 3145 15712 3179
rect 15660 3136 15712 3145
rect 17408 3179 17460 3188
rect 17408 3145 17417 3179
rect 17417 3145 17451 3179
rect 17451 3145 17460 3179
rect 17408 3136 17460 3145
rect 18880 3136 18932 3188
rect 23480 3136 23532 3188
rect 26884 3136 26936 3188
rect 30840 3179 30892 3188
rect 30840 3145 30849 3179
rect 30849 3145 30883 3179
rect 30883 3145 30892 3179
rect 30840 3136 30892 3145
rect 31300 3179 31352 3188
rect 31300 3145 31309 3179
rect 31309 3145 31343 3179
rect 31343 3145 31352 3179
rect 31300 3136 31352 3145
rect 32220 3136 32272 3188
rect 17316 3068 17368 3120
rect 19248 3068 19300 3120
rect 24032 3068 24084 3120
rect 9128 3000 9180 3052
rect 16488 3043 16540 3052
rect 16488 3009 16497 3043
rect 16497 3009 16531 3043
rect 16531 3009 16540 3043
rect 16488 3000 16540 3009
rect 11520 2932 11572 2984
rect 17316 2932 17368 2984
rect 18328 2975 18380 2984
rect 18328 2941 18337 2975
rect 18337 2941 18371 2975
rect 18371 2941 18380 2975
rect 18328 2932 18380 2941
rect 18420 2932 18472 2984
rect 18880 2975 18932 2984
rect 18880 2941 18889 2975
rect 18889 2941 18923 2975
rect 18923 2941 18932 2975
rect 18880 2932 18932 2941
rect 19248 2975 19300 2984
rect 19248 2941 19257 2975
rect 19257 2941 19291 2975
rect 19291 2941 19300 2975
rect 19248 2932 19300 2941
rect 19340 2932 19392 2984
rect 25228 3000 25280 3052
rect 5908 2864 5960 2916
rect 8208 2864 8260 2916
rect 8392 2907 8444 2916
rect 8392 2873 8401 2907
rect 8401 2873 8435 2907
rect 8435 2873 8444 2907
rect 8392 2864 8444 2873
rect 9036 2907 9088 2916
rect 9036 2873 9045 2907
rect 9045 2873 9079 2907
rect 9079 2873 9088 2907
rect 9036 2864 9088 2873
rect 9404 2907 9456 2916
rect 9404 2873 9413 2907
rect 9413 2873 9447 2907
rect 9447 2873 9456 2907
rect 9404 2864 9456 2873
rect 10876 2907 10928 2916
rect 10876 2873 10885 2907
rect 10885 2873 10919 2907
rect 10919 2873 10928 2907
rect 10876 2864 10928 2873
rect 10968 2907 11020 2916
rect 10968 2873 10977 2907
rect 10977 2873 11011 2907
rect 11011 2873 11020 2907
rect 10968 2864 11020 2873
rect 2412 2839 2464 2848
rect 2412 2805 2421 2839
rect 2421 2805 2455 2839
rect 2455 2805 2464 2839
rect 2412 2796 2464 2805
rect 3056 2796 3108 2848
rect 7196 2839 7248 2848
rect 7196 2805 7205 2839
rect 7205 2805 7239 2839
rect 7239 2805 7248 2839
rect 7196 2796 7248 2805
rect 7472 2839 7524 2848
rect 7472 2805 7481 2839
rect 7481 2805 7515 2839
rect 7515 2805 7524 2839
rect 7472 2796 7524 2805
rect 12716 2907 12768 2916
rect 12716 2873 12725 2907
rect 12725 2873 12759 2907
rect 12759 2873 12768 2907
rect 14188 2907 14240 2916
rect 12716 2864 12768 2873
rect 12808 2796 12860 2848
rect 14188 2873 14197 2907
rect 14197 2873 14231 2907
rect 14231 2873 14240 2907
rect 14188 2864 14240 2873
rect 16948 2864 17000 2916
rect 19064 2864 19116 2916
rect 20352 2907 20404 2916
rect 20352 2873 20361 2907
rect 20361 2873 20395 2907
rect 20395 2873 20404 2907
rect 20352 2864 20404 2873
rect 26884 2932 26936 2984
rect 30840 2932 30892 2984
rect 32312 2932 32364 2984
rect 33232 3068 33284 3120
rect 34704 3068 34756 3120
rect 24584 2864 24636 2916
rect 25136 2864 25188 2916
rect 17868 2796 17920 2848
rect 18420 2796 18472 2848
rect 21456 2839 21508 2848
rect 21456 2805 21465 2839
rect 21465 2805 21499 2839
rect 21499 2805 21508 2839
rect 21456 2796 21508 2805
rect 22284 2796 22336 2848
rect 29920 2796 29972 2848
rect 14315 2694 14367 2746
rect 14379 2694 14431 2746
rect 14443 2694 14495 2746
rect 14507 2694 14559 2746
rect 27648 2694 27700 2746
rect 27712 2694 27764 2746
rect 27776 2694 27828 2746
rect 27840 2694 27892 2746
rect 3700 2592 3752 2644
rect 3884 2635 3936 2644
rect 3884 2601 3893 2635
rect 3893 2601 3927 2635
rect 3927 2601 3936 2635
rect 3884 2592 3936 2601
rect 5356 2592 5408 2644
rect 7104 2635 7156 2644
rect 7104 2601 7113 2635
rect 7113 2601 7147 2635
rect 7147 2601 7156 2635
rect 7104 2592 7156 2601
rect 10692 2592 10744 2644
rect 2412 2567 2464 2576
rect 2412 2533 2421 2567
rect 2421 2533 2455 2567
rect 2455 2533 2464 2567
rect 2412 2524 2464 2533
rect 1400 2499 1452 2508
rect 1400 2465 1409 2499
rect 1409 2465 1443 2499
rect 1443 2465 1452 2499
rect 1400 2456 1452 2465
rect 3056 2499 3108 2508
rect 3056 2465 3065 2499
rect 3065 2465 3099 2499
rect 3099 2465 3108 2499
rect 3056 2456 3108 2465
rect 6920 2499 6972 2508
rect 1308 2388 1360 2440
rect 6920 2465 6929 2499
rect 6929 2465 6963 2499
rect 6963 2465 6972 2499
rect 6920 2456 6972 2465
rect 7932 2499 7984 2508
rect 7932 2465 7941 2499
rect 7941 2465 7975 2499
rect 7975 2465 7984 2499
rect 7932 2456 7984 2465
rect 8300 2524 8352 2576
rect 10600 2567 10652 2576
rect 10600 2533 10609 2567
rect 10609 2533 10643 2567
rect 10643 2533 10652 2567
rect 10600 2524 10652 2533
rect 8392 2456 8444 2508
rect 11244 2592 11296 2644
rect 12440 2635 12492 2644
rect 12440 2601 12449 2635
rect 12449 2601 12483 2635
rect 12483 2601 12492 2635
rect 12440 2592 12492 2601
rect 12808 2592 12860 2644
rect 16304 2635 16356 2644
rect 16304 2601 16313 2635
rect 16313 2601 16347 2635
rect 16347 2601 16356 2635
rect 16304 2592 16356 2601
rect 11888 2524 11940 2576
rect 12992 2567 13044 2576
rect 12992 2533 13001 2567
rect 13001 2533 13035 2567
rect 13035 2533 13044 2567
rect 12992 2524 13044 2533
rect 14740 2524 14792 2576
rect 16948 2592 17000 2644
rect 19340 2592 19392 2644
rect 25136 2635 25188 2644
rect 11704 2499 11756 2508
rect 11704 2465 11713 2499
rect 11713 2465 11747 2499
rect 11747 2465 11756 2499
rect 11704 2456 11756 2465
rect 15200 2456 15252 2508
rect 17132 2524 17184 2576
rect 20352 2524 20404 2576
rect 25136 2601 25145 2635
rect 25145 2601 25179 2635
rect 25179 2601 25188 2635
rect 25136 2592 25188 2601
rect 32220 2635 32272 2644
rect 32220 2601 32229 2635
rect 32229 2601 32263 2635
rect 32263 2601 32272 2635
rect 32220 2592 32272 2601
rect 33232 2635 33284 2644
rect 33232 2601 33241 2635
rect 33241 2601 33275 2635
rect 33275 2601 33284 2635
rect 33232 2592 33284 2601
rect 21456 2524 21508 2576
rect 17868 2456 17920 2508
rect 19064 2499 19116 2508
rect 19064 2465 19073 2499
rect 19073 2465 19107 2499
rect 19107 2465 19116 2499
rect 19064 2456 19116 2465
rect 20076 2456 20128 2508
rect 21272 2499 21324 2508
rect 21272 2465 21281 2499
rect 21281 2465 21315 2499
rect 21315 2465 21324 2499
rect 21272 2456 21324 2465
rect 25504 2456 25556 2508
rect 5632 2320 5684 2372
rect 7196 2252 7248 2304
rect 8668 2431 8720 2440
rect 8668 2397 8677 2431
rect 8677 2397 8711 2431
rect 8711 2397 8720 2431
rect 8668 2388 8720 2397
rect 11060 2388 11112 2440
rect 14924 2388 14976 2440
rect 16948 2388 17000 2440
rect 8208 2363 8260 2372
rect 8208 2329 8217 2363
rect 8217 2329 8251 2363
rect 8251 2329 8260 2363
rect 8208 2320 8260 2329
rect 10876 2320 10928 2372
rect 11980 2320 12032 2372
rect 18880 2320 18932 2372
rect 22376 2320 22428 2372
rect 31760 2320 31812 2372
rect 34152 2320 34204 2372
rect 11520 2252 11572 2304
rect 18236 2252 18288 2304
rect 7648 2150 7700 2202
rect 7712 2150 7764 2202
rect 7776 2150 7828 2202
rect 7840 2150 7892 2202
rect 20982 2150 21034 2202
rect 21046 2150 21098 2202
rect 21110 2150 21162 2202
rect 21174 2150 21226 2202
rect 34315 2150 34367 2202
rect 34379 2150 34431 2202
rect 34443 2150 34495 2202
rect 34507 2150 34559 2202
rect 8116 76 8168 128
rect 12164 76 12216 128
<< metal2 >>
rect 2226 15586 2282 16000
rect 2056 15558 2282 15586
rect 1490 14784 1546 14793
rect 1490 14719 1546 14728
rect 1398 9344 1454 9353
rect 1398 9279 1454 9288
rect 1412 7342 1440 9279
rect 1504 8090 1532 14719
rect 1582 13696 1638 13705
rect 1582 13631 1638 13640
rect 1596 12986 1624 13631
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 1860 12640 1912 12646
rect 1860 12582 1912 12588
rect 1872 8945 1900 12582
rect 1858 8936 1914 8945
rect 1858 8871 1914 8880
rect 1492 8084 1544 8090
rect 1492 8026 1544 8032
rect 1400 7336 1452 7342
rect 110 7304 166 7313
rect 1400 7278 1452 7284
rect 110 7239 166 7248
rect 124 7206 152 7239
rect 112 7200 164 7206
rect 112 7142 164 7148
rect 1584 6792 1636 6798
rect 1584 6734 1636 6740
rect 1030 5536 1086 5545
rect 1030 5471 1086 5480
rect 1044 5370 1072 5471
rect 1032 5364 1084 5370
rect 1032 5306 1084 5312
rect 1400 3936 1452 3942
rect 1400 3878 1452 3884
rect 112 3392 164 3398
rect 112 3334 164 3340
rect 124 3233 152 3334
rect 110 3224 166 3233
rect 110 3159 166 3168
rect 1412 2990 1440 3878
rect 1596 3670 1624 6734
rect 1676 6180 1728 6186
rect 1676 6122 1728 6128
rect 1688 4826 1716 6122
rect 1872 5137 1900 8871
rect 2056 6866 2084 15558
rect 2226 15520 2282 15558
rect 5632 15564 5684 15570
rect 6642 15564 6698 16000
rect 6642 15520 6644 15564
rect 5632 15506 5684 15512
rect 6696 15520 6698 15564
rect 11058 15564 11114 16000
rect 15566 15586 15622 16000
rect 19982 15586 20038 16000
rect 24398 15586 24454 16000
rect 28906 15586 28962 16000
rect 33322 15586 33378 16000
rect 11058 15520 11060 15564
rect 6644 15506 6696 15512
rect 11112 15520 11114 15564
rect 15488 15558 15622 15586
rect 11060 15506 11112 15512
rect 2688 8288 2740 8294
rect 2688 8230 2740 8236
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 2516 7002 2544 7686
rect 2504 6996 2556 7002
rect 2504 6938 2556 6944
rect 2044 6860 2096 6866
rect 2044 6802 2096 6808
rect 2056 6458 2084 6802
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 2044 6452 2096 6458
rect 1964 6412 2044 6440
rect 1858 5128 1914 5137
rect 1858 5063 1914 5072
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1688 4486 1716 4762
rect 1858 4720 1914 4729
rect 1964 4690 1992 6412
rect 2044 6394 2096 6400
rect 2332 6322 2360 6598
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2044 5160 2096 5166
rect 2042 5128 2044 5137
rect 2096 5128 2098 5137
rect 2042 5063 2098 5072
rect 2056 5030 2084 5063
rect 2044 5024 2096 5030
rect 2044 4966 2096 4972
rect 2516 4690 2544 6938
rect 1858 4655 1914 4664
rect 1952 4684 2004 4690
rect 1676 4480 1728 4486
rect 1676 4422 1728 4428
rect 1872 4282 1900 4655
rect 1952 4626 2004 4632
rect 2504 4684 2556 4690
rect 2504 4626 2556 4632
rect 1860 4276 1912 4282
rect 1860 4218 1912 4224
rect 1964 3738 1992 4626
rect 2700 4214 2728 8230
rect 5644 8022 5672 15506
rect 6656 15475 6684 15506
rect 11072 15475 11100 15506
rect 14289 13628 14585 13648
rect 14345 13626 14369 13628
rect 14425 13626 14449 13628
rect 14505 13626 14529 13628
rect 14367 13574 14369 13626
rect 14431 13574 14443 13626
rect 14505 13574 14507 13626
rect 14345 13572 14369 13574
rect 14425 13572 14449 13574
rect 14505 13572 14529 13574
rect 14289 13552 14585 13572
rect 7622 13084 7918 13104
rect 7678 13082 7702 13084
rect 7758 13082 7782 13084
rect 7838 13082 7862 13084
rect 7700 13030 7702 13082
rect 7764 13030 7776 13082
rect 7838 13030 7840 13082
rect 7678 13028 7702 13030
rect 7758 13028 7782 13030
rect 7838 13028 7862 13030
rect 7622 13008 7918 13028
rect 14289 12540 14585 12560
rect 14345 12538 14369 12540
rect 14425 12538 14449 12540
rect 14505 12538 14529 12540
rect 14367 12486 14369 12538
rect 14431 12486 14443 12538
rect 14505 12486 14507 12538
rect 14345 12484 14369 12486
rect 14425 12484 14449 12486
rect 14505 12484 14529 12486
rect 14289 12464 14585 12484
rect 7010 12064 7066 12073
rect 7010 11999 7066 12008
rect 7024 11898 7052 11999
rect 7622 11996 7918 12016
rect 7678 11994 7702 11996
rect 7758 11994 7782 11996
rect 7838 11994 7862 11996
rect 7700 11942 7702 11994
rect 7764 11942 7776 11994
rect 7838 11942 7840 11994
rect 7678 11940 7702 11942
rect 7758 11940 7782 11942
rect 7838 11940 7862 11942
rect 7622 11920 7918 11940
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 7380 11552 7432 11558
rect 7380 11494 7432 11500
rect 4620 8016 4672 8022
rect 4620 7958 4672 7964
rect 5632 8016 5684 8022
rect 5632 7958 5684 7964
rect 3332 7948 3384 7954
rect 3332 7890 3384 7896
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2792 7546 2820 7822
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 2780 6112 2832 6118
rect 2780 6054 2832 6060
rect 2792 5846 2820 6054
rect 2780 5840 2832 5846
rect 2780 5782 2832 5788
rect 2792 5030 2820 5782
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 2780 5024 2832 5030
rect 2780 4966 2832 4972
rect 2688 4208 2740 4214
rect 2688 4150 2740 4156
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 1584 3664 1636 3670
rect 2504 3664 2556 3670
rect 1584 3606 1636 3612
rect 2424 3624 2504 3652
rect 2136 3392 2188 3398
rect 2136 3334 2188 3340
rect 2148 3058 2176 3334
rect 2136 3052 2188 3058
rect 2136 2994 2188 3000
rect 1400 2984 1452 2990
rect 1400 2926 1452 2932
rect 1412 2514 1440 2926
rect 2424 2854 2452 3624
rect 2504 3606 2556 3612
rect 2700 3466 2728 4150
rect 2688 3460 2740 3466
rect 2688 3402 2740 3408
rect 2792 2922 2820 4966
rect 2884 4826 2912 5102
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2872 4684 2924 4690
rect 2872 4626 2924 4632
rect 2884 4010 2912 4626
rect 2872 4004 2924 4010
rect 2872 3946 2924 3952
rect 2976 3942 3004 7686
rect 3344 7410 3372 7890
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 3148 7268 3200 7274
rect 3148 7210 3200 7216
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 3068 6254 3096 6598
rect 3056 6248 3108 6254
rect 3056 6190 3108 6196
rect 3068 5148 3096 6190
rect 3160 5914 3188 7210
rect 4632 7206 4660 7958
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 4724 7478 4752 7822
rect 4712 7472 4764 7478
rect 4712 7414 4764 7420
rect 4908 7410 4936 7822
rect 5264 7812 5316 7818
rect 5264 7754 5316 7760
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 5276 7274 5304 7754
rect 5264 7268 5316 7274
rect 5264 7210 5316 7216
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 3528 6390 3556 6598
rect 3516 6384 3568 6390
rect 3516 6326 3568 6332
rect 3424 6248 3476 6254
rect 3424 6190 3476 6196
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 3332 5908 3384 5914
rect 3332 5850 3384 5856
rect 3344 5234 3372 5850
rect 3436 5846 3464 6190
rect 3424 5840 3476 5846
rect 3424 5782 3476 5788
rect 3436 5710 3464 5782
rect 3528 5778 3556 6326
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 3792 5840 3844 5846
rect 3792 5782 3844 5788
rect 3516 5772 3568 5778
rect 3516 5714 3568 5720
rect 3424 5704 3476 5710
rect 3424 5646 3476 5652
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 3148 5160 3200 5166
rect 3068 5120 3148 5148
rect 3068 4554 3096 5120
rect 3148 5102 3200 5108
rect 3344 4554 3372 5170
rect 3804 5166 3832 5782
rect 4080 5234 4108 6190
rect 4264 5778 4292 6258
rect 4252 5772 4304 5778
rect 4252 5714 4304 5720
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 4264 5030 4292 5714
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 3056 4548 3108 4554
rect 3332 4548 3384 4554
rect 3108 4508 3188 4536
rect 3056 4490 3108 4496
rect 3160 4146 3188 4508
rect 3332 4490 3384 4496
rect 3344 4282 3372 4490
rect 3332 4276 3384 4282
rect 3332 4218 3384 4224
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 3056 4004 3108 4010
rect 3056 3946 3108 3952
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 2780 2916 2832 2922
rect 2780 2858 2832 2864
rect 2412 2848 2464 2854
rect 2412 2790 2464 2796
rect 2424 2582 2452 2790
rect 2412 2576 2464 2582
rect 2412 2518 2464 2524
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 1308 2440 1360 2446
rect 1308 2382 1360 2388
rect 1122 82 1178 480
rect 1320 82 1348 2382
rect 1412 1193 1440 2450
rect 2976 1737 3004 3878
rect 3068 2854 3096 3946
rect 3528 3602 3556 4762
rect 3700 4684 3752 4690
rect 3700 4626 3752 4632
rect 3712 4282 3740 4626
rect 4264 4554 4292 4966
rect 4356 4593 4384 6598
rect 4632 6458 4660 7142
rect 5552 7002 5580 7142
rect 4988 6996 5040 7002
rect 4988 6938 5040 6944
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 5000 6186 5028 6938
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 4988 6180 5040 6186
rect 4988 6122 5040 6128
rect 5552 6118 5580 6734
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 4342 4584 4398 4593
rect 4252 4548 4304 4554
rect 4342 4519 4398 4528
rect 4252 4490 4304 4496
rect 3700 4276 3752 4282
rect 3700 4218 3752 4224
rect 4264 4214 4292 4490
rect 4252 4208 4304 4214
rect 4252 4150 4304 4156
rect 4264 4078 4292 4150
rect 4252 4072 4304 4078
rect 4252 4014 4304 4020
rect 3700 3936 3752 3942
rect 3700 3878 3752 3884
rect 3516 3596 3568 3602
rect 3516 3538 3568 3544
rect 3516 2916 3568 2922
rect 3516 2858 3568 2864
rect 3056 2848 3108 2854
rect 3056 2790 3108 2796
rect 3068 2514 3096 2790
rect 3056 2508 3108 2514
rect 3056 2450 3108 2456
rect 2962 1728 3018 1737
rect 2962 1663 3018 1672
rect 1398 1184 1454 1193
rect 1398 1119 1454 1128
rect 1122 54 1348 82
rect 3422 82 3478 480
rect 3528 82 3556 2858
rect 3712 2650 3740 3878
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3896 3194 3924 3334
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 3896 2650 3924 3130
rect 4356 3058 4384 4519
rect 4540 4486 4568 5714
rect 5092 5302 5120 5850
rect 5552 5846 5580 6054
rect 5540 5840 5592 5846
rect 5540 5782 5592 5788
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 5080 5296 5132 5302
rect 5080 5238 5132 5244
rect 5092 4690 5120 5238
rect 5368 4690 5396 5646
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5080 4684 5132 4690
rect 5080 4626 5132 4632
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 4528 4480 4580 4486
rect 4528 4422 4580 4428
rect 4540 4185 4568 4422
rect 4526 4176 4582 4185
rect 5092 4154 5120 4626
rect 5092 4126 5304 4154
rect 4526 4111 4582 4120
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 4816 3602 4844 4014
rect 5276 4010 5304 4126
rect 5264 4004 5316 4010
rect 5264 3946 5316 3952
rect 5368 3602 5396 4626
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 4804 3460 4856 3466
rect 4804 3402 4856 3408
rect 4816 3058 4844 3402
rect 4344 3052 4396 3058
rect 4344 2994 4396 3000
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 5368 2650 5396 3538
rect 5552 3466 5580 5510
rect 5644 5166 5672 7958
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7300 7546 7328 7890
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 6840 7002 6868 7346
rect 7300 7206 7328 7482
rect 7288 7200 7340 7206
rect 7288 7142 7340 7148
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6460 6860 6512 6866
rect 6460 6802 6512 6808
rect 6472 6390 6500 6802
rect 6644 6724 6696 6730
rect 6644 6666 6696 6672
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 6656 5914 6684 6666
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7208 6254 7236 6598
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 6184 5772 6236 5778
rect 6184 5714 6236 5720
rect 6196 5370 6224 5714
rect 6656 5642 6684 5850
rect 6644 5636 6696 5642
rect 6644 5578 6696 5584
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 6184 5364 6236 5370
rect 6184 5306 6236 5312
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 5908 5092 5960 5098
rect 5908 5034 5960 5040
rect 5724 4684 5776 4690
rect 5644 4644 5724 4672
rect 5644 4078 5672 4644
rect 5724 4626 5776 4632
rect 5632 4072 5684 4078
rect 5632 4014 5684 4020
rect 5644 3602 5672 4014
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 5540 3460 5592 3466
rect 5540 3402 5592 3408
rect 5644 3194 5672 3538
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 3700 2644 3752 2650
rect 3700 2586 3752 2592
rect 3884 2644 3936 2650
rect 3884 2586 3936 2592
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 5644 2378 5672 2994
rect 5920 2922 5948 5034
rect 6368 4616 6420 4622
rect 6368 4558 6420 4564
rect 6380 3602 6408 4558
rect 6472 4078 6500 5510
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6656 4282 6684 4558
rect 6748 4486 6776 6054
rect 7208 5914 7236 6190
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7300 5817 7328 7142
rect 7392 6390 7420 11494
rect 14289 11452 14585 11472
rect 14345 11450 14369 11452
rect 14425 11450 14449 11452
rect 14505 11450 14529 11452
rect 14367 11398 14369 11450
rect 14431 11398 14443 11450
rect 14505 11398 14507 11450
rect 14345 11396 14369 11398
rect 14425 11396 14449 11398
rect 14505 11396 14529 11398
rect 14289 11376 14585 11396
rect 11150 11112 11206 11121
rect 11150 11047 11206 11056
rect 7622 10908 7918 10928
rect 7678 10906 7702 10908
rect 7758 10906 7782 10908
rect 7838 10906 7862 10908
rect 7700 10854 7702 10906
rect 7764 10854 7776 10906
rect 7838 10854 7840 10906
rect 7678 10852 7702 10854
rect 7758 10852 7782 10854
rect 7838 10852 7862 10854
rect 7622 10832 7918 10852
rect 7622 9820 7918 9840
rect 7678 9818 7702 9820
rect 7758 9818 7782 9820
rect 7838 9818 7862 9820
rect 7700 9766 7702 9818
rect 7764 9766 7776 9818
rect 7838 9766 7840 9818
rect 7678 9764 7702 9766
rect 7758 9764 7782 9766
rect 7838 9764 7862 9766
rect 7622 9744 7918 9764
rect 7622 8732 7918 8752
rect 7678 8730 7702 8732
rect 7758 8730 7782 8732
rect 7838 8730 7862 8732
rect 7700 8678 7702 8730
rect 7764 8678 7776 8730
rect 7838 8678 7840 8730
rect 7678 8676 7702 8678
rect 7758 8676 7782 8678
rect 7838 8676 7862 8678
rect 7622 8656 7918 8676
rect 11164 8634 11192 11047
rect 15488 10713 15516 15558
rect 15566 15520 15622 15558
rect 16488 15564 16540 15570
rect 16488 15506 16540 15512
rect 19720 15558 20038 15586
rect 16212 12708 16264 12714
rect 16212 12650 16264 12656
rect 15474 10704 15530 10713
rect 15474 10639 15530 10648
rect 14289 10364 14585 10384
rect 14345 10362 14369 10364
rect 14425 10362 14449 10364
rect 14505 10362 14529 10364
rect 14367 10310 14369 10362
rect 14431 10310 14443 10362
rect 14505 10310 14507 10362
rect 14345 10308 14369 10310
rect 14425 10308 14449 10310
rect 14505 10308 14529 10310
rect 14289 10288 14585 10308
rect 14289 9276 14585 9296
rect 14345 9274 14369 9276
rect 14425 9274 14449 9276
rect 14505 9274 14529 9276
rect 14367 9222 14369 9274
rect 14431 9222 14443 9274
rect 14505 9222 14507 9274
rect 14345 9220 14369 9222
rect 14425 9220 14449 9222
rect 14505 9220 14529 9222
rect 14289 9200 14585 9220
rect 12072 8968 12124 8974
rect 12072 8910 12124 8916
rect 12898 8936 12954 8945
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11164 8430 11192 8570
rect 9864 8424 9916 8430
rect 11152 8424 11204 8430
rect 9864 8366 9916 8372
rect 11058 8392 11114 8401
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 9588 7948 9640 7954
rect 9588 7890 9640 7896
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7484 6798 7512 7686
rect 7622 7644 7918 7664
rect 7678 7642 7702 7644
rect 7758 7642 7782 7644
rect 7838 7642 7862 7644
rect 7700 7590 7702 7642
rect 7764 7590 7776 7642
rect 7838 7590 7840 7642
rect 7678 7588 7702 7590
rect 7758 7588 7782 7590
rect 7838 7588 7862 7590
rect 7622 7568 7918 7588
rect 8036 7274 8064 7822
rect 8300 7812 8352 7818
rect 8300 7754 8352 7760
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 8128 7410 8156 7686
rect 8116 7404 8168 7410
rect 8116 7346 8168 7352
rect 8024 7268 8076 7274
rect 8024 7210 8076 7216
rect 8036 6934 8064 7210
rect 8312 6934 8340 7754
rect 8588 7546 8616 7890
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 9600 7206 9628 7890
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 8024 6928 8076 6934
rect 8024 6870 8076 6876
rect 8300 6928 8352 6934
rect 8300 6870 8352 6876
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7622 6556 7918 6576
rect 7678 6554 7702 6556
rect 7758 6554 7782 6556
rect 7838 6554 7862 6556
rect 7700 6502 7702 6554
rect 7764 6502 7776 6554
rect 7838 6502 7840 6554
rect 7678 6500 7702 6502
rect 7758 6500 7782 6502
rect 7838 6500 7862 6502
rect 7622 6480 7918 6500
rect 8036 6458 8064 6870
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 7380 6384 7432 6390
rect 7380 6326 7432 6332
rect 8956 6118 8984 6598
rect 8944 6112 8996 6118
rect 8944 6054 8996 6060
rect 7286 5808 7342 5817
rect 7196 5772 7248 5778
rect 7286 5743 7342 5752
rect 7380 5772 7432 5778
rect 7196 5714 7248 5720
rect 7380 5714 7432 5720
rect 7104 5704 7156 5710
rect 7104 5646 7156 5652
rect 7116 5370 7144 5646
rect 7104 5364 7156 5370
rect 7104 5306 7156 5312
rect 7116 4758 7144 5306
rect 7208 4826 7236 5714
rect 7392 5642 7420 5714
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 7380 5636 7432 5642
rect 7380 5578 7432 5584
rect 7622 5468 7918 5488
rect 7678 5466 7702 5468
rect 7758 5466 7782 5468
rect 7838 5466 7862 5468
rect 7700 5414 7702 5466
rect 7764 5414 7776 5466
rect 7838 5414 7840 5466
rect 7678 5412 7702 5414
rect 7758 5412 7782 5414
rect 7838 5412 7862 5414
rect 7622 5392 7918 5412
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 7104 4752 7156 4758
rect 7208 4729 7236 4762
rect 7104 4694 7156 4700
rect 7194 4720 7250 4729
rect 7012 4684 7064 4690
rect 7194 4655 7250 4664
rect 7012 4626 7064 4632
rect 6920 4548 6972 4554
rect 6920 4490 6972 4496
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 6644 4276 6696 4282
rect 6644 4218 6696 4224
rect 6460 4072 6512 4078
rect 6460 4014 6512 4020
rect 6748 3777 6776 4422
rect 6734 3768 6790 3777
rect 6734 3703 6736 3712
rect 6788 3703 6790 3712
rect 6736 3674 6788 3680
rect 6368 3596 6420 3602
rect 6368 3538 6420 3544
rect 6092 3392 6144 3398
rect 6092 3334 6144 3340
rect 6104 3194 6132 3334
rect 6748 3194 6776 3674
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 5908 2916 5960 2922
rect 5908 2858 5960 2864
rect 6932 2514 6960 4490
rect 7024 4154 7052 4626
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 7024 4126 7144 4154
rect 7116 2650 7144 4126
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 7208 3777 7236 3878
rect 7194 3768 7250 3777
rect 7194 3703 7250 3712
rect 7300 3126 7328 4558
rect 7484 4486 7512 5102
rect 8116 5092 8168 5098
rect 8116 5034 8168 5040
rect 8300 5092 8352 5098
rect 8300 5034 8352 5040
rect 8024 4684 8076 4690
rect 8024 4626 8076 4632
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 7288 3120 7340 3126
rect 7288 3062 7340 3068
rect 7484 3058 7512 4422
rect 7622 4380 7918 4400
rect 7678 4378 7702 4380
rect 7758 4378 7782 4380
rect 7838 4378 7862 4380
rect 7700 4326 7702 4378
rect 7764 4326 7776 4378
rect 7838 4326 7840 4378
rect 7678 4324 7702 4326
rect 7758 4324 7782 4326
rect 7838 4324 7862 4326
rect 7622 4304 7918 4324
rect 7746 4040 7802 4049
rect 8036 4010 8064 4626
rect 8128 4486 8156 5034
rect 8312 4622 8340 5034
rect 8772 5030 8800 5646
rect 8956 5234 8984 6054
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8116 4480 8168 4486
rect 8116 4422 8168 4428
rect 7746 3975 7802 3984
rect 8024 4004 8076 4010
rect 7760 3942 7788 3975
rect 8024 3946 8076 3952
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 8036 3670 8064 3946
rect 8128 3738 8156 4422
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 8116 3732 8168 3738
rect 8116 3674 8168 3680
rect 8024 3664 8076 3670
rect 8024 3606 8076 3612
rect 7622 3292 7918 3312
rect 7678 3290 7702 3292
rect 7758 3290 7782 3292
rect 7838 3290 7862 3292
rect 7700 3238 7702 3290
rect 7764 3238 7776 3290
rect 7838 3238 7840 3290
rect 7678 3236 7702 3238
rect 7758 3236 7782 3238
rect 7838 3236 7862 3238
rect 7622 3216 7918 3236
rect 7932 3120 7984 3126
rect 8036 3108 8064 3606
rect 8220 3602 8248 3878
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 7984 3080 8064 3108
rect 7932 3062 7984 3068
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 7484 2854 7512 2994
rect 7196 2848 7248 2854
rect 7196 2790 7248 2796
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 5632 2372 5684 2378
rect 5632 2314 5684 2320
rect 3422 54 3556 82
rect 5644 82 5672 2314
rect 7208 2310 7236 2790
rect 7484 2417 7512 2790
rect 7944 2514 7972 3062
rect 8220 3058 8248 3538
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 8208 2916 8260 2922
rect 8208 2858 8260 2864
rect 7932 2508 7984 2514
rect 7932 2450 7984 2456
rect 7470 2408 7526 2417
rect 8220 2378 8248 2858
rect 8312 2582 8340 4558
rect 8772 4486 8800 4966
rect 8760 4480 8812 4486
rect 8760 4422 8812 4428
rect 8772 4214 8800 4422
rect 8760 4208 8812 4214
rect 8760 4150 8812 4156
rect 8956 4146 8984 5170
rect 9036 4276 9088 4282
rect 9036 4218 9088 4224
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 8484 4004 8536 4010
rect 8484 3946 8536 3952
rect 8496 3913 8524 3946
rect 8482 3904 8538 3913
rect 8482 3839 8538 3848
rect 8956 3738 8984 4082
rect 9048 4078 9076 4218
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 9034 3904 9090 3913
rect 9034 3839 9090 3848
rect 8944 3732 8996 3738
rect 8944 3674 8996 3680
rect 9048 2922 9076 3839
rect 9140 3058 9168 5850
rect 9600 4826 9628 7142
rect 9692 5914 9720 7142
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9784 6186 9812 6802
rect 9772 6180 9824 6186
rect 9772 6122 9824 6128
rect 9876 6066 9904 8366
rect 11152 8366 11204 8372
rect 11058 8327 11114 8336
rect 11072 8022 11100 8327
rect 12084 8294 12112 8910
rect 12898 8871 12954 8880
rect 12912 8634 12940 8871
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 12900 8628 12952 8634
rect 12952 8588 13032 8616
rect 12900 8570 12952 8576
rect 12256 8560 12308 8566
rect 12256 8502 12308 8508
rect 12348 8560 12400 8566
rect 12348 8502 12400 8508
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 12072 8288 12124 8294
rect 12072 8230 12124 8236
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 10508 7744 10560 7750
rect 10508 7686 10560 7692
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10048 6724 10100 6730
rect 10048 6666 10100 6672
rect 10060 6322 10088 6666
rect 10140 6656 10192 6662
rect 10192 6616 10272 6644
rect 10140 6598 10192 6604
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 9784 6038 9904 6066
rect 9680 5908 9732 5914
rect 9680 5850 9732 5856
rect 9588 4820 9640 4826
rect 9588 4762 9640 4768
rect 9218 4176 9274 4185
rect 9218 4111 9274 4120
rect 9232 3602 9260 4111
rect 9784 3602 9812 6038
rect 9864 5160 9916 5166
rect 9968 5148 9996 6190
rect 10060 5302 10088 6258
rect 10244 6254 10272 6616
rect 10232 6248 10284 6254
rect 10232 6190 10284 6196
rect 10324 6180 10376 6186
rect 10376 6140 10456 6168
rect 10324 6122 10376 6128
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10244 5574 10272 6054
rect 10324 5772 10376 5778
rect 10324 5714 10376 5720
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10048 5296 10100 5302
rect 10048 5238 10100 5244
rect 10060 5166 10088 5238
rect 9916 5120 9996 5148
rect 10048 5160 10100 5166
rect 9864 5102 9916 5108
rect 10048 5102 10100 5108
rect 10140 5160 10192 5166
rect 10140 5102 10192 5108
rect 9876 5001 9904 5102
rect 9862 4992 9918 5001
rect 9862 4927 9918 4936
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 9968 4282 9996 4626
rect 9956 4276 10008 4282
rect 9956 4218 10008 4224
rect 9968 4146 9996 4218
rect 10060 4185 10088 4626
rect 10046 4176 10102 4185
rect 9956 4140 10008 4146
rect 10152 4146 10180 5102
rect 10244 4758 10272 5510
rect 10232 4752 10284 4758
rect 10232 4694 10284 4700
rect 10046 4111 10102 4120
rect 10140 4140 10192 4146
rect 9956 4082 10008 4088
rect 10140 4082 10192 4088
rect 10244 4078 10272 4694
rect 10336 4554 10364 5714
rect 10324 4548 10376 4554
rect 10324 4490 10376 4496
rect 10324 4208 10376 4214
rect 10324 4150 10376 4156
rect 10232 4072 10284 4078
rect 10232 4014 10284 4020
rect 9220 3596 9272 3602
rect 9220 3538 9272 3544
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 9128 3052 9180 3058
rect 9128 2994 9180 3000
rect 9416 2922 9444 3334
rect 9784 3194 9812 3538
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 8392 2916 8444 2922
rect 8392 2858 8444 2864
rect 9036 2916 9088 2922
rect 9036 2858 9088 2864
rect 9404 2916 9456 2922
rect 9404 2858 9456 2864
rect 8300 2576 8352 2582
rect 8300 2518 8352 2524
rect 8404 2514 8432 2858
rect 8666 2544 8722 2553
rect 8392 2508 8444 2514
rect 8666 2479 8722 2488
rect 8392 2450 8444 2456
rect 8680 2446 8708 2479
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 7470 2343 7526 2352
rect 8208 2372 8260 2378
rect 8208 2314 8260 2320
rect 7196 2304 7248 2310
rect 7196 2246 7248 2252
rect 7622 2204 7918 2224
rect 7678 2202 7702 2204
rect 7758 2202 7782 2204
rect 7838 2202 7862 2204
rect 7700 2150 7702 2202
rect 7764 2150 7776 2202
rect 7838 2150 7840 2202
rect 7678 2148 7702 2150
rect 7758 2148 7782 2150
rect 7838 2148 7862 2150
rect 7622 2128 7918 2148
rect 5814 82 5870 480
rect 5644 54 5870 82
rect 1122 0 1178 54
rect 3422 0 3478 54
rect 5814 0 5870 54
rect 8114 128 8170 480
rect 8114 76 8116 128
rect 8168 76 8170 128
rect 8114 0 8170 76
rect 10336 82 10364 4150
rect 10428 4078 10456 6140
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 10428 3602 10456 4014
rect 10520 3738 10548 7686
rect 10888 7410 10916 7686
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 10600 7336 10652 7342
rect 10600 7278 10652 7284
rect 10612 6390 10640 7278
rect 10888 7002 10916 7346
rect 10980 7274 11008 7482
rect 11072 7478 11100 7958
rect 11704 7812 11756 7818
rect 11704 7754 11756 7760
rect 11060 7472 11112 7478
rect 11060 7414 11112 7420
rect 10968 7268 11020 7274
rect 10968 7210 11020 7216
rect 11612 7268 11664 7274
rect 11612 7210 11664 7216
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 11336 6928 11388 6934
rect 11336 6870 11388 6876
rect 10600 6384 10652 6390
rect 10600 6326 10652 6332
rect 10612 4214 10640 6326
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 10968 6112 11020 6118
rect 10968 6054 11020 6060
rect 10784 5840 10836 5846
rect 10784 5782 10836 5788
rect 10692 5772 10744 5778
rect 10692 5714 10744 5720
rect 10704 5098 10732 5714
rect 10796 5642 10824 5782
rect 10980 5710 11008 6054
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 10784 5636 10836 5642
rect 10784 5578 10836 5584
rect 10796 5166 10824 5578
rect 11072 5234 11100 6190
rect 11348 6118 11376 6870
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11532 6118 11560 6734
rect 11624 6730 11652 7210
rect 11612 6724 11664 6730
rect 11612 6666 11664 6672
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10692 5092 10744 5098
rect 10692 5034 10744 5040
rect 10704 4690 10732 5034
rect 10692 4684 10744 4690
rect 10692 4626 10744 4632
rect 10600 4208 10652 4214
rect 10600 4150 10652 4156
rect 10598 3768 10654 3777
rect 10508 3732 10560 3738
rect 10598 3703 10654 3712
rect 10508 3674 10560 3680
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 10612 2582 10640 3703
rect 10692 2644 10744 2650
rect 10796 2632 10824 5102
rect 11242 4176 11298 4185
rect 11242 4111 11298 4120
rect 11256 3942 11284 4111
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 11256 3466 11284 3878
rect 11348 3777 11376 6054
rect 11532 5846 11560 6054
rect 11520 5840 11572 5846
rect 11520 5782 11572 5788
rect 11520 4548 11572 4554
rect 11520 4490 11572 4496
rect 11532 4457 11560 4490
rect 11518 4448 11574 4457
rect 11518 4383 11574 4392
rect 11334 3768 11390 3777
rect 11334 3703 11390 3712
rect 11520 3596 11572 3602
rect 11716 3584 11744 7754
rect 11900 7750 11928 8230
rect 11888 7744 11940 7750
rect 11888 7686 11940 7692
rect 11900 7410 11928 7686
rect 11888 7404 11940 7410
rect 11888 7346 11940 7352
rect 12268 6304 12296 8502
rect 12360 8022 12388 8502
rect 12900 8424 12952 8430
rect 12900 8366 12952 8372
rect 12532 8288 12584 8294
rect 12532 8230 12584 8236
rect 12348 8016 12400 8022
rect 12348 7958 12400 7964
rect 12440 8016 12492 8022
rect 12440 7958 12492 7964
rect 12452 7546 12480 7958
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12452 7002 12480 7482
rect 12440 6996 12492 7002
rect 12440 6938 12492 6944
rect 12268 6276 12388 6304
rect 12254 6216 12310 6225
rect 12254 6151 12310 6160
rect 12268 5778 12296 6151
rect 12256 5772 12308 5778
rect 12256 5714 12308 5720
rect 11796 5636 11848 5642
rect 11796 5578 11848 5584
rect 11808 4729 11836 5578
rect 11888 5568 11940 5574
rect 11888 5510 11940 5516
rect 11794 4720 11850 4729
rect 11794 4655 11850 4664
rect 11808 4554 11836 4655
rect 11796 4548 11848 4554
rect 11796 4490 11848 4496
rect 11900 3720 11928 5510
rect 12268 5370 12296 5714
rect 12256 5364 12308 5370
rect 12256 5306 12308 5312
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 11992 4078 12020 4626
rect 12268 4154 12296 5306
rect 12176 4126 12296 4154
rect 11980 4072 12032 4078
rect 11980 4014 12032 4020
rect 11992 3913 12020 4014
rect 11978 3904 12034 3913
rect 11978 3839 12034 3848
rect 12072 3732 12124 3738
rect 11900 3692 12020 3720
rect 11888 3596 11940 3602
rect 11716 3556 11888 3584
rect 11520 3538 11572 3544
rect 11888 3538 11940 3544
rect 11244 3460 11296 3466
rect 11244 3402 11296 3408
rect 11532 2990 11560 3538
rect 11704 3392 11756 3398
rect 11900 3369 11928 3538
rect 11704 3334 11756 3340
rect 11886 3360 11942 3369
rect 11520 2984 11572 2990
rect 11520 2926 11572 2932
rect 10876 2916 10928 2922
rect 10876 2858 10928 2864
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 10744 2604 10824 2632
rect 10692 2586 10744 2592
rect 10600 2576 10652 2582
rect 10600 2518 10652 2524
rect 10888 2378 10916 2858
rect 10876 2372 10928 2378
rect 10876 2314 10928 2320
rect 10980 2145 11008 2858
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 11060 2440 11112 2446
rect 11256 2428 11284 2586
rect 11112 2400 11284 2428
rect 11060 2382 11112 2388
rect 11532 2310 11560 2926
rect 11716 2514 11744 3334
rect 11886 3295 11942 3304
rect 11900 2582 11928 3295
rect 11888 2576 11940 2582
rect 11888 2518 11940 2524
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 11716 2417 11744 2450
rect 11702 2408 11758 2417
rect 11992 2378 12020 3692
rect 12072 3674 12124 3680
rect 12084 3602 12112 3674
rect 12072 3596 12124 3602
rect 12072 3538 12124 3544
rect 11702 2343 11758 2352
rect 11980 2372 12032 2378
rect 11980 2314 12032 2320
rect 11520 2304 11572 2310
rect 11520 2246 11572 2252
rect 10966 2136 11022 2145
rect 10966 2071 11022 2080
rect 10506 82 10562 480
rect 12176 134 12204 4126
rect 12360 3942 12388 6276
rect 12348 3936 12400 3942
rect 12348 3878 12400 3884
rect 12256 3596 12308 3602
rect 12360 3584 12388 3878
rect 12308 3556 12388 3584
rect 12256 3538 12308 3544
rect 12268 3194 12296 3538
rect 12440 3460 12492 3466
rect 12440 3402 12492 3408
rect 12256 3188 12308 3194
rect 12256 3130 12308 3136
rect 12452 2650 12480 3402
rect 12544 3233 12572 8230
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12820 7410 12848 7822
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 12624 7268 12676 7274
rect 12624 7210 12676 7216
rect 12636 6934 12664 7210
rect 12624 6928 12676 6934
rect 12624 6870 12676 6876
rect 12820 6866 12848 7346
rect 12808 6860 12860 6866
rect 12808 6802 12860 6808
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 12636 6254 12664 6598
rect 12624 6248 12676 6254
rect 12624 6190 12676 6196
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 12728 5234 12756 5850
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 12820 5098 12848 5510
rect 12808 5092 12860 5098
rect 12728 5052 12808 5080
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 12636 4146 12664 4558
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12728 4049 12756 5052
rect 12808 5034 12860 5040
rect 12912 4978 12940 8366
rect 13004 7410 13032 8588
rect 13464 7546 13492 8774
rect 16224 8634 16252 12650
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16028 8424 16080 8430
rect 16028 8366 16080 8372
rect 15292 8356 15344 8362
rect 15292 8298 15344 8304
rect 14289 8188 14585 8208
rect 14345 8186 14369 8188
rect 14425 8186 14449 8188
rect 14505 8186 14529 8188
rect 14367 8134 14369 8186
rect 14431 8134 14443 8186
rect 14505 8134 14507 8186
rect 14345 8132 14369 8134
rect 14425 8132 14449 8134
rect 14505 8132 14529 8134
rect 14289 8112 14585 8132
rect 13912 7948 13964 7954
rect 13912 7890 13964 7896
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 13176 6928 13228 6934
rect 13176 6870 13228 6876
rect 13188 6458 13216 6870
rect 13464 6798 13492 7482
rect 13924 7449 13952 7890
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 14004 7472 14056 7478
rect 13910 7440 13966 7449
rect 14004 7414 14056 7420
rect 13910 7375 13966 7384
rect 13924 7342 13952 7375
rect 13912 7336 13964 7342
rect 13912 7278 13964 7284
rect 13912 7200 13964 7206
rect 13912 7142 13964 7148
rect 13452 6792 13504 6798
rect 13452 6734 13504 6740
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 13084 6180 13136 6186
rect 13084 6122 13136 6128
rect 13176 6180 13228 6186
rect 13176 6122 13228 6128
rect 13096 5846 13124 6122
rect 13084 5840 13136 5846
rect 13084 5782 13136 5788
rect 12992 5636 13044 5642
rect 12992 5578 13044 5584
rect 12820 4950 12940 4978
rect 12714 4040 12770 4049
rect 12714 3975 12770 3984
rect 12624 3664 12676 3670
rect 12624 3606 12676 3612
rect 12636 3505 12664 3606
rect 12622 3496 12678 3505
rect 12622 3431 12678 3440
rect 12716 3460 12768 3466
rect 12716 3402 12768 3408
rect 12530 3224 12586 3233
rect 12530 3159 12586 3168
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 10336 54 10562 82
rect 12164 128 12216 134
rect 12164 70 12216 76
rect 12544 82 12572 3159
rect 12728 3126 12756 3402
rect 12716 3120 12768 3126
rect 12716 3062 12768 3068
rect 12728 2922 12756 3062
rect 12716 2916 12768 2922
rect 12716 2858 12768 2864
rect 12820 2854 12848 4950
rect 13004 4154 13032 5578
rect 13096 5370 13124 5782
rect 13084 5364 13136 5370
rect 13084 5306 13136 5312
rect 13188 5234 13216 6122
rect 13924 5914 13952 7142
rect 13912 5908 13964 5914
rect 13912 5850 13964 5856
rect 13268 5704 13320 5710
rect 13268 5646 13320 5652
rect 13176 5228 13228 5234
rect 13176 5170 13228 5176
rect 12912 4146 13032 4154
rect 13188 4146 13216 5170
rect 13280 4826 13308 5646
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13728 5160 13780 5166
rect 13728 5102 13780 5108
rect 13268 4820 13320 4826
rect 13268 4762 13320 4768
rect 13740 4758 13768 5102
rect 13832 5098 13860 5306
rect 13820 5092 13872 5098
rect 13820 5034 13872 5040
rect 13832 4826 13860 5034
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13728 4752 13780 4758
rect 13728 4694 13780 4700
rect 13832 4146 13860 4762
rect 12900 4140 13032 4146
rect 12952 4126 13032 4140
rect 13176 4140 13228 4146
rect 12900 4082 12952 4088
rect 13176 4082 13228 4088
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 12990 4040 13046 4049
rect 12900 4004 12952 4010
rect 12990 3975 13046 3984
rect 12900 3946 12952 3952
rect 12912 3534 12940 3946
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 12808 2848 12860 2854
rect 12808 2790 12860 2796
rect 12820 2650 12848 2790
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 13004 2582 13032 3975
rect 13188 3126 13216 4082
rect 14016 4078 14044 7414
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 14289 7100 14585 7120
rect 14345 7098 14369 7100
rect 14425 7098 14449 7100
rect 14505 7098 14529 7100
rect 14367 7046 14369 7098
rect 14431 7046 14443 7098
rect 14505 7046 14507 7098
rect 14345 7044 14369 7046
rect 14425 7044 14449 7046
rect 14505 7044 14529 7046
rect 14289 7024 14585 7044
rect 14372 6656 14424 6662
rect 14372 6598 14424 6604
rect 14384 6322 14412 6598
rect 14372 6316 14424 6322
rect 14372 6258 14424 6264
rect 14188 6112 14240 6118
rect 14188 6054 14240 6060
rect 14200 5914 14228 6054
rect 14289 6012 14585 6032
rect 14345 6010 14369 6012
rect 14425 6010 14449 6012
rect 14505 6010 14529 6012
rect 14367 5958 14369 6010
rect 14431 5958 14443 6010
rect 14505 5958 14507 6010
rect 14345 5956 14369 5958
rect 14425 5956 14449 5958
rect 14505 5956 14529 5958
rect 14289 5936 14585 5956
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 14648 5568 14700 5574
rect 14648 5510 14700 5516
rect 14096 5296 14148 5302
rect 14096 5238 14148 5244
rect 14108 5001 14136 5238
rect 14094 4992 14150 5001
rect 14094 4927 14150 4936
rect 14289 4924 14585 4944
rect 14345 4922 14369 4924
rect 14425 4922 14449 4924
rect 14505 4922 14529 4924
rect 14367 4870 14369 4922
rect 14431 4870 14443 4922
rect 14505 4870 14507 4922
rect 14345 4868 14369 4870
rect 14425 4868 14449 4870
rect 14505 4868 14529 4870
rect 14289 4848 14585 4868
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 14004 4072 14056 4078
rect 14004 4014 14056 4020
rect 14200 3738 14228 4422
rect 14289 3836 14585 3856
rect 14345 3834 14369 3836
rect 14425 3834 14449 3836
rect 14505 3834 14529 3836
rect 14367 3782 14369 3834
rect 14431 3782 14443 3834
rect 14505 3782 14507 3834
rect 14345 3780 14369 3782
rect 14425 3780 14449 3782
rect 14505 3780 14529 3782
rect 14289 3760 14585 3780
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 13636 3664 13688 3670
rect 13636 3606 13688 3612
rect 14554 3632 14610 3641
rect 13648 3194 13676 3606
rect 14554 3567 14610 3576
rect 14188 3460 14240 3466
rect 14188 3402 14240 3408
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 13176 3120 13228 3126
rect 13176 3062 13228 3068
rect 14200 2922 14228 3402
rect 14568 3398 14596 3567
rect 14660 3398 14688 5510
rect 14752 5137 14780 7142
rect 14738 5128 14794 5137
rect 14738 5063 14794 5072
rect 14936 4690 14964 7686
rect 15106 7440 15162 7449
rect 15106 7375 15162 7384
rect 15016 4820 15068 4826
rect 15016 4762 15068 4768
rect 14924 4684 14976 4690
rect 14924 4626 14976 4632
rect 14830 4040 14886 4049
rect 14830 3975 14886 3984
rect 14844 3942 14872 3975
rect 14832 3936 14884 3942
rect 14832 3878 14884 3884
rect 14740 3664 14792 3670
rect 14740 3606 14792 3612
rect 14556 3392 14608 3398
rect 14556 3334 14608 3340
rect 14648 3392 14700 3398
rect 14648 3334 14700 3340
rect 14752 3126 14780 3606
rect 14740 3120 14792 3126
rect 14740 3062 14792 3068
rect 14188 2916 14240 2922
rect 14188 2858 14240 2864
rect 14289 2748 14585 2768
rect 14345 2746 14369 2748
rect 14425 2746 14449 2748
rect 14505 2746 14529 2748
rect 14367 2694 14369 2746
rect 14431 2694 14443 2746
rect 14505 2694 14507 2746
rect 14345 2692 14369 2694
rect 14425 2692 14449 2694
rect 14505 2692 14529 2694
rect 14289 2672 14585 2692
rect 14752 2582 14780 3062
rect 12992 2576 13044 2582
rect 12992 2518 13044 2524
rect 14740 2576 14792 2582
rect 14740 2518 14792 2524
rect 14936 2446 14964 4626
rect 15028 3738 15056 4762
rect 15016 3732 15068 3738
rect 15016 3674 15068 3680
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 12806 82 12862 480
rect 12544 54 12862 82
rect 15120 82 15148 7375
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 15212 5370 15240 6054
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 15200 3936 15252 3942
rect 15200 3878 15252 3884
rect 15212 2514 15240 3878
rect 15304 3602 15332 8298
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 15396 6934 15424 7822
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 15384 6928 15436 6934
rect 15384 6870 15436 6876
rect 15476 6928 15528 6934
rect 15476 6870 15528 6876
rect 15396 6458 15424 6870
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15488 6118 15516 6870
rect 15476 6112 15528 6118
rect 15476 6054 15528 6060
rect 15580 5846 15608 7142
rect 16040 6934 16068 8366
rect 16500 8090 16528 15506
rect 19720 12306 19748 15558
rect 19982 15520 20038 15558
rect 24136 15558 24454 15586
rect 20956 13084 21252 13104
rect 21012 13082 21036 13084
rect 21092 13082 21116 13084
rect 21172 13082 21196 13084
rect 21034 13030 21036 13082
rect 21098 13030 21110 13082
rect 21172 13030 21174 13082
rect 21012 13028 21036 13030
rect 21092 13028 21116 13030
rect 21172 13028 21196 13030
rect 20956 13008 21252 13028
rect 24136 12986 24164 15558
rect 24398 15520 24454 15558
rect 28552 15558 28962 15586
rect 27622 13628 27918 13648
rect 27678 13626 27702 13628
rect 27758 13626 27782 13628
rect 27838 13626 27862 13628
rect 27700 13574 27702 13626
rect 27764 13574 27776 13626
rect 27838 13574 27840 13626
rect 27678 13572 27702 13574
rect 27758 13572 27782 13574
rect 27838 13572 27862 13574
rect 27622 13552 27918 13572
rect 28552 12986 28580 15558
rect 28906 15520 28962 15558
rect 33152 15558 33378 15586
rect 24124 12980 24176 12986
rect 24124 12922 24176 12928
rect 28540 12980 28592 12986
rect 28540 12922 28592 12928
rect 24308 12776 24360 12782
rect 24308 12718 24360 12724
rect 26792 12776 26844 12782
rect 26792 12718 26844 12724
rect 24320 12646 24348 12718
rect 26804 12646 26832 12718
rect 24308 12640 24360 12646
rect 24308 12582 24360 12588
rect 26792 12640 26844 12646
rect 26792 12582 26844 12588
rect 19708 12300 19760 12306
rect 19708 12242 19760 12248
rect 19720 11898 19748 12242
rect 20956 11996 21252 12016
rect 21012 11994 21036 11996
rect 21092 11994 21116 11996
rect 21172 11994 21196 11996
rect 21034 11942 21036 11994
rect 21098 11942 21110 11994
rect 21172 11942 21174 11994
rect 21012 11940 21036 11942
rect 21092 11940 21116 11942
rect 21172 11940 21196 11942
rect 20956 11920 21252 11940
rect 19708 11892 19760 11898
rect 19708 11834 19760 11840
rect 19720 8634 19748 11834
rect 24320 11665 24348 12582
rect 24306 11656 24362 11665
rect 24306 11591 24362 11600
rect 20956 10908 21252 10928
rect 21012 10906 21036 10908
rect 21092 10906 21116 10908
rect 21172 10906 21196 10908
rect 21034 10854 21036 10906
rect 21098 10854 21110 10906
rect 21172 10854 21174 10906
rect 21012 10852 21036 10854
rect 21092 10852 21116 10854
rect 21172 10852 21196 10854
rect 20956 10832 21252 10852
rect 20956 9820 21252 9840
rect 21012 9818 21036 9820
rect 21092 9818 21116 9820
rect 21172 9818 21196 9820
rect 21034 9766 21036 9818
rect 21098 9766 21110 9818
rect 21172 9766 21174 9818
rect 21012 9764 21036 9766
rect 21092 9764 21116 9766
rect 21172 9764 21196 9766
rect 20956 9744 21252 9764
rect 20956 8732 21252 8752
rect 21012 8730 21036 8732
rect 21092 8730 21116 8732
rect 21172 8730 21196 8732
rect 21034 8678 21036 8730
rect 21098 8678 21110 8730
rect 21172 8678 21174 8730
rect 21012 8676 21036 8678
rect 21092 8676 21116 8678
rect 21172 8676 21196 8678
rect 20956 8656 21252 8676
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 24320 8090 24348 11591
rect 24674 10568 24730 10577
rect 24674 10503 24730 10512
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 24308 8084 24360 8090
rect 24308 8026 24360 8032
rect 16672 7948 16724 7954
rect 16672 7890 16724 7896
rect 16684 7206 16712 7890
rect 20956 7644 21252 7664
rect 21012 7642 21036 7644
rect 21092 7642 21116 7644
rect 21172 7642 21196 7644
rect 21034 7590 21036 7642
rect 21098 7590 21110 7642
rect 21172 7590 21174 7642
rect 21012 7588 21036 7590
rect 21092 7588 21116 7590
rect 21172 7588 21196 7590
rect 20956 7568 21252 7588
rect 24320 7342 24348 8026
rect 24688 7954 24716 10503
rect 24676 7948 24728 7954
rect 24676 7890 24728 7896
rect 24688 7546 24716 7890
rect 25136 7812 25188 7818
rect 25136 7754 25188 7760
rect 25044 7744 25096 7750
rect 25044 7686 25096 7692
rect 24676 7540 24728 7546
rect 24676 7482 24728 7488
rect 18236 7336 18288 7342
rect 18236 7278 18288 7284
rect 24308 7336 24360 7342
rect 24308 7278 24360 7284
rect 17592 7268 17644 7274
rect 17592 7210 17644 7216
rect 16672 7200 16724 7206
rect 16672 7142 16724 7148
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 16028 6928 16080 6934
rect 16028 6870 16080 6876
rect 16040 6322 16068 6870
rect 16684 6730 16712 7142
rect 16776 7002 16804 7142
rect 16764 6996 16816 7002
rect 16764 6938 16816 6944
rect 16672 6724 16724 6730
rect 16672 6666 16724 6672
rect 16776 6322 16804 6938
rect 17604 6934 17632 7210
rect 17592 6928 17644 6934
rect 17592 6870 17644 6876
rect 17604 6458 17632 6870
rect 17868 6792 17920 6798
rect 17868 6734 17920 6740
rect 17880 6458 17908 6734
rect 17592 6452 17644 6458
rect 17592 6394 17644 6400
rect 17868 6452 17920 6458
rect 17868 6394 17920 6400
rect 16028 6316 16080 6322
rect 16028 6258 16080 6264
rect 16764 6316 16816 6322
rect 16764 6258 16816 6264
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 15568 5840 15620 5846
rect 15568 5782 15620 5788
rect 15844 5840 15896 5846
rect 15844 5782 15896 5788
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 15396 4758 15424 5510
rect 15856 5234 15884 5782
rect 15844 5228 15896 5234
rect 15844 5170 15896 5176
rect 16040 4758 16068 6258
rect 16868 5846 16896 6258
rect 18248 6186 18276 7278
rect 25056 7274 25084 7686
rect 25148 7410 25176 7754
rect 25136 7404 25188 7410
rect 25136 7346 25188 7352
rect 24400 7268 24452 7274
rect 24400 7210 24452 7216
rect 25044 7268 25096 7274
rect 25044 7210 25096 7216
rect 25780 7268 25832 7274
rect 25780 7210 25832 7216
rect 18328 7200 18380 7206
rect 18328 7142 18380 7148
rect 17224 6180 17276 6186
rect 17224 6122 17276 6128
rect 18236 6180 18288 6186
rect 18236 6122 18288 6128
rect 16856 5840 16908 5846
rect 16856 5782 16908 5788
rect 16764 5772 16816 5778
rect 16764 5714 16816 5720
rect 16304 5364 16356 5370
rect 16304 5306 16356 5312
rect 16316 5098 16344 5306
rect 16776 5166 16804 5714
rect 17132 5568 17184 5574
rect 17132 5510 17184 5516
rect 16764 5160 16816 5166
rect 16764 5102 16816 5108
rect 16304 5092 16356 5098
rect 16304 5034 16356 5040
rect 16856 5092 16908 5098
rect 16856 5034 16908 5040
rect 15384 4752 15436 4758
rect 15384 4694 15436 4700
rect 16028 4752 16080 4758
rect 16028 4694 16080 4700
rect 15396 3670 15424 4694
rect 15566 4448 15622 4457
rect 15566 4383 15622 4392
rect 15580 4282 15608 4383
rect 15568 4276 15620 4282
rect 15568 4218 15620 4224
rect 15936 4072 15988 4078
rect 15936 4014 15988 4020
rect 15844 4004 15896 4010
rect 15844 3946 15896 3952
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 15384 3664 15436 3670
rect 15384 3606 15436 3612
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 15304 3194 15332 3538
rect 15672 3505 15700 3878
rect 15856 3602 15884 3946
rect 15948 3670 15976 4014
rect 15936 3664 15988 3670
rect 15936 3606 15988 3612
rect 15844 3596 15896 3602
rect 15844 3538 15896 3544
rect 15658 3496 15714 3505
rect 15658 3431 15714 3440
rect 15672 3194 15700 3431
rect 15856 3398 15884 3538
rect 15844 3392 15896 3398
rect 15842 3360 15844 3369
rect 15896 3360 15898 3369
rect 15842 3295 15898 3304
rect 15856 3269 15884 3295
rect 15292 3188 15344 3194
rect 15292 3130 15344 3136
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 16316 2650 16344 5034
rect 16580 4752 16632 4758
rect 16500 4729 16580 4740
rect 16486 4720 16580 4729
rect 16542 4712 16580 4720
rect 16580 4694 16632 4700
rect 16486 4655 16542 4664
rect 16488 4548 16540 4554
rect 16488 4490 16540 4496
rect 16500 3058 16528 4490
rect 16488 3052 16540 3058
rect 16488 2994 16540 3000
rect 16304 2644 16356 2650
rect 16304 2586 16356 2592
rect 16868 2553 16896 5034
rect 17040 4820 17092 4826
rect 17040 4762 17092 4768
rect 17052 4593 17080 4762
rect 17038 4584 17094 4593
rect 17038 4519 17094 4528
rect 17144 4146 17172 5510
rect 17236 5234 17264 6122
rect 18248 5914 18276 6122
rect 17592 5908 17644 5914
rect 17592 5850 17644 5856
rect 18236 5908 18288 5914
rect 18236 5850 18288 5856
rect 17604 5370 17632 5850
rect 18144 5772 18196 5778
rect 18144 5714 18196 5720
rect 17592 5364 17644 5370
rect 17592 5306 17644 5312
rect 17224 5228 17276 5234
rect 17224 5170 17276 5176
rect 17224 4684 17276 4690
rect 17224 4626 17276 4632
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 17776 4684 17828 4690
rect 17776 4626 17828 4632
rect 17236 4146 17264 4626
rect 17132 4140 17184 4146
rect 17132 4082 17184 4088
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17132 3936 17184 3942
rect 17132 3878 17184 3884
rect 17144 3398 17172 3878
rect 17236 3670 17264 4082
rect 17328 3942 17356 4626
rect 17500 4616 17552 4622
rect 17420 4576 17500 4604
rect 17420 4078 17448 4576
rect 17500 4558 17552 4564
rect 17788 4486 17816 4626
rect 17776 4480 17828 4486
rect 17776 4422 17828 4428
rect 17500 4208 17552 4214
rect 17500 4150 17552 4156
rect 17408 4072 17460 4078
rect 17408 4014 17460 4020
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 17224 3664 17276 3670
rect 17224 3606 17276 3612
rect 17316 3596 17368 3602
rect 17316 3538 17368 3544
rect 17132 3392 17184 3398
rect 17132 3334 17184 3340
rect 16948 2916 17000 2922
rect 16948 2858 17000 2864
rect 16960 2650 16988 2858
rect 16948 2644 17000 2650
rect 16948 2586 17000 2592
rect 16854 2544 16910 2553
rect 15200 2508 15252 2514
rect 16854 2479 16910 2488
rect 15200 2450 15252 2456
rect 16960 2446 16988 2586
rect 17144 2582 17172 3334
rect 17328 3126 17356 3538
rect 17420 3194 17448 4014
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 17316 3120 17368 3126
rect 17316 3062 17368 3068
rect 17328 2990 17356 3062
rect 17316 2984 17368 2990
rect 17316 2926 17368 2932
rect 17132 2576 17184 2582
rect 17132 2518 17184 2524
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 15198 82 15254 480
rect 15120 54 15254 82
rect 17512 82 17540 4150
rect 17682 4040 17738 4049
rect 17682 3975 17738 3984
rect 17696 3942 17724 3975
rect 17684 3936 17736 3942
rect 17684 3878 17736 3884
rect 17696 3602 17724 3878
rect 17788 3670 17816 4422
rect 18156 3942 18184 5714
rect 18340 4690 18368 7142
rect 20168 6860 20220 6866
rect 20168 6802 20220 6808
rect 21364 6860 21416 6866
rect 21364 6802 21416 6808
rect 21916 6860 21968 6866
rect 21916 6802 21968 6808
rect 22100 6860 22152 6866
rect 22100 6802 22152 6808
rect 23296 6860 23348 6866
rect 23296 6802 23348 6808
rect 18512 6724 18564 6730
rect 18512 6666 18564 6672
rect 18420 6656 18472 6662
rect 18420 6598 18472 6604
rect 18432 6322 18460 6598
rect 18524 6322 18552 6666
rect 20180 6662 20208 6802
rect 20168 6656 20220 6662
rect 20168 6598 20220 6604
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 18420 6316 18472 6322
rect 18420 6258 18472 6264
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 20180 6254 20208 6598
rect 20640 6304 20668 6598
rect 20956 6556 21252 6576
rect 21012 6554 21036 6556
rect 21092 6554 21116 6556
rect 21172 6554 21196 6556
rect 21034 6502 21036 6554
rect 21098 6502 21110 6554
rect 21172 6502 21174 6554
rect 21012 6500 21036 6502
rect 21092 6500 21116 6502
rect 21172 6500 21196 6502
rect 20956 6480 21252 6500
rect 20720 6316 20772 6322
rect 20640 6276 20720 6304
rect 19432 6248 19484 6254
rect 19432 6190 19484 6196
rect 20168 6248 20220 6254
rect 20168 6190 20220 6196
rect 18328 4684 18380 4690
rect 18328 4626 18380 4632
rect 18420 4480 18472 4486
rect 18420 4422 18472 4428
rect 19156 4480 19208 4486
rect 19156 4422 19208 4428
rect 19248 4480 19300 4486
rect 19248 4422 19300 4428
rect 18432 4078 18460 4422
rect 18880 4208 18932 4214
rect 18880 4150 18932 4156
rect 18236 4072 18288 4078
rect 18236 4014 18288 4020
rect 18420 4072 18472 4078
rect 18892 4049 18920 4150
rect 19168 4146 19196 4422
rect 19156 4140 19208 4146
rect 19156 4082 19208 4088
rect 19064 4072 19116 4078
rect 18420 4014 18472 4020
rect 18878 4040 18934 4049
rect 18144 3936 18196 3942
rect 18144 3878 18196 3884
rect 17776 3664 17828 3670
rect 17776 3606 17828 3612
rect 18248 3602 18276 4014
rect 18432 3602 18460 4014
rect 19064 4014 19116 4020
rect 18878 3975 18934 3984
rect 18892 3720 18920 3975
rect 18892 3692 19012 3720
rect 18984 3602 19012 3692
rect 19076 3670 19104 4014
rect 19064 3664 19116 3670
rect 19064 3606 19116 3612
rect 17684 3596 17736 3602
rect 17684 3538 17736 3544
rect 18236 3596 18288 3602
rect 18236 3538 18288 3544
rect 18420 3596 18472 3602
rect 18420 3538 18472 3544
rect 18880 3596 18932 3602
rect 18880 3538 18932 3544
rect 18972 3596 19024 3602
rect 18972 3538 19024 3544
rect 17868 2848 17920 2854
rect 17868 2790 17920 2796
rect 17880 2514 17908 2790
rect 17868 2508 17920 2514
rect 17868 2450 17920 2456
rect 18248 2310 18276 3538
rect 18432 3398 18460 3538
rect 18420 3392 18472 3398
rect 18420 3334 18472 3340
rect 18432 2990 18460 3334
rect 18892 3194 18920 3538
rect 19260 3534 19288 4422
rect 19444 4282 19472 6190
rect 19708 6112 19760 6118
rect 19708 6054 19760 6060
rect 19524 5568 19576 5574
rect 19524 5510 19576 5516
rect 19536 5030 19564 5510
rect 19524 5024 19576 5030
rect 19524 4966 19576 4972
rect 19536 4622 19564 4966
rect 19720 4758 19748 6054
rect 20640 5914 20668 6276
rect 20720 6258 20772 6264
rect 21272 6248 21324 6254
rect 21272 6190 21324 6196
rect 20628 5908 20680 5914
rect 20628 5850 20680 5856
rect 19800 5772 19852 5778
rect 19800 5714 19852 5720
rect 20444 5772 20496 5778
rect 20444 5714 20496 5720
rect 19812 5098 19840 5714
rect 20456 5302 20484 5714
rect 20628 5704 20680 5710
rect 20628 5646 20680 5652
rect 20444 5296 20496 5302
rect 20444 5238 20496 5244
rect 20456 5166 20484 5238
rect 20640 5166 20668 5646
rect 20956 5468 21252 5488
rect 21012 5466 21036 5468
rect 21092 5466 21116 5468
rect 21172 5466 21196 5468
rect 21034 5414 21036 5466
rect 21098 5414 21110 5466
rect 21172 5414 21174 5466
rect 21012 5412 21036 5414
rect 21092 5412 21116 5414
rect 21172 5412 21196 5414
rect 20956 5392 21252 5412
rect 20444 5160 20496 5166
rect 20444 5102 20496 5108
rect 20628 5160 20680 5166
rect 20628 5102 20680 5108
rect 19800 5092 19852 5098
rect 19800 5034 19852 5040
rect 20640 4758 20668 5102
rect 21284 5030 21312 6190
rect 21376 6118 21404 6802
rect 21928 6254 21956 6802
rect 22112 6322 22140 6802
rect 22100 6316 22152 6322
rect 22100 6258 22152 6264
rect 21916 6248 21968 6254
rect 21916 6190 21968 6196
rect 21640 6180 21692 6186
rect 21640 6122 21692 6128
rect 21364 6112 21416 6118
rect 21364 6054 21416 6060
rect 21652 5234 21680 6122
rect 21928 5778 21956 6190
rect 22112 5778 22140 6258
rect 23308 6118 23336 6802
rect 23572 6792 23624 6798
rect 23572 6734 23624 6740
rect 23584 6322 23612 6734
rect 23572 6316 23624 6322
rect 23572 6258 23624 6264
rect 24412 6118 24440 7210
rect 24492 7200 24544 7206
rect 24492 7142 24544 7148
rect 24504 6934 24532 7142
rect 24492 6928 24544 6934
rect 24492 6870 24544 6876
rect 25044 6928 25096 6934
rect 25044 6870 25096 6876
rect 22192 6112 22244 6118
rect 22192 6054 22244 6060
rect 23020 6112 23072 6118
rect 23020 6054 23072 6060
rect 23296 6112 23348 6118
rect 23296 6054 23348 6060
rect 24032 6112 24084 6118
rect 24032 6054 24084 6060
rect 24400 6112 24452 6118
rect 24400 6054 24452 6060
rect 21916 5772 21968 5778
rect 21916 5714 21968 5720
rect 22100 5772 22152 5778
rect 22100 5714 22152 5720
rect 21640 5228 21692 5234
rect 21640 5170 21692 5176
rect 21272 5024 21324 5030
rect 21272 4966 21324 4972
rect 19708 4752 19760 4758
rect 19708 4694 19760 4700
rect 20628 4752 20680 4758
rect 20628 4694 20680 4700
rect 19892 4684 19944 4690
rect 19892 4626 19944 4632
rect 20720 4684 20772 4690
rect 20720 4626 20772 4632
rect 19524 4616 19576 4622
rect 19524 4558 19576 4564
rect 19432 4276 19484 4282
rect 19432 4218 19484 4224
rect 19444 4078 19472 4218
rect 19904 4214 19932 4626
rect 19892 4208 19944 4214
rect 19892 4150 19944 4156
rect 20732 4078 20760 4626
rect 20956 4380 21252 4400
rect 21012 4378 21036 4380
rect 21092 4378 21116 4380
rect 21172 4378 21196 4380
rect 21034 4326 21036 4378
rect 21098 4326 21110 4378
rect 21172 4326 21174 4378
rect 21012 4324 21036 4326
rect 21092 4324 21116 4326
rect 21172 4324 21196 4326
rect 20956 4304 21252 4324
rect 21284 4078 21312 4966
rect 21928 4826 21956 5714
rect 22112 5166 22140 5714
rect 22204 5370 22232 6054
rect 23032 5846 23060 6054
rect 23020 5840 23072 5846
rect 23308 5817 23336 6054
rect 23020 5782 23072 5788
rect 23294 5808 23350 5817
rect 23032 5370 23060 5782
rect 23294 5743 23350 5752
rect 23204 5704 23256 5710
rect 23204 5646 23256 5652
rect 22192 5364 22244 5370
rect 22192 5306 22244 5312
rect 23020 5364 23072 5370
rect 23020 5306 23072 5312
rect 22100 5160 22152 5166
rect 22100 5102 22152 5108
rect 21916 4820 21968 4826
rect 21916 4762 21968 4768
rect 22112 4690 22140 5102
rect 23216 4826 23244 5646
rect 24044 5370 24072 6054
rect 24412 5914 24440 6054
rect 24504 5914 24532 6870
rect 25056 6458 25084 6870
rect 25792 6730 25820 7210
rect 26700 6928 26752 6934
rect 26700 6870 26752 6876
rect 26056 6792 26108 6798
rect 26056 6734 26108 6740
rect 26608 6792 26660 6798
rect 26608 6734 26660 6740
rect 25780 6724 25832 6730
rect 25780 6666 25832 6672
rect 25136 6656 25188 6662
rect 25136 6598 25188 6604
rect 25044 6452 25096 6458
rect 25044 6394 25096 6400
rect 25148 6322 25176 6598
rect 25792 6322 25820 6666
rect 26068 6390 26096 6734
rect 26424 6724 26476 6730
rect 26424 6666 26476 6672
rect 26056 6384 26108 6390
rect 26056 6326 26108 6332
rect 25136 6316 25188 6322
rect 25136 6258 25188 6264
rect 25780 6316 25832 6322
rect 25780 6258 25832 6264
rect 24400 5908 24452 5914
rect 24400 5850 24452 5856
rect 24492 5908 24544 5914
rect 24492 5850 24544 5856
rect 25148 5710 25176 6258
rect 25596 6180 25648 6186
rect 25596 6122 25648 6128
rect 25608 5846 25636 6122
rect 25596 5840 25648 5846
rect 25596 5782 25648 5788
rect 25504 5772 25556 5778
rect 25504 5714 25556 5720
rect 25136 5704 25188 5710
rect 25136 5646 25188 5652
rect 24032 5364 24084 5370
rect 24032 5306 24084 5312
rect 24044 5166 24072 5306
rect 24216 5228 24268 5234
rect 24216 5170 24268 5176
rect 24032 5160 24084 5166
rect 24032 5102 24084 5108
rect 22560 4820 22612 4826
rect 22560 4762 22612 4768
rect 23204 4820 23256 4826
rect 23204 4762 23256 4768
rect 21364 4684 21416 4690
rect 21364 4626 21416 4632
rect 21732 4684 21784 4690
rect 21732 4626 21784 4632
rect 22100 4684 22152 4690
rect 22100 4626 22152 4632
rect 19432 4072 19484 4078
rect 19432 4014 19484 4020
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 21272 4072 21324 4078
rect 21272 4014 21324 4020
rect 20444 3936 20496 3942
rect 20444 3878 20496 3884
rect 19984 3732 20036 3738
rect 19984 3674 20036 3680
rect 19340 3596 19392 3602
rect 19340 3538 19392 3544
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 19352 3233 19380 3538
rect 19338 3224 19394 3233
rect 18880 3188 18932 3194
rect 19338 3159 19394 3168
rect 18880 3130 18932 3136
rect 18892 2990 18920 3130
rect 19248 3120 19300 3126
rect 19248 3062 19300 3068
rect 19260 2990 19288 3062
rect 18328 2984 18380 2990
rect 18328 2926 18380 2932
rect 18420 2984 18472 2990
rect 18420 2926 18472 2932
rect 18880 2984 18932 2990
rect 18880 2926 18932 2932
rect 19248 2984 19300 2990
rect 19248 2926 19300 2932
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 18236 2304 18288 2310
rect 18236 2246 18288 2252
rect 18340 1873 18368 2926
rect 18432 2854 18460 2926
rect 18420 2848 18472 2854
rect 18420 2790 18472 2796
rect 18892 2378 18920 2926
rect 19064 2916 19116 2922
rect 19064 2858 19116 2864
rect 19076 2514 19104 2858
rect 19352 2650 19380 2926
rect 19340 2644 19392 2650
rect 19340 2586 19392 2592
rect 19064 2508 19116 2514
rect 19064 2450 19116 2456
rect 18880 2372 18932 2378
rect 18880 2314 18932 2320
rect 18326 1864 18382 1873
rect 18326 1799 18382 1808
rect 17590 82 17646 480
rect 17512 54 17646 82
rect 10506 0 10562 54
rect 12806 0 12862 54
rect 15198 0 15254 54
rect 17590 0 17646 54
rect 19890 82 19946 480
rect 19996 82 20024 3674
rect 20456 3641 20484 3878
rect 20732 3670 20760 4014
rect 21376 4010 21404 4626
rect 21640 4616 21692 4622
rect 21640 4558 21692 4564
rect 21652 4078 21680 4558
rect 21640 4072 21692 4078
rect 21744 4049 21772 4626
rect 22572 4282 22600 4762
rect 23664 4480 23716 4486
rect 23664 4422 23716 4428
rect 22560 4276 22612 4282
rect 22560 4218 22612 4224
rect 23676 4146 23704 4422
rect 24044 4282 24072 5102
rect 24228 4826 24256 5170
rect 24400 5092 24452 5098
rect 24400 5034 24452 5040
rect 24768 5092 24820 5098
rect 24768 5034 24820 5040
rect 24216 4820 24268 4826
rect 24216 4762 24268 4768
rect 24412 4758 24440 5034
rect 24780 4826 24808 5034
rect 25516 5030 25544 5714
rect 25608 5370 25636 5782
rect 26068 5642 26096 6326
rect 26056 5636 26108 5642
rect 26056 5578 26108 5584
rect 25596 5364 25648 5370
rect 25596 5306 25648 5312
rect 26068 5234 26096 5578
rect 26056 5228 26108 5234
rect 26056 5170 26108 5176
rect 25504 5024 25556 5030
rect 25504 4966 25556 4972
rect 25780 5024 25832 5030
rect 25780 4966 25832 4972
rect 24768 4820 24820 4826
rect 24768 4762 24820 4768
rect 24400 4752 24452 4758
rect 24400 4694 24452 4700
rect 24676 4616 24728 4622
rect 24676 4558 24728 4564
rect 24032 4276 24084 4282
rect 24032 4218 24084 4224
rect 23664 4140 23716 4146
rect 23664 4082 23716 4088
rect 21640 4014 21692 4020
rect 21730 4040 21786 4049
rect 21364 4004 21416 4010
rect 21364 3946 21416 3952
rect 21652 3738 21680 4014
rect 21730 3975 21786 3984
rect 24044 3942 24072 4218
rect 24032 3936 24084 3942
rect 24032 3878 24084 3884
rect 24584 3936 24636 3942
rect 24584 3878 24636 3884
rect 21640 3732 21692 3738
rect 21640 3674 21692 3680
rect 24044 3670 24072 3878
rect 20720 3664 20772 3670
rect 20442 3632 20498 3641
rect 20720 3606 20772 3612
rect 24032 3664 24084 3670
rect 24032 3606 24084 3612
rect 20442 3567 20498 3576
rect 21456 3596 21508 3602
rect 20456 3534 20484 3567
rect 21456 3538 21508 3544
rect 23480 3596 23532 3602
rect 23480 3538 23532 3544
rect 20444 3528 20496 3534
rect 20444 3470 20496 3476
rect 20994 3496 21050 3505
rect 20904 3460 20956 3466
rect 20956 3440 20994 3448
rect 20956 3431 21050 3440
rect 20956 3420 21036 3431
rect 20904 3402 20956 3408
rect 20956 3292 21252 3312
rect 21012 3290 21036 3292
rect 21092 3290 21116 3292
rect 21172 3290 21196 3292
rect 21034 3238 21036 3290
rect 21098 3238 21110 3290
rect 21172 3238 21174 3290
rect 21012 3236 21036 3238
rect 21092 3236 21116 3238
rect 21172 3236 21196 3238
rect 20956 3216 21252 3236
rect 20352 2916 20404 2922
rect 20352 2858 20404 2864
rect 20364 2582 20392 2858
rect 21468 2854 21496 3538
rect 23492 3505 23520 3538
rect 23478 3496 23534 3505
rect 23478 3431 23534 3440
rect 23492 3194 23520 3431
rect 23480 3188 23532 3194
rect 23480 3130 23532 3136
rect 24044 3126 24072 3606
rect 24032 3120 24084 3126
rect 24032 3062 24084 3068
rect 24596 2922 24624 3878
rect 24688 3738 24716 4558
rect 24780 4214 24808 4762
rect 25412 4752 25464 4758
rect 25412 4694 25464 4700
rect 24768 4208 24820 4214
rect 24768 4150 24820 4156
rect 25424 4146 25452 4694
rect 25412 4140 25464 4146
rect 25412 4082 25464 4088
rect 24676 3732 24728 3738
rect 24676 3674 24728 3680
rect 25516 3602 25544 4966
rect 25792 4826 25820 4966
rect 26068 4826 26096 5170
rect 25780 4820 25832 4826
rect 25780 4762 25832 4768
rect 26056 4820 26108 4826
rect 26056 4762 26108 4768
rect 26436 4622 26464 6666
rect 26620 5914 26648 6734
rect 26712 6458 26740 6870
rect 26700 6452 26752 6458
rect 26700 6394 26752 6400
rect 26608 5908 26660 5914
rect 26608 5850 26660 5856
rect 26608 5704 26660 5710
rect 26608 5646 26660 5652
rect 26620 5370 26648 5646
rect 26608 5364 26660 5370
rect 26608 5306 26660 5312
rect 26700 4752 26752 4758
rect 26700 4694 26752 4700
rect 26424 4616 26476 4622
rect 26424 4558 26476 4564
rect 26436 4214 26464 4558
rect 26712 4282 26740 4694
rect 26700 4276 26752 4282
rect 26700 4218 26752 4224
rect 26424 4208 26476 4214
rect 26424 4150 26476 4156
rect 26804 4146 26832 12582
rect 27622 12540 27918 12560
rect 27678 12538 27702 12540
rect 27758 12538 27782 12540
rect 27838 12538 27862 12540
rect 27700 12486 27702 12538
rect 27764 12486 27776 12538
rect 27838 12486 27840 12538
rect 27678 12484 27702 12486
rect 27758 12484 27782 12486
rect 27838 12484 27862 12486
rect 27622 12464 27918 12484
rect 27622 11452 27918 11472
rect 27678 11450 27702 11452
rect 27758 11450 27782 11452
rect 27838 11450 27862 11452
rect 27700 11398 27702 11450
rect 27764 11398 27776 11450
rect 27838 11398 27840 11450
rect 27678 11396 27702 11398
rect 27758 11396 27782 11398
rect 27838 11396 27862 11398
rect 27622 11376 27918 11396
rect 27622 10364 27918 10384
rect 27678 10362 27702 10364
rect 27758 10362 27782 10364
rect 27838 10362 27862 10364
rect 27700 10310 27702 10362
rect 27764 10310 27776 10362
rect 27838 10310 27840 10362
rect 27678 10308 27702 10310
rect 27758 10308 27782 10310
rect 27838 10308 27862 10310
rect 27622 10288 27918 10308
rect 27622 9276 27918 9296
rect 27678 9274 27702 9276
rect 27758 9274 27782 9276
rect 27838 9274 27862 9276
rect 27700 9222 27702 9274
rect 27764 9222 27776 9274
rect 27838 9222 27840 9274
rect 27678 9220 27702 9222
rect 27758 9220 27782 9222
rect 27838 9220 27862 9222
rect 27622 9200 27918 9220
rect 27622 8188 27918 8208
rect 27678 8186 27702 8188
rect 27758 8186 27782 8188
rect 27838 8186 27862 8188
rect 27700 8134 27702 8186
rect 27764 8134 27776 8186
rect 27838 8134 27840 8186
rect 27678 8132 27702 8134
rect 27758 8132 27782 8134
rect 27838 8132 27862 8134
rect 27622 8112 27918 8132
rect 33152 8090 33180 15558
rect 33322 15520 33378 15558
rect 37738 15586 37794 16000
rect 37738 15558 37872 15586
rect 37738 15520 37794 15558
rect 35622 13696 35678 13705
rect 35622 13631 35678 13640
rect 34289 13084 34585 13104
rect 34345 13082 34369 13084
rect 34425 13082 34449 13084
rect 34505 13082 34529 13084
rect 34367 13030 34369 13082
rect 34431 13030 34443 13082
rect 34505 13030 34507 13082
rect 34345 13028 34369 13030
rect 34425 13028 34449 13030
rect 34505 13028 34529 13030
rect 34289 13008 34585 13028
rect 35636 12986 35664 13631
rect 35624 12980 35676 12986
rect 35624 12922 35676 12928
rect 35256 12776 35308 12782
rect 35256 12718 35308 12724
rect 34289 11996 34585 12016
rect 34345 11994 34369 11996
rect 34425 11994 34449 11996
rect 34505 11994 34529 11996
rect 34367 11942 34369 11994
rect 34431 11942 34443 11994
rect 34505 11942 34507 11994
rect 34345 11940 34369 11942
rect 34425 11940 34449 11942
rect 34505 11940 34529 11942
rect 34289 11920 34585 11940
rect 34289 10908 34585 10928
rect 34345 10906 34369 10908
rect 34425 10906 34449 10908
rect 34505 10906 34529 10908
rect 34367 10854 34369 10906
rect 34431 10854 34443 10906
rect 34505 10854 34507 10906
rect 34345 10852 34369 10854
rect 34425 10852 34449 10854
rect 34505 10852 34529 10854
rect 34289 10832 34585 10852
rect 34289 9820 34585 9840
rect 34345 9818 34369 9820
rect 34425 9818 34449 9820
rect 34505 9818 34529 9820
rect 34367 9766 34369 9818
rect 34431 9766 34443 9818
rect 34505 9766 34507 9818
rect 34345 9764 34369 9766
rect 34425 9764 34449 9766
rect 34505 9764 34529 9766
rect 34289 9744 34585 9764
rect 34289 8732 34585 8752
rect 34345 8730 34369 8732
rect 34425 8730 34449 8732
rect 34505 8730 34529 8732
rect 34367 8678 34369 8730
rect 34431 8678 34443 8730
rect 34505 8678 34507 8730
rect 34345 8676 34369 8678
rect 34425 8676 34449 8678
rect 34505 8676 34529 8678
rect 34289 8656 34585 8676
rect 33140 8084 33192 8090
rect 33140 8026 33192 8032
rect 32220 7948 32272 7954
rect 32220 7890 32272 7896
rect 32232 7313 32260 7890
rect 34289 7644 34585 7664
rect 34345 7642 34369 7644
rect 34425 7642 34449 7644
rect 34505 7642 34529 7644
rect 34367 7590 34369 7642
rect 34431 7590 34443 7642
rect 34505 7590 34507 7642
rect 34345 7588 34369 7590
rect 34425 7588 34449 7590
rect 34505 7588 34529 7590
rect 34289 7568 34585 7588
rect 35268 7449 35296 12718
rect 37844 11665 37872 15558
rect 39578 15328 39634 15337
rect 39578 15263 39634 15272
rect 39592 12714 39620 15263
rect 39580 12708 39632 12714
rect 39580 12650 39632 12656
rect 39578 12608 39634 12617
rect 39578 12543 39634 12552
rect 39592 12102 39620 12543
rect 39580 12096 39632 12102
rect 39580 12038 39632 12044
rect 37830 11656 37886 11665
rect 37830 11591 37886 11600
rect 39580 11348 39632 11354
rect 39580 11290 39632 11296
rect 39592 11257 39620 11290
rect 39578 11248 39634 11257
rect 35440 11212 35492 11218
rect 39578 11183 39634 11192
rect 35440 11154 35492 11160
rect 35452 10674 35480 11154
rect 35440 10668 35492 10674
rect 35440 10610 35492 10616
rect 35452 10577 35480 10610
rect 35438 10568 35494 10577
rect 35438 10503 35494 10512
rect 35622 9344 35678 9353
rect 35622 9279 35678 9288
rect 35636 9178 35664 9279
rect 35624 9172 35676 9178
rect 35624 9114 35676 9120
rect 35440 9036 35492 9042
rect 35440 8978 35492 8984
rect 35452 8294 35480 8978
rect 35440 8288 35492 8294
rect 35440 8230 35492 8236
rect 35254 7440 35310 7449
rect 35254 7375 35310 7384
rect 32218 7304 32274 7313
rect 32218 7239 32274 7248
rect 32232 7206 32260 7239
rect 32220 7200 32272 7206
rect 32220 7142 32272 7148
rect 27622 7100 27918 7120
rect 27678 7098 27702 7100
rect 27758 7098 27782 7100
rect 27838 7098 27862 7100
rect 27700 7046 27702 7098
rect 27764 7046 27776 7098
rect 27838 7046 27840 7098
rect 27678 7044 27702 7046
rect 27758 7044 27782 7046
rect 27838 7044 27862 7046
rect 27622 7024 27918 7044
rect 27988 6656 28040 6662
rect 27988 6598 28040 6604
rect 28000 6322 28028 6598
rect 32232 6458 32260 7142
rect 34612 6860 34664 6866
rect 34612 6802 34664 6808
rect 34289 6556 34585 6576
rect 34345 6554 34369 6556
rect 34425 6554 34449 6556
rect 34505 6554 34529 6556
rect 34367 6502 34369 6554
rect 34431 6502 34443 6554
rect 34505 6502 34507 6554
rect 34345 6500 34369 6502
rect 34425 6500 34449 6502
rect 34505 6500 34529 6502
rect 34289 6480 34585 6500
rect 32220 6452 32272 6458
rect 32220 6394 32272 6400
rect 27988 6316 28040 6322
rect 27988 6258 28040 6264
rect 27622 6012 27918 6032
rect 27678 6010 27702 6012
rect 27758 6010 27782 6012
rect 27838 6010 27862 6012
rect 27700 5958 27702 6010
rect 27764 5958 27776 6010
rect 27838 5958 27840 6010
rect 27678 5956 27702 5958
rect 27758 5956 27782 5958
rect 27838 5956 27862 5958
rect 27622 5936 27918 5956
rect 28000 5914 28028 6258
rect 34624 6254 34652 6802
rect 34612 6248 34664 6254
rect 35452 6225 35480 8230
rect 36082 8120 36138 8129
rect 36082 8055 36138 8064
rect 36096 6458 36124 8055
rect 36084 6452 36136 6458
rect 36084 6394 36136 6400
rect 36096 6254 36124 6394
rect 39580 6384 39632 6390
rect 39580 6326 39632 6332
rect 36084 6248 36136 6254
rect 34612 6190 34664 6196
rect 35438 6216 35494 6225
rect 36084 6190 36136 6196
rect 35438 6151 35494 6160
rect 31392 6112 31444 6118
rect 31392 6054 31444 6060
rect 27988 5908 28040 5914
rect 27988 5850 28040 5856
rect 26976 5840 27028 5846
rect 26976 5782 27028 5788
rect 26988 5302 27016 5782
rect 27436 5364 27488 5370
rect 27436 5306 27488 5312
rect 26976 5296 27028 5302
rect 26976 5238 27028 5244
rect 26884 5092 26936 5098
rect 26884 5034 26936 5040
rect 26896 4622 26924 5034
rect 26884 4616 26936 4622
rect 26884 4558 26936 4564
rect 26792 4140 26844 4146
rect 26792 4082 26844 4088
rect 25504 3596 25556 3602
rect 25504 3538 25556 3544
rect 25228 3528 25280 3534
rect 25228 3470 25280 3476
rect 25240 3058 25268 3470
rect 25228 3052 25280 3058
rect 25228 2994 25280 3000
rect 24584 2916 24636 2922
rect 24584 2858 24636 2864
rect 25136 2916 25188 2922
rect 25136 2858 25188 2864
rect 21456 2848 21508 2854
rect 21456 2790 21508 2796
rect 22284 2848 22336 2854
rect 22284 2790 22336 2796
rect 21468 2582 21496 2790
rect 20352 2576 20404 2582
rect 20352 2518 20404 2524
rect 21456 2576 21508 2582
rect 22296 2553 22324 2790
rect 25148 2650 25176 2858
rect 25136 2644 25188 2650
rect 25136 2586 25188 2592
rect 21456 2518 21508 2524
rect 22282 2544 22338 2553
rect 20076 2508 20128 2514
rect 20076 2450 20128 2456
rect 21272 2508 21324 2514
rect 21272 2450 21324 2456
rect 20088 2145 20116 2450
rect 21284 2417 21312 2450
rect 21270 2408 21326 2417
rect 21270 2343 21326 2352
rect 20956 2204 21252 2224
rect 21012 2202 21036 2204
rect 21092 2202 21116 2204
rect 21172 2202 21196 2204
rect 21034 2150 21036 2202
rect 21098 2150 21110 2202
rect 21172 2150 21174 2202
rect 21012 2148 21036 2150
rect 21092 2148 21116 2150
rect 21172 2148 21196 2150
rect 20074 2136 20130 2145
rect 20956 2128 21252 2148
rect 20074 2071 20130 2080
rect 21468 1465 21496 2518
rect 25516 2514 25544 3538
rect 22282 2479 22338 2488
rect 25504 2508 25556 2514
rect 25504 2450 25556 2456
rect 22376 2372 22428 2378
rect 22376 2314 22428 2320
rect 21454 1456 21510 1465
rect 21454 1391 21510 1400
rect 19890 54 20024 82
rect 22282 82 22338 480
rect 22388 82 22416 2314
rect 22282 54 22416 82
rect 24582 96 24638 480
rect 19890 0 19946 54
rect 22282 0 22338 54
rect 26804 82 26832 4082
rect 26896 3194 26924 4558
rect 27448 4282 27476 5306
rect 27622 4924 27918 4944
rect 27678 4922 27702 4924
rect 27758 4922 27782 4924
rect 27838 4922 27862 4924
rect 27700 4870 27702 4922
rect 27764 4870 27776 4922
rect 27838 4870 27840 4922
rect 27678 4868 27702 4870
rect 27758 4868 27782 4870
rect 27838 4868 27862 4870
rect 27622 4848 27918 4868
rect 27436 4276 27488 4282
rect 27436 4218 27488 4224
rect 31404 4146 31432 6054
rect 39592 5953 39620 6326
rect 39578 5944 39634 5953
rect 39578 5879 39634 5888
rect 34289 5468 34585 5488
rect 34345 5466 34369 5468
rect 34425 5466 34449 5468
rect 34505 5466 34529 5468
rect 34367 5414 34369 5466
rect 34431 5414 34443 5466
rect 34505 5414 34507 5466
rect 34345 5412 34369 5414
rect 34425 5412 34449 5414
rect 34505 5412 34529 5414
rect 34289 5392 34585 5412
rect 34289 4380 34585 4400
rect 34345 4378 34369 4380
rect 34425 4378 34449 4380
rect 34505 4378 34529 4380
rect 34367 4326 34369 4378
rect 34431 4326 34443 4378
rect 34505 4326 34507 4378
rect 34345 4324 34369 4326
rect 34425 4324 34449 4326
rect 34505 4324 34529 4326
rect 34289 4304 34585 4324
rect 35530 4312 35586 4321
rect 35530 4247 35586 4256
rect 35544 4146 35572 4247
rect 36084 4208 36136 4214
rect 36084 4150 36136 4156
rect 31392 4140 31444 4146
rect 31392 4082 31444 4088
rect 31668 4140 31720 4146
rect 31668 4082 31720 4088
rect 35532 4140 35584 4146
rect 35532 4082 35584 4088
rect 31300 3936 31352 3942
rect 31300 3878 31352 3884
rect 27622 3836 27918 3856
rect 27678 3834 27702 3836
rect 27758 3834 27782 3836
rect 27838 3834 27862 3836
rect 27700 3782 27702 3834
rect 27764 3782 27776 3834
rect 27838 3782 27840 3834
rect 27678 3780 27702 3782
rect 27758 3780 27782 3782
rect 27838 3780 27862 3782
rect 27622 3760 27918 3780
rect 31312 3618 31340 3878
rect 31404 3738 31432 4082
rect 31484 4004 31536 4010
rect 31484 3946 31536 3952
rect 31392 3732 31444 3738
rect 31392 3674 31444 3680
rect 31496 3618 31524 3946
rect 31312 3590 31524 3618
rect 30840 3392 30892 3398
rect 30840 3334 30892 3340
rect 30852 3194 30880 3334
rect 31312 3194 31340 3590
rect 31680 3466 31708 4082
rect 32312 3664 32364 3670
rect 32312 3606 32364 3612
rect 32220 3528 32272 3534
rect 32220 3470 32272 3476
rect 31668 3460 31720 3466
rect 31668 3402 31720 3408
rect 26884 3188 26936 3194
rect 26884 3130 26936 3136
rect 30840 3188 30892 3194
rect 30840 3130 30892 3136
rect 31300 3188 31352 3194
rect 31300 3130 31352 3136
rect 26896 2990 26924 3130
rect 30852 2990 30880 3130
rect 26884 2984 26936 2990
rect 26884 2926 26936 2932
rect 30840 2984 30892 2990
rect 30840 2926 30892 2932
rect 29920 2848 29972 2854
rect 29920 2790 29972 2796
rect 27622 2748 27918 2768
rect 27678 2746 27702 2748
rect 27758 2746 27782 2748
rect 27838 2746 27862 2748
rect 27700 2694 27702 2746
rect 27764 2694 27776 2746
rect 27838 2694 27840 2746
rect 27678 2692 27702 2694
rect 27758 2692 27782 2694
rect 27838 2692 27862 2694
rect 27622 2672 27918 2692
rect 29932 1601 29960 2790
rect 31680 2417 31708 3402
rect 32232 3194 32260 3470
rect 32220 3188 32272 3194
rect 32220 3130 32272 3136
rect 32232 2650 32260 3130
rect 32324 2990 32352 3606
rect 34289 3292 34585 3312
rect 34345 3290 34369 3292
rect 34425 3290 34449 3292
rect 34505 3290 34529 3292
rect 34367 3238 34369 3290
rect 34431 3238 34443 3290
rect 34505 3238 34507 3290
rect 34345 3236 34369 3238
rect 34425 3236 34449 3238
rect 34505 3236 34529 3238
rect 34289 3216 34585 3236
rect 34702 3224 34758 3233
rect 34702 3159 34758 3168
rect 34716 3126 34744 3159
rect 33232 3120 33284 3126
rect 33232 3062 33284 3068
rect 34704 3120 34756 3126
rect 34704 3062 34756 3068
rect 32312 2984 32364 2990
rect 32312 2926 32364 2932
rect 33244 2650 33272 3062
rect 32220 2644 32272 2650
rect 32220 2586 32272 2592
rect 33232 2644 33284 2650
rect 33232 2586 33284 2592
rect 31666 2408 31722 2417
rect 31666 2343 31722 2352
rect 31760 2372 31812 2378
rect 31760 2314 31812 2320
rect 34152 2372 34204 2378
rect 34152 2314 34204 2320
rect 29918 1592 29974 1601
rect 29918 1527 29974 1536
rect 29090 1456 29146 1465
rect 29090 1391 29146 1400
rect 26974 82 27030 480
rect 26804 54 27030 82
rect 29104 82 29132 1391
rect 29366 82 29422 480
rect 29104 54 29422 82
rect 24582 0 24638 40
rect 26974 0 27030 54
rect 29366 0 29422 54
rect 31666 82 31722 480
rect 31772 82 31800 2314
rect 31666 54 31800 82
rect 34058 82 34114 480
rect 34164 82 34192 2314
rect 34289 2204 34585 2224
rect 34345 2202 34369 2204
rect 34425 2202 34449 2204
rect 34505 2202 34529 2204
rect 34367 2150 34369 2202
rect 34431 2150 34443 2202
rect 34505 2150 34507 2202
rect 34345 2148 34369 2150
rect 34425 2148 34449 2150
rect 34505 2148 34529 2150
rect 34289 2128 34585 2148
rect 34058 54 34192 82
rect 36096 82 36124 4150
rect 38474 2544 38530 2553
rect 38474 2479 38530 2488
rect 36358 82 36414 480
rect 36096 54 36414 82
rect 38488 82 38516 2479
rect 39394 1864 39450 1873
rect 39450 1822 39620 1850
rect 39394 1799 39450 1808
rect 39592 649 39620 1822
rect 39578 640 39634 649
rect 39578 575 39634 584
rect 38750 82 38806 480
rect 38488 54 38806 82
rect 31666 0 31722 54
rect 34058 0 34114 54
rect 36358 0 36414 54
rect 38750 0 38806 54
<< via2 >>
rect 1490 14728 1546 14784
rect 1398 9288 1454 9344
rect 1582 13640 1638 13696
rect 1858 8880 1914 8936
rect 110 7248 166 7304
rect 1030 5480 1086 5536
rect 110 3168 166 3224
rect 1858 5072 1914 5128
rect 1858 4664 1914 4720
rect 2042 5108 2044 5128
rect 2044 5108 2096 5128
rect 2096 5108 2098 5128
rect 2042 5072 2098 5108
rect 14289 13626 14345 13628
rect 14369 13626 14425 13628
rect 14449 13626 14505 13628
rect 14529 13626 14585 13628
rect 14289 13574 14315 13626
rect 14315 13574 14345 13626
rect 14369 13574 14379 13626
rect 14379 13574 14425 13626
rect 14449 13574 14495 13626
rect 14495 13574 14505 13626
rect 14529 13574 14559 13626
rect 14559 13574 14585 13626
rect 14289 13572 14345 13574
rect 14369 13572 14425 13574
rect 14449 13572 14505 13574
rect 14529 13572 14585 13574
rect 7622 13082 7678 13084
rect 7702 13082 7758 13084
rect 7782 13082 7838 13084
rect 7862 13082 7918 13084
rect 7622 13030 7648 13082
rect 7648 13030 7678 13082
rect 7702 13030 7712 13082
rect 7712 13030 7758 13082
rect 7782 13030 7828 13082
rect 7828 13030 7838 13082
rect 7862 13030 7892 13082
rect 7892 13030 7918 13082
rect 7622 13028 7678 13030
rect 7702 13028 7758 13030
rect 7782 13028 7838 13030
rect 7862 13028 7918 13030
rect 14289 12538 14345 12540
rect 14369 12538 14425 12540
rect 14449 12538 14505 12540
rect 14529 12538 14585 12540
rect 14289 12486 14315 12538
rect 14315 12486 14345 12538
rect 14369 12486 14379 12538
rect 14379 12486 14425 12538
rect 14449 12486 14495 12538
rect 14495 12486 14505 12538
rect 14529 12486 14559 12538
rect 14559 12486 14585 12538
rect 14289 12484 14345 12486
rect 14369 12484 14425 12486
rect 14449 12484 14505 12486
rect 14529 12484 14585 12486
rect 7010 12008 7066 12064
rect 7622 11994 7678 11996
rect 7702 11994 7758 11996
rect 7782 11994 7838 11996
rect 7862 11994 7918 11996
rect 7622 11942 7648 11994
rect 7648 11942 7678 11994
rect 7702 11942 7712 11994
rect 7712 11942 7758 11994
rect 7782 11942 7828 11994
rect 7828 11942 7838 11994
rect 7862 11942 7892 11994
rect 7892 11942 7918 11994
rect 7622 11940 7678 11942
rect 7702 11940 7758 11942
rect 7782 11940 7838 11942
rect 7862 11940 7918 11942
rect 4342 4528 4398 4584
rect 2962 1672 3018 1728
rect 1398 1128 1454 1184
rect 4526 4120 4582 4176
rect 14289 11450 14345 11452
rect 14369 11450 14425 11452
rect 14449 11450 14505 11452
rect 14529 11450 14585 11452
rect 14289 11398 14315 11450
rect 14315 11398 14345 11450
rect 14369 11398 14379 11450
rect 14379 11398 14425 11450
rect 14449 11398 14495 11450
rect 14495 11398 14505 11450
rect 14529 11398 14559 11450
rect 14559 11398 14585 11450
rect 14289 11396 14345 11398
rect 14369 11396 14425 11398
rect 14449 11396 14505 11398
rect 14529 11396 14585 11398
rect 11150 11056 11206 11112
rect 7622 10906 7678 10908
rect 7702 10906 7758 10908
rect 7782 10906 7838 10908
rect 7862 10906 7918 10908
rect 7622 10854 7648 10906
rect 7648 10854 7678 10906
rect 7702 10854 7712 10906
rect 7712 10854 7758 10906
rect 7782 10854 7828 10906
rect 7828 10854 7838 10906
rect 7862 10854 7892 10906
rect 7892 10854 7918 10906
rect 7622 10852 7678 10854
rect 7702 10852 7758 10854
rect 7782 10852 7838 10854
rect 7862 10852 7918 10854
rect 7622 9818 7678 9820
rect 7702 9818 7758 9820
rect 7782 9818 7838 9820
rect 7862 9818 7918 9820
rect 7622 9766 7648 9818
rect 7648 9766 7678 9818
rect 7702 9766 7712 9818
rect 7712 9766 7758 9818
rect 7782 9766 7828 9818
rect 7828 9766 7838 9818
rect 7862 9766 7892 9818
rect 7892 9766 7918 9818
rect 7622 9764 7678 9766
rect 7702 9764 7758 9766
rect 7782 9764 7838 9766
rect 7862 9764 7918 9766
rect 7622 8730 7678 8732
rect 7702 8730 7758 8732
rect 7782 8730 7838 8732
rect 7862 8730 7918 8732
rect 7622 8678 7648 8730
rect 7648 8678 7678 8730
rect 7702 8678 7712 8730
rect 7712 8678 7758 8730
rect 7782 8678 7828 8730
rect 7828 8678 7838 8730
rect 7862 8678 7892 8730
rect 7892 8678 7918 8730
rect 7622 8676 7678 8678
rect 7702 8676 7758 8678
rect 7782 8676 7838 8678
rect 7862 8676 7918 8678
rect 15474 10648 15530 10704
rect 14289 10362 14345 10364
rect 14369 10362 14425 10364
rect 14449 10362 14505 10364
rect 14529 10362 14585 10364
rect 14289 10310 14315 10362
rect 14315 10310 14345 10362
rect 14369 10310 14379 10362
rect 14379 10310 14425 10362
rect 14449 10310 14495 10362
rect 14495 10310 14505 10362
rect 14529 10310 14559 10362
rect 14559 10310 14585 10362
rect 14289 10308 14345 10310
rect 14369 10308 14425 10310
rect 14449 10308 14505 10310
rect 14529 10308 14585 10310
rect 14289 9274 14345 9276
rect 14369 9274 14425 9276
rect 14449 9274 14505 9276
rect 14529 9274 14585 9276
rect 14289 9222 14315 9274
rect 14315 9222 14345 9274
rect 14369 9222 14379 9274
rect 14379 9222 14425 9274
rect 14449 9222 14495 9274
rect 14495 9222 14505 9274
rect 14529 9222 14559 9274
rect 14559 9222 14585 9274
rect 14289 9220 14345 9222
rect 14369 9220 14425 9222
rect 14449 9220 14505 9222
rect 14529 9220 14585 9222
rect 7622 7642 7678 7644
rect 7702 7642 7758 7644
rect 7782 7642 7838 7644
rect 7862 7642 7918 7644
rect 7622 7590 7648 7642
rect 7648 7590 7678 7642
rect 7702 7590 7712 7642
rect 7712 7590 7758 7642
rect 7782 7590 7828 7642
rect 7828 7590 7838 7642
rect 7862 7590 7892 7642
rect 7892 7590 7918 7642
rect 7622 7588 7678 7590
rect 7702 7588 7758 7590
rect 7782 7588 7838 7590
rect 7862 7588 7918 7590
rect 7622 6554 7678 6556
rect 7702 6554 7758 6556
rect 7782 6554 7838 6556
rect 7862 6554 7918 6556
rect 7622 6502 7648 6554
rect 7648 6502 7678 6554
rect 7702 6502 7712 6554
rect 7712 6502 7758 6554
rect 7782 6502 7828 6554
rect 7828 6502 7838 6554
rect 7862 6502 7892 6554
rect 7892 6502 7918 6554
rect 7622 6500 7678 6502
rect 7702 6500 7758 6502
rect 7782 6500 7838 6502
rect 7862 6500 7918 6502
rect 7286 5752 7342 5808
rect 7622 5466 7678 5468
rect 7702 5466 7758 5468
rect 7782 5466 7838 5468
rect 7862 5466 7918 5468
rect 7622 5414 7648 5466
rect 7648 5414 7678 5466
rect 7702 5414 7712 5466
rect 7712 5414 7758 5466
rect 7782 5414 7828 5466
rect 7828 5414 7838 5466
rect 7862 5414 7892 5466
rect 7892 5414 7918 5466
rect 7622 5412 7678 5414
rect 7702 5412 7758 5414
rect 7782 5412 7838 5414
rect 7862 5412 7918 5414
rect 7194 4664 7250 4720
rect 6734 3732 6790 3768
rect 6734 3712 6736 3732
rect 6736 3712 6788 3732
rect 6788 3712 6790 3732
rect 7194 3712 7250 3768
rect 7622 4378 7678 4380
rect 7702 4378 7758 4380
rect 7782 4378 7838 4380
rect 7862 4378 7918 4380
rect 7622 4326 7648 4378
rect 7648 4326 7678 4378
rect 7702 4326 7712 4378
rect 7712 4326 7758 4378
rect 7782 4326 7828 4378
rect 7828 4326 7838 4378
rect 7862 4326 7892 4378
rect 7892 4326 7918 4378
rect 7622 4324 7678 4326
rect 7702 4324 7758 4326
rect 7782 4324 7838 4326
rect 7862 4324 7918 4326
rect 7746 3984 7802 4040
rect 7622 3290 7678 3292
rect 7702 3290 7758 3292
rect 7782 3290 7838 3292
rect 7862 3290 7918 3292
rect 7622 3238 7648 3290
rect 7648 3238 7678 3290
rect 7702 3238 7712 3290
rect 7712 3238 7758 3290
rect 7782 3238 7828 3290
rect 7828 3238 7838 3290
rect 7862 3238 7892 3290
rect 7892 3238 7918 3290
rect 7622 3236 7678 3238
rect 7702 3236 7758 3238
rect 7782 3236 7838 3238
rect 7862 3236 7918 3238
rect 7470 2352 7526 2408
rect 8482 3848 8538 3904
rect 9034 3848 9090 3904
rect 11058 8336 11114 8392
rect 12898 8880 12954 8936
rect 9218 4120 9274 4176
rect 9862 4936 9918 4992
rect 10046 4120 10102 4176
rect 8666 2488 8722 2544
rect 7622 2202 7678 2204
rect 7702 2202 7758 2204
rect 7782 2202 7838 2204
rect 7862 2202 7918 2204
rect 7622 2150 7648 2202
rect 7648 2150 7678 2202
rect 7702 2150 7712 2202
rect 7712 2150 7758 2202
rect 7782 2150 7828 2202
rect 7828 2150 7838 2202
rect 7862 2150 7892 2202
rect 7892 2150 7918 2202
rect 7622 2148 7678 2150
rect 7702 2148 7758 2150
rect 7782 2148 7838 2150
rect 7862 2148 7918 2150
rect 10598 3712 10654 3768
rect 11242 4120 11298 4176
rect 11518 4392 11574 4448
rect 11334 3712 11390 3768
rect 12254 6160 12310 6216
rect 11794 4664 11850 4720
rect 11978 3848 12034 3904
rect 11886 3304 11942 3360
rect 11702 2352 11758 2408
rect 10966 2080 11022 2136
rect 14289 8186 14345 8188
rect 14369 8186 14425 8188
rect 14449 8186 14505 8188
rect 14529 8186 14585 8188
rect 14289 8134 14315 8186
rect 14315 8134 14345 8186
rect 14369 8134 14379 8186
rect 14379 8134 14425 8186
rect 14449 8134 14495 8186
rect 14495 8134 14505 8186
rect 14529 8134 14559 8186
rect 14559 8134 14585 8186
rect 14289 8132 14345 8134
rect 14369 8132 14425 8134
rect 14449 8132 14505 8134
rect 14529 8132 14585 8134
rect 13910 7384 13966 7440
rect 12714 3984 12770 4040
rect 12622 3440 12678 3496
rect 12530 3168 12586 3224
rect 12990 3984 13046 4040
rect 14289 7098 14345 7100
rect 14369 7098 14425 7100
rect 14449 7098 14505 7100
rect 14529 7098 14585 7100
rect 14289 7046 14315 7098
rect 14315 7046 14345 7098
rect 14369 7046 14379 7098
rect 14379 7046 14425 7098
rect 14449 7046 14495 7098
rect 14495 7046 14505 7098
rect 14529 7046 14559 7098
rect 14559 7046 14585 7098
rect 14289 7044 14345 7046
rect 14369 7044 14425 7046
rect 14449 7044 14505 7046
rect 14529 7044 14585 7046
rect 14289 6010 14345 6012
rect 14369 6010 14425 6012
rect 14449 6010 14505 6012
rect 14529 6010 14585 6012
rect 14289 5958 14315 6010
rect 14315 5958 14345 6010
rect 14369 5958 14379 6010
rect 14379 5958 14425 6010
rect 14449 5958 14495 6010
rect 14495 5958 14505 6010
rect 14529 5958 14559 6010
rect 14559 5958 14585 6010
rect 14289 5956 14345 5958
rect 14369 5956 14425 5958
rect 14449 5956 14505 5958
rect 14529 5956 14585 5958
rect 14094 4936 14150 4992
rect 14289 4922 14345 4924
rect 14369 4922 14425 4924
rect 14449 4922 14505 4924
rect 14529 4922 14585 4924
rect 14289 4870 14315 4922
rect 14315 4870 14345 4922
rect 14369 4870 14379 4922
rect 14379 4870 14425 4922
rect 14449 4870 14495 4922
rect 14495 4870 14505 4922
rect 14529 4870 14559 4922
rect 14559 4870 14585 4922
rect 14289 4868 14345 4870
rect 14369 4868 14425 4870
rect 14449 4868 14505 4870
rect 14529 4868 14585 4870
rect 14289 3834 14345 3836
rect 14369 3834 14425 3836
rect 14449 3834 14505 3836
rect 14529 3834 14585 3836
rect 14289 3782 14315 3834
rect 14315 3782 14345 3834
rect 14369 3782 14379 3834
rect 14379 3782 14425 3834
rect 14449 3782 14495 3834
rect 14495 3782 14505 3834
rect 14529 3782 14559 3834
rect 14559 3782 14585 3834
rect 14289 3780 14345 3782
rect 14369 3780 14425 3782
rect 14449 3780 14505 3782
rect 14529 3780 14585 3782
rect 14554 3576 14610 3632
rect 14738 5072 14794 5128
rect 15106 7384 15162 7440
rect 14830 3984 14886 4040
rect 14289 2746 14345 2748
rect 14369 2746 14425 2748
rect 14449 2746 14505 2748
rect 14529 2746 14585 2748
rect 14289 2694 14315 2746
rect 14315 2694 14345 2746
rect 14369 2694 14379 2746
rect 14379 2694 14425 2746
rect 14449 2694 14495 2746
rect 14495 2694 14505 2746
rect 14529 2694 14559 2746
rect 14559 2694 14585 2746
rect 14289 2692 14345 2694
rect 14369 2692 14425 2694
rect 14449 2692 14505 2694
rect 14529 2692 14585 2694
rect 20956 13082 21012 13084
rect 21036 13082 21092 13084
rect 21116 13082 21172 13084
rect 21196 13082 21252 13084
rect 20956 13030 20982 13082
rect 20982 13030 21012 13082
rect 21036 13030 21046 13082
rect 21046 13030 21092 13082
rect 21116 13030 21162 13082
rect 21162 13030 21172 13082
rect 21196 13030 21226 13082
rect 21226 13030 21252 13082
rect 20956 13028 21012 13030
rect 21036 13028 21092 13030
rect 21116 13028 21172 13030
rect 21196 13028 21252 13030
rect 27622 13626 27678 13628
rect 27702 13626 27758 13628
rect 27782 13626 27838 13628
rect 27862 13626 27918 13628
rect 27622 13574 27648 13626
rect 27648 13574 27678 13626
rect 27702 13574 27712 13626
rect 27712 13574 27758 13626
rect 27782 13574 27828 13626
rect 27828 13574 27838 13626
rect 27862 13574 27892 13626
rect 27892 13574 27918 13626
rect 27622 13572 27678 13574
rect 27702 13572 27758 13574
rect 27782 13572 27838 13574
rect 27862 13572 27918 13574
rect 20956 11994 21012 11996
rect 21036 11994 21092 11996
rect 21116 11994 21172 11996
rect 21196 11994 21252 11996
rect 20956 11942 20982 11994
rect 20982 11942 21012 11994
rect 21036 11942 21046 11994
rect 21046 11942 21092 11994
rect 21116 11942 21162 11994
rect 21162 11942 21172 11994
rect 21196 11942 21226 11994
rect 21226 11942 21252 11994
rect 20956 11940 21012 11942
rect 21036 11940 21092 11942
rect 21116 11940 21172 11942
rect 21196 11940 21252 11942
rect 24306 11600 24362 11656
rect 20956 10906 21012 10908
rect 21036 10906 21092 10908
rect 21116 10906 21172 10908
rect 21196 10906 21252 10908
rect 20956 10854 20982 10906
rect 20982 10854 21012 10906
rect 21036 10854 21046 10906
rect 21046 10854 21092 10906
rect 21116 10854 21162 10906
rect 21162 10854 21172 10906
rect 21196 10854 21226 10906
rect 21226 10854 21252 10906
rect 20956 10852 21012 10854
rect 21036 10852 21092 10854
rect 21116 10852 21172 10854
rect 21196 10852 21252 10854
rect 20956 9818 21012 9820
rect 21036 9818 21092 9820
rect 21116 9818 21172 9820
rect 21196 9818 21252 9820
rect 20956 9766 20982 9818
rect 20982 9766 21012 9818
rect 21036 9766 21046 9818
rect 21046 9766 21092 9818
rect 21116 9766 21162 9818
rect 21162 9766 21172 9818
rect 21196 9766 21226 9818
rect 21226 9766 21252 9818
rect 20956 9764 21012 9766
rect 21036 9764 21092 9766
rect 21116 9764 21172 9766
rect 21196 9764 21252 9766
rect 20956 8730 21012 8732
rect 21036 8730 21092 8732
rect 21116 8730 21172 8732
rect 21196 8730 21252 8732
rect 20956 8678 20982 8730
rect 20982 8678 21012 8730
rect 21036 8678 21046 8730
rect 21046 8678 21092 8730
rect 21116 8678 21162 8730
rect 21162 8678 21172 8730
rect 21196 8678 21226 8730
rect 21226 8678 21252 8730
rect 20956 8676 21012 8678
rect 21036 8676 21092 8678
rect 21116 8676 21172 8678
rect 21196 8676 21252 8678
rect 24674 10512 24730 10568
rect 20956 7642 21012 7644
rect 21036 7642 21092 7644
rect 21116 7642 21172 7644
rect 21196 7642 21252 7644
rect 20956 7590 20982 7642
rect 20982 7590 21012 7642
rect 21036 7590 21046 7642
rect 21046 7590 21092 7642
rect 21116 7590 21162 7642
rect 21162 7590 21172 7642
rect 21196 7590 21226 7642
rect 21226 7590 21252 7642
rect 20956 7588 21012 7590
rect 21036 7588 21092 7590
rect 21116 7588 21172 7590
rect 21196 7588 21252 7590
rect 15566 4392 15622 4448
rect 15658 3440 15714 3496
rect 15842 3340 15844 3360
rect 15844 3340 15896 3360
rect 15896 3340 15898 3360
rect 15842 3304 15898 3340
rect 16486 4664 16542 4720
rect 17038 4528 17094 4584
rect 16854 2488 16910 2544
rect 17682 3984 17738 4040
rect 20956 6554 21012 6556
rect 21036 6554 21092 6556
rect 21116 6554 21172 6556
rect 21196 6554 21252 6556
rect 20956 6502 20982 6554
rect 20982 6502 21012 6554
rect 21036 6502 21046 6554
rect 21046 6502 21092 6554
rect 21116 6502 21162 6554
rect 21162 6502 21172 6554
rect 21196 6502 21226 6554
rect 21226 6502 21252 6554
rect 20956 6500 21012 6502
rect 21036 6500 21092 6502
rect 21116 6500 21172 6502
rect 21196 6500 21252 6502
rect 18878 3984 18934 4040
rect 20956 5466 21012 5468
rect 21036 5466 21092 5468
rect 21116 5466 21172 5468
rect 21196 5466 21252 5468
rect 20956 5414 20982 5466
rect 20982 5414 21012 5466
rect 21036 5414 21046 5466
rect 21046 5414 21092 5466
rect 21116 5414 21162 5466
rect 21162 5414 21172 5466
rect 21196 5414 21226 5466
rect 21226 5414 21252 5466
rect 20956 5412 21012 5414
rect 21036 5412 21092 5414
rect 21116 5412 21172 5414
rect 21196 5412 21252 5414
rect 20956 4378 21012 4380
rect 21036 4378 21092 4380
rect 21116 4378 21172 4380
rect 21196 4378 21252 4380
rect 20956 4326 20982 4378
rect 20982 4326 21012 4378
rect 21036 4326 21046 4378
rect 21046 4326 21092 4378
rect 21116 4326 21162 4378
rect 21162 4326 21172 4378
rect 21196 4326 21226 4378
rect 21226 4326 21252 4378
rect 20956 4324 21012 4326
rect 21036 4324 21092 4326
rect 21116 4324 21172 4326
rect 21196 4324 21252 4326
rect 23294 5752 23350 5808
rect 19338 3168 19394 3224
rect 18326 1808 18382 1864
rect 21730 3984 21786 4040
rect 20442 3576 20498 3632
rect 20994 3440 21050 3496
rect 20956 3290 21012 3292
rect 21036 3290 21092 3292
rect 21116 3290 21172 3292
rect 21196 3290 21252 3292
rect 20956 3238 20982 3290
rect 20982 3238 21012 3290
rect 21036 3238 21046 3290
rect 21046 3238 21092 3290
rect 21116 3238 21162 3290
rect 21162 3238 21172 3290
rect 21196 3238 21226 3290
rect 21226 3238 21252 3290
rect 20956 3236 21012 3238
rect 21036 3236 21092 3238
rect 21116 3236 21172 3238
rect 21196 3236 21252 3238
rect 23478 3440 23534 3496
rect 27622 12538 27678 12540
rect 27702 12538 27758 12540
rect 27782 12538 27838 12540
rect 27862 12538 27918 12540
rect 27622 12486 27648 12538
rect 27648 12486 27678 12538
rect 27702 12486 27712 12538
rect 27712 12486 27758 12538
rect 27782 12486 27828 12538
rect 27828 12486 27838 12538
rect 27862 12486 27892 12538
rect 27892 12486 27918 12538
rect 27622 12484 27678 12486
rect 27702 12484 27758 12486
rect 27782 12484 27838 12486
rect 27862 12484 27918 12486
rect 27622 11450 27678 11452
rect 27702 11450 27758 11452
rect 27782 11450 27838 11452
rect 27862 11450 27918 11452
rect 27622 11398 27648 11450
rect 27648 11398 27678 11450
rect 27702 11398 27712 11450
rect 27712 11398 27758 11450
rect 27782 11398 27828 11450
rect 27828 11398 27838 11450
rect 27862 11398 27892 11450
rect 27892 11398 27918 11450
rect 27622 11396 27678 11398
rect 27702 11396 27758 11398
rect 27782 11396 27838 11398
rect 27862 11396 27918 11398
rect 27622 10362 27678 10364
rect 27702 10362 27758 10364
rect 27782 10362 27838 10364
rect 27862 10362 27918 10364
rect 27622 10310 27648 10362
rect 27648 10310 27678 10362
rect 27702 10310 27712 10362
rect 27712 10310 27758 10362
rect 27782 10310 27828 10362
rect 27828 10310 27838 10362
rect 27862 10310 27892 10362
rect 27892 10310 27918 10362
rect 27622 10308 27678 10310
rect 27702 10308 27758 10310
rect 27782 10308 27838 10310
rect 27862 10308 27918 10310
rect 27622 9274 27678 9276
rect 27702 9274 27758 9276
rect 27782 9274 27838 9276
rect 27862 9274 27918 9276
rect 27622 9222 27648 9274
rect 27648 9222 27678 9274
rect 27702 9222 27712 9274
rect 27712 9222 27758 9274
rect 27782 9222 27828 9274
rect 27828 9222 27838 9274
rect 27862 9222 27892 9274
rect 27892 9222 27918 9274
rect 27622 9220 27678 9222
rect 27702 9220 27758 9222
rect 27782 9220 27838 9222
rect 27862 9220 27918 9222
rect 27622 8186 27678 8188
rect 27702 8186 27758 8188
rect 27782 8186 27838 8188
rect 27862 8186 27918 8188
rect 27622 8134 27648 8186
rect 27648 8134 27678 8186
rect 27702 8134 27712 8186
rect 27712 8134 27758 8186
rect 27782 8134 27828 8186
rect 27828 8134 27838 8186
rect 27862 8134 27892 8186
rect 27892 8134 27918 8186
rect 27622 8132 27678 8134
rect 27702 8132 27758 8134
rect 27782 8132 27838 8134
rect 27862 8132 27918 8134
rect 35622 13640 35678 13696
rect 34289 13082 34345 13084
rect 34369 13082 34425 13084
rect 34449 13082 34505 13084
rect 34529 13082 34585 13084
rect 34289 13030 34315 13082
rect 34315 13030 34345 13082
rect 34369 13030 34379 13082
rect 34379 13030 34425 13082
rect 34449 13030 34495 13082
rect 34495 13030 34505 13082
rect 34529 13030 34559 13082
rect 34559 13030 34585 13082
rect 34289 13028 34345 13030
rect 34369 13028 34425 13030
rect 34449 13028 34505 13030
rect 34529 13028 34585 13030
rect 34289 11994 34345 11996
rect 34369 11994 34425 11996
rect 34449 11994 34505 11996
rect 34529 11994 34585 11996
rect 34289 11942 34315 11994
rect 34315 11942 34345 11994
rect 34369 11942 34379 11994
rect 34379 11942 34425 11994
rect 34449 11942 34495 11994
rect 34495 11942 34505 11994
rect 34529 11942 34559 11994
rect 34559 11942 34585 11994
rect 34289 11940 34345 11942
rect 34369 11940 34425 11942
rect 34449 11940 34505 11942
rect 34529 11940 34585 11942
rect 34289 10906 34345 10908
rect 34369 10906 34425 10908
rect 34449 10906 34505 10908
rect 34529 10906 34585 10908
rect 34289 10854 34315 10906
rect 34315 10854 34345 10906
rect 34369 10854 34379 10906
rect 34379 10854 34425 10906
rect 34449 10854 34495 10906
rect 34495 10854 34505 10906
rect 34529 10854 34559 10906
rect 34559 10854 34585 10906
rect 34289 10852 34345 10854
rect 34369 10852 34425 10854
rect 34449 10852 34505 10854
rect 34529 10852 34585 10854
rect 34289 9818 34345 9820
rect 34369 9818 34425 9820
rect 34449 9818 34505 9820
rect 34529 9818 34585 9820
rect 34289 9766 34315 9818
rect 34315 9766 34345 9818
rect 34369 9766 34379 9818
rect 34379 9766 34425 9818
rect 34449 9766 34495 9818
rect 34495 9766 34505 9818
rect 34529 9766 34559 9818
rect 34559 9766 34585 9818
rect 34289 9764 34345 9766
rect 34369 9764 34425 9766
rect 34449 9764 34505 9766
rect 34529 9764 34585 9766
rect 34289 8730 34345 8732
rect 34369 8730 34425 8732
rect 34449 8730 34505 8732
rect 34529 8730 34585 8732
rect 34289 8678 34315 8730
rect 34315 8678 34345 8730
rect 34369 8678 34379 8730
rect 34379 8678 34425 8730
rect 34449 8678 34495 8730
rect 34495 8678 34505 8730
rect 34529 8678 34559 8730
rect 34559 8678 34585 8730
rect 34289 8676 34345 8678
rect 34369 8676 34425 8678
rect 34449 8676 34505 8678
rect 34529 8676 34585 8678
rect 34289 7642 34345 7644
rect 34369 7642 34425 7644
rect 34449 7642 34505 7644
rect 34529 7642 34585 7644
rect 34289 7590 34315 7642
rect 34315 7590 34345 7642
rect 34369 7590 34379 7642
rect 34379 7590 34425 7642
rect 34449 7590 34495 7642
rect 34495 7590 34505 7642
rect 34529 7590 34559 7642
rect 34559 7590 34585 7642
rect 34289 7588 34345 7590
rect 34369 7588 34425 7590
rect 34449 7588 34505 7590
rect 34529 7588 34585 7590
rect 39578 15272 39634 15328
rect 39578 12552 39634 12608
rect 37830 11600 37886 11656
rect 39578 11192 39634 11248
rect 35438 10512 35494 10568
rect 35622 9288 35678 9344
rect 35254 7384 35310 7440
rect 32218 7248 32274 7304
rect 27622 7098 27678 7100
rect 27702 7098 27758 7100
rect 27782 7098 27838 7100
rect 27862 7098 27918 7100
rect 27622 7046 27648 7098
rect 27648 7046 27678 7098
rect 27702 7046 27712 7098
rect 27712 7046 27758 7098
rect 27782 7046 27828 7098
rect 27828 7046 27838 7098
rect 27862 7046 27892 7098
rect 27892 7046 27918 7098
rect 27622 7044 27678 7046
rect 27702 7044 27758 7046
rect 27782 7044 27838 7046
rect 27862 7044 27918 7046
rect 34289 6554 34345 6556
rect 34369 6554 34425 6556
rect 34449 6554 34505 6556
rect 34529 6554 34585 6556
rect 34289 6502 34315 6554
rect 34315 6502 34345 6554
rect 34369 6502 34379 6554
rect 34379 6502 34425 6554
rect 34449 6502 34495 6554
rect 34495 6502 34505 6554
rect 34529 6502 34559 6554
rect 34559 6502 34585 6554
rect 34289 6500 34345 6502
rect 34369 6500 34425 6502
rect 34449 6500 34505 6502
rect 34529 6500 34585 6502
rect 27622 6010 27678 6012
rect 27702 6010 27758 6012
rect 27782 6010 27838 6012
rect 27862 6010 27918 6012
rect 27622 5958 27648 6010
rect 27648 5958 27678 6010
rect 27702 5958 27712 6010
rect 27712 5958 27758 6010
rect 27782 5958 27828 6010
rect 27828 5958 27838 6010
rect 27862 5958 27892 6010
rect 27892 5958 27918 6010
rect 27622 5956 27678 5958
rect 27702 5956 27758 5958
rect 27782 5956 27838 5958
rect 27862 5956 27918 5958
rect 36082 8064 36138 8120
rect 35438 6160 35494 6216
rect 21270 2352 21326 2408
rect 20956 2202 21012 2204
rect 21036 2202 21092 2204
rect 21116 2202 21172 2204
rect 21196 2202 21252 2204
rect 20956 2150 20982 2202
rect 20982 2150 21012 2202
rect 21036 2150 21046 2202
rect 21046 2150 21092 2202
rect 21116 2150 21162 2202
rect 21162 2150 21172 2202
rect 21196 2150 21226 2202
rect 21226 2150 21252 2202
rect 20956 2148 21012 2150
rect 21036 2148 21092 2150
rect 21116 2148 21172 2150
rect 21196 2148 21252 2150
rect 20074 2080 20130 2136
rect 22282 2488 22338 2544
rect 21454 1400 21510 1456
rect 24582 40 24638 96
rect 27622 4922 27678 4924
rect 27702 4922 27758 4924
rect 27782 4922 27838 4924
rect 27862 4922 27918 4924
rect 27622 4870 27648 4922
rect 27648 4870 27678 4922
rect 27702 4870 27712 4922
rect 27712 4870 27758 4922
rect 27782 4870 27828 4922
rect 27828 4870 27838 4922
rect 27862 4870 27892 4922
rect 27892 4870 27918 4922
rect 27622 4868 27678 4870
rect 27702 4868 27758 4870
rect 27782 4868 27838 4870
rect 27862 4868 27918 4870
rect 39578 5888 39634 5944
rect 34289 5466 34345 5468
rect 34369 5466 34425 5468
rect 34449 5466 34505 5468
rect 34529 5466 34585 5468
rect 34289 5414 34315 5466
rect 34315 5414 34345 5466
rect 34369 5414 34379 5466
rect 34379 5414 34425 5466
rect 34449 5414 34495 5466
rect 34495 5414 34505 5466
rect 34529 5414 34559 5466
rect 34559 5414 34585 5466
rect 34289 5412 34345 5414
rect 34369 5412 34425 5414
rect 34449 5412 34505 5414
rect 34529 5412 34585 5414
rect 34289 4378 34345 4380
rect 34369 4378 34425 4380
rect 34449 4378 34505 4380
rect 34529 4378 34585 4380
rect 34289 4326 34315 4378
rect 34315 4326 34345 4378
rect 34369 4326 34379 4378
rect 34379 4326 34425 4378
rect 34449 4326 34495 4378
rect 34495 4326 34505 4378
rect 34529 4326 34559 4378
rect 34559 4326 34585 4378
rect 34289 4324 34345 4326
rect 34369 4324 34425 4326
rect 34449 4324 34505 4326
rect 34529 4324 34585 4326
rect 35530 4256 35586 4312
rect 27622 3834 27678 3836
rect 27702 3834 27758 3836
rect 27782 3834 27838 3836
rect 27862 3834 27918 3836
rect 27622 3782 27648 3834
rect 27648 3782 27678 3834
rect 27702 3782 27712 3834
rect 27712 3782 27758 3834
rect 27782 3782 27828 3834
rect 27828 3782 27838 3834
rect 27862 3782 27892 3834
rect 27892 3782 27918 3834
rect 27622 3780 27678 3782
rect 27702 3780 27758 3782
rect 27782 3780 27838 3782
rect 27862 3780 27918 3782
rect 27622 2746 27678 2748
rect 27702 2746 27758 2748
rect 27782 2746 27838 2748
rect 27862 2746 27918 2748
rect 27622 2694 27648 2746
rect 27648 2694 27678 2746
rect 27702 2694 27712 2746
rect 27712 2694 27758 2746
rect 27782 2694 27828 2746
rect 27828 2694 27838 2746
rect 27862 2694 27892 2746
rect 27892 2694 27918 2746
rect 27622 2692 27678 2694
rect 27702 2692 27758 2694
rect 27782 2692 27838 2694
rect 27862 2692 27918 2694
rect 34289 3290 34345 3292
rect 34369 3290 34425 3292
rect 34449 3290 34505 3292
rect 34529 3290 34585 3292
rect 34289 3238 34315 3290
rect 34315 3238 34345 3290
rect 34369 3238 34379 3290
rect 34379 3238 34425 3290
rect 34449 3238 34495 3290
rect 34495 3238 34505 3290
rect 34529 3238 34559 3290
rect 34559 3238 34585 3290
rect 34289 3236 34345 3238
rect 34369 3236 34425 3238
rect 34449 3236 34505 3238
rect 34529 3236 34585 3238
rect 34702 3168 34758 3224
rect 31666 2352 31722 2408
rect 29918 1536 29974 1592
rect 29090 1400 29146 1456
rect 34289 2202 34345 2204
rect 34369 2202 34425 2204
rect 34449 2202 34505 2204
rect 34529 2202 34585 2204
rect 34289 2150 34315 2202
rect 34315 2150 34345 2202
rect 34369 2150 34379 2202
rect 34379 2150 34425 2202
rect 34449 2150 34495 2202
rect 34495 2150 34505 2202
rect 34529 2150 34559 2202
rect 34559 2150 34585 2202
rect 34289 2148 34345 2150
rect 34369 2148 34425 2150
rect 34449 2148 34505 2150
rect 34529 2148 34585 2150
rect 38474 2488 38530 2544
rect 39394 1808 39450 1864
rect 39578 584 39634 640
<< metal3 >>
rect 0 15240 480 15360
rect 39520 15330 40000 15360
rect 39492 15328 40000 15330
rect 39492 15272 39578 15328
rect 39634 15272 40000 15328
rect 39492 15270 40000 15272
rect 39520 15240 40000 15270
rect 62 14786 122 15240
rect 1485 14786 1551 14789
rect 62 14784 1551 14786
rect 62 14728 1490 14784
rect 1546 14728 1551 14784
rect 62 14726 1551 14728
rect 1485 14723 1551 14726
rect 0 13880 480 14000
rect 39520 13880 40000 14000
rect 62 13698 122 13880
rect 1577 13698 1643 13701
rect 62 13696 1643 13698
rect 62 13640 1582 13696
rect 1638 13640 1643 13696
rect 62 13638 1643 13640
rect 1577 13635 1643 13638
rect 35617 13698 35683 13701
rect 39622 13698 39682 13880
rect 35617 13696 39682 13698
rect 35617 13640 35622 13696
rect 35678 13640 39682 13696
rect 35617 13638 39682 13640
rect 35617 13635 35683 13638
rect 14277 13632 14597 13633
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 13567 14597 13568
rect 27610 13632 27930 13633
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 13567 27930 13568
rect 7610 13088 7930 13089
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7930 13088
rect 7610 13023 7930 13024
rect 20944 13088 21264 13089
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 13023 21264 13024
rect 34277 13088 34597 13089
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 34277 13023 34597 13024
rect 0 12520 480 12640
rect 39520 12610 40000 12640
rect 39492 12608 40000 12610
rect 39492 12552 39578 12608
rect 39634 12552 40000 12608
rect 39492 12550 40000 12552
rect 14277 12544 14597 12545
rect 62 12066 122 12520
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 12479 14597 12480
rect 27610 12544 27930 12545
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 39520 12520 40000 12550
rect 27610 12479 27930 12480
rect 7005 12066 7071 12069
rect 62 12064 7071 12066
rect 62 12008 7010 12064
rect 7066 12008 7071 12064
rect 62 12006 7071 12008
rect 7005 12003 7071 12006
rect 7610 12000 7930 12001
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7930 12000
rect 7610 11935 7930 11936
rect 20944 12000 21264 12001
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 11935 21264 11936
rect 34277 12000 34597 12001
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 34277 11935 34597 11936
rect 24301 11658 24367 11661
rect 37825 11658 37891 11661
rect 24301 11656 37891 11658
rect 24301 11600 24306 11656
rect 24362 11600 37830 11656
rect 37886 11600 37891 11656
rect 24301 11598 37891 11600
rect 24301 11595 24367 11598
rect 37825 11595 37891 11598
rect 14277 11456 14597 11457
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 11391 14597 11392
rect 27610 11456 27930 11457
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 27610 11391 27930 11392
rect 0 11252 480 11280
rect 0 11188 60 11252
rect 124 11188 480 11252
rect 39520 11250 40000 11280
rect 39492 11248 40000 11250
rect 39492 11192 39578 11248
rect 39634 11192 40000 11248
rect 39492 11190 40000 11192
rect 0 11160 480 11188
rect 39520 11160 40000 11190
rect 11145 11114 11211 11117
rect 614 11112 11211 11114
rect 614 11056 11150 11112
rect 11206 11056 11211 11112
rect 614 11054 11211 11056
rect 54 10916 60 10980
rect 124 10978 130 10980
rect 614 10978 674 11054
rect 11145 11051 11211 11054
rect 124 10918 674 10978
rect 124 10916 130 10918
rect 7610 10912 7930 10913
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7930 10912
rect 7610 10847 7930 10848
rect 20944 10912 21264 10913
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 10847 21264 10848
rect 34277 10912 34597 10913
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 34277 10847 34597 10848
rect 15469 10706 15535 10709
rect 15469 10704 23490 10706
rect 15469 10648 15474 10704
rect 15530 10648 23490 10704
rect 15469 10646 23490 10648
rect 15469 10643 15535 10646
rect 23430 10570 23490 10646
rect 24669 10570 24735 10573
rect 35433 10570 35499 10573
rect 23430 10568 35499 10570
rect 23430 10512 24674 10568
rect 24730 10512 35438 10568
rect 35494 10512 35499 10568
rect 23430 10510 35499 10512
rect 24669 10507 24735 10510
rect 35433 10507 35499 10510
rect 14277 10368 14597 10369
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 10303 14597 10304
rect 27610 10368 27930 10369
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 10303 27930 10304
rect 0 9800 480 9920
rect 7610 9824 7930 9825
rect 62 9346 122 9800
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7930 9824
rect 7610 9759 7930 9760
rect 20944 9824 21264 9825
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 9759 21264 9760
rect 34277 9824 34597 9825
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 39520 9800 40000 9920
rect 34277 9759 34597 9760
rect 1393 9346 1459 9349
rect 62 9344 1459 9346
rect 62 9288 1398 9344
rect 1454 9288 1459 9344
rect 62 9286 1459 9288
rect 1393 9283 1459 9286
rect 35617 9346 35683 9349
rect 39622 9346 39682 9800
rect 35617 9344 39682 9346
rect 35617 9288 35622 9344
rect 35678 9288 39682 9344
rect 35617 9286 39682 9288
rect 35617 9283 35683 9286
rect 14277 9280 14597 9281
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 9215 14597 9216
rect 27610 9280 27930 9281
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 27610 9215 27930 9216
rect 1853 8938 1919 8941
rect 12893 8938 12959 8941
rect 1853 8936 12959 8938
rect 1853 8880 1858 8936
rect 1914 8880 12898 8936
rect 12954 8880 12959 8936
rect 1853 8878 12959 8880
rect 1853 8875 1919 8878
rect 12893 8875 12959 8878
rect 7610 8736 7930 8737
rect 0 8576 480 8696
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7930 8736
rect 7610 8671 7930 8672
rect 20944 8736 21264 8737
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 8671 21264 8672
rect 34277 8736 34597 8737
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 8671 34597 8672
rect 39520 8576 40000 8696
rect 62 8394 122 8576
rect 11053 8394 11119 8397
rect 62 8392 11119 8394
rect 62 8336 11058 8392
rect 11114 8336 11119 8392
rect 62 8334 11119 8336
rect 11053 8331 11119 8334
rect 14277 8192 14597 8193
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 8127 14597 8128
rect 27610 8192 27930 8193
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 8127 27930 8128
rect 36077 8122 36143 8125
rect 39622 8122 39682 8576
rect 36077 8120 39682 8122
rect 36077 8064 36082 8120
rect 36138 8064 39682 8120
rect 36077 8062 39682 8064
rect 36077 8059 36143 8062
rect 7610 7648 7930 7649
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7930 7648
rect 7610 7583 7930 7584
rect 20944 7648 21264 7649
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 7583 21264 7584
rect 34277 7648 34597 7649
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 7583 34597 7584
rect 13905 7442 13971 7445
rect 15101 7442 15167 7445
rect 35249 7442 35315 7445
rect 13905 7440 35315 7442
rect 13905 7384 13910 7440
rect 13966 7384 15106 7440
rect 15162 7384 35254 7440
rect 35310 7384 35315 7440
rect 13905 7382 35315 7384
rect 13905 7379 13971 7382
rect 15101 7379 15167 7382
rect 35249 7379 35315 7382
rect 0 7304 480 7336
rect 0 7248 110 7304
rect 166 7248 480 7304
rect 0 7216 480 7248
rect 32213 7306 32279 7309
rect 39520 7306 40000 7336
rect 32213 7304 40000 7306
rect 32213 7248 32218 7304
rect 32274 7248 40000 7304
rect 32213 7246 40000 7248
rect 32213 7243 32279 7246
rect 39520 7216 40000 7246
rect 14277 7104 14597 7105
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 7039 14597 7040
rect 27610 7104 27930 7105
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 7039 27930 7040
rect 7610 6560 7930 6561
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7930 6560
rect 7610 6495 7930 6496
rect 20944 6560 21264 6561
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 6495 21264 6496
rect 34277 6560 34597 6561
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 34277 6495 34597 6496
rect 12249 6218 12315 6221
rect 35433 6218 35499 6221
rect 12249 6216 35499 6218
rect 12249 6160 12254 6216
rect 12310 6160 35438 6216
rect 35494 6160 35499 6216
rect 12249 6158 35499 6160
rect 12249 6155 12315 6158
rect 35433 6155 35499 6158
rect 14277 6016 14597 6017
rect 0 5856 480 5976
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 5951 14597 5952
rect 27610 6016 27930 6017
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 5951 27930 5952
rect 39520 5946 40000 5976
rect 39492 5944 40000 5946
rect 39492 5888 39578 5944
rect 39634 5888 40000 5944
rect 39492 5886 40000 5888
rect 39520 5856 40000 5886
rect 62 5538 122 5856
rect 7281 5810 7347 5813
rect 23289 5810 23355 5813
rect 7281 5808 23355 5810
rect 7281 5752 7286 5808
rect 7342 5752 23294 5808
rect 23350 5752 23355 5808
rect 7281 5750 23355 5752
rect 7281 5747 7347 5750
rect 23289 5747 23355 5750
rect 1025 5538 1091 5541
rect 62 5536 1091 5538
rect 62 5480 1030 5536
rect 1086 5480 1091 5536
rect 62 5478 1091 5480
rect 1025 5475 1091 5478
rect 7610 5472 7930 5473
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7930 5472
rect 7610 5407 7930 5408
rect 20944 5472 21264 5473
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 5407 21264 5408
rect 34277 5472 34597 5473
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 34277 5407 34597 5408
rect 1853 5130 1919 5133
rect 62 5128 1919 5130
rect 62 5072 1858 5128
rect 1914 5072 1919 5128
rect 62 5070 1919 5072
rect 62 4616 122 5070
rect 1853 5067 1919 5070
rect 2037 5130 2103 5133
rect 14733 5132 14799 5133
rect 14733 5130 14780 5132
rect 2037 5128 14780 5130
rect 2037 5072 2042 5128
rect 2098 5072 14738 5128
rect 2037 5070 14780 5072
rect 2037 5067 2103 5070
rect 14733 5068 14780 5070
rect 14844 5068 14850 5132
rect 14733 5067 14799 5068
rect 9857 4994 9923 4997
rect 14089 4994 14155 4997
rect 9857 4992 14155 4994
rect 9857 4936 9862 4992
rect 9918 4936 14094 4992
rect 14150 4936 14155 4992
rect 9857 4934 14155 4936
rect 9857 4931 9923 4934
rect 14089 4931 14155 4934
rect 14277 4928 14597 4929
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 4863 14597 4864
rect 27610 4928 27930 4929
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 4863 27930 4864
rect 1853 4722 1919 4725
rect 7189 4722 7255 4725
rect 1853 4720 7255 4722
rect 1853 4664 1858 4720
rect 1914 4664 7194 4720
rect 7250 4664 7255 4720
rect 1853 4662 7255 4664
rect 1853 4659 1919 4662
rect 7189 4659 7255 4662
rect 11789 4722 11855 4725
rect 16481 4722 16547 4725
rect 11789 4720 16547 4722
rect 11789 4664 11794 4720
rect 11850 4664 16486 4720
rect 16542 4664 16547 4720
rect 11789 4662 16547 4664
rect 11789 4659 11855 4662
rect 16481 4659 16547 4662
rect 0 4496 480 4616
rect 4337 4586 4403 4589
rect 17033 4586 17099 4589
rect 4337 4584 17099 4586
rect 4337 4528 4342 4584
rect 4398 4528 17038 4584
rect 17094 4528 17099 4584
rect 4337 4526 17099 4528
rect 4337 4523 4403 4526
rect 17033 4523 17099 4526
rect 39520 4496 40000 4616
rect 11513 4450 11579 4453
rect 15561 4450 15627 4453
rect 11513 4448 15627 4450
rect 11513 4392 11518 4448
rect 11574 4392 15566 4448
rect 15622 4392 15627 4448
rect 11513 4390 15627 4392
rect 11513 4387 11579 4390
rect 15561 4387 15627 4390
rect 7610 4384 7930 4385
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7930 4384
rect 7610 4319 7930 4320
rect 20944 4384 21264 4385
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 4319 21264 4320
rect 34277 4384 34597 4385
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 34277 4319 34597 4320
rect 35525 4314 35591 4317
rect 39622 4314 39682 4496
rect 35525 4312 39682 4314
rect 35525 4256 35530 4312
rect 35586 4256 39682 4312
rect 35525 4254 39682 4256
rect 35525 4251 35591 4254
rect 4521 4178 4587 4181
rect 9213 4178 9279 4181
rect 10041 4178 10107 4181
rect 11237 4178 11303 4181
rect 4521 4176 11303 4178
rect 4521 4120 4526 4176
rect 4582 4120 9218 4176
rect 9274 4120 10046 4176
rect 10102 4120 11242 4176
rect 11298 4120 11303 4176
rect 4521 4118 11303 4120
rect 4521 4115 4587 4118
rect 9213 4115 9279 4118
rect 10041 4115 10107 4118
rect 11237 4115 11303 4118
rect 7741 4042 7807 4045
rect 12709 4042 12775 4045
rect 12985 4042 13051 4045
rect 7741 4040 13051 4042
rect 7741 3984 7746 4040
rect 7802 3984 12714 4040
rect 12770 3984 12990 4040
rect 13046 3984 13051 4040
rect 7741 3982 13051 3984
rect 7741 3979 7807 3982
rect 12709 3979 12775 3982
rect 12985 3979 13051 3982
rect 14825 4042 14891 4045
rect 17677 4042 17743 4045
rect 18873 4042 18939 4045
rect 21725 4042 21791 4045
rect 14825 4040 21791 4042
rect 14825 3984 14830 4040
rect 14886 3984 17682 4040
rect 17738 3984 18878 4040
rect 18934 3984 21730 4040
rect 21786 3984 21791 4040
rect 14825 3982 21791 3984
rect 14825 3979 14891 3982
rect 17677 3979 17743 3982
rect 18873 3979 18939 3982
rect 21725 3979 21791 3982
rect 8477 3906 8543 3909
rect 9029 3906 9095 3909
rect 11973 3906 12039 3909
rect 8477 3904 12039 3906
rect 8477 3848 8482 3904
rect 8538 3848 9034 3904
rect 9090 3848 11978 3904
rect 12034 3848 12039 3904
rect 8477 3846 12039 3848
rect 8477 3843 8543 3846
rect 9029 3843 9095 3846
rect 11973 3843 12039 3846
rect 14277 3840 14597 3841
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 3775 14597 3776
rect 27610 3840 27930 3841
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 27610 3775 27930 3776
rect 6729 3770 6795 3773
rect 7189 3770 7255 3773
rect 10593 3770 10659 3773
rect 11329 3770 11395 3773
rect 6729 3768 11395 3770
rect 6729 3712 6734 3768
rect 6790 3712 7194 3768
rect 7250 3712 10598 3768
rect 10654 3712 11334 3768
rect 11390 3712 11395 3768
rect 6729 3710 11395 3712
rect 6729 3707 6795 3710
rect 7189 3707 7255 3710
rect 10593 3707 10659 3710
rect 11329 3707 11395 3710
rect 14549 3634 14615 3637
rect 20437 3634 20503 3637
rect 14549 3632 20503 3634
rect 14549 3576 14554 3632
rect 14610 3576 20442 3632
rect 20498 3576 20503 3632
rect 14549 3574 20503 3576
rect 14549 3571 14615 3574
rect 20437 3571 20503 3574
rect 12617 3498 12683 3501
rect 15653 3498 15719 3501
rect 12617 3496 15719 3498
rect 12617 3440 12622 3496
rect 12678 3440 15658 3496
rect 15714 3440 15719 3496
rect 12617 3438 15719 3440
rect 12617 3435 12683 3438
rect 15653 3435 15719 3438
rect 20989 3498 21055 3501
rect 23473 3498 23539 3501
rect 20989 3496 23539 3498
rect 20989 3440 20994 3496
rect 21050 3440 23478 3496
rect 23534 3440 23539 3496
rect 20989 3438 23539 3440
rect 20989 3435 21055 3438
rect 23473 3435 23539 3438
rect 11881 3362 11947 3365
rect 15837 3362 15903 3365
rect 11881 3360 15903 3362
rect 11881 3304 11886 3360
rect 11942 3304 15842 3360
rect 15898 3304 15903 3360
rect 11881 3302 15903 3304
rect 11881 3299 11947 3302
rect 15837 3299 15903 3302
rect 7610 3296 7930 3297
rect 0 3224 480 3256
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7930 3296
rect 7610 3231 7930 3232
rect 20944 3296 21264 3297
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 3231 21264 3232
rect 34277 3296 34597 3297
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 3231 34597 3232
rect 0 3168 110 3224
rect 166 3168 480 3224
rect 0 3136 480 3168
rect 12525 3226 12591 3229
rect 19333 3226 19399 3229
rect 12525 3224 19399 3226
rect 12525 3168 12530 3224
rect 12586 3168 19338 3224
rect 19394 3168 19399 3224
rect 12525 3166 19399 3168
rect 12525 3163 12591 3166
rect 19333 3163 19399 3166
rect 34697 3226 34763 3229
rect 39520 3226 40000 3256
rect 34697 3224 40000 3226
rect 34697 3168 34702 3224
rect 34758 3168 40000 3224
rect 34697 3166 40000 3168
rect 34697 3163 34763 3166
rect 39520 3136 40000 3166
rect 14277 2752 14597 2753
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2687 14597 2688
rect 27610 2752 27930 2753
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 27610 2687 27930 2688
rect 8661 2546 8727 2549
rect 16849 2546 16915 2549
rect 8661 2544 16915 2546
rect 8661 2488 8666 2544
rect 8722 2488 16854 2544
rect 16910 2488 16915 2544
rect 8661 2486 16915 2488
rect 8661 2483 8727 2486
rect 16849 2483 16915 2486
rect 22277 2546 22343 2549
rect 38469 2546 38535 2549
rect 22277 2544 38535 2546
rect 22277 2488 22282 2544
rect 22338 2488 38474 2544
rect 38530 2488 38535 2544
rect 22277 2486 38535 2488
rect 22277 2483 22343 2486
rect 38469 2483 38535 2486
rect 7465 2410 7531 2413
rect 62 2408 7531 2410
rect 62 2352 7470 2408
rect 7526 2352 7531 2408
rect 62 2350 7531 2352
rect 62 1896 122 2350
rect 7465 2347 7531 2350
rect 11697 2410 11763 2413
rect 21265 2410 21331 2413
rect 11697 2408 21331 2410
rect 11697 2352 11702 2408
rect 11758 2352 21270 2408
rect 21326 2352 21331 2408
rect 11697 2350 21331 2352
rect 11697 2347 11763 2350
rect 21265 2347 21331 2350
rect 31518 2348 31524 2412
rect 31588 2410 31594 2412
rect 31661 2410 31727 2413
rect 31588 2408 31727 2410
rect 31588 2352 31666 2408
rect 31722 2352 31727 2408
rect 31588 2350 31727 2352
rect 31588 2348 31594 2350
rect 31661 2347 31727 2350
rect 7610 2208 7930 2209
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7930 2208
rect 7610 2143 7930 2144
rect 20944 2208 21264 2209
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2143 21264 2144
rect 34277 2208 34597 2209
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 34277 2143 34597 2144
rect 10961 2138 11027 2141
rect 20069 2138 20135 2141
rect 10961 2136 20135 2138
rect 10961 2080 10966 2136
rect 11022 2080 20074 2136
rect 20130 2080 20135 2136
rect 10961 2078 20135 2080
rect 10961 2075 11027 2078
rect 20069 2075 20135 2078
rect 0 1776 480 1896
rect 18321 1866 18387 1869
rect 39389 1866 39455 1869
rect 18321 1864 39455 1866
rect 18321 1808 18326 1864
rect 18382 1808 39394 1864
rect 39450 1808 39455 1864
rect 18321 1806 39455 1808
rect 18321 1803 18387 1806
rect 39389 1803 39455 1806
rect 39520 1776 40000 1896
rect 2957 1730 3023 1733
rect 4102 1730 4108 1732
rect 2957 1728 4108 1730
rect 2957 1672 2962 1728
rect 3018 1672 4108 1728
rect 2957 1670 4108 1672
rect 2957 1667 3023 1670
rect 4102 1668 4108 1670
rect 4172 1668 4178 1732
rect 29913 1594 29979 1597
rect 39622 1594 39682 1776
rect 29913 1592 39682 1594
rect 29913 1536 29918 1592
rect 29974 1536 39682 1592
rect 29913 1534 39682 1536
rect 29913 1531 29979 1534
rect 21449 1458 21515 1461
rect 29085 1458 29151 1461
rect 21449 1456 29151 1458
rect 21449 1400 21454 1456
rect 21510 1400 29090 1456
rect 29146 1400 29151 1456
rect 21449 1398 29151 1400
rect 21449 1395 21515 1398
rect 29085 1395 29151 1398
rect 1393 1186 1459 1189
rect 62 1184 1459 1186
rect 62 1128 1398 1184
rect 1454 1128 1459 1184
rect 62 1126 1459 1128
rect 62 672 122 1126
rect 1393 1123 1459 1126
rect 0 552 480 672
rect 39520 642 40000 672
rect 39492 640 40000 642
rect 39492 584 39578 640
rect 39634 584 40000 640
rect 39492 582 40000 584
rect 39520 552 40000 582
rect 23422 36 23428 100
rect 23492 98 23498 100
rect 24577 98 24643 101
rect 23492 96 24643 98
rect 23492 40 24582 96
rect 24638 40 24643 96
rect 23492 38 24643 40
rect 23492 36 23498 38
rect 24577 35 24643 38
<< via3 >>
rect 14285 13628 14349 13632
rect 14285 13572 14289 13628
rect 14289 13572 14345 13628
rect 14345 13572 14349 13628
rect 14285 13568 14349 13572
rect 14365 13628 14429 13632
rect 14365 13572 14369 13628
rect 14369 13572 14425 13628
rect 14425 13572 14429 13628
rect 14365 13568 14429 13572
rect 14445 13628 14509 13632
rect 14445 13572 14449 13628
rect 14449 13572 14505 13628
rect 14505 13572 14509 13628
rect 14445 13568 14509 13572
rect 14525 13628 14589 13632
rect 14525 13572 14529 13628
rect 14529 13572 14585 13628
rect 14585 13572 14589 13628
rect 14525 13568 14589 13572
rect 27618 13628 27682 13632
rect 27618 13572 27622 13628
rect 27622 13572 27678 13628
rect 27678 13572 27682 13628
rect 27618 13568 27682 13572
rect 27698 13628 27762 13632
rect 27698 13572 27702 13628
rect 27702 13572 27758 13628
rect 27758 13572 27762 13628
rect 27698 13568 27762 13572
rect 27778 13628 27842 13632
rect 27778 13572 27782 13628
rect 27782 13572 27838 13628
rect 27838 13572 27842 13628
rect 27778 13568 27842 13572
rect 27858 13628 27922 13632
rect 27858 13572 27862 13628
rect 27862 13572 27918 13628
rect 27918 13572 27922 13628
rect 27858 13568 27922 13572
rect 7618 13084 7682 13088
rect 7618 13028 7622 13084
rect 7622 13028 7678 13084
rect 7678 13028 7682 13084
rect 7618 13024 7682 13028
rect 7698 13084 7762 13088
rect 7698 13028 7702 13084
rect 7702 13028 7758 13084
rect 7758 13028 7762 13084
rect 7698 13024 7762 13028
rect 7778 13084 7842 13088
rect 7778 13028 7782 13084
rect 7782 13028 7838 13084
rect 7838 13028 7842 13084
rect 7778 13024 7842 13028
rect 7858 13084 7922 13088
rect 7858 13028 7862 13084
rect 7862 13028 7918 13084
rect 7918 13028 7922 13084
rect 7858 13024 7922 13028
rect 20952 13084 21016 13088
rect 20952 13028 20956 13084
rect 20956 13028 21012 13084
rect 21012 13028 21016 13084
rect 20952 13024 21016 13028
rect 21032 13084 21096 13088
rect 21032 13028 21036 13084
rect 21036 13028 21092 13084
rect 21092 13028 21096 13084
rect 21032 13024 21096 13028
rect 21112 13084 21176 13088
rect 21112 13028 21116 13084
rect 21116 13028 21172 13084
rect 21172 13028 21176 13084
rect 21112 13024 21176 13028
rect 21192 13084 21256 13088
rect 21192 13028 21196 13084
rect 21196 13028 21252 13084
rect 21252 13028 21256 13084
rect 21192 13024 21256 13028
rect 34285 13084 34349 13088
rect 34285 13028 34289 13084
rect 34289 13028 34345 13084
rect 34345 13028 34349 13084
rect 34285 13024 34349 13028
rect 34365 13084 34429 13088
rect 34365 13028 34369 13084
rect 34369 13028 34425 13084
rect 34425 13028 34429 13084
rect 34365 13024 34429 13028
rect 34445 13084 34509 13088
rect 34445 13028 34449 13084
rect 34449 13028 34505 13084
rect 34505 13028 34509 13084
rect 34445 13024 34509 13028
rect 34525 13084 34589 13088
rect 34525 13028 34529 13084
rect 34529 13028 34585 13084
rect 34585 13028 34589 13084
rect 34525 13024 34589 13028
rect 14285 12540 14349 12544
rect 14285 12484 14289 12540
rect 14289 12484 14345 12540
rect 14345 12484 14349 12540
rect 14285 12480 14349 12484
rect 14365 12540 14429 12544
rect 14365 12484 14369 12540
rect 14369 12484 14425 12540
rect 14425 12484 14429 12540
rect 14365 12480 14429 12484
rect 14445 12540 14509 12544
rect 14445 12484 14449 12540
rect 14449 12484 14505 12540
rect 14505 12484 14509 12540
rect 14445 12480 14509 12484
rect 14525 12540 14589 12544
rect 14525 12484 14529 12540
rect 14529 12484 14585 12540
rect 14585 12484 14589 12540
rect 14525 12480 14589 12484
rect 27618 12540 27682 12544
rect 27618 12484 27622 12540
rect 27622 12484 27678 12540
rect 27678 12484 27682 12540
rect 27618 12480 27682 12484
rect 27698 12540 27762 12544
rect 27698 12484 27702 12540
rect 27702 12484 27758 12540
rect 27758 12484 27762 12540
rect 27698 12480 27762 12484
rect 27778 12540 27842 12544
rect 27778 12484 27782 12540
rect 27782 12484 27838 12540
rect 27838 12484 27842 12540
rect 27778 12480 27842 12484
rect 27858 12540 27922 12544
rect 27858 12484 27862 12540
rect 27862 12484 27918 12540
rect 27918 12484 27922 12540
rect 27858 12480 27922 12484
rect 7618 11996 7682 12000
rect 7618 11940 7622 11996
rect 7622 11940 7678 11996
rect 7678 11940 7682 11996
rect 7618 11936 7682 11940
rect 7698 11996 7762 12000
rect 7698 11940 7702 11996
rect 7702 11940 7758 11996
rect 7758 11940 7762 11996
rect 7698 11936 7762 11940
rect 7778 11996 7842 12000
rect 7778 11940 7782 11996
rect 7782 11940 7838 11996
rect 7838 11940 7842 11996
rect 7778 11936 7842 11940
rect 7858 11996 7922 12000
rect 7858 11940 7862 11996
rect 7862 11940 7918 11996
rect 7918 11940 7922 11996
rect 7858 11936 7922 11940
rect 20952 11996 21016 12000
rect 20952 11940 20956 11996
rect 20956 11940 21012 11996
rect 21012 11940 21016 11996
rect 20952 11936 21016 11940
rect 21032 11996 21096 12000
rect 21032 11940 21036 11996
rect 21036 11940 21092 11996
rect 21092 11940 21096 11996
rect 21032 11936 21096 11940
rect 21112 11996 21176 12000
rect 21112 11940 21116 11996
rect 21116 11940 21172 11996
rect 21172 11940 21176 11996
rect 21112 11936 21176 11940
rect 21192 11996 21256 12000
rect 21192 11940 21196 11996
rect 21196 11940 21252 11996
rect 21252 11940 21256 11996
rect 21192 11936 21256 11940
rect 34285 11996 34349 12000
rect 34285 11940 34289 11996
rect 34289 11940 34345 11996
rect 34345 11940 34349 11996
rect 34285 11936 34349 11940
rect 34365 11996 34429 12000
rect 34365 11940 34369 11996
rect 34369 11940 34425 11996
rect 34425 11940 34429 11996
rect 34365 11936 34429 11940
rect 34445 11996 34509 12000
rect 34445 11940 34449 11996
rect 34449 11940 34505 11996
rect 34505 11940 34509 11996
rect 34445 11936 34509 11940
rect 34525 11996 34589 12000
rect 34525 11940 34529 11996
rect 34529 11940 34585 11996
rect 34585 11940 34589 11996
rect 34525 11936 34589 11940
rect 14285 11452 14349 11456
rect 14285 11396 14289 11452
rect 14289 11396 14345 11452
rect 14345 11396 14349 11452
rect 14285 11392 14349 11396
rect 14365 11452 14429 11456
rect 14365 11396 14369 11452
rect 14369 11396 14425 11452
rect 14425 11396 14429 11452
rect 14365 11392 14429 11396
rect 14445 11452 14509 11456
rect 14445 11396 14449 11452
rect 14449 11396 14505 11452
rect 14505 11396 14509 11452
rect 14445 11392 14509 11396
rect 14525 11452 14589 11456
rect 14525 11396 14529 11452
rect 14529 11396 14585 11452
rect 14585 11396 14589 11452
rect 14525 11392 14589 11396
rect 27618 11452 27682 11456
rect 27618 11396 27622 11452
rect 27622 11396 27678 11452
rect 27678 11396 27682 11452
rect 27618 11392 27682 11396
rect 27698 11452 27762 11456
rect 27698 11396 27702 11452
rect 27702 11396 27758 11452
rect 27758 11396 27762 11452
rect 27698 11392 27762 11396
rect 27778 11452 27842 11456
rect 27778 11396 27782 11452
rect 27782 11396 27838 11452
rect 27838 11396 27842 11452
rect 27778 11392 27842 11396
rect 27858 11452 27922 11456
rect 27858 11396 27862 11452
rect 27862 11396 27918 11452
rect 27918 11396 27922 11452
rect 27858 11392 27922 11396
rect 60 11188 124 11252
rect 60 10916 124 10980
rect 7618 10908 7682 10912
rect 7618 10852 7622 10908
rect 7622 10852 7678 10908
rect 7678 10852 7682 10908
rect 7618 10848 7682 10852
rect 7698 10908 7762 10912
rect 7698 10852 7702 10908
rect 7702 10852 7758 10908
rect 7758 10852 7762 10908
rect 7698 10848 7762 10852
rect 7778 10908 7842 10912
rect 7778 10852 7782 10908
rect 7782 10852 7838 10908
rect 7838 10852 7842 10908
rect 7778 10848 7842 10852
rect 7858 10908 7922 10912
rect 7858 10852 7862 10908
rect 7862 10852 7918 10908
rect 7918 10852 7922 10908
rect 7858 10848 7922 10852
rect 20952 10908 21016 10912
rect 20952 10852 20956 10908
rect 20956 10852 21012 10908
rect 21012 10852 21016 10908
rect 20952 10848 21016 10852
rect 21032 10908 21096 10912
rect 21032 10852 21036 10908
rect 21036 10852 21092 10908
rect 21092 10852 21096 10908
rect 21032 10848 21096 10852
rect 21112 10908 21176 10912
rect 21112 10852 21116 10908
rect 21116 10852 21172 10908
rect 21172 10852 21176 10908
rect 21112 10848 21176 10852
rect 21192 10908 21256 10912
rect 21192 10852 21196 10908
rect 21196 10852 21252 10908
rect 21252 10852 21256 10908
rect 21192 10848 21256 10852
rect 34285 10908 34349 10912
rect 34285 10852 34289 10908
rect 34289 10852 34345 10908
rect 34345 10852 34349 10908
rect 34285 10848 34349 10852
rect 34365 10908 34429 10912
rect 34365 10852 34369 10908
rect 34369 10852 34425 10908
rect 34425 10852 34429 10908
rect 34365 10848 34429 10852
rect 34445 10908 34509 10912
rect 34445 10852 34449 10908
rect 34449 10852 34505 10908
rect 34505 10852 34509 10908
rect 34445 10848 34509 10852
rect 34525 10908 34589 10912
rect 34525 10852 34529 10908
rect 34529 10852 34585 10908
rect 34585 10852 34589 10908
rect 34525 10848 34589 10852
rect 14285 10364 14349 10368
rect 14285 10308 14289 10364
rect 14289 10308 14345 10364
rect 14345 10308 14349 10364
rect 14285 10304 14349 10308
rect 14365 10364 14429 10368
rect 14365 10308 14369 10364
rect 14369 10308 14425 10364
rect 14425 10308 14429 10364
rect 14365 10304 14429 10308
rect 14445 10364 14509 10368
rect 14445 10308 14449 10364
rect 14449 10308 14505 10364
rect 14505 10308 14509 10364
rect 14445 10304 14509 10308
rect 14525 10364 14589 10368
rect 14525 10308 14529 10364
rect 14529 10308 14585 10364
rect 14585 10308 14589 10364
rect 14525 10304 14589 10308
rect 27618 10364 27682 10368
rect 27618 10308 27622 10364
rect 27622 10308 27678 10364
rect 27678 10308 27682 10364
rect 27618 10304 27682 10308
rect 27698 10364 27762 10368
rect 27698 10308 27702 10364
rect 27702 10308 27758 10364
rect 27758 10308 27762 10364
rect 27698 10304 27762 10308
rect 27778 10364 27842 10368
rect 27778 10308 27782 10364
rect 27782 10308 27838 10364
rect 27838 10308 27842 10364
rect 27778 10304 27842 10308
rect 27858 10364 27922 10368
rect 27858 10308 27862 10364
rect 27862 10308 27918 10364
rect 27918 10308 27922 10364
rect 27858 10304 27922 10308
rect 7618 9820 7682 9824
rect 7618 9764 7622 9820
rect 7622 9764 7678 9820
rect 7678 9764 7682 9820
rect 7618 9760 7682 9764
rect 7698 9820 7762 9824
rect 7698 9764 7702 9820
rect 7702 9764 7758 9820
rect 7758 9764 7762 9820
rect 7698 9760 7762 9764
rect 7778 9820 7842 9824
rect 7778 9764 7782 9820
rect 7782 9764 7838 9820
rect 7838 9764 7842 9820
rect 7778 9760 7842 9764
rect 7858 9820 7922 9824
rect 7858 9764 7862 9820
rect 7862 9764 7918 9820
rect 7918 9764 7922 9820
rect 7858 9760 7922 9764
rect 20952 9820 21016 9824
rect 20952 9764 20956 9820
rect 20956 9764 21012 9820
rect 21012 9764 21016 9820
rect 20952 9760 21016 9764
rect 21032 9820 21096 9824
rect 21032 9764 21036 9820
rect 21036 9764 21092 9820
rect 21092 9764 21096 9820
rect 21032 9760 21096 9764
rect 21112 9820 21176 9824
rect 21112 9764 21116 9820
rect 21116 9764 21172 9820
rect 21172 9764 21176 9820
rect 21112 9760 21176 9764
rect 21192 9820 21256 9824
rect 21192 9764 21196 9820
rect 21196 9764 21252 9820
rect 21252 9764 21256 9820
rect 21192 9760 21256 9764
rect 34285 9820 34349 9824
rect 34285 9764 34289 9820
rect 34289 9764 34345 9820
rect 34345 9764 34349 9820
rect 34285 9760 34349 9764
rect 34365 9820 34429 9824
rect 34365 9764 34369 9820
rect 34369 9764 34425 9820
rect 34425 9764 34429 9820
rect 34365 9760 34429 9764
rect 34445 9820 34509 9824
rect 34445 9764 34449 9820
rect 34449 9764 34505 9820
rect 34505 9764 34509 9820
rect 34445 9760 34509 9764
rect 34525 9820 34589 9824
rect 34525 9764 34529 9820
rect 34529 9764 34585 9820
rect 34585 9764 34589 9820
rect 34525 9760 34589 9764
rect 14285 9276 14349 9280
rect 14285 9220 14289 9276
rect 14289 9220 14345 9276
rect 14345 9220 14349 9276
rect 14285 9216 14349 9220
rect 14365 9276 14429 9280
rect 14365 9220 14369 9276
rect 14369 9220 14425 9276
rect 14425 9220 14429 9276
rect 14365 9216 14429 9220
rect 14445 9276 14509 9280
rect 14445 9220 14449 9276
rect 14449 9220 14505 9276
rect 14505 9220 14509 9276
rect 14445 9216 14509 9220
rect 14525 9276 14589 9280
rect 14525 9220 14529 9276
rect 14529 9220 14585 9276
rect 14585 9220 14589 9276
rect 14525 9216 14589 9220
rect 27618 9276 27682 9280
rect 27618 9220 27622 9276
rect 27622 9220 27678 9276
rect 27678 9220 27682 9276
rect 27618 9216 27682 9220
rect 27698 9276 27762 9280
rect 27698 9220 27702 9276
rect 27702 9220 27758 9276
rect 27758 9220 27762 9276
rect 27698 9216 27762 9220
rect 27778 9276 27842 9280
rect 27778 9220 27782 9276
rect 27782 9220 27838 9276
rect 27838 9220 27842 9276
rect 27778 9216 27842 9220
rect 27858 9276 27922 9280
rect 27858 9220 27862 9276
rect 27862 9220 27918 9276
rect 27918 9220 27922 9276
rect 27858 9216 27922 9220
rect 7618 8732 7682 8736
rect 7618 8676 7622 8732
rect 7622 8676 7678 8732
rect 7678 8676 7682 8732
rect 7618 8672 7682 8676
rect 7698 8732 7762 8736
rect 7698 8676 7702 8732
rect 7702 8676 7758 8732
rect 7758 8676 7762 8732
rect 7698 8672 7762 8676
rect 7778 8732 7842 8736
rect 7778 8676 7782 8732
rect 7782 8676 7838 8732
rect 7838 8676 7842 8732
rect 7778 8672 7842 8676
rect 7858 8732 7922 8736
rect 7858 8676 7862 8732
rect 7862 8676 7918 8732
rect 7918 8676 7922 8732
rect 7858 8672 7922 8676
rect 20952 8732 21016 8736
rect 20952 8676 20956 8732
rect 20956 8676 21012 8732
rect 21012 8676 21016 8732
rect 20952 8672 21016 8676
rect 21032 8732 21096 8736
rect 21032 8676 21036 8732
rect 21036 8676 21092 8732
rect 21092 8676 21096 8732
rect 21032 8672 21096 8676
rect 21112 8732 21176 8736
rect 21112 8676 21116 8732
rect 21116 8676 21172 8732
rect 21172 8676 21176 8732
rect 21112 8672 21176 8676
rect 21192 8732 21256 8736
rect 21192 8676 21196 8732
rect 21196 8676 21252 8732
rect 21252 8676 21256 8732
rect 21192 8672 21256 8676
rect 34285 8732 34349 8736
rect 34285 8676 34289 8732
rect 34289 8676 34345 8732
rect 34345 8676 34349 8732
rect 34285 8672 34349 8676
rect 34365 8732 34429 8736
rect 34365 8676 34369 8732
rect 34369 8676 34425 8732
rect 34425 8676 34429 8732
rect 34365 8672 34429 8676
rect 34445 8732 34509 8736
rect 34445 8676 34449 8732
rect 34449 8676 34505 8732
rect 34505 8676 34509 8732
rect 34445 8672 34509 8676
rect 34525 8732 34589 8736
rect 34525 8676 34529 8732
rect 34529 8676 34585 8732
rect 34585 8676 34589 8732
rect 34525 8672 34589 8676
rect 14285 8188 14349 8192
rect 14285 8132 14289 8188
rect 14289 8132 14345 8188
rect 14345 8132 14349 8188
rect 14285 8128 14349 8132
rect 14365 8188 14429 8192
rect 14365 8132 14369 8188
rect 14369 8132 14425 8188
rect 14425 8132 14429 8188
rect 14365 8128 14429 8132
rect 14445 8188 14509 8192
rect 14445 8132 14449 8188
rect 14449 8132 14505 8188
rect 14505 8132 14509 8188
rect 14445 8128 14509 8132
rect 14525 8188 14589 8192
rect 14525 8132 14529 8188
rect 14529 8132 14585 8188
rect 14585 8132 14589 8188
rect 14525 8128 14589 8132
rect 27618 8188 27682 8192
rect 27618 8132 27622 8188
rect 27622 8132 27678 8188
rect 27678 8132 27682 8188
rect 27618 8128 27682 8132
rect 27698 8188 27762 8192
rect 27698 8132 27702 8188
rect 27702 8132 27758 8188
rect 27758 8132 27762 8188
rect 27698 8128 27762 8132
rect 27778 8188 27842 8192
rect 27778 8132 27782 8188
rect 27782 8132 27838 8188
rect 27838 8132 27842 8188
rect 27778 8128 27842 8132
rect 27858 8188 27922 8192
rect 27858 8132 27862 8188
rect 27862 8132 27918 8188
rect 27918 8132 27922 8188
rect 27858 8128 27922 8132
rect 7618 7644 7682 7648
rect 7618 7588 7622 7644
rect 7622 7588 7678 7644
rect 7678 7588 7682 7644
rect 7618 7584 7682 7588
rect 7698 7644 7762 7648
rect 7698 7588 7702 7644
rect 7702 7588 7758 7644
rect 7758 7588 7762 7644
rect 7698 7584 7762 7588
rect 7778 7644 7842 7648
rect 7778 7588 7782 7644
rect 7782 7588 7838 7644
rect 7838 7588 7842 7644
rect 7778 7584 7842 7588
rect 7858 7644 7922 7648
rect 7858 7588 7862 7644
rect 7862 7588 7918 7644
rect 7918 7588 7922 7644
rect 7858 7584 7922 7588
rect 20952 7644 21016 7648
rect 20952 7588 20956 7644
rect 20956 7588 21012 7644
rect 21012 7588 21016 7644
rect 20952 7584 21016 7588
rect 21032 7644 21096 7648
rect 21032 7588 21036 7644
rect 21036 7588 21092 7644
rect 21092 7588 21096 7644
rect 21032 7584 21096 7588
rect 21112 7644 21176 7648
rect 21112 7588 21116 7644
rect 21116 7588 21172 7644
rect 21172 7588 21176 7644
rect 21112 7584 21176 7588
rect 21192 7644 21256 7648
rect 21192 7588 21196 7644
rect 21196 7588 21252 7644
rect 21252 7588 21256 7644
rect 21192 7584 21256 7588
rect 34285 7644 34349 7648
rect 34285 7588 34289 7644
rect 34289 7588 34345 7644
rect 34345 7588 34349 7644
rect 34285 7584 34349 7588
rect 34365 7644 34429 7648
rect 34365 7588 34369 7644
rect 34369 7588 34425 7644
rect 34425 7588 34429 7644
rect 34365 7584 34429 7588
rect 34445 7644 34509 7648
rect 34445 7588 34449 7644
rect 34449 7588 34505 7644
rect 34505 7588 34509 7644
rect 34445 7584 34509 7588
rect 34525 7644 34589 7648
rect 34525 7588 34529 7644
rect 34529 7588 34585 7644
rect 34585 7588 34589 7644
rect 34525 7584 34589 7588
rect 14285 7100 14349 7104
rect 14285 7044 14289 7100
rect 14289 7044 14345 7100
rect 14345 7044 14349 7100
rect 14285 7040 14349 7044
rect 14365 7100 14429 7104
rect 14365 7044 14369 7100
rect 14369 7044 14425 7100
rect 14425 7044 14429 7100
rect 14365 7040 14429 7044
rect 14445 7100 14509 7104
rect 14445 7044 14449 7100
rect 14449 7044 14505 7100
rect 14505 7044 14509 7100
rect 14445 7040 14509 7044
rect 14525 7100 14589 7104
rect 14525 7044 14529 7100
rect 14529 7044 14585 7100
rect 14585 7044 14589 7100
rect 14525 7040 14589 7044
rect 27618 7100 27682 7104
rect 27618 7044 27622 7100
rect 27622 7044 27678 7100
rect 27678 7044 27682 7100
rect 27618 7040 27682 7044
rect 27698 7100 27762 7104
rect 27698 7044 27702 7100
rect 27702 7044 27758 7100
rect 27758 7044 27762 7100
rect 27698 7040 27762 7044
rect 27778 7100 27842 7104
rect 27778 7044 27782 7100
rect 27782 7044 27838 7100
rect 27838 7044 27842 7100
rect 27778 7040 27842 7044
rect 27858 7100 27922 7104
rect 27858 7044 27862 7100
rect 27862 7044 27918 7100
rect 27918 7044 27922 7100
rect 27858 7040 27922 7044
rect 7618 6556 7682 6560
rect 7618 6500 7622 6556
rect 7622 6500 7678 6556
rect 7678 6500 7682 6556
rect 7618 6496 7682 6500
rect 7698 6556 7762 6560
rect 7698 6500 7702 6556
rect 7702 6500 7758 6556
rect 7758 6500 7762 6556
rect 7698 6496 7762 6500
rect 7778 6556 7842 6560
rect 7778 6500 7782 6556
rect 7782 6500 7838 6556
rect 7838 6500 7842 6556
rect 7778 6496 7842 6500
rect 7858 6556 7922 6560
rect 7858 6500 7862 6556
rect 7862 6500 7918 6556
rect 7918 6500 7922 6556
rect 7858 6496 7922 6500
rect 20952 6556 21016 6560
rect 20952 6500 20956 6556
rect 20956 6500 21012 6556
rect 21012 6500 21016 6556
rect 20952 6496 21016 6500
rect 21032 6556 21096 6560
rect 21032 6500 21036 6556
rect 21036 6500 21092 6556
rect 21092 6500 21096 6556
rect 21032 6496 21096 6500
rect 21112 6556 21176 6560
rect 21112 6500 21116 6556
rect 21116 6500 21172 6556
rect 21172 6500 21176 6556
rect 21112 6496 21176 6500
rect 21192 6556 21256 6560
rect 21192 6500 21196 6556
rect 21196 6500 21252 6556
rect 21252 6500 21256 6556
rect 21192 6496 21256 6500
rect 34285 6556 34349 6560
rect 34285 6500 34289 6556
rect 34289 6500 34345 6556
rect 34345 6500 34349 6556
rect 34285 6496 34349 6500
rect 34365 6556 34429 6560
rect 34365 6500 34369 6556
rect 34369 6500 34425 6556
rect 34425 6500 34429 6556
rect 34365 6496 34429 6500
rect 34445 6556 34509 6560
rect 34445 6500 34449 6556
rect 34449 6500 34505 6556
rect 34505 6500 34509 6556
rect 34445 6496 34509 6500
rect 34525 6556 34589 6560
rect 34525 6500 34529 6556
rect 34529 6500 34585 6556
rect 34585 6500 34589 6556
rect 34525 6496 34589 6500
rect 14285 6012 14349 6016
rect 14285 5956 14289 6012
rect 14289 5956 14345 6012
rect 14345 5956 14349 6012
rect 14285 5952 14349 5956
rect 14365 6012 14429 6016
rect 14365 5956 14369 6012
rect 14369 5956 14425 6012
rect 14425 5956 14429 6012
rect 14365 5952 14429 5956
rect 14445 6012 14509 6016
rect 14445 5956 14449 6012
rect 14449 5956 14505 6012
rect 14505 5956 14509 6012
rect 14445 5952 14509 5956
rect 14525 6012 14589 6016
rect 14525 5956 14529 6012
rect 14529 5956 14585 6012
rect 14585 5956 14589 6012
rect 14525 5952 14589 5956
rect 27618 6012 27682 6016
rect 27618 5956 27622 6012
rect 27622 5956 27678 6012
rect 27678 5956 27682 6012
rect 27618 5952 27682 5956
rect 27698 6012 27762 6016
rect 27698 5956 27702 6012
rect 27702 5956 27758 6012
rect 27758 5956 27762 6012
rect 27698 5952 27762 5956
rect 27778 6012 27842 6016
rect 27778 5956 27782 6012
rect 27782 5956 27838 6012
rect 27838 5956 27842 6012
rect 27778 5952 27842 5956
rect 27858 6012 27922 6016
rect 27858 5956 27862 6012
rect 27862 5956 27918 6012
rect 27918 5956 27922 6012
rect 27858 5952 27922 5956
rect 7618 5468 7682 5472
rect 7618 5412 7622 5468
rect 7622 5412 7678 5468
rect 7678 5412 7682 5468
rect 7618 5408 7682 5412
rect 7698 5468 7762 5472
rect 7698 5412 7702 5468
rect 7702 5412 7758 5468
rect 7758 5412 7762 5468
rect 7698 5408 7762 5412
rect 7778 5468 7842 5472
rect 7778 5412 7782 5468
rect 7782 5412 7838 5468
rect 7838 5412 7842 5468
rect 7778 5408 7842 5412
rect 7858 5468 7922 5472
rect 7858 5412 7862 5468
rect 7862 5412 7918 5468
rect 7918 5412 7922 5468
rect 7858 5408 7922 5412
rect 20952 5468 21016 5472
rect 20952 5412 20956 5468
rect 20956 5412 21012 5468
rect 21012 5412 21016 5468
rect 20952 5408 21016 5412
rect 21032 5468 21096 5472
rect 21032 5412 21036 5468
rect 21036 5412 21092 5468
rect 21092 5412 21096 5468
rect 21032 5408 21096 5412
rect 21112 5468 21176 5472
rect 21112 5412 21116 5468
rect 21116 5412 21172 5468
rect 21172 5412 21176 5468
rect 21112 5408 21176 5412
rect 21192 5468 21256 5472
rect 21192 5412 21196 5468
rect 21196 5412 21252 5468
rect 21252 5412 21256 5468
rect 21192 5408 21256 5412
rect 34285 5468 34349 5472
rect 34285 5412 34289 5468
rect 34289 5412 34345 5468
rect 34345 5412 34349 5468
rect 34285 5408 34349 5412
rect 34365 5468 34429 5472
rect 34365 5412 34369 5468
rect 34369 5412 34425 5468
rect 34425 5412 34429 5468
rect 34365 5408 34429 5412
rect 34445 5468 34509 5472
rect 34445 5412 34449 5468
rect 34449 5412 34505 5468
rect 34505 5412 34509 5468
rect 34445 5408 34509 5412
rect 34525 5468 34589 5472
rect 34525 5412 34529 5468
rect 34529 5412 34585 5468
rect 34585 5412 34589 5468
rect 34525 5408 34589 5412
rect 14780 5128 14844 5132
rect 14780 5072 14794 5128
rect 14794 5072 14844 5128
rect 14780 5068 14844 5072
rect 14285 4924 14349 4928
rect 14285 4868 14289 4924
rect 14289 4868 14345 4924
rect 14345 4868 14349 4924
rect 14285 4864 14349 4868
rect 14365 4924 14429 4928
rect 14365 4868 14369 4924
rect 14369 4868 14425 4924
rect 14425 4868 14429 4924
rect 14365 4864 14429 4868
rect 14445 4924 14509 4928
rect 14445 4868 14449 4924
rect 14449 4868 14505 4924
rect 14505 4868 14509 4924
rect 14445 4864 14509 4868
rect 14525 4924 14589 4928
rect 14525 4868 14529 4924
rect 14529 4868 14585 4924
rect 14585 4868 14589 4924
rect 14525 4864 14589 4868
rect 27618 4924 27682 4928
rect 27618 4868 27622 4924
rect 27622 4868 27678 4924
rect 27678 4868 27682 4924
rect 27618 4864 27682 4868
rect 27698 4924 27762 4928
rect 27698 4868 27702 4924
rect 27702 4868 27758 4924
rect 27758 4868 27762 4924
rect 27698 4864 27762 4868
rect 27778 4924 27842 4928
rect 27778 4868 27782 4924
rect 27782 4868 27838 4924
rect 27838 4868 27842 4924
rect 27778 4864 27842 4868
rect 27858 4924 27922 4928
rect 27858 4868 27862 4924
rect 27862 4868 27918 4924
rect 27918 4868 27922 4924
rect 27858 4864 27922 4868
rect 7618 4380 7682 4384
rect 7618 4324 7622 4380
rect 7622 4324 7678 4380
rect 7678 4324 7682 4380
rect 7618 4320 7682 4324
rect 7698 4380 7762 4384
rect 7698 4324 7702 4380
rect 7702 4324 7758 4380
rect 7758 4324 7762 4380
rect 7698 4320 7762 4324
rect 7778 4380 7842 4384
rect 7778 4324 7782 4380
rect 7782 4324 7838 4380
rect 7838 4324 7842 4380
rect 7778 4320 7842 4324
rect 7858 4380 7922 4384
rect 7858 4324 7862 4380
rect 7862 4324 7918 4380
rect 7918 4324 7922 4380
rect 7858 4320 7922 4324
rect 20952 4380 21016 4384
rect 20952 4324 20956 4380
rect 20956 4324 21012 4380
rect 21012 4324 21016 4380
rect 20952 4320 21016 4324
rect 21032 4380 21096 4384
rect 21032 4324 21036 4380
rect 21036 4324 21092 4380
rect 21092 4324 21096 4380
rect 21032 4320 21096 4324
rect 21112 4380 21176 4384
rect 21112 4324 21116 4380
rect 21116 4324 21172 4380
rect 21172 4324 21176 4380
rect 21112 4320 21176 4324
rect 21192 4380 21256 4384
rect 21192 4324 21196 4380
rect 21196 4324 21252 4380
rect 21252 4324 21256 4380
rect 21192 4320 21256 4324
rect 34285 4380 34349 4384
rect 34285 4324 34289 4380
rect 34289 4324 34345 4380
rect 34345 4324 34349 4380
rect 34285 4320 34349 4324
rect 34365 4380 34429 4384
rect 34365 4324 34369 4380
rect 34369 4324 34425 4380
rect 34425 4324 34429 4380
rect 34365 4320 34429 4324
rect 34445 4380 34509 4384
rect 34445 4324 34449 4380
rect 34449 4324 34505 4380
rect 34505 4324 34509 4380
rect 34445 4320 34509 4324
rect 34525 4380 34589 4384
rect 34525 4324 34529 4380
rect 34529 4324 34585 4380
rect 34585 4324 34589 4380
rect 34525 4320 34589 4324
rect 14285 3836 14349 3840
rect 14285 3780 14289 3836
rect 14289 3780 14345 3836
rect 14345 3780 14349 3836
rect 14285 3776 14349 3780
rect 14365 3836 14429 3840
rect 14365 3780 14369 3836
rect 14369 3780 14425 3836
rect 14425 3780 14429 3836
rect 14365 3776 14429 3780
rect 14445 3836 14509 3840
rect 14445 3780 14449 3836
rect 14449 3780 14505 3836
rect 14505 3780 14509 3836
rect 14445 3776 14509 3780
rect 14525 3836 14589 3840
rect 14525 3780 14529 3836
rect 14529 3780 14585 3836
rect 14585 3780 14589 3836
rect 14525 3776 14589 3780
rect 27618 3836 27682 3840
rect 27618 3780 27622 3836
rect 27622 3780 27678 3836
rect 27678 3780 27682 3836
rect 27618 3776 27682 3780
rect 27698 3836 27762 3840
rect 27698 3780 27702 3836
rect 27702 3780 27758 3836
rect 27758 3780 27762 3836
rect 27698 3776 27762 3780
rect 27778 3836 27842 3840
rect 27778 3780 27782 3836
rect 27782 3780 27838 3836
rect 27838 3780 27842 3836
rect 27778 3776 27842 3780
rect 27858 3836 27922 3840
rect 27858 3780 27862 3836
rect 27862 3780 27918 3836
rect 27918 3780 27922 3836
rect 27858 3776 27922 3780
rect 7618 3292 7682 3296
rect 7618 3236 7622 3292
rect 7622 3236 7678 3292
rect 7678 3236 7682 3292
rect 7618 3232 7682 3236
rect 7698 3292 7762 3296
rect 7698 3236 7702 3292
rect 7702 3236 7758 3292
rect 7758 3236 7762 3292
rect 7698 3232 7762 3236
rect 7778 3292 7842 3296
rect 7778 3236 7782 3292
rect 7782 3236 7838 3292
rect 7838 3236 7842 3292
rect 7778 3232 7842 3236
rect 7858 3292 7922 3296
rect 7858 3236 7862 3292
rect 7862 3236 7918 3292
rect 7918 3236 7922 3292
rect 7858 3232 7922 3236
rect 20952 3292 21016 3296
rect 20952 3236 20956 3292
rect 20956 3236 21012 3292
rect 21012 3236 21016 3292
rect 20952 3232 21016 3236
rect 21032 3292 21096 3296
rect 21032 3236 21036 3292
rect 21036 3236 21092 3292
rect 21092 3236 21096 3292
rect 21032 3232 21096 3236
rect 21112 3292 21176 3296
rect 21112 3236 21116 3292
rect 21116 3236 21172 3292
rect 21172 3236 21176 3292
rect 21112 3232 21176 3236
rect 21192 3292 21256 3296
rect 21192 3236 21196 3292
rect 21196 3236 21252 3292
rect 21252 3236 21256 3292
rect 21192 3232 21256 3236
rect 34285 3292 34349 3296
rect 34285 3236 34289 3292
rect 34289 3236 34345 3292
rect 34345 3236 34349 3292
rect 34285 3232 34349 3236
rect 34365 3292 34429 3296
rect 34365 3236 34369 3292
rect 34369 3236 34425 3292
rect 34425 3236 34429 3292
rect 34365 3232 34429 3236
rect 34445 3292 34509 3296
rect 34445 3236 34449 3292
rect 34449 3236 34505 3292
rect 34505 3236 34509 3292
rect 34445 3232 34509 3236
rect 34525 3292 34589 3296
rect 34525 3236 34529 3292
rect 34529 3236 34585 3292
rect 34585 3236 34589 3292
rect 34525 3232 34589 3236
rect 14285 2748 14349 2752
rect 14285 2692 14289 2748
rect 14289 2692 14345 2748
rect 14345 2692 14349 2748
rect 14285 2688 14349 2692
rect 14365 2748 14429 2752
rect 14365 2692 14369 2748
rect 14369 2692 14425 2748
rect 14425 2692 14429 2748
rect 14365 2688 14429 2692
rect 14445 2748 14509 2752
rect 14445 2692 14449 2748
rect 14449 2692 14505 2748
rect 14505 2692 14509 2748
rect 14445 2688 14509 2692
rect 14525 2748 14589 2752
rect 14525 2692 14529 2748
rect 14529 2692 14585 2748
rect 14585 2692 14589 2748
rect 14525 2688 14589 2692
rect 27618 2748 27682 2752
rect 27618 2692 27622 2748
rect 27622 2692 27678 2748
rect 27678 2692 27682 2748
rect 27618 2688 27682 2692
rect 27698 2748 27762 2752
rect 27698 2692 27702 2748
rect 27702 2692 27758 2748
rect 27758 2692 27762 2748
rect 27698 2688 27762 2692
rect 27778 2748 27842 2752
rect 27778 2692 27782 2748
rect 27782 2692 27838 2748
rect 27838 2692 27842 2748
rect 27778 2688 27842 2692
rect 27858 2748 27922 2752
rect 27858 2692 27862 2748
rect 27862 2692 27918 2748
rect 27918 2692 27922 2748
rect 27858 2688 27922 2692
rect 31524 2348 31588 2412
rect 7618 2204 7682 2208
rect 7618 2148 7622 2204
rect 7622 2148 7678 2204
rect 7678 2148 7682 2204
rect 7618 2144 7682 2148
rect 7698 2204 7762 2208
rect 7698 2148 7702 2204
rect 7702 2148 7758 2204
rect 7758 2148 7762 2204
rect 7698 2144 7762 2148
rect 7778 2204 7842 2208
rect 7778 2148 7782 2204
rect 7782 2148 7838 2204
rect 7838 2148 7842 2204
rect 7778 2144 7842 2148
rect 7858 2204 7922 2208
rect 7858 2148 7862 2204
rect 7862 2148 7918 2204
rect 7918 2148 7922 2204
rect 7858 2144 7922 2148
rect 20952 2204 21016 2208
rect 20952 2148 20956 2204
rect 20956 2148 21012 2204
rect 21012 2148 21016 2204
rect 20952 2144 21016 2148
rect 21032 2204 21096 2208
rect 21032 2148 21036 2204
rect 21036 2148 21092 2204
rect 21092 2148 21096 2204
rect 21032 2144 21096 2148
rect 21112 2204 21176 2208
rect 21112 2148 21116 2204
rect 21116 2148 21172 2204
rect 21172 2148 21176 2204
rect 21112 2144 21176 2148
rect 21192 2204 21256 2208
rect 21192 2148 21196 2204
rect 21196 2148 21252 2204
rect 21252 2148 21256 2204
rect 21192 2144 21256 2148
rect 34285 2204 34349 2208
rect 34285 2148 34289 2204
rect 34289 2148 34345 2204
rect 34345 2148 34349 2204
rect 34285 2144 34349 2148
rect 34365 2204 34429 2208
rect 34365 2148 34369 2204
rect 34369 2148 34425 2204
rect 34425 2148 34429 2204
rect 34365 2144 34429 2148
rect 34445 2204 34509 2208
rect 34445 2148 34449 2204
rect 34449 2148 34505 2204
rect 34505 2148 34509 2204
rect 34445 2144 34509 2148
rect 34525 2204 34589 2208
rect 34525 2148 34529 2204
rect 34529 2148 34585 2204
rect 34585 2148 34589 2204
rect 34525 2144 34589 2148
rect 4108 1668 4172 1732
rect 23428 36 23492 100
<< metal4 >>
rect 7610 13088 7931 13648
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7931 13088
rect 7610 12000 7931 13024
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7931 12000
rect 59 11252 125 11253
rect 59 11188 60 11252
rect 124 11188 125 11252
rect 59 11187 125 11188
rect 62 10981 122 11187
rect 59 10980 125 10981
rect 59 10916 60 10980
rect 124 10916 125 10980
rect 59 10915 125 10916
rect 7610 10912 7931 11936
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7931 10912
rect 7610 9824 7931 10848
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7931 9824
rect 7610 8736 7931 9760
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7931 8736
rect 7610 7648 7931 8672
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7931 7648
rect 7610 6560 7931 7584
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7931 6560
rect 7610 5472 7931 6496
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7931 5472
rect 7610 4384 7931 5408
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7931 4384
rect 7610 3296 7931 4320
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7931 3296
rect 4110 1733 4170 2262
rect 7610 2208 7931 3232
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7931 2208
rect 7610 2128 7931 2144
rect 14277 13632 14597 13648
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 12544 14597 13568
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 11456 14597 12480
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 10368 14597 11392
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 9280 14597 10304
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 8192 14597 9216
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 7104 14597 8128
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 6016 14597 7040
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 4928 14597 5952
rect 20944 13088 21264 13648
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 12000 21264 13024
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 10912 21264 11936
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 9824 21264 10848
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 8736 21264 9760
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 7648 21264 8672
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 6560 21264 7584
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 5472 21264 6496
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 14779 5132 14845 5133
rect 14779 5068 14780 5132
rect 14844 5068 14845 5132
rect 14779 5067 14845 5068
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 3840 14597 4864
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 2752 14597 3776
rect 14782 3178 14842 5067
rect 20944 4384 21264 5408
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 3296 21264 4320
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2128 14597 2688
rect 20944 2208 21264 3232
rect 27610 13632 27930 13648
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 12544 27930 13568
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 27610 11456 27930 12480
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 27610 10368 27930 11392
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 9280 27930 10304
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 27610 8192 27930 9216
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 7104 27930 8128
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 6016 27930 7040
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 4928 27930 5952
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 3840 27930 4864
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2128 21264 2144
rect 4107 1732 4173 1733
rect 4107 1668 4108 1732
rect 4172 1668 4173 1732
rect 4107 1667 4173 1668
rect 23430 101 23490 2942
rect 27610 2752 27930 3776
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 27610 2128 27930 2688
rect 34277 13088 34597 13648
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 34277 12000 34597 13024
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 34277 10912 34597 11936
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 34277 9824 34597 10848
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 34277 8736 34597 9760
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 7648 34597 8672
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 6560 34597 7584
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 34277 5472 34597 6496
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 34277 4384 34597 5408
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 34277 3296 34597 4320
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 2208 34597 3232
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 34277 2128 34597 2144
rect 23427 100 23493 101
rect 23427 36 23428 100
rect 23492 36 23493 100
rect 23427 35 23493 36
<< via4 >>
rect 4022 2262 4258 2498
rect 14694 2942 14930 3178
rect 23342 2942 23578 3178
rect 31438 2412 31674 2498
rect 31438 2348 31524 2412
rect 31524 2348 31588 2412
rect 31588 2348 31674 2412
rect 31438 2262 31674 2348
<< metal5 >>
rect 14652 3178 23620 3220
rect 14652 2942 14694 3178
rect 14930 2942 23342 3178
rect 23578 2942 23620 3178
rect 14652 2900 23620 2942
rect 3980 2498 31716 2540
rect 3980 2262 4022 2498
rect 4258 2262 31438 2498
rect 31674 2262 31716 2498
rect 3980 2220 31716 2262
use scs8hd_fill_2  FILLER_0_6 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__047__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_buf_1  _037_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_1_16
timestamp 1586364061
transform 1 0 2576 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_12
timestamp 1586364061
transform 1 0 2208 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_10
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__037__A
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_8  _090_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use scs8hd_inv_8  _047_
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__050__C
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2852 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_32
timestamp 1586364061
transform 1 0 4048 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__050__D
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__051__D
timestamp 1586364061
transform 1 0 4232 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_42 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_1  _045_
timestamp 1586364061
transform 1 0 4232 0 -1 2720
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_1_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3036 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_36
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_41
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_37
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__041__A
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__045__A
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_51
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__050__B
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 1050 592
use scs8hd_inv_8  _041_
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__C
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_55
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_55
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__043__A
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_59
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_43
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_67
timestamp 1586364061
transform 1 0 7268 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_70
timestamp 1586364061
transform 1 0 7544 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_66
timestamp 1586364061
transform 1 0 7176 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__D
timestamp 1586364061
transform 1 0 7360 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__C
timestamp 1586364061
transform 1 0 7084 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__A
timestamp 1586364061
transform 1 0 7452 0 1 2720
box -38 -48 222 592
use scs8hd_buf_1  _043_
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use scs8hd_or4_4  _054_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_80
timestamp 1586364061
transform 1 0 8464 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_84
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_87
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_83
timestamp 1586364061
transform 1 0 8740 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__D
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__B
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__B
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 8648 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9200 0 1 2720
box -38 -48 866 592
use scs8hd_or4_4  _066_
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_97
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_97
timestamp 1586364061
transform 1 0 10028 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_91
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_44
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_1  _055_
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_101
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_101
timestamp 1586364061
transform 1 0 10396 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__055__A
timestamp 1586364061
transform 1 0 10212 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__039__A
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__B
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__D
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_45
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_56
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_123 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12512 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_133
timestamp 1586364061
transform 1 0 13340 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_125 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_137
timestamp 1586364061
transform 1 0 13708 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_140
timestamp 1586364061
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13892 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14076 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 -1 2720
box -38 -48 866 592
use scs8hd_decap_4  FILLER_0_144
timestamp 1586364061
transform 1 0 14352 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_150
timestamp 1586364061
transform 1 0 14904 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_148
timestamp 1586364061
transform 1 0 14720 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_156
timestamp 1586364061
transform 1 0 15456 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 15272 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_46
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_160
timestamp 1586364061
transform 1 0 15824 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_159
timestamp 1586364061
transform 1 0 15732 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__C
timestamp 1586364061
transform 1 0 15640 0 1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16468 0 -1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 16192 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15916 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__D
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_163
timestamp 1586364061
transform 1 0 16100 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_178
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_57
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_47
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use scs8hd_nor4_4  _078_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_1_205
timestamp 1586364061
transform 1 0 19964 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_201
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_204
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_200
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 19688 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__C
timestamp 1586364061
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 19780 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _098_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19964 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_209
timestamp 1586364061
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__C
timestamp 1586364061
transform 1 0 20148 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_8  _086_
timestamp 1586364061
transform 1 0 20332 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_222
timestamp 1586364061
transform 1 0 21528 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_218
timestamp 1586364061
transform 1 0 21160 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_48
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_229
timestamp 1586364061
transform 1 0 22172 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_231
timestamp 1586364061
transform 1 0 22356 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_227
timestamp 1586364061
transform 1 0 21988 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22356 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 21712 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 22172 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21896 0 1 2720
box -38 -48 314 592
use scs8hd_inv_8  _087_
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 866 592
use scs8hd_decap_8  FILLER_1_233 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 22540 0 1 2720
box -38 -48 774 592
use scs8hd_decap_8  FILLER_0_238
timestamp 1586364061
transform 1 0 23000 0 -1 2720
box -38 -48 774 592
use scs8hd_conb_1  _093_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 22724 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_249
timestamp 1586364061
transform 1 0 24012 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_241
timestamp 1586364061
transform 1 0 23276 0 1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_246
timestamp 1586364061
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 23828 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_58
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_49
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25024 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24840 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24196 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_257
timestamp 1586364061
transform 1 0 24748 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_262 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25208 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_253
timestamp 1586364061
transform 1 0 24380 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26588 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_50
timestamp 1586364061
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27048 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_274
timestamp 1586364061
transform 1 0 26312 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_278
timestamp 1586364061
transform 1 0 26680 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_280
timestamp 1586364061
transform 1 0 26864 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_280
timestamp 1586364061
transform 1 0 26864 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_284
timestamp 1586364061
transform 1 0 27232 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_292
timestamp 1586364061
transform 1 0 27968 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_296
timestamp 1586364061
transform 1 0 28336 0 1 2720
box -38 -48 774 592
use scs8hd_fill_1  FILLER_1_304
timestamp 1586364061
transform 1 0 29072 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_304 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 29072 0 -1 2720
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_59
timestamp 1586364061
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_51
timestamp 1586364061
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _113_
timestamp 1586364061
transform 1 0 29716 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_318
timestamp 1586364061
transform 1 0 30360 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_315
timestamp 1586364061
transform 1 0 30084 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 30268 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_306
timestamp 1586364061
transform 1 0 29256 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_319
timestamp 1586364061
transform 1 0 30452 0 -1 2720
box -38 -48 1142 592
use scs8hd_inv_8  _091_
timestamp 1586364061
transform 1 0 31004 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32108 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 30820 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32108 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_331
timestamp 1586364061
transform 1 0 31556 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_1_322
timestamp 1586364061
transform 1 0 30728 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_334
timestamp 1586364061
transform 1 0 31832 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_345
timestamp 1586364061
transform 1 0 32844 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_339
timestamp 1586364061
transform 1 0 32292 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_346
timestamp 1586364061
transform 1 0 32936 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_339
timestamp 1586364061
transform 1 0 32292 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33028 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_52
timestamp 1586364061
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32568 0 1 2720
box -38 -48 314 592
use scs8hd_buf_2  _110_
timestamp 1586364061
transform 1 0 32568 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 33120 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_349
timestamp 1586364061
transform 1 0 33212 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_350
timestamp 1586364061
transform 1 0 33304 0 -1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_53
timestamp 1586364061
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_60
timestamp 1586364061
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_362
timestamp 1586364061
transform 1 0 34408 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_370
timestamp 1586364061
transform 1 0 35144 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_373
timestamp 1586364061
transform 1 0 35420 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_361
timestamp 1586364061
transform 1 0 34316 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_365
timestamp 1586364061
transform 1 0 34684 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_367
timestamp 1586364061
transform 1 0 34868 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_385
timestamp 1586364061
transform 1 0 36524 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_379
timestamp 1586364061
transform 1 0 35972 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_391
timestamp 1586364061
transform 1 0 37076 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 38824 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 38824 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_54
timestamp 1586364061
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_397
timestamp 1586364061
transform 1 0 37628 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_3  FILLER_0_404
timestamp 1586364061
transform 1 0 38272 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_403
timestamp 1586364061
transform 1 0 38180 0 1 2720
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 3808
box -38 -48 866 592
use scs8hd_inv_1  mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__038__A
timestamp 1586364061
transform 1 0 1840 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_6
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_10
timestamp 1586364061
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _050_
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_61
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__052__D
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__050__A
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__052__C
timestamp 1586364061
transform 1 0 5796 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_49
timestamp 1586364061
transform 1 0 5612 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_53
timestamp 1586364061
transform 1 0 5980 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6348 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__042__B
timestamp 1586364061
transform 1 0 7544 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__052__B
timestamp 1586364061
transform 1 0 6164 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 222 592
use scs8hd_or2_4  _081_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8096 0 -1 3808
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__046__B
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__B
timestamp 1586364061
transform 1 0 7912 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_72
timestamp 1586364061
transform 1 0 7728 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_83
timestamp 1586364061
transform 1 0 8740 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_8  _039_
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_62
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__044__C
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_106
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _079_
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__079__C
timestamp 1586364061
transform 1 0 11040 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13340 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_127
timestamp 1586364061
transform 1 0 12788 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_131
timestamp 1586364061
transform 1 0 13156 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _100_
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_63
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 15824 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_144
timestamp 1586364061
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_148
timestamp 1586364061
transform 1 0 14720 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_158
timestamp 1586364061
transform 1 0 15640 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_8  _080_
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__084__B
timestamp 1586364061
transform 1 0 17388 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 16192 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_162
timestamp 1586364061
transform 1 0 16008 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_175
timestamp 1586364061
transform 1 0 17204 0 -1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _085_
timestamp 1586364061
transform 1 0 17940 0 -1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__085__D
timestamp 1586364061
transform 1 0 17756 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_179
timestamp 1586364061
transform 1 0 17572 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_64
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__068__B
timestamp 1586364061
transform 1 0 20424 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__D
timestamp 1586364061
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__C
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_200
timestamp 1586364061
transform 1 0 19504 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_204
timestamp 1586364061
transform 1 0 19872 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_208
timestamp 1586364061
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_212
timestamp 1586364061
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 21344 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__D
timestamp 1586364061
transform 1 0 21712 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_218
timestamp 1586364061
transform 1 0 21160 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_222
timestamp 1586364061
transform 1 0 21528 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_226
timestamp 1586364061
transform 1 0 21896 0 -1 3808
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 23460 0 -1 3808
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_2_238
timestamp 1586364061
transform 1 0 23000 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_242
timestamp 1586364061
transform 1 0 23368 0 -1 3808
box -38 -48 130 592
use scs8hd_conb_1  _095_
timestamp 1586364061
transform 1 0 25208 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24656 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_254
timestamp 1586364061
transform 1 0 24472 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_258
timestamp 1586364061
transform 1 0 24840 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_2_265
timestamp 1586364061
transform 1 0 25484 0 -1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_65
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_273
timestamp 1586364061
transform 1 0 26220 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_288
timestamp 1586364061
transform 1 0 27600 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_300
timestamp 1586364061
transform 1 0 28704 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_312
timestamp 1586364061
transform 1 0 29808 0 -1 3808
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32108 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_66
timestamp 1586364061
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31280 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_324
timestamp 1586364061
transform 1 0 30912 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_6  FILLER_2_330
timestamp 1586364061
transform 1 0 31464 0 -1 3808
box -38 -48 590 592
use scs8hd_decap_12  FILLER_2_346
timestamp 1586364061
transform 1 0 32936 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_358
timestamp 1586364061
transform 1 0 34040 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_370
timestamp 1586364061
transform 1 0 35144 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_382
timestamp 1586364061
transform 1 0 36248 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 38824 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_67
timestamp 1586364061
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_394
timestamp 1586364061
transform 1 0 37352 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_398
timestamp 1586364061
transform 1 0 37720 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_406
timestamp 1586364061
transform 1 0 38456 0 -1 3808
box -38 -48 130 592
use scs8hd_buf_1  _060_
timestamp 1586364061
transform 1 0 1656 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2668 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__060__A
timestamp 1586364061
transform 1 0 2116 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__051__B
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_9
timestamp 1586364061
transform 1 0 1932 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_13
timestamp 1586364061
transform 1 0 2300 0 1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _051_
timestamp 1586364061
transform 1 0 4232 0 1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__048__A
timestamp 1586364061
transform 1 0 3680 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__052__A
timestamp 1586364061
transform 1 0 4048 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_26
timestamp 1586364061
transform 1 0 3496 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_30
timestamp 1586364061
transform 1 0 3864 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__051__C
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_68
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__042__A
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_55
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 406 592
use scs8hd_nor4_4  _046_
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__042__C
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__046__A
timestamp 1586364061
transform 1 0 8832 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__042__D
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_73
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_77
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_81
timestamp 1586364061
transform 1 0 8556 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__044__A
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_103
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_107
timestamp 1586364061
transform 1 0 10948 0 1 3808
box -38 -48 222 592
use scs8hd_buf_1  _064_
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_69
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__044__B
timestamp 1586364061
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 13708 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14076 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_139
timestamp 1586364061
transform 1 0 13892 0 1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _082_
timestamp 1586364061
transform 1 0 15640 0 1 3808
box -38 -48 1602 592
use scs8hd_buf_2  _105_
timestamp 1586364061
transform 1 0 14260 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 14812 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__D
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_151
timestamp 1586364061
transform 1 0 14996 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_155
timestamp 1586364061
transform 1 0 15364 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__084__D
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_175
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _083_
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_70
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__083__D
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _068_
timestamp 1586364061
transform 1 0 20424 0 1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19780 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__B
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_201
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_205
timestamp 1586364061
transform 1 0 19964 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__068__C
timestamp 1586364061
transform 1 0 22172 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_227
timestamp 1586364061
transform 1 0 21988 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_231
timestamp 1586364061
transform 1 0 22356 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_71
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__C
timestamp 1586364061
transform 1 0 22540 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_235
timestamp 1586364061
transform 1 0 22724 0 1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_241
timestamp 1586364061
transform 1 0 23276 0 1 3808
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 25392 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 24840 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 25208 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_256
timestamp 1586364061
transform 1 0 24656 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_260
timestamp 1586364061
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 27140 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26588 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26956 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_275
timestamp 1586364061
transform 1 0 26404 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_279
timestamp 1586364061
transform 1 0 26772 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27600 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_286
timestamp 1586364061
transform 1 0 27416 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_290
timestamp 1586364061
transform 1 0 27784 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_3_302
timestamp 1586364061
transform 1 0 28888 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_72
timestamp 1586364061
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_306
timestamp 1586364061
transform 1 0 29256 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_318
timestamp 1586364061
transform 1 0 30360 0 1 3808
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 31280 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31096 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_337
timestamp 1586364061
transform 1 0 32108 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_349
timestamp 1586364061
transform 1 0 33212 0 1 3808
box -38 -48 1142 592
use scs8hd_buf_2  _108_
timestamp 1586364061
transform 1 0 34868 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 35420 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_361
timestamp 1586364061
transform 1 0 34316 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_365
timestamp 1586364061
transform 1 0 34684 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_371
timestamp 1586364061
transform 1 0 35236 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_375
timestamp 1586364061
transform 1 0 35604 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_387
timestamp 1586364061
transform 1 0 36708 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 38824 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_399
timestamp 1586364061
transform 1 0 37812 0 1 3808
box -38 -48 774 592
use scs8hd_inv_8  _038_
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__058__C
timestamp 1586364061
transform 1 0 2576 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_12
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 406 592
use scs8hd_buf_1  _048_
timestamp 1586364061
transform 1 0 2944 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__051__A
timestamp 1586364061
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__B
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__A
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_18
timestamp 1586364061
transform 1 0 2760 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use scs8hd_nor4_4  _052_
timestamp 1586364061
transform 1 0 4600 0 -1 4896
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_4_36
timestamp 1586364061
transform 1 0 4416 0 -1 4896
box -38 -48 222 592
use scs8hd_or4_4  _042_
timestamp 1586364061
transform 1 0 7452 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6348 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_55
timestamp 1586364061
transform 1 0 6164 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_59
timestamp 1586364061
transform 1 0 6532 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_64
timestamp 1586364061
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__046__D
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__046__C
timestamp 1586364061
transform 1 0 8648 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_78
timestamp 1586364061
transform 1 0 8280 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_88
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use scs8hd_nor4_4  _044_
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__044__D
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_or2_4  _076_
timestamp 1586364061
transform 1 0 11960 0 -1 4896
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 11408 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__B
timestamp 1586364061
transform 1 0 11776 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_110
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_114
timestamp 1586364061
transform 1 0 11592 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 12788 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13248 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_125
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use scs8hd_nor4_4  _084_
timestamp 1586364061
transform 1 0 16928 0 -1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__084__C
timestamp 1586364061
transform 1 0 16744 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_163
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_168
timestamp 1586364061
transform 1 0 16560 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 18676 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 19044 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_189
timestamp 1586364061
transform 1 0 18492 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_193
timestamp 1586364061
transform 1 0 18860 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19228 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__B
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_200
timestamp 1586364061
transform 1 0 19504 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_204
timestamp 1586364061
transform 1 0 19872 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_208
timestamp 1586364061
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_212
timestamp 1586364061
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use scs8hd_nor4_4  _070_
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__072__C
timestamp 1586364061
transform 1 0 22632 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23184 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23644 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_232
timestamp 1586364061
transform 1 0 22448 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_236
timestamp 1586364061
transform 1 0 22816 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_3  FILLER_4_242
timestamp 1586364061
transform 1 0 23368 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_4_247
timestamp 1586364061
transform 1 0 23828 0 -1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 24380 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25576 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_264
timestamp 1586364061
transform 1 0 25392 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25944 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_268
timestamp 1586364061
transform 1 0 25760 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_272
timestamp 1586364061
transform 1 0 26128 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_285
timestamp 1586364061
transform 1 0 27324 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_297
timestamp 1586364061
transform 1 0 28428 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_309
timestamp 1586364061
transform 1 0 29532 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_321
timestamp 1586364061
transform 1 0 30636 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_333
timestamp 1586364061
transform 1 0 31740 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_337
timestamp 1586364061
transform 1 0 32108 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_349
timestamp 1586364061
transform 1 0 33212 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_361
timestamp 1586364061
transform 1 0 34316 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_373
timestamp 1586364061
transform 1 0 35420 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_385
timestamp 1586364061
transform 1 0 36524 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 38824 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_398
timestamp 1586364061
transform 1 0 37720 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_406
timestamp 1586364061
transform 1 0 38456 0 -1 4896
box -38 -48 130 592
use scs8hd_nor4_4  _058_
timestamp 1586364061
transform 1 0 2576 0 1 4896
box -38 -48 1602 592
use scs8hd_buf_2  _106_
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 2300 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_7
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_11
timestamp 1586364061
transform 1 0 2116 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__057__A
timestamp 1586364061
transform 1 0 4324 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_33
timestamp 1586364061
transform 1 0 4140 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _053_
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__053__A
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_37
timestamp 1586364061
transform 1 0 4508 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_41
timestamp 1586364061
transform 1 0 4876 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _065_
timestamp 1586364061
transform 1 0 7544 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__C
timestamp 1586364061
transform 1 0 6992 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__D
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__D
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_66
timestamp 1586364061
transform 1 0 7176 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__C
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__A
timestamp 1586364061
transform 1 0 8648 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_79
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_84
timestamp 1586364061
transform 1 0 8832 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_88
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 222 592
use scs8hd_nor4_4  _059_
timestamp 1586364061
transform 1 0 9568 0 1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__062__C
timestamp 1586364061
transform 1 0 9384 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__B
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__D
timestamp 1586364061
transform 1 0 11684 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_109
timestamp 1586364061
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_113
timestamp 1586364061
transform 1 0 11500 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_117
timestamp 1586364061
transform 1 0 11868 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 14076 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_134
timestamp 1586364061
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_138
timestamp 1586364061
transform 1 0 13800 0 1 4896
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_154
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_160
timestamp 1586364061
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16192 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_175
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _089_
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_193
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 314 592
use scs8hd_nor4_4  _071_
timestamp 1586364061
transform 1 0 20056 0 1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 19872 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__C
timestamp 1586364061
transform 1 0 19504 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_198
timestamp 1586364061
transform 1 0 19320 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_202
timestamp 1586364061
transform 1 0 19688 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 21804 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__B
timestamp 1586364061
transform 1 0 22172 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_223
timestamp 1586364061
transform 1 0 21620 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_227
timestamp 1586364061
transform 1 0 21988 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_231
timestamp 1586364061
transform 1 0 22356 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 24012 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__D
timestamp 1586364061
transform 1 0 22540 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_235
timestamp 1586364061
transform 1 0 22724 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_239
timestamp 1586364061
transform 1 0 23092 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_242
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 24196 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_262
timestamp 1586364061
transform 1 0 25208 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_266
timestamp 1586364061
transform 1 0 25576 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25944 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26956 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25760 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27324 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_279
timestamp 1586364061
transform 1 0 26772 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_283
timestamp 1586364061
transform 1 0 27140 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_287
timestamp 1586364061
transform 1 0 27508 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_5_299
timestamp 1586364061
transform 1 0 28612 0 1 4896
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_306
timestamp 1586364061
transform 1 0 29256 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_318
timestamp 1586364061
transform 1 0 30360 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_330
timestamp 1586364061
transform 1 0 31464 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_342
timestamp 1586364061
transform 1 0 32568 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_354
timestamp 1586364061
transform 1 0 33672 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_367
timestamp 1586364061
transform 1 0 34868 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_379
timestamp 1586364061
transform 1 0 35972 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_391
timestamp 1586364061
transform 1 0 37076 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 38824 0 1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_5_403
timestamp 1586364061
transform 1 0 38180 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_8
timestamp 1586364061
transform 1 0 1840 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_8
timestamp 1586364061
transform 1 0 1840 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__056__D
timestamp 1586364061
transform 1 0 1656 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__056__B
timestamp 1586364061
transform 1 0 1656 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__058__D
timestamp 1586364061
transform 1 0 2024 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__061__A
timestamp 1586364061
transform 1 0 2024 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 5984
box -38 -48 1050 592
use scs8hd_nor4_4  _056_
timestamp 1586364061
transform 1 0 2208 0 1 5984
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__B
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_33
timestamp 1586364061
transform 1 0 4140 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_29
timestamp 1586364061
transform 1 0 3772 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__C
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 3956 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4324 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_nor4_4  _057_
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1602 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 4508 0 1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5796 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5704 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_49
timestamp 1586364061
transform 1 0 5612 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_53
timestamp 1586364061
transform 1 0 5980 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_48
timestamp 1586364061
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_52
timestamp 1586364061
transform 1 0 5888 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_56
timestamp 1586364061
transform 1 0 6256 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_59
timestamp 1586364061
transform 1 0 6532 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6348 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__B
timestamp 1586364061
transform 1 0 6716 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6992 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7176 0 1 5984
box -38 -48 1050 592
use scs8hd_nor4_4  _063_
timestamp 1586364061
transform 1 0 6900 0 -1 5984
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__049__C
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__049__A
timestamp 1586364061
transform 1 0 8648 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_6_88
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_77
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_81
timestamp 1586364061
transform 1 0 8556 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_84
timestamp 1586364061
transform 1 0 8832 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_88
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 222 592
use scs8hd_nor4_4  _049_
timestamp 1586364061
transform 1 0 9568 0 1 5984
box -38 -48 1602 592
use scs8hd_nor4_4  _062_
timestamp 1586364061
transform 1 0 10028 0 -1 5984
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__040__A
timestamp 1586364061
transform 1 0 9384 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__049__D
timestamp 1586364061
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__D
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_113
timestamp 1586364061
transform 1 0 11500 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_109
timestamp 1586364061
transform 1 0 11132 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_114
timestamp 1586364061
transform 1 0 11592 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11684 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11316 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_117
timestamp 1586364061
transform 1 0 11868 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_118
timestamp 1586364061
transform 1 0 11960 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12328 0 -1 5984
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_6_133
timestamp 1586364061
transform 1 0 13340 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_125
timestamp 1586364061
transform 1 0 12604 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13156 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_138
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_134
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 5984
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_160
timestamp 1586364061
transform 1 0 15824 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_156
timestamp 1586364061
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_152
timestamp 1586364061
transform 1 0 15088 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15456 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15272 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 17204 0 -1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16652 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17020 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_167
timestamp 1586364061
transform 1 0 16468 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_171
timestamp 1586364061
transform 1 0 16836 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18400 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_186
timestamp 1586364061
transform 1 0 18216 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_193
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_203
timestamp 1586364061
transform 1 0 19780 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__073__B
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 19964 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  _067_
timestamp 1586364061
transform 1 0 19780 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_210
timestamp 1586364061
transform 1 0 20424 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_206
timestamp 1586364061
transform 1 0 20056 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__D
timestamp 1586364061
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__C
timestamp 1586364061
transform 1 0 20240 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_nor4_4  _073_
timestamp 1586364061
transform 1 0 20148 0 1 5984
box -38 -48 1602 592
use scs8hd_nor4_4  _072_
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__074__B
timestamp 1586364061
transform 1 0 21896 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__D
timestamp 1586364061
transform 1 0 22264 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_224
timestamp 1586364061
transform 1 0 21712 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_228
timestamp 1586364061
transform 1 0 22080 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_240
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_236
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_232
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_232
timestamp 1586364061
transform 1 0 22448 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__074__C
timestamp 1586364061
transform 1 0 22632 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 23184 0 -1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_7_256
timestamp 1586364061
transform 1 0 24656 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24748 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24840 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_260
timestamp 1586364061
transform 1 0 25024 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_266
timestamp 1586364061
transform 1 0 25576 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_6_262
timestamp 1586364061
transform 1 0 25208 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25392 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25208 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24932 0 -1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25392 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26956 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26496 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_272
timestamp 1586364061
transform 1 0 26128 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_285
timestamp 1586364061
transform 1 0 27324 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_273
timestamp 1586364061
transform 1 0 26220 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_278
timestamp 1586364061
transform 1 0 26680 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27968 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27508 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_289
timestamp 1586364061
transform 1 0 27692 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_301
timestamp 1586364061
transform 1 0 28796 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_290
timestamp 1586364061
transform 1 0 27784 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_294
timestamp 1586364061
transform 1 0 28152 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_302
timestamp 1586364061
transform 1 0 28888 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_313
timestamp 1586364061
transform 1 0 29900 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_306
timestamp 1586364061
transform 1 0 29256 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_318
timestamp 1586364061
transform 1 0 30360 0 1 5984
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31464 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31924 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_325
timestamp 1586364061
transform 1 0 31004 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_6_333
timestamp 1586364061
transform 1 0 31740 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_337
timestamp 1586364061
transform 1 0 32108 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_333
timestamp 1586364061
transform 1 0 31740 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_337
timestamp 1586364061
transform 1 0 32108 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_349
timestamp 1586364061
transform 1 0 33212 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_349
timestamp 1586364061
transform 1 0 33212 0 1 5984
box -38 -48 1142 592
use scs8hd_buf_2  _099_
timestamp 1586364061
transform 1 0 35420 0 1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34592 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_361
timestamp 1586364061
transform 1 0 34316 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_373
timestamp 1586364061
transform 1 0 35420 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_7_361
timestamp 1586364061
transform 1 0 34316 0 1 5984
box -38 -48 314 592
use scs8hd_decap_6  FILLER_7_367
timestamp 1586364061
transform 1 0 34868 0 1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 35972 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_385
timestamp 1586364061
transform 1 0 36524 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_377
timestamp 1586364061
transform 1 0 35788 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_381
timestamp 1586364061
transform 1 0 36156 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 38824 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 38824 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_398
timestamp 1586364061
transform 1 0 37720 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_406
timestamp 1586364061
transform 1 0 38456 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_393
timestamp 1586364061
transform 1 0 37260 0 1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_405
timestamp 1586364061
transform 1 0 38364 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  _061_
timestamp 1586364061
transform 1 0 2576 0 -1 7072
box -38 -48 314 592
use scs8hd_conb_1  _097_
timestamp 1586364061
transform 1 0 1564 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__056__A
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_8
timestamp 1586364061
transform 1 0 1840 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_14
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__056__C
timestamp 1586364061
transform 1 0 3036 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_19
timestamp 1586364061
transform 1 0 2852 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4600 0 -1 7072
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_8_36
timestamp 1586364061
transform 1 0 4416 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_49
timestamp 1586364061
transform 1 0 5612 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6532 0 -1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_57
timestamp 1586364061
transform 1 0 6348 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_62
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_66
timestamp 1586364061
transform 1 0 7176 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_79
timestamp 1586364061
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_83
timestamp 1586364061
transform 1 0 8740 0 -1 7072
box -38 -48 774 592
use scs8hd_buf_1  _040_
timestamp 1586364061
transform 1 0 9752 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__049__B
timestamp 1586364061
transform 1 0 10212 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_91
timestamp 1586364061
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_97
timestamp 1586364061
transform 1 0 10028 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_101
timestamp 1586364061
transform 1 0 10396 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  FILLER_8_107
timestamp 1586364061
transform 1 0 10948 0 -1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_121
timestamp 1586364061
transform 1 0 12236 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12788 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_125
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_138
timestamp 1586364061
transform 1 0 13800 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_142
timestamp 1586364061
transform 1 0 14168 0 -1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17388 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_163
timestamp 1586364061
transform 1 0 16100 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_168
timestamp 1586364061
transform 1 0 16560 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_176
timestamp 1586364061
transform 1 0 17296 0 -1 7072
box -38 -48 130 592
use scs8hd_conb_1  _096_
timestamp 1586364061
transform 1 0 18952 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18400 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_186
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 20148 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__D
timestamp 1586364061
transform 1 0 20516 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_197
timestamp 1586364061
transform 1 0 19228 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_205
timestamp 1586364061
transform 1 0 19964 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_209
timestamp 1586364061
transform 1 0 20332 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_213
timestamp 1586364061
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use scs8hd_nor4_4  _074_
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1602 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23736 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_232
timestamp 1586364061
transform 1 0 22448 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_8_244
timestamp 1586364061
transform 1 0 23552 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_249
timestamp 1586364061
transform 1 0 24012 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_253
timestamp 1586364061
transform 1 0 24380 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_257
timestamp 1586364061
transform 1 0 24748 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_267
timestamp 1586364061
transform 1 0 25668 0 -1 7072
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_285
timestamp 1586364061
transform 1 0 27324 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_297
timestamp 1586364061
transform 1 0 28428 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_309
timestamp 1586364061
transform 1 0 29532 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_321
timestamp 1586364061
transform 1 0 30636 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_333
timestamp 1586364061
transform 1 0 31740 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_337
timestamp 1586364061
transform 1 0 32108 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_349
timestamp 1586364061
transform 1 0 33212 0 -1 7072
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34592 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_361
timestamp 1586364061
transform 1 0 34316 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_367
timestamp 1586364061
transform 1 0 34868 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_379
timestamp 1586364061
transform 1 0 35972 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_8_391
timestamp 1586364061
transform 1 0 37076 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 38824 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_398
timestamp 1586364061
transform 1 0 37720 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_406
timestamp 1586364061
transform 1 0 38456 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_2  _104_
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_7
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_11
timestamp 1586364061
transform 1 0 2116 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_16
timestamp 1586364061
transform 1 0 2576 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2944 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2760 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_29
timestamp 1586364061
transform 1 0 3772 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_35
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7544 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7176 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_68
timestamp 1586364061
transform 1 0 7360 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_79
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_83
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 9568 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_91
timestamp 1586364061
transform 1 0 9476 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_97
timestamp 1586364061
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_101
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_132
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_136
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15548 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14444 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_143
timestamp 1586364061
transform 1 0 14260 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_155
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_160
timestamp 1586364061
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16652 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_164
timestamp 1586364061
transform 1 0 16192 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_168
timestamp 1586364061
transform 1 0 16560 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_171
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_inv_8  _088_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_193
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_205
timestamp 1586364061
transform 1 0 19964 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_217
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_229
timestamp 1586364061
transform 1 0 22172 0 1 7072
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23920 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_9_241
timestamp 1586364061
transform 1 0 23276 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24932 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_251
timestamp 1586364061
transform 1 0 24196 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_268
timestamp 1586364061
transform 1 0 25760 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_280
timestamp 1586364061
transform 1 0 26864 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_292
timestamp 1586364061
transform 1 0 27968 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_304
timestamp 1586364061
transform 1 0 29072 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_306
timestamp 1586364061
transform 1 0 29256 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_318
timestamp 1586364061
transform 1 0 30360 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 32108 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_330
timestamp 1586364061
transform 1 0 31464 0 1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_9_336
timestamp 1586364061
transform 1 0 32016 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_339
timestamp 1586364061
transform 1 0 32292 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_351
timestamp 1586364061
transform 1 0 33396 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_9_363
timestamp 1586364061
transform 1 0 34500 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_367
timestamp 1586364061
transform 1 0 34868 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_379
timestamp 1586364061
transform 1 0 35972 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_391
timestamp 1586364061
transform 1 0 37076 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 38824 0 1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_9_403
timestamp 1586364061
transform 1 0 38180 0 1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_6
timestamp 1586364061
transform 1 0 1656 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_10
timestamp 1586364061
transform 1 0 2024 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_16
timestamp 1586364061
transform 1 0 2576 0 -1 8160
box -38 -48 222 592
use scs8hd_conb_1  _094_
timestamp 1586364061
transform 1 0 2760 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_21
timestamp 1586364061
transform 1 0 3036 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_25
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_4  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4508 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5520 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_36
timestamp 1586364061
transform 1 0 4416 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_46
timestamp 1586364061
transform 1 0 5336 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_50
timestamp 1586364061
transform 1 0 5704 0 -1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7176 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_62
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_69
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_1  _075_
timestamp 1586364061
transform 1 0 8556 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_73
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_77
timestamp 1586364061
transform 1 0 8188 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_8  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use scs8hd_buf_1  _077_
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_96
timestamp 1586364061
transform 1 0 9936 0 -1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12236 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_108
timestamp 1586364061
transform 1 0 11040 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_113
timestamp 1586364061
transform 1 0 11500 0 -1 8160
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13800 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13248 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_130
timestamp 1586364061
transform 1 0 13064 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_134
timestamp 1586364061
transform 1 0 13432 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_141
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use scs8hd_conb_1  _092_
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_157
timestamp 1586364061
transform 1 0 15548 0 -1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16652 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_172
timestamp 1586364061
transform 1 0 16928 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_184
timestamp 1586364061
transform 1 0 18032 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_196
timestamp 1586364061
transform 1 0 19136 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_6  FILLER_10_208
timestamp 1586364061
transform 1 0 20240 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23920 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_247
timestamp 1586364061
transform 1 0 23828 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25024 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25392 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_250
timestamp 1586364061
transform 1 0 24104 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_254
timestamp 1586364061
transform 1 0 24472 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_258
timestamp 1586364061
transform 1 0 24840 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_262
timestamp 1586364061
transform 1 0 25208 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_266
timestamp 1586364061
transform 1 0 25576 0 -1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_274
timestamp 1586364061
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_288
timestamp 1586364061
transform 1 0 27600 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_300
timestamp 1586364061
transform 1 0 28704 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_312
timestamp 1586364061
transform 1 0 29808 0 -1 8160
box -38 -48 1142 592
use scs8hd_buf_2  _101_
timestamp 1586364061
transform 1 0 32108 0 -1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_324
timestamp 1586364061
transform 1 0 30912 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_341
timestamp 1586364061
transform 1 0 32476 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_353
timestamp 1586364061
transform 1 0 33580 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_365
timestamp 1586364061
transform 1 0 34684 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_377
timestamp 1586364061
transform 1 0 35788 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_389
timestamp 1586364061
transform 1 0 36892 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 38824 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_398
timestamp 1586364061
transform 1 0 37720 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_406
timestamp 1586364061
transform 1 0 38456 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_19
timestamp 1586364061
transform 1 0 2852 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_31
timestamp 1586364061
transform 1 0 3956 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_43
timestamp 1586364061
transform 1 0 5060 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_decap_6  FILLER_11_55
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 590 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use scs8hd_buf_1  _069_
timestamp 1586364061
transform 1 0 10304 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_98
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_103
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_107
timestamp 1586364061
transform 1 0 10948 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_120
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_126
timestamp 1586364061
transform 1 0 12696 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_130
timestamp 1586364061
transform 1 0 13064 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_142
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_11_154
timestamp 1586364061
transform 1 0 15272 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_160
timestamp 1586364061
transform 1 0 15824 0 1 8160
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15916 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16376 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_164
timestamp 1586364061
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_168
timestamp 1586364061
transform 1 0 16560 0 1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_180
timestamp 1586364061
transform 1 0 17664 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_187
timestamp 1586364061
transform 1 0 18308 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_191
timestamp 1586364061
transform 1 0 18676 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_203
timestamp 1586364061
transform 1 0 19780 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_215
timestamp 1586364061
transform 1 0 20884 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_227
timestamp 1586364061
transform 1 0 21988 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_11_239
timestamp 1586364061
transform 1 0 23092 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_243
timestamp 1586364061
transform 1 0 23460 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_281
timestamp 1586364061
transform 1 0 26956 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_293
timestamp 1586364061
transform 1 0 28060 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_306
timestamp 1586364061
transform 1 0 29256 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_318
timestamp 1586364061
transform 1 0 30360 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_330
timestamp 1586364061
transform 1 0 31464 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_342
timestamp 1586364061
transform 1 0 32568 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_354
timestamp 1586364061
transform 1 0 33672 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 35420 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_367
timestamp 1586364061
transform 1 0 34868 0 1 8160
box -38 -48 590 592
use scs8hd_decap_12  FILLER_11_375
timestamp 1586364061
transform 1 0 35604 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_387
timestamp 1586364061
transform 1 0 36708 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 38824 0 1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_11_399
timestamp 1586364061
transform 1 0 37812 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11960 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_121
timestamp 1586364061
transform 1 0 12236 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_133
timestamp 1586364061
transform 1 0 13340 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_166
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_178
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_190
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_202
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_263
timestamp 1586364061
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_288
timestamp 1586364061
transform 1 0 27600 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_300
timestamp 1586364061
transform 1 0 28704 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_312
timestamp 1586364061
transform 1 0 29808 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_324
timestamp 1586364061
transform 1 0 30912 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_337
timestamp 1586364061
transform 1 0 32108 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_349
timestamp 1586364061
transform 1 0 33212 0 -1 9248
box -38 -48 1142 592
use scs8hd_buf_2  _115_
timestamp 1586364061
transform 1 0 35420 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_361
timestamp 1586364061
transform 1 0 34316 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_377
timestamp 1586364061
transform 1 0 35788 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_12_389
timestamp 1586364061
transform 1 0 36892 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 38824 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_398
timestamp 1586364061
transform 1 0 37720 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_406
timestamp 1586364061
transform 1 0 38456 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_98
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_110
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_117
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_129
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_147
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_159
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_171
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_178
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_196
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_202
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_281
timestamp 1586364061
transform 1 0 26956 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_293
timestamp 1586364061
transform 1 0 28060 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_288
timestamp 1586364061
transform 1 0 27600 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_300
timestamp 1586364061
transform 1 0 28704 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_306
timestamp 1586364061
transform 1 0 29256 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_318
timestamp 1586364061
transform 1 0 30360 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_312
timestamp 1586364061
transform 1 0 29808 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_330
timestamp 1586364061
transform 1 0 31464 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_324
timestamp 1586364061
transform 1 0 30912 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_337
timestamp 1586364061
transform 1 0 32108 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_342
timestamp 1586364061
transform 1 0 32568 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_354
timestamp 1586364061
transform 1 0 33672 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_349
timestamp 1586364061
transform 1 0 33212 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_367
timestamp 1586364061
transform 1 0 34868 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_361
timestamp 1586364061
transform 1 0 34316 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_373
timestamp 1586364061
transform 1 0 35420 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_379
timestamp 1586364061
transform 1 0 35972 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_391
timestamp 1586364061
transform 1 0 37076 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_385
timestamp 1586364061
transform 1 0 36524 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 38824 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 38824 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_403
timestamp 1586364061
transform 1 0 38180 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_398
timestamp 1586364061
transform 1 0 37720 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_406
timestamp 1586364061
transform 1 0 38456 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_110
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_159
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_220
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_281
timestamp 1586364061
transform 1 0 26956 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_293
timestamp 1586364061
transform 1 0 28060 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_306
timestamp 1586364061
transform 1 0 29256 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_318
timestamp 1586364061
transform 1 0 30360 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_330
timestamp 1586364061
transform 1 0 31464 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_342
timestamp 1586364061
transform 1 0 32568 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_354
timestamp 1586364061
transform 1 0 33672 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 35420 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_367
timestamp 1586364061
transform 1 0 34868 0 1 10336
box -38 -48 590 592
use scs8hd_decap_12  FILLER_15_375
timestamp 1586364061
transform 1 0 35604 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_387
timestamp 1586364061
transform 1 0 36708 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 38824 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_399
timestamp 1586364061
transform 1 0 37812 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_117
timestamp 1586364061
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_129
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_166
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_178
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_190
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_202
timestamp 1586364061
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_288
timestamp 1586364061
transform 1 0 27600 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_300
timestamp 1586364061
transform 1 0 28704 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_312
timestamp 1586364061
transform 1 0 29808 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_324
timestamp 1586364061
transform 1 0 30912 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_337
timestamp 1586364061
transform 1 0 32108 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_349
timestamp 1586364061
transform 1 0 33212 0 -1 11424
box -38 -48 1142 592
use scs8hd_buf_2  _112_
timestamp 1586364061
transform 1 0 35420 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_361
timestamp 1586364061
transform 1 0 34316 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_377
timestamp 1586364061
transform 1 0 35788 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_389
timestamp 1586364061
transform 1 0 36892 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 38824 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_398
timestamp 1586364061
transform 1 0 37720 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_406
timestamp 1586364061
transform 1 0 38456 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use scs8hd_buf_2  _114_
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 7360 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_66
timestamp 1586364061
transform 1 0 7176 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_70
timestamp 1586364061
transform 1 0 7544 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_82
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_94
timestamp 1586364061
transform 1 0 9752 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_106
timestamp 1586364061
transform 1 0 10856 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_147
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_159
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_171
timestamp 1586364061
transform 1 0 16836 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 19320 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_200
timestamp 1586364061
transform 1 0 19504 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_212
timestamp 1586364061
transform 1 0 20608 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_224
timestamp 1586364061
transform 1 0 21712 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_17_236
timestamp 1586364061
transform 1 0 22816 0 1 11424
box -38 -48 774 592
use scs8hd_decap_12  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_281
timestamp 1586364061
transform 1 0 26956 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_293
timestamp 1586364061
transform 1 0 28060 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_306
timestamp 1586364061
transform 1 0 29256 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_318
timestamp 1586364061
transform 1 0 30360 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_330
timestamp 1586364061
transform 1 0 31464 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_342
timestamp 1586364061
transform 1 0 32568 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_354
timestamp 1586364061
transform 1 0 33672 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_367
timestamp 1586364061
transform 1 0 34868 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_379
timestamp 1586364061
transform 1 0 35972 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_391
timestamp 1586364061
transform 1 0 37076 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 38824 0 1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_17_403
timestamp 1586364061
transform 1 0 38180 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_117
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_129
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 774 592
use scs8hd_buf_2  _109_
timestamp 1586364061
transform 1 0 19320 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_288
timestamp 1586364061
transform 1 0 27600 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_300
timestamp 1586364061
transform 1 0 28704 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_312
timestamp 1586364061
transform 1 0 29808 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_324
timestamp 1586364061
transform 1 0 30912 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_337
timestamp 1586364061
transform 1 0 32108 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_349
timestamp 1586364061
transform 1 0 33212 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_361
timestamp 1586364061
transform 1 0 34316 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_373
timestamp 1586364061
transform 1 0 35420 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_385
timestamp 1586364061
transform 1 0 36524 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 38824 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_398
timestamp 1586364061
transform 1 0 37720 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_406
timestamp 1586364061
transform 1 0 38456 0 -1 12512
box -38 -48 130 592
use scs8hd_buf_2  _111_
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 1932 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_11
timestamp 1586364061
transform 1 0 2116 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_23
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_35
timestamp 1586364061
transform 1 0 4324 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_47
timestamp 1586364061
transform 1 0 5428 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_63
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_75
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_87
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_94
timestamp 1586364061
transform 1 0 9752 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_118
timestamp 1586364061
transform 1 0 11960 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_137
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 15364 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_156
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_171
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_168
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_180
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_187
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_199
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_211
timestamp 1586364061
transform 1 0 20516 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_218
timestamp 1586364061
transform 1 0 21160 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_230
timestamp 1586364061
transform 1 0 22264 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_2  _103_
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 23920 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_19_249
timestamp 1586364061
transform 1 0 24012 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_242
timestamp 1586364061
transform 1 0 23368 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_249
timestamp 1586364061
transform 1 0 24012 0 -1 13600
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 24196 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_253
timestamp 1586364061
transform 1 0 24380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_265
timestamp 1586364061
transform 1 0 25484 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_261
timestamp 1586364061
transform 1 0 25116 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_2  _102_
timestamp 1586364061
transform 1 0 26220 0 1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 26772 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 26772 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_277
timestamp 1586364061
transform 1 0 26588 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_281
timestamp 1586364061
transform 1 0 26956 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_273
timestamp 1586364061
transform 1 0 26220 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_280
timestamp 1586364061
transform 1 0 26864 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_293
timestamp 1586364061
transform 1 0 28060 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_292
timestamp 1586364061
transform 1 0 27968 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 29624 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_306
timestamp 1586364061
transform 1 0 29256 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_318
timestamp 1586364061
transform 1 0 30360 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_304
timestamp 1586364061
transform 1 0 29072 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_311
timestamp 1586364061
transform 1 0 29716 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_330
timestamp 1586364061
transform 1 0 31464 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_323
timestamp 1586364061
transform 1 0 30820 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_335
timestamp 1586364061
transform 1 0 31924 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 32476 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_342
timestamp 1586364061
transform 1 0 32568 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_354
timestamp 1586364061
transform 1 0 33672 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_342
timestamp 1586364061
transform 1 0 32568 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_354
timestamp 1586364061
transform 1 0 33672 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_2  _107_
timestamp 1586364061
transform 1 0 35420 0 1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 35328 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_19_367
timestamp 1586364061
transform 1 0 34868 0 1 12512
box -38 -48 590 592
use scs8hd_decap_6  FILLER_20_366
timestamp 1586364061
transform 1 0 34776 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_373
timestamp 1586364061
transform 1 0 35420 0 -1 13600
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 35972 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_377
timestamp 1586364061
transform 1 0 35788 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_381
timestamp 1586364061
transform 1 0 36156 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_385
timestamp 1586364061
transform 1 0 36524 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 38824 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 38824 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 38180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_393
timestamp 1586364061
transform 1 0 37260 0 1 12512
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_19_405
timestamp 1586364061
transform 1 0 38364 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_397
timestamp 1586364061
transform 1 0 37628 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_3  FILLER_20_404
timestamp 1586364061
transform 1 0 38272 0 -1 13600
box -38 -48 314 592
<< labels >>
rlabel metal2 s 5814 0 5870 480 6 address[0]
port 0 nsew default input
rlabel metal3 s 0 552 480 672 6 address[1]
port 1 nsew default input
rlabel metal2 s 2226 15520 2282 16000 6 address[2]
port 2 nsew default input
rlabel metal3 s 0 1776 480 1896 6 address[3]
port 3 nsew default input
rlabel metal2 s 6642 15520 6698 16000 6 address[4]
port 4 nsew default input
rlabel metal3 s 39520 552 40000 672 6 address[5]
port 5 nsew default input
rlabel metal3 s 39520 1776 40000 1896 6 bottom_grid_pin_0_
port 6 nsew default tristate
rlabel metal2 s 11058 15520 11114 16000 6 bottom_grid_pin_4_
port 7 nsew default tristate
rlabel metal3 s 0 3136 480 3256 6 bottom_grid_pin_8_
port 8 nsew default tristate
rlabel metal2 s 8114 0 8170 480 6 chanx_left_in[0]
port 9 nsew default input
rlabel metal2 s 10506 0 10562 480 6 chanx_left_in[1]
port 10 nsew default input
rlabel metal2 s 12806 0 12862 480 6 chanx_left_in[2]
port 11 nsew default input
rlabel metal2 s 15566 15520 15622 16000 6 chanx_left_in[3]
port 12 nsew default input
rlabel metal3 s 0 4496 480 4616 6 chanx_left_in[4]
port 13 nsew default input
rlabel metal3 s 39520 3136 40000 3256 6 chanx_left_in[5]
port 14 nsew default input
rlabel metal2 s 19982 15520 20038 16000 6 chanx_left_in[6]
port 15 nsew default input
rlabel metal3 s 39520 4496 40000 4616 6 chanx_left_in[7]
port 16 nsew default input
rlabel metal2 s 15198 0 15254 480 6 chanx_left_in[8]
port 17 nsew default input
rlabel metal3 s 0 5856 480 5976 6 chanx_left_out[0]
port 18 nsew default tristate
rlabel metal2 s 17590 0 17646 480 6 chanx_left_out[1]
port 19 nsew default tristate
rlabel metal3 s 0 7216 480 7336 6 chanx_left_out[2]
port 20 nsew default tristate
rlabel metal2 s 24398 15520 24454 16000 6 chanx_left_out[3]
port 21 nsew default tristate
rlabel metal2 s 28906 15520 28962 16000 6 chanx_left_out[4]
port 22 nsew default tristate
rlabel metal2 s 33322 15520 33378 16000 6 chanx_left_out[5]
port 23 nsew default tristate
rlabel metal2 s 19890 0 19946 480 6 chanx_left_out[6]
port 24 nsew default tristate
rlabel metal3 s 39520 5856 40000 5976 6 chanx_left_out[7]
port 25 nsew default tristate
rlabel metal2 s 22282 0 22338 480 6 chanx_left_out[8]
port 26 nsew default tristate
rlabel metal2 s 24582 0 24638 480 6 chanx_right_in[0]
port 27 nsew default input
rlabel metal3 s 0 8576 480 8696 6 chanx_right_in[1]
port 28 nsew default input
rlabel metal3 s 0 9800 480 9920 6 chanx_right_in[2]
port 29 nsew default input
rlabel metal2 s 37738 15520 37794 16000 6 chanx_right_in[3]
port 30 nsew default input
rlabel metal2 s 26974 0 27030 480 6 chanx_right_in[4]
port 31 nsew default input
rlabel metal3 s 39520 7216 40000 7336 6 chanx_right_in[5]
port 32 nsew default input
rlabel metal3 s 0 11160 480 11280 6 chanx_right_in[6]
port 33 nsew default input
rlabel metal3 s 39520 8576 40000 8696 6 chanx_right_in[7]
port 34 nsew default input
rlabel metal2 s 29366 0 29422 480 6 chanx_right_in[8]
port 35 nsew default input
rlabel metal3 s 39520 9800 40000 9920 6 chanx_right_out[0]
port 36 nsew default tristate
rlabel metal3 s 0 12520 480 12640 6 chanx_right_out[1]
port 37 nsew default tristate
rlabel metal2 s 31666 0 31722 480 6 chanx_right_out[2]
port 38 nsew default tristate
rlabel metal3 s 39520 11160 40000 11280 6 chanx_right_out[3]
port 39 nsew default tristate
rlabel metal3 s 0 13880 480 14000 6 chanx_right_out[4]
port 40 nsew default tristate
rlabel metal2 s 34058 0 34114 480 6 chanx_right_out[5]
port 41 nsew default tristate
rlabel metal3 s 39520 12520 40000 12640 6 chanx_right_out[6]
port 42 nsew default tristate
rlabel metal2 s 36358 0 36414 480 6 chanx_right_out[7]
port 43 nsew default tristate
rlabel metal3 s 39520 13880 40000 14000 6 chanx_right_out[8]
port 44 nsew default tristate
rlabel metal2 s 3422 0 3478 480 6 data_in
port 45 nsew default input
rlabel metal2 s 1122 0 1178 480 6 enable
port 46 nsew default input
rlabel metal3 s 0 15240 480 15360 6 top_grid_pin_14_
port 47 nsew default tristate
rlabel metal3 s 39520 15240 40000 15360 6 top_grid_pin_2_
port 48 nsew default tristate
rlabel metal2 s 38750 0 38806 480 6 top_grid_pin_6_
port 49 nsew default tristate
rlabel metal4 s 7611 2128 7931 13648 6 vpwr
port 50 nsew default input
rlabel metal4 s 14277 2128 14597 13648 6 vgnd
port 51 nsew default input
<< end >>
