magic
tech sky130A
magscale 1 2
timestamp 1606236403
<< viali >>
rect 11751 4641 11785 4675
rect 12119 4641 12153 4675
rect 12211 4437 12245 4471
rect 12763 3689 12797 3723
rect 8690 3553 8724 3587
rect 11650 3553 11684 3587
rect 11383 3485 11417 3519
rect 8761 3349 8795 3383
rect 7795 3009 7829 3043
rect 6415 2941 6449 2975
rect 7887 2873 7921 2907
rect 8807 2873 8841 2907
rect 6599 2805 6633 2839
rect 6691 2533 6725 2567
rect 7611 2533 7645 2567
rect 6599 2397 6633 2431
<< metal1 >>
rect 38 6554 14758 6576
rect 38 6502 2381 6554
rect 2433 6502 2445 6554
rect 2497 6502 2509 6554
rect 2561 6502 2573 6554
rect 2625 6502 7312 6554
rect 7364 6502 7376 6554
rect 7428 6502 7440 6554
rect 7492 6502 7504 6554
rect 7556 6502 12242 6554
rect 12294 6502 12306 6554
rect 12358 6502 12370 6554
rect 12422 6502 12434 6554
rect 12486 6502 14758 6554
rect 38 6480 14758 6502
rect 38 6010 14758 6032
rect 38 5958 4846 6010
rect 4898 5958 4910 6010
rect 4962 5958 4974 6010
rect 5026 5958 5038 6010
rect 5090 5958 9777 6010
rect 9829 5958 9841 6010
rect 9893 5958 9905 6010
rect 9957 5958 9969 6010
rect 10021 5958 14758 6010
rect 38 5936 14758 5958
rect 38 5466 14758 5488
rect 38 5414 2381 5466
rect 2433 5414 2445 5466
rect 2497 5414 2509 5466
rect 2561 5414 2573 5466
rect 2625 5414 7312 5466
rect 7364 5414 7376 5466
rect 7428 5414 7440 5466
rect 7492 5414 7504 5466
rect 7556 5414 12242 5466
rect 12294 5414 12306 5466
rect 12358 5414 12370 5466
rect 12422 5414 12434 5466
rect 12486 5414 14758 5466
rect 38 5392 14758 5414
rect 38 4922 14758 4944
rect 38 4870 4846 4922
rect 4898 4870 4910 4922
rect 4962 4870 4974 4922
rect 5026 4870 5038 4922
rect 5090 4870 9777 4922
rect 9829 4870 9841 4922
rect 9893 4870 9905 4922
rect 9957 4870 9969 4922
rect 10021 4870 14758 4922
rect 38 4848 14758 4870
rect 11736 4672 11742 4684
rect 11697 4644 11742 4672
rect 11736 4632 11742 4644
rect 11794 4632 11800 4684
rect 12104 4672 12110 4684
rect 12065 4644 12110 4672
rect 12104 4632 12110 4644
rect 12162 4632 12168 4684
rect 11460 4428 11466 4480
rect 11518 4468 11524 4480
rect 12199 4471 12257 4477
rect 12199 4468 12211 4471
rect 11518 4440 12211 4468
rect 11518 4428 11524 4440
rect 12199 4437 12211 4440
rect 12245 4437 12257 4471
rect 12199 4431 12257 4437
rect 38 4378 14758 4400
rect 38 4326 2381 4378
rect 2433 4326 2445 4378
rect 2497 4326 2509 4378
rect 2561 4326 2573 4378
rect 2625 4326 7312 4378
rect 7364 4326 7376 4378
rect 7428 4326 7440 4378
rect 7492 4326 7504 4378
rect 7556 4326 12242 4378
rect 12294 4326 12306 4378
rect 12358 4326 12370 4378
rect 12422 4326 12434 4378
rect 12486 4326 14758 4378
rect 38 4304 14758 4326
rect 38 3834 14758 3856
rect 38 3782 4846 3834
rect 4898 3782 4910 3834
rect 4962 3782 4974 3834
rect 5026 3782 5038 3834
rect 5090 3782 9777 3834
rect 9829 3782 9841 3834
rect 9893 3782 9905 3834
rect 9957 3782 9969 3834
rect 10021 3782 14758 3834
rect 38 3760 14758 3782
rect 12104 3680 12110 3732
rect 12162 3720 12168 3732
rect 12751 3723 12809 3729
rect 12751 3720 12763 3723
rect 12162 3692 12763 3720
rect 12162 3680 12168 3692
rect 12751 3689 12763 3692
rect 12797 3689 12809 3723
rect 12751 3683 12809 3689
rect 7780 3544 7786 3596
rect 7838 3584 7844 3596
rect 8678 3587 8736 3593
rect 8678 3584 8690 3587
rect 7838 3556 8690 3584
rect 7838 3544 7844 3556
rect 8678 3553 8690 3556
rect 8724 3584 8736 3587
rect 10816 3584 10822 3596
rect 8724 3556 10822 3584
rect 8724 3553 8736 3556
rect 8678 3547 8736 3553
rect 10816 3544 10822 3556
rect 10874 3584 10880 3596
rect 11460 3584 11466 3596
rect 10874 3556 11466 3584
rect 10874 3544 10880 3556
rect 11460 3544 11466 3556
rect 11518 3544 11524 3596
rect 11638 3587 11696 3593
rect 11638 3553 11650 3587
rect 11684 3584 11696 3587
rect 12656 3584 12662 3596
rect 11684 3556 12662 3584
rect 11684 3553 11696 3556
rect 11638 3547 11696 3553
rect 12656 3544 12662 3556
rect 12714 3544 12720 3596
rect 11368 3516 11374 3528
rect 11329 3488 11374 3516
rect 11368 3476 11374 3488
rect 11426 3476 11432 3528
rect 7872 3340 7878 3392
rect 7930 3380 7936 3392
rect 8749 3383 8807 3389
rect 8749 3380 8761 3383
rect 7930 3352 8761 3380
rect 7930 3340 7936 3352
rect 8749 3349 8761 3352
rect 8795 3349 8807 3383
rect 8749 3343 8807 3349
rect 38 3290 14758 3312
rect 38 3238 2381 3290
rect 2433 3238 2445 3290
rect 2497 3238 2509 3290
rect 2561 3238 2573 3290
rect 2625 3238 7312 3290
rect 7364 3238 7376 3290
rect 7428 3238 7440 3290
rect 7492 3238 7504 3290
rect 7556 3238 12242 3290
rect 12294 3238 12306 3290
rect 12358 3238 12370 3290
rect 12422 3238 12434 3290
rect 12486 3238 14758 3290
rect 38 3216 14758 3238
rect 7783 3043 7841 3049
rect 7783 3009 7795 3043
rect 7829 3040 7841 3043
rect 14220 3040 14226 3052
rect 7829 3012 14226 3040
rect 7829 3009 7841 3012
rect 7783 3003 7841 3009
rect 14220 3000 14226 3012
rect 14278 3000 14284 3052
rect 6403 2975 6461 2981
rect 6403 2941 6415 2975
rect 6449 2972 6461 2975
rect 6449 2944 6722 2972
rect 6449 2941 6461 2944
rect 6403 2935 6461 2941
rect 604 2796 610 2848
rect 662 2836 668 2848
rect 6587 2839 6645 2845
rect 6587 2836 6599 2839
rect 662 2808 6599 2836
rect 662 2796 668 2808
rect 6587 2805 6599 2808
rect 6633 2805 6645 2839
rect 6694 2836 6722 2944
rect 7872 2864 7878 2916
rect 7930 2904 7936 2916
rect 8795 2907 8853 2913
rect 7930 2876 7975 2904
rect 7930 2864 7936 2876
rect 8795 2873 8807 2907
rect 8841 2873 8853 2907
rect 8795 2867 8853 2873
rect 7688 2836 7694 2848
rect 6694 2808 7694 2836
rect 6587 2799 6645 2805
rect 7688 2796 7694 2808
rect 7746 2836 7752 2848
rect 8810 2836 8838 2867
rect 7746 2808 8838 2836
rect 7746 2796 7752 2808
rect 38 2746 14758 2768
rect 38 2694 4846 2746
rect 4898 2694 4910 2746
rect 4962 2694 4974 2746
rect 5026 2694 5038 2746
rect 5090 2694 9777 2746
rect 9829 2694 9841 2746
rect 9893 2694 9905 2746
rect 9957 2694 9969 2746
rect 10021 2694 14758 2746
rect 38 2672 14758 2694
rect 7780 2632 7786 2644
rect 6694 2604 7786 2632
rect 6694 2573 6722 2604
rect 7780 2592 7786 2604
rect 7838 2592 7844 2644
rect 6679 2567 6737 2573
rect 6679 2533 6691 2567
rect 6725 2533 6737 2567
rect 6679 2527 6737 2533
rect 7599 2567 7657 2573
rect 7599 2533 7611 2567
rect 7645 2564 7657 2567
rect 7964 2564 7970 2576
rect 7645 2536 7970 2564
rect 7645 2533 7657 2536
rect 7599 2527 7657 2533
rect 7964 2524 7970 2536
rect 8022 2524 8028 2576
rect 4008 2388 4014 2440
rect 4066 2428 4072 2440
rect 6587 2431 6645 2437
rect 6587 2428 6599 2431
rect 4066 2400 6599 2428
rect 4066 2388 4072 2400
rect 6587 2397 6599 2400
rect 6633 2397 6645 2431
rect 6587 2391 6645 2397
rect 38 2202 14758 2224
rect 38 2150 2381 2202
rect 2433 2150 2445 2202
rect 2497 2150 2509 2202
rect 2561 2150 2573 2202
rect 2625 2150 7312 2202
rect 7364 2150 7376 2202
rect 7428 2150 7440 2202
rect 7492 2150 7504 2202
rect 7556 2150 12242 2202
rect 12294 2150 12306 2202
rect 12358 2150 12370 2202
rect 12422 2150 12434 2202
rect 12486 2150 14758 2202
rect 38 2128 14758 2150
<< via1 >>
rect 2381 6502 2433 6554
rect 2445 6502 2497 6554
rect 2509 6502 2561 6554
rect 2573 6502 2625 6554
rect 7312 6502 7364 6554
rect 7376 6502 7428 6554
rect 7440 6502 7492 6554
rect 7504 6502 7556 6554
rect 12242 6502 12294 6554
rect 12306 6502 12358 6554
rect 12370 6502 12422 6554
rect 12434 6502 12486 6554
rect 4846 5958 4898 6010
rect 4910 5958 4962 6010
rect 4974 5958 5026 6010
rect 5038 5958 5090 6010
rect 9777 5958 9829 6010
rect 9841 5958 9893 6010
rect 9905 5958 9957 6010
rect 9969 5958 10021 6010
rect 2381 5414 2433 5466
rect 2445 5414 2497 5466
rect 2509 5414 2561 5466
rect 2573 5414 2625 5466
rect 7312 5414 7364 5466
rect 7376 5414 7428 5466
rect 7440 5414 7492 5466
rect 7504 5414 7556 5466
rect 12242 5414 12294 5466
rect 12306 5414 12358 5466
rect 12370 5414 12422 5466
rect 12434 5414 12486 5466
rect 4846 4870 4898 4922
rect 4910 4870 4962 4922
rect 4974 4870 5026 4922
rect 5038 4870 5090 4922
rect 9777 4870 9829 4922
rect 9841 4870 9893 4922
rect 9905 4870 9957 4922
rect 9969 4870 10021 4922
rect 11742 4675 11794 4684
rect 11742 4641 11751 4675
rect 11751 4641 11785 4675
rect 11785 4641 11794 4675
rect 11742 4632 11794 4641
rect 12110 4675 12162 4684
rect 12110 4641 12119 4675
rect 12119 4641 12153 4675
rect 12153 4641 12162 4675
rect 12110 4632 12162 4641
rect 11466 4428 11518 4480
rect 2381 4326 2433 4378
rect 2445 4326 2497 4378
rect 2509 4326 2561 4378
rect 2573 4326 2625 4378
rect 7312 4326 7364 4378
rect 7376 4326 7428 4378
rect 7440 4326 7492 4378
rect 7504 4326 7556 4378
rect 12242 4326 12294 4378
rect 12306 4326 12358 4378
rect 12370 4326 12422 4378
rect 12434 4326 12486 4378
rect 4846 3782 4898 3834
rect 4910 3782 4962 3834
rect 4974 3782 5026 3834
rect 5038 3782 5090 3834
rect 9777 3782 9829 3834
rect 9841 3782 9893 3834
rect 9905 3782 9957 3834
rect 9969 3782 10021 3834
rect 12110 3680 12162 3732
rect 7786 3544 7838 3596
rect 10822 3544 10874 3596
rect 11466 3544 11518 3596
rect 12662 3544 12714 3596
rect 11374 3519 11426 3528
rect 11374 3485 11383 3519
rect 11383 3485 11417 3519
rect 11417 3485 11426 3519
rect 11374 3476 11426 3485
rect 7878 3340 7930 3392
rect 2381 3238 2433 3290
rect 2445 3238 2497 3290
rect 2509 3238 2561 3290
rect 2573 3238 2625 3290
rect 7312 3238 7364 3290
rect 7376 3238 7428 3290
rect 7440 3238 7492 3290
rect 7504 3238 7556 3290
rect 12242 3238 12294 3290
rect 12306 3238 12358 3290
rect 12370 3238 12422 3290
rect 12434 3238 12486 3290
rect 14226 3000 14278 3052
rect 610 2796 662 2848
rect 7878 2907 7930 2916
rect 7878 2873 7887 2907
rect 7887 2873 7921 2907
rect 7921 2873 7930 2907
rect 7878 2864 7930 2873
rect 7694 2796 7746 2848
rect 4846 2694 4898 2746
rect 4910 2694 4962 2746
rect 4974 2694 5026 2746
rect 5038 2694 5090 2746
rect 9777 2694 9829 2746
rect 9841 2694 9893 2746
rect 9905 2694 9957 2746
rect 9969 2694 10021 2746
rect 7786 2592 7838 2644
rect 7970 2524 8022 2576
rect 4014 2388 4066 2440
rect 2381 2150 2433 2202
rect 2445 2150 2497 2202
rect 2509 2150 2561 2202
rect 2573 2150 2625 2202
rect 7312 2150 7364 2202
rect 7376 2150 7428 2202
rect 7440 2150 7492 2202
rect 7504 2150 7556 2202
rect 12242 2150 12294 2202
rect 12306 2150 12358 2202
rect 12370 2150 12422 2202
rect 12434 2150 12486 2202
<< metal2 >>
rect 7416 8520 7472 9000
rect 7430 6882 7458 8520
rect 11740 7848 11796 7857
rect 11740 7783 11796 7792
rect 7430 6854 8010 6882
rect 2355 6556 2651 6576
rect 2411 6554 2435 6556
rect 2491 6554 2515 6556
rect 2571 6554 2595 6556
rect 2433 6502 2435 6554
rect 2497 6502 2509 6554
rect 2571 6502 2573 6554
rect 2411 6500 2435 6502
rect 2491 6500 2515 6502
rect 2571 6500 2595 6502
rect 2355 6480 2651 6500
rect 7286 6556 7582 6576
rect 7342 6554 7366 6556
rect 7422 6554 7446 6556
rect 7502 6554 7526 6556
rect 7364 6502 7366 6554
rect 7428 6502 7440 6554
rect 7502 6502 7504 6554
rect 7342 6500 7366 6502
rect 7422 6500 7446 6502
rect 7502 6500 7526 6502
rect 7286 6480 7582 6500
rect 4820 6012 5116 6032
rect 4876 6010 4900 6012
rect 4956 6010 4980 6012
rect 5036 6010 5060 6012
rect 4898 5958 4900 6010
rect 4962 5958 4974 6010
rect 5036 5958 5038 6010
rect 4876 5956 4900 5958
rect 4956 5956 4980 5958
rect 5036 5956 5060 5958
rect 4820 5936 5116 5956
rect 2355 5468 2651 5488
rect 2411 5466 2435 5468
rect 2491 5466 2515 5468
rect 2571 5466 2595 5468
rect 2433 5414 2435 5466
rect 2497 5414 2509 5466
rect 2571 5414 2573 5466
rect 2411 5412 2435 5414
rect 2491 5412 2515 5414
rect 2571 5412 2595 5414
rect 2355 5392 2651 5412
rect 7286 5468 7582 5488
rect 7342 5466 7366 5468
rect 7422 5466 7446 5468
rect 7502 5466 7526 5468
rect 7364 5414 7366 5466
rect 7428 5414 7440 5466
rect 7502 5414 7504 5466
rect 7342 5412 7366 5414
rect 7422 5412 7446 5414
rect 7502 5412 7526 5414
rect 7286 5392 7582 5412
rect 4820 4924 5116 4944
rect 4876 4922 4900 4924
rect 4956 4922 4980 4924
rect 5036 4922 5060 4924
rect 4898 4870 4900 4922
rect 4962 4870 4974 4922
rect 5036 4870 5038 4922
rect 4876 4868 4900 4870
rect 4956 4868 4980 4870
rect 5036 4868 5060 4870
rect 4820 4848 5116 4868
rect 2355 4380 2651 4400
rect 2411 4378 2435 4380
rect 2491 4378 2515 4380
rect 2571 4378 2595 4380
rect 2433 4326 2435 4378
rect 2497 4326 2509 4378
rect 2571 4326 2573 4378
rect 2411 4324 2435 4326
rect 2491 4324 2515 4326
rect 2571 4324 2595 4326
rect 2355 4304 2651 4324
rect 7286 4380 7582 4400
rect 7342 4378 7366 4380
rect 7422 4378 7446 4380
rect 7502 4378 7526 4380
rect 7364 4326 7366 4378
rect 7428 4326 7440 4378
rect 7502 4326 7504 4378
rect 7342 4324 7366 4326
rect 7422 4324 7446 4326
rect 7502 4324 7526 4326
rect 7286 4304 7582 4324
rect 4820 3836 5116 3856
rect 4876 3834 4900 3836
rect 4956 3834 4980 3836
rect 5036 3834 5060 3836
rect 4898 3782 4900 3834
rect 4962 3782 4974 3834
rect 5036 3782 5038 3834
rect 4876 3780 4900 3782
rect 4956 3780 4980 3782
rect 5036 3780 5060 3782
rect 4820 3760 5116 3780
rect 7786 3596 7838 3602
rect 7786 3538 7838 3544
rect 2355 3292 2651 3312
rect 2411 3290 2435 3292
rect 2491 3290 2515 3292
rect 2571 3290 2595 3292
rect 2433 3238 2435 3290
rect 2497 3238 2509 3290
rect 2571 3238 2573 3290
rect 2411 3236 2435 3238
rect 2491 3236 2515 3238
rect 2571 3236 2595 3238
rect 2355 3216 2651 3236
rect 7286 3292 7582 3312
rect 7342 3290 7366 3292
rect 7422 3290 7446 3292
rect 7502 3290 7526 3292
rect 7364 3238 7366 3290
rect 7428 3238 7440 3290
rect 7502 3238 7504 3290
rect 7342 3236 7366 3238
rect 7422 3236 7446 3238
rect 7502 3236 7526 3238
rect 7286 3216 7582 3236
rect 610 2848 662 2854
rect 610 2790 662 2796
rect 7694 2848 7746 2854
rect 7694 2790 7746 2796
rect 622 480 650 2790
rect 4820 2748 5116 2768
rect 4876 2746 4900 2748
rect 4956 2746 4980 2748
rect 5036 2746 5060 2748
rect 4898 2694 4900 2746
rect 4962 2694 4974 2746
rect 5036 2694 5038 2746
rect 4876 2692 4900 2694
rect 4956 2692 4980 2694
rect 5036 2692 5060 2694
rect 4820 2672 5116 2692
rect 4014 2440 4066 2446
rect 4014 2382 4066 2388
rect 2355 2204 2651 2224
rect 2411 2202 2435 2204
rect 2491 2202 2515 2204
rect 2571 2202 2595 2204
rect 2433 2150 2435 2202
rect 2497 2150 2509 2202
rect 2571 2150 2573 2202
rect 2411 2148 2435 2150
rect 2491 2148 2515 2150
rect 2571 2148 2595 2150
rect 2355 2128 2651 2148
rect 4026 480 4054 2382
rect 7286 2204 7582 2224
rect 7342 2202 7366 2204
rect 7422 2202 7446 2204
rect 7502 2202 7526 2204
rect 7364 2150 7366 2202
rect 7428 2150 7440 2202
rect 7502 2150 7504 2202
rect 7342 2148 7366 2150
rect 7422 2148 7446 2150
rect 7502 2148 7526 2150
rect 7286 2128 7582 2148
rect 7706 1986 7734 2790
rect 7798 2650 7826 3538
rect 7878 3392 7930 3398
rect 7878 3334 7930 3340
rect 7890 2922 7918 3334
rect 7878 2916 7930 2922
rect 7878 2858 7930 2864
rect 7786 2644 7838 2650
rect 7786 2586 7838 2592
rect 7982 2582 8010 6854
rect 9751 6012 10047 6032
rect 9807 6010 9831 6012
rect 9887 6010 9911 6012
rect 9967 6010 9991 6012
rect 9829 5958 9831 6010
rect 9893 5958 9905 6010
rect 9967 5958 9969 6010
rect 9807 5956 9831 5958
rect 9887 5956 9911 5958
rect 9967 5956 9991 5958
rect 9751 5936 10047 5956
rect 9751 4924 10047 4944
rect 9807 4922 9831 4924
rect 9887 4922 9911 4924
rect 9967 4922 9991 4924
rect 9829 4870 9831 4922
rect 9893 4870 9905 4922
rect 9967 4870 9969 4922
rect 9807 4868 9831 4870
rect 9887 4868 9911 4870
rect 9967 4868 9991 4870
rect 9751 4848 10047 4868
rect 11754 4690 11782 7783
rect 12216 6556 12512 6576
rect 12272 6554 12296 6556
rect 12352 6554 12376 6556
rect 12432 6554 12456 6556
rect 12294 6502 12296 6554
rect 12358 6502 12370 6554
rect 12432 6502 12434 6554
rect 12272 6500 12296 6502
rect 12352 6500 12376 6502
rect 12432 6500 12456 6502
rect 12216 6480 12512 6500
rect 12108 5672 12164 5681
rect 12108 5607 12164 5616
rect 12122 4690 12150 5607
rect 12216 5468 12512 5488
rect 12272 5466 12296 5468
rect 12352 5466 12376 5468
rect 12432 5466 12456 5468
rect 12294 5414 12296 5466
rect 12358 5414 12370 5466
rect 12432 5414 12434 5466
rect 12272 5412 12296 5414
rect 12352 5412 12376 5414
rect 12432 5412 12456 5414
rect 12216 5392 12512 5412
rect 11742 4684 11794 4690
rect 11742 4626 11794 4632
rect 12110 4684 12162 4690
rect 12110 4626 12162 4632
rect 11466 4480 11518 4486
rect 11466 4422 11518 4428
rect 9751 3836 10047 3856
rect 9807 3834 9831 3836
rect 9887 3834 9911 3836
rect 9967 3834 9991 3836
rect 9829 3782 9831 3834
rect 9893 3782 9905 3834
rect 9967 3782 9969 3834
rect 9807 3780 9831 3782
rect 9887 3780 9911 3782
rect 9967 3780 9991 3782
rect 9751 3760 10047 3780
rect 11478 3602 11506 4422
rect 12122 3738 12150 4626
rect 12216 4380 12512 4400
rect 12272 4378 12296 4380
rect 12352 4378 12376 4380
rect 12432 4378 12456 4380
rect 12294 4326 12296 4378
rect 12358 4326 12370 4378
rect 12432 4326 12434 4378
rect 12272 4324 12296 4326
rect 12352 4324 12376 4326
rect 12432 4324 12456 4326
rect 12216 4304 12512 4324
rect 12110 3732 12162 3738
rect 12110 3674 12162 3680
rect 10822 3596 10874 3602
rect 10822 3538 10874 3544
rect 11466 3596 11518 3602
rect 11466 3538 11518 3544
rect 12662 3596 12714 3602
rect 12662 3538 12714 3544
rect 9751 2748 10047 2768
rect 9807 2746 9831 2748
rect 9887 2746 9911 2748
rect 9967 2746 9991 2748
rect 9829 2694 9831 2746
rect 9893 2694 9905 2746
rect 9967 2694 9969 2746
rect 9807 2692 9831 2694
rect 9887 2692 9911 2694
rect 9967 2692 9991 2694
rect 9751 2672 10047 2692
rect 7970 2576 8022 2582
rect 7970 2518 8022 2524
rect 7430 1958 7734 1986
rect 7430 480 7458 1958
rect 10834 480 10862 3538
rect 11374 3528 11426 3534
rect 11374 3470 11426 3476
rect 11386 1193 11414 3470
rect 12674 3369 12702 3538
rect 12660 3360 12716 3369
rect 12216 3292 12512 3312
rect 12660 3295 12716 3304
rect 12272 3290 12296 3292
rect 12352 3290 12376 3292
rect 12432 3290 12456 3292
rect 12294 3238 12296 3290
rect 12358 3238 12370 3290
rect 12432 3238 12434 3290
rect 12272 3236 12296 3238
rect 12352 3236 12376 3238
rect 12432 3236 12456 3238
rect 12216 3216 12512 3236
rect 14226 3052 14278 3058
rect 14226 2994 14278 3000
rect 12216 2204 12512 2224
rect 12272 2202 12296 2204
rect 12352 2202 12376 2204
rect 12432 2202 12456 2204
rect 12294 2150 12296 2202
rect 12358 2150 12370 2202
rect 12432 2150 12434 2202
rect 12272 2148 12296 2150
rect 12352 2148 12376 2150
rect 12432 2148 12456 2150
rect 12216 2128 12512 2148
rect 11372 1184 11428 1193
rect 11372 1119 11428 1128
rect 14238 480 14266 2994
rect 608 0 664 480
rect 4012 0 4068 480
rect 7416 0 7472 480
rect 10820 0 10876 480
rect 14224 0 14280 480
<< via2 >>
rect 11740 7792 11796 7848
rect 2355 6554 2411 6556
rect 2435 6554 2491 6556
rect 2515 6554 2571 6556
rect 2595 6554 2651 6556
rect 2355 6502 2381 6554
rect 2381 6502 2411 6554
rect 2435 6502 2445 6554
rect 2445 6502 2491 6554
rect 2515 6502 2561 6554
rect 2561 6502 2571 6554
rect 2595 6502 2625 6554
rect 2625 6502 2651 6554
rect 2355 6500 2411 6502
rect 2435 6500 2491 6502
rect 2515 6500 2571 6502
rect 2595 6500 2651 6502
rect 7286 6554 7342 6556
rect 7366 6554 7422 6556
rect 7446 6554 7502 6556
rect 7526 6554 7582 6556
rect 7286 6502 7312 6554
rect 7312 6502 7342 6554
rect 7366 6502 7376 6554
rect 7376 6502 7422 6554
rect 7446 6502 7492 6554
rect 7492 6502 7502 6554
rect 7526 6502 7556 6554
rect 7556 6502 7582 6554
rect 7286 6500 7342 6502
rect 7366 6500 7422 6502
rect 7446 6500 7502 6502
rect 7526 6500 7582 6502
rect 4820 6010 4876 6012
rect 4900 6010 4956 6012
rect 4980 6010 5036 6012
rect 5060 6010 5116 6012
rect 4820 5958 4846 6010
rect 4846 5958 4876 6010
rect 4900 5958 4910 6010
rect 4910 5958 4956 6010
rect 4980 5958 5026 6010
rect 5026 5958 5036 6010
rect 5060 5958 5090 6010
rect 5090 5958 5116 6010
rect 4820 5956 4876 5958
rect 4900 5956 4956 5958
rect 4980 5956 5036 5958
rect 5060 5956 5116 5958
rect 2355 5466 2411 5468
rect 2435 5466 2491 5468
rect 2515 5466 2571 5468
rect 2595 5466 2651 5468
rect 2355 5414 2381 5466
rect 2381 5414 2411 5466
rect 2435 5414 2445 5466
rect 2445 5414 2491 5466
rect 2515 5414 2561 5466
rect 2561 5414 2571 5466
rect 2595 5414 2625 5466
rect 2625 5414 2651 5466
rect 2355 5412 2411 5414
rect 2435 5412 2491 5414
rect 2515 5412 2571 5414
rect 2595 5412 2651 5414
rect 7286 5466 7342 5468
rect 7366 5466 7422 5468
rect 7446 5466 7502 5468
rect 7526 5466 7582 5468
rect 7286 5414 7312 5466
rect 7312 5414 7342 5466
rect 7366 5414 7376 5466
rect 7376 5414 7422 5466
rect 7446 5414 7492 5466
rect 7492 5414 7502 5466
rect 7526 5414 7556 5466
rect 7556 5414 7582 5466
rect 7286 5412 7342 5414
rect 7366 5412 7422 5414
rect 7446 5412 7502 5414
rect 7526 5412 7582 5414
rect 4820 4922 4876 4924
rect 4900 4922 4956 4924
rect 4980 4922 5036 4924
rect 5060 4922 5116 4924
rect 4820 4870 4846 4922
rect 4846 4870 4876 4922
rect 4900 4870 4910 4922
rect 4910 4870 4956 4922
rect 4980 4870 5026 4922
rect 5026 4870 5036 4922
rect 5060 4870 5090 4922
rect 5090 4870 5116 4922
rect 4820 4868 4876 4870
rect 4900 4868 4956 4870
rect 4980 4868 5036 4870
rect 5060 4868 5116 4870
rect 2355 4378 2411 4380
rect 2435 4378 2491 4380
rect 2515 4378 2571 4380
rect 2595 4378 2651 4380
rect 2355 4326 2381 4378
rect 2381 4326 2411 4378
rect 2435 4326 2445 4378
rect 2445 4326 2491 4378
rect 2515 4326 2561 4378
rect 2561 4326 2571 4378
rect 2595 4326 2625 4378
rect 2625 4326 2651 4378
rect 2355 4324 2411 4326
rect 2435 4324 2491 4326
rect 2515 4324 2571 4326
rect 2595 4324 2651 4326
rect 7286 4378 7342 4380
rect 7366 4378 7422 4380
rect 7446 4378 7502 4380
rect 7526 4378 7582 4380
rect 7286 4326 7312 4378
rect 7312 4326 7342 4378
rect 7366 4326 7376 4378
rect 7376 4326 7422 4378
rect 7446 4326 7492 4378
rect 7492 4326 7502 4378
rect 7526 4326 7556 4378
rect 7556 4326 7582 4378
rect 7286 4324 7342 4326
rect 7366 4324 7422 4326
rect 7446 4324 7502 4326
rect 7526 4324 7582 4326
rect 4820 3834 4876 3836
rect 4900 3834 4956 3836
rect 4980 3834 5036 3836
rect 5060 3834 5116 3836
rect 4820 3782 4846 3834
rect 4846 3782 4876 3834
rect 4900 3782 4910 3834
rect 4910 3782 4956 3834
rect 4980 3782 5026 3834
rect 5026 3782 5036 3834
rect 5060 3782 5090 3834
rect 5090 3782 5116 3834
rect 4820 3780 4876 3782
rect 4900 3780 4956 3782
rect 4980 3780 5036 3782
rect 5060 3780 5116 3782
rect 2355 3290 2411 3292
rect 2435 3290 2491 3292
rect 2515 3290 2571 3292
rect 2595 3290 2651 3292
rect 2355 3238 2381 3290
rect 2381 3238 2411 3290
rect 2435 3238 2445 3290
rect 2445 3238 2491 3290
rect 2515 3238 2561 3290
rect 2561 3238 2571 3290
rect 2595 3238 2625 3290
rect 2625 3238 2651 3290
rect 2355 3236 2411 3238
rect 2435 3236 2491 3238
rect 2515 3236 2571 3238
rect 2595 3236 2651 3238
rect 7286 3290 7342 3292
rect 7366 3290 7422 3292
rect 7446 3290 7502 3292
rect 7526 3290 7582 3292
rect 7286 3238 7312 3290
rect 7312 3238 7342 3290
rect 7366 3238 7376 3290
rect 7376 3238 7422 3290
rect 7446 3238 7492 3290
rect 7492 3238 7502 3290
rect 7526 3238 7556 3290
rect 7556 3238 7582 3290
rect 7286 3236 7342 3238
rect 7366 3236 7422 3238
rect 7446 3236 7502 3238
rect 7526 3236 7582 3238
rect 4820 2746 4876 2748
rect 4900 2746 4956 2748
rect 4980 2746 5036 2748
rect 5060 2746 5116 2748
rect 4820 2694 4846 2746
rect 4846 2694 4876 2746
rect 4900 2694 4910 2746
rect 4910 2694 4956 2746
rect 4980 2694 5026 2746
rect 5026 2694 5036 2746
rect 5060 2694 5090 2746
rect 5090 2694 5116 2746
rect 4820 2692 4876 2694
rect 4900 2692 4956 2694
rect 4980 2692 5036 2694
rect 5060 2692 5116 2694
rect 2355 2202 2411 2204
rect 2435 2202 2491 2204
rect 2515 2202 2571 2204
rect 2595 2202 2651 2204
rect 2355 2150 2381 2202
rect 2381 2150 2411 2202
rect 2435 2150 2445 2202
rect 2445 2150 2491 2202
rect 2515 2150 2561 2202
rect 2561 2150 2571 2202
rect 2595 2150 2625 2202
rect 2625 2150 2651 2202
rect 2355 2148 2411 2150
rect 2435 2148 2491 2150
rect 2515 2148 2571 2150
rect 2595 2148 2651 2150
rect 7286 2202 7342 2204
rect 7366 2202 7422 2204
rect 7446 2202 7502 2204
rect 7526 2202 7582 2204
rect 7286 2150 7312 2202
rect 7312 2150 7342 2202
rect 7366 2150 7376 2202
rect 7376 2150 7422 2202
rect 7446 2150 7492 2202
rect 7492 2150 7502 2202
rect 7526 2150 7556 2202
rect 7556 2150 7582 2202
rect 7286 2148 7342 2150
rect 7366 2148 7422 2150
rect 7446 2148 7502 2150
rect 7526 2148 7582 2150
rect 9751 6010 9807 6012
rect 9831 6010 9887 6012
rect 9911 6010 9967 6012
rect 9991 6010 10047 6012
rect 9751 5958 9777 6010
rect 9777 5958 9807 6010
rect 9831 5958 9841 6010
rect 9841 5958 9887 6010
rect 9911 5958 9957 6010
rect 9957 5958 9967 6010
rect 9991 5958 10021 6010
rect 10021 5958 10047 6010
rect 9751 5956 9807 5958
rect 9831 5956 9887 5958
rect 9911 5956 9967 5958
rect 9991 5956 10047 5958
rect 9751 4922 9807 4924
rect 9831 4922 9887 4924
rect 9911 4922 9967 4924
rect 9991 4922 10047 4924
rect 9751 4870 9777 4922
rect 9777 4870 9807 4922
rect 9831 4870 9841 4922
rect 9841 4870 9887 4922
rect 9911 4870 9957 4922
rect 9957 4870 9967 4922
rect 9991 4870 10021 4922
rect 10021 4870 10047 4922
rect 9751 4868 9807 4870
rect 9831 4868 9887 4870
rect 9911 4868 9967 4870
rect 9991 4868 10047 4870
rect 12216 6554 12272 6556
rect 12296 6554 12352 6556
rect 12376 6554 12432 6556
rect 12456 6554 12512 6556
rect 12216 6502 12242 6554
rect 12242 6502 12272 6554
rect 12296 6502 12306 6554
rect 12306 6502 12352 6554
rect 12376 6502 12422 6554
rect 12422 6502 12432 6554
rect 12456 6502 12486 6554
rect 12486 6502 12512 6554
rect 12216 6500 12272 6502
rect 12296 6500 12352 6502
rect 12376 6500 12432 6502
rect 12456 6500 12512 6502
rect 12108 5616 12164 5672
rect 12216 5466 12272 5468
rect 12296 5466 12352 5468
rect 12376 5466 12432 5468
rect 12456 5466 12512 5468
rect 12216 5414 12242 5466
rect 12242 5414 12272 5466
rect 12296 5414 12306 5466
rect 12306 5414 12352 5466
rect 12376 5414 12422 5466
rect 12422 5414 12432 5466
rect 12456 5414 12486 5466
rect 12486 5414 12512 5466
rect 12216 5412 12272 5414
rect 12296 5412 12352 5414
rect 12376 5412 12432 5414
rect 12456 5412 12512 5414
rect 9751 3834 9807 3836
rect 9831 3834 9887 3836
rect 9911 3834 9967 3836
rect 9991 3834 10047 3836
rect 9751 3782 9777 3834
rect 9777 3782 9807 3834
rect 9831 3782 9841 3834
rect 9841 3782 9887 3834
rect 9911 3782 9957 3834
rect 9957 3782 9967 3834
rect 9991 3782 10021 3834
rect 10021 3782 10047 3834
rect 9751 3780 9807 3782
rect 9831 3780 9887 3782
rect 9911 3780 9967 3782
rect 9991 3780 10047 3782
rect 12216 4378 12272 4380
rect 12296 4378 12352 4380
rect 12376 4378 12432 4380
rect 12456 4378 12512 4380
rect 12216 4326 12242 4378
rect 12242 4326 12272 4378
rect 12296 4326 12306 4378
rect 12306 4326 12352 4378
rect 12376 4326 12422 4378
rect 12422 4326 12432 4378
rect 12456 4326 12486 4378
rect 12486 4326 12512 4378
rect 12216 4324 12272 4326
rect 12296 4324 12352 4326
rect 12376 4324 12432 4326
rect 12456 4324 12512 4326
rect 9751 2746 9807 2748
rect 9831 2746 9887 2748
rect 9911 2746 9967 2748
rect 9991 2746 10047 2748
rect 9751 2694 9777 2746
rect 9777 2694 9807 2746
rect 9831 2694 9841 2746
rect 9841 2694 9887 2746
rect 9911 2694 9957 2746
rect 9957 2694 9967 2746
rect 9991 2694 10021 2746
rect 10021 2694 10047 2746
rect 9751 2692 9807 2694
rect 9831 2692 9887 2694
rect 9911 2692 9967 2694
rect 9991 2692 10047 2694
rect 12660 3304 12716 3360
rect 12216 3290 12272 3292
rect 12296 3290 12352 3292
rect 12376 3290 12432 3292
rect 12456 3290 12512 3292
rect 12216 3238 12242 3290
rect 12242 3238 12272 3290
rect 12296 3238 12306 3290
rect 12306 3238 12352 3290
rect 12376 3238 12422 3290
rect 12422 3238 12432 3290
rect 12456 3238 12486 3290
rect 12486 3238 12512 3290
rect 12216 3236 12272 3238
rect 12296 3236 12352 3238
rect 12376 3236 12432 3238
rect 12456 3236 12512 3238
rect 12216 2202 12272 2204
rect 12296 2202 12352 2204
rect 12376 2202 12432 2204
rect 12456 2202 12512 2204
rect 12216 2150 12242 2202
rect 12242 2150 12272 2202
rect 12296 2150 12306 2202
rect 12306 2150 12352 2202
rect 12376 2150 12422 2202
rect 12422 2150 12432 2202
rect 12456 2150 12486 2202
rect 12486 2150 12512 2202
rect 12216 2148 12272 2150
rect 12296 2148 12352 2150
rect 12376 2148 12432 2150
rect 12456 2148 12512 2150
rect 11372 1128 11428 1184
<< metal3 >>
rect 11735 7850 11801 7853
rect 15454 7850 15934 7880
rect 11735 7848 15934 7850
rect 11735 7792 11740 7848
rect 11796 7792 15934 7848
rect 11735 7790 15934 7792
rect 11735 7787 11801 7790
rect 15454 7760 15934 7790
rect 2343 6560 2663 6561
rect 2343 6496 2351 6560
rect 2415 6496 2431 6560
rect 2495 6496 2511 6560
rect 2575 6496 2591 6560
rect 2655 6496 2663 6560
rect 2343 6495 2663 6496
rect 7274 6560 7594 6561
rect 7274 6496 7282 6560
rect 7346 6496 7362 6560
rect 7426 6496 7442 6560
rect 7506 6496 7522 6560
rect 7586 6496 7594 6560
rect 7274 6495 7594 6496
rect 12204 6560 12524 6561
rect 12204 6496 12212 6560
rect 12276 6496 12292 6560
rect 12356 6496 12372 6560
rect 12436 6496 12452 6560
rect 12516 6496 12524 6560
rect 12204 6495 12524 6496
rect 4808 6016 5128 6017
rect 4808 5952 4816 6016
rect 4880 5952 4896 6016
rect 4960 5952 4976 6016
rect 5040 5952 5056 6016
rect 5120 5952 5128 6016
rect 4808 5951 5128 5952
rect 9739 6016 10059 6017
rect 9739 5952 9747 6016
rect 9811 5952 9827 6016
rect 9891 5952 9907 6016
rect 9971 5952 9987 6016
rect 10051 5952 10059 6016
rect 9739 5951 10059 5952
rect 12103 5674 12169 5677
rect 15454 5674 15934 5704
rect 12103 5672 15934 5674
rect 12103 5616 12108 5672
rect 12164 5616 15934 5672
rect 12103 5614 15934 5616
rect 12103 5611 12169 5614
rect 15454 5584 15934 5614
rect 2343 5472 2663 5473
rect 2343 5408 2351 5472
rect 2415 5408 2431 5472
rect 2495 5408 2511 5472
rect 2575 5408 2591 5472
rect 2655 5408 2663 5472
rect 2343 5407 2663 5408
rect 7274 5472 7594 5473
rect 7274 5408 7282 5472
rect 7346 5408 7362 5472
rect 7426 5408 7442 5472
rect 7506 5408 7522 5472
rect 7586 5408 7594 5472
rect 7274 5407 7594 5408
rect 12204 5472 12524 5473
rect 12204 5408 12212 5472
rect 12276 5408 12292 5472
rect 12356 5408 12372 5472
rect 12436 5408 12452 5472
rect 12516 5408 12524 5472
rect 12204 5407 12524 5408
rect 4808 4928 5128 4929
rect 4808 4864 4816 4928
rect 4880 4864 4896 4928
rect 4960 4864 4976 4928
rect 5040 4864 5056 4928
rect 5120 4864 5128 4928
rect 4808 4863 5128 4864
rect 9739 4928 10059 4929
rect 9739 4864 9747 4928
rect 9811 4864 9827 4928
rect 9891 4864 9907 4928
rect 9971 4864 9987 4928
rect 10051 4864 10059 4928
rect 9739 4863 10059 4864
rect 2343 4384 2663 4385
rect 2343 4320 2351 4384
rect 2415 4320 2431 4384
rect 2495 4320 2511 4384
rect 2575 4320 2591 4384
rect 2655 4320 2663 4384
rect 2343 4319 2663 4320
rect 7274 4384 7594 4385
rect 7274 4320 7282 4384
rect 7346 4320 7362 4384
rect 7426 4320 7442 4384
rect 7506 4320 7522 4384
rect 7586 4320 7594 4384
rect 7274 4319 7594 4320
rect 12204 4384 12524 4385
rect 12204 4320 12212 4384
rect 12276 4320 12292 4384
rect 12356 4320 12372 4384
rect 12436 4320 12452 4384
rect 12516 4320 12524 4384
rect 12204 4319 12524 4320
rect 4808 3840 5128 3841
rect 4808 3776 4816 3840
rect 4880 3776 4896 3840
rect 4960 3776 4976 3840
rect 5040 3776 5056 3840
rect 5120 3776 5128 3840
rect 4808 3775 5128 3776
rect 9739 3840 10059 3841
rect 9739 3776 9747 3840
rect 9811 3776 9827 3840
rect 9891 3776 9907 3840
rect 9971 3776 9987 3840
rect 10051 3776 10059 3840
rect 9739 3775 10059 3776
rect 12655 3362 12721 3365
rect 15454 3362 15934 3392
rect 12655 3360 15934 3362
rect 12655 3304 12660 3360
rect 12716 3304 15934 3360
rect 12655 3302 15934 3304
rect 12655 3299 12721 3302
rect 2343 3296 2663 3297
rect 2343 3232 2351 3296
rect 2415 3232 2431 3296
rect 2495 3232 2511 3296
rect 2575 3232 2591 3296
rect 2655 3232 2663 3296
rect 2343 3231 2663 3232
rect 7274 3296 7594 3297
rect 7274 3232 7282 3296
rect 7346 3232 7362 3296
rect 7426 3232 7442 3296
rect 7506 3232 7522 3296
rect 7586 3232 7594 3296
rect 7274 3231 7594 3232
rect 12204 3296 12524 3297
rect 12204 3232 12212 3296
rect 12276 3232 12292 3296
rect 12356 3232 12372 3296
rect 12436 3232 12452 3296
rect 12516 3232 12524 3296
rect 15454 3272 15934 3302
rect 12204 3231 12524 3232
rect 4808 2752 5128 2753
rect 4808 2688 4816 2752
rect 4880 2688 4896 2752
rect 4960 2688 4976 2752
rect 5040 2688 5056 2752
rect 5120 2688 5128 2752
rect 4808 2687 5128 2688
rect 9739 2752 10059 2753
rect 9739 2688 9747 2752
rect 9811 2688 9827 2752
rect 9891 2688 9907 2752
rect 9971 2688 9987 2752
rect 10051 2688 10059 2752
rect 9739 2687 10059 2688
rect 2343 2208 2663 2209
rect 2343 2144 2351 2208
rect 2415 2144 2431 2208
rect 2495 2144 2511 2208
rect 2575 2144 2591 2208
rect 2655 2144 2663 2208
rect 2343 2143 2663 2144
rect 7274 2208 7594 2209
rect 7274 2144 7282 2208
rect 7346 2144 7362 2208
rect 7426 2144 7442 2208
rect 7506 2144 7522 2208
rect 7586 2144 7594 2208
rect 7274 2143 7594 2144
rect 12204 2208 12524 2209
rect 12204 2144 12212 2208
rect 12276 2144 12292 2208
rect 12356 2144 12372 2208
rect 12436 2144 12452 2208
rect 12516 2144 12524 2208
rect 12204 2143 12524 2144
rect 11367 1186 11433 1189
rect 15454 1186 15934 1216
rect 11367 1184 15934 1186
rect 11367 1128 11372 1184
rect 11428 1128 15934 1184
rect 11367 1126 15934 1128
rect 11367 1123 11433 1126
rect 15454 1096 15934 1126
<< via3 >>
rect 2351 6556 2415 6560
rect 2351 6500 2355 6556
rect 2355 6500 2411 6556
rect 2411 6500 2415 6556
rect 2351 6496 2415 6500
rect 2431 6556 2495 6560
rect 2431 6500 2435 6556
rect 2435 6500 2491 6556
rect 2491 6500 2495 6556
rect 2431 6496 2495 6500
rect 2511 6556 2575 6560
rect 2511 6500 2515 6556
rect 2515 6500 2571 6556
rect 2571 6500 2575 6556
rect 2511 6496 2575 6500
rect 2591 6556 2655 6560
rect 2591 6500 2595 6556
rect 2595 6500 2651 6556
rect 2651 6500 2655 6556
rect 2591 6496 2655 6500
rect 7282 6556 7346 6560
rect 7282 6500 7286 6556
rect 7286 6500 7342 6556
rect 7342 6500 7346 6556
rect 7282 6496 7346 6500
rect 7362 6556 7426 6560
rect 7362 6500 7366 6556
rect 7366 6500 7422 6556
rect 7422 6500 7426 6556
rect 7362 6496 7426 6500
rect 7442 6556 7506 6560
rect 7442 6500 7446 6556
rect 7446 6500 7502 6556
rect 7502 6500 7506 6556
rect 7442 6496 7506 6500
rect 7522 6556 7586 6560
rect 7522 6500 7526 6556
rect 7526 6500 7582 6556
rect 7582 6500 7586 6556
rect 7522 6496 7586 6500
rect 12212 6556 12276 6560
rect 12212 6500 12216 6556
rect 12216 6500 12272 6556
rect 12272 6500 12276 6556
rect 12212 6496 12276 6500
rect 12292 6556 12356 6560
rect 12292 6500 12296 6556
rect 12296 6500 12352 6556
rect 12352 6500 12356 6556
rect 12292 6496 12356 6500
rect 12372 6556 12436 6560
rect 12372 6500 12376 6556
rect 12376 6500 12432 6556
rect 12432 6500 12436 6556
rect 12372 6496 12436 6500
rect 12452 6556 12516 6560
rect 12452 6500 12456 6556
rect 12456 6500 12512 6556
rect 12512 6500 12516 6556
rect 12452 6496 12516 6500
rect 4816 6012 4880 6016
rect 4816 5956 4820 6012
rect 4820 5956 4876 6012
rect 4876 5956 4880 6012
rect 4816 5952 4880 5956
rect 4896 6012 4960 6016
rect 4896 5956 4900 6012
rect 4900 5956 4956 6012
rect 4956 5956 4960 6012
rect 4896 5952 4960 5956
rect 4976 6012 5040 6016
rect 4976 5956 4980 6012
rect 4980 5956 5036 6012
rect 5036 5956 5040 6012
rect 4976 5952 5040 5956
rect 5056 6012 5120 6016
rect 5056 5956 5060 6012
rect 5060 5956 5116 6012
rect 5116 5956 5120 6012
rect 5056 5952 5120 5956
rect 9747 6012 9811 6016
rect 9747 5956 9751 6012
rect 9751 5956 9807 6012
rect 9807 5956 9811 6012
rect 9747 5952 9811 5956
rect 9827 6012 9891 6016
rect 9827 5956 9831 6012
rect 9831 5956 9887 6012
rect 9887 5956 9891 6012
rect 9827 5952 9891 5956
rect 9907 6012 9971 6016
rect 9907 5956 9911 6012
rect 9911 5956 9967 6012
rect 9967 5956 9971 6012
rect 9907 5952 9971 5956
rect 9987 6012 10051 6016
rect 9987 5956 9991 6012
rect 9991 5956 10047 6012
rect 10047 5956 10051 6012
rect 9987 5952 10051 5956
rect 2351 5468 2415 5472
rect 2351 5412 2355 5468
rect 2355 5412 2411 5468
rect 2411 5412 2415 5468
rect 2351 5408 2415 5412
rect 2431 5468 2495 5472
rect 2431 5412 2435 5468
rect 2435 5412 2491 5468
rect 2491 5412 2495 5468
rect 2431 5408 2495 5412
rect 2511 5468 2575 5472
rect 2511 5412 2515 5468
rect 2515 5412 2571 5468
rect 2571 5412 2575 5468
rect 2511 5408 2575 5412
rect 2591 5468 2655 5472
rect 2591 5412 2595 5468
rect 2595 5412 2651 5468
rect 2651 5412 2655 5468
rect 2591 5408 2655 5412
rect 7282 5468 7346 5472
rect 7282 5412 7286 5468
rect 7286 5412 7342 5468
rect 7342 5412 7346 5468
rect 7282 5408 7346 5412
rect 7362 5468 7426 5472
rect 7362 5412 7366 5468
rect 7366 5412 7422 5468
rect 7422 5412 7426 5468
rect 7362 5408 7426 5412
rect 7442 5468 7506 5472
rect 7442 5412 7446 5468
rect 7446 5412 7502 5468
rect 7502 5412 7506 5468
rect 7442 5408 7506 5412
rect 7522 5468 7586 5472
rect 7522 5412 7526 5468
rect 7526 5412 7582 5468
rect 7582 5412 7586 5468
rect 7522 5408 7586 5412
rect 12212 5468 12276 5472
rect 12212 5412 12216 5468
rect 12216 5412 12272 5468
rect 12272 5412 12276 5468
rect 12212 5408 12276 5412
rect 12292 5468 12356 5472
rect 12292 5412 12296 5468
rect 12296 5412 12352 5468
rect 12352 5412 12356 5468
rect 12292 5408 12356 5412
rect 12372 5468 12436 5472
rect 12372 5412 12376 5468
rect 12376 5412 12432 5468
rect 12432 5412 12436 5468
rect 12372 5408 12436 5412
rect 12452 5468 12516 5472
rect 12452 5412 12456 5468
rect 12456 5412 12512 5468
rect 12512 5412 12516 5468
rect 12452 5408 12516 5412
rect 4816 4924 4880 4928
rect 4816 4868 4820 4924
rect 4820 4868 4876 4924
rect 4876 4868 4880 4924
rect 4816 4864 4880 4868
rect 4896 4924 4960 4928
rect 4896 4868 4900 4924
rect 4900 4868 4956 4924
rect 4956 4868 4960 4924
rect 4896 4864 4960 4868
rect 4976 4924 5040 4928
rect 4976 4868 4980 4924
rect 4980 4868 5036 4924
rect 5036 4868 5040 4924
rect 4976 4864 5040 4868
rect 5056 4924 5120 4928
rect 5056 4868 5060 4924
rect 5060 4868 5116 4924
rect 5116 4868 5120 4924
rect 5056 4864 5120 4868
rect 9747 4924 9811 4928
rect 9747 4868 9751 4924
rect 9751 4868 9807 4924
rect 9807 4868 9811 4924
rect 9747 4864 9811 4868
rect 9827 4924 9891 4928
rect 9827 4868 9831 4924
rect 9831 4868 9887 4924
rect 9887 4868 9891 4924
rect 9827 4864 9891 4868
rect 9907 4924 9971 4928
rect 9907 4868 9911 4924
rect 9911 4868 9967 4924
rect 9967 4868 9971 4924
rect 9907 4864 9971 4868
rect 9987 4924 10051 4928
rect 9987 4868 9991 4924
rect 9991 4868 10047 4924
rect 10047 4868 10051 4924
rect 9987 4864 10051 4868
rect 2351 4380 2415 4384
rect 2351 4324 2355 4380
rect 2355 4324 2411 4380
rect 2411 4324 2415 4380
rect 2351 4320 2415 4324
rect 2431 4380 2495 4384
rect 2431 4324 2435 4380
rect 2435 4324 2491 4380
rect 2491 4324 2495 4380
rect 2431 4320 2495 4324
rect 2511 4380 2575 4384
rect 2511 4324 2515 4380
rect 2515 4324 2571 4380
rect 2571 4324 2575 4380
rect 2511 4320 2575 4324
rect 2591 4380 2655 4384
rect 2591 4324 2595 4380
rect 2595 4324 2651 4380
rect 2651 4324 2655 4380
rect 2591 4320 2655 4324
rect 7282 4380 7346 4384
rect 7282 4324 7286 4380
rect 7286 4324 7342 4380
rect 7342 4324 7346 4380
rect 7282 4320 7346 4324
rect 7362 4380 7426 4384
rect 7362 4324 7366 4380
rect 7366 4324 7422 4380
rect 7422 4324 7426 4380
rect 7362 4320 7426 4324
rect 7442 4380 7506 4384
rect 7442 4324 7446 4380
rect 7446 4324 7502 4380
rect 7502 4324 7506 4380
rect 7442 4320 7506 4324
rect 7522 4380 7586 4384
rect 7522 4324 7526 4380
rect 7526 4324 7582 4380
rect 7582 4324 7586 4380
rect 7522 4320 7586 4324
rect 12212 4380 12276 4384
rect 12212 4324 12216 4380
rect 12216 4324 12272 4380
rect 12272 4324 12276 4380
rect 12212 4320 12276 4324
rect 12292 4380 12356 4384
rect 12292 4324 12296 4380
rect 12296 4324 12352 4380
rect 12352 4324 12356 4380
rect 12292 4320 12356 4324
rect 12372 4380 12436 4384
rect 12372 4324 12376 4380
rect 12376 4324 12432 4380
rect 12432 4324 12436 4380
rect 12372 4320 12436 4324
rect 12452 4380 12516 4384
rect 12452 4324 12456 4380
rect 12456 4324 12512 4380
rect 12512 4324 12516 4380
rect 12452 4320 12516 4324
rect 4816 3836 4880 3840
rect 4816 3780 4820 3836
rect 4820 3780 4876 3836
rect 4876 3780 4880 3836
rect 4816 3776 4880 3780
rect 4896 3836 4960 3840
rect 4896 3780 4900 3836
rect 4900 3780 4956 3836
rect 4956 3780 4960 3836
rect 4896 3776 4960 3780
rect 4976 3836 5040 3840
rect 4976 3780 4980 3836
rect 4980 3780 5036 3836
rect 5036 3780 5040 3836
rect 4976 3776 5040 3780
rect 5056 3836 5120 3840
rect 5056 3780 5060 3836
rect 5060 3780 5116 3836
rect 5116 3780 5120 3836
rect 5056 3776 5120 3780
rect 9747 3836 9811 3840
rect 9747 3780 9751 3836
rect 9751 3780 9807 3836
rect 9807 3780 9811 3836
rect 9747 3776 9811 3780
rect 9827 3836 9891 3840
rect 9827 3780 9831 3836
rect 9831 3780 9887 3836
rect 9887 3780 9891 3836
rect 9827 3776 9891 3780
rect 9907 3836 9971 3840
rect 9907 3780 9911 3836
rect 9911 3780 9967 3836
rect 9967 3780 9971 3836
rect 9907 3776 9971 3780
rect 9987 3836 10051 3840
rect 9987 3780 9991 3836
rect 9991 3780 10047 3836
rect 10047 3780 10051 3836
rect 9987 3776 10051 3780
rect 2351 3292 2415 3296
rect 2351 3236 2355 3292
rect 2355 3236 2411 3292
rect 2411 3236 2415 3292
rect 2351 3232 2415 3236
rect 2431 3292 2495 3296
rect 2431 3236 2435 3292
rect 2435 3236 2491 3292
rect 2491 3236 2495 3292
rect 2431 3232 2495 3236
rect 2511 3292 2575 3296
rect 2511 3236 2515 3292
rect 2515 3236 2571 3292
rect 2571 3236 2575 3292
rect 2511 3232 2575 3236
rect 2591 3292 2655 3296
rect 2591 3236 2595 3292
rect 2595 3236 2651 3292
rect 2651 3236 2655 3292
rect 2591 3232 2655 3236
rect 7282 3292 7346 3296
rect 7282 3236 7286 3292
rect 7286 3236 7342 3292
rect 7342 3236 7346 3292
rect 7282 3232 7346 3236
rect 7362 3292 7426 3296
rect 7362 3236 7366 3292
rect 7366 3236 7422 3292
rect 7422 3236 7426 3292
rect 7362 3232 7426 3236
rect 7442 3292 7506 3296
rect 7442 3236 7446 3292
rect 7446 3236 7502 3292
rect 7502 3236 7506 3292
rect 7442 3232 7506 3236
rect 7522 3292 7586 3296
rect 7522 3236 7526 3292
rect 7526 3236 7582 3292
rect 7582 3236 7586 3292
rect 7522 3232 7586 3236
rect 12212 3292 12276 3296
rect 12212 3236 12216 3292
rect 12216 3236 12272 3292
rect 12272 3236 12276 3292
rect 12212 3232 12276 3236
rect 12292 3292 12356 3296
rect 12292 3236 12296 3292
rect 12296 3236 12352 3292
rect 12352 3236 12356 3292
rect 12292 3232 12356 3236
rect 12372 3292 12436 3296
rect 12372 3236 12376 3292
rect 12376 3236 12432 3292
rect 12432 3236 12436 3292
rect 12372 3232 12436 3236
rect 12452 3292 12516 3296
rect 12452 3236 12456 3292
rect 12456 3236 12512 3292
rect 12512 3236 12516 3292
rect 12452 3232 12516 3236
rect 4816 2748 4880 2752
rect 4816 2692 4820 2748
rect 4820 2692 4876 2748
rect 4876 2692 4880 2748
rect 4816 2688 4880 2692
rect 4896 2748 4960 2752
rect 4896 2692 4900 2748
rect 4900 2692 4956 2748
rect 4956 2692 4960 2748
rect 4896 2688 4960 2692
rect 4976 2748 5040 2752
rect 4976 2692 4980 2748
rect 4980 2692 5036 2748
rect 5036 2692 5040 2748
rect 4976 2688 5040 2692
rect 5056 2748 5120 2752
rect 5056 2692 5060 2748
rect 5060 2692 5116 2748
rect 5116 2692 5120 2748
rect 5056 2688 5120 2692
rect 9747 2748 9811 2752
rect 9747 2692 9751 2748
rect 9751 2692 9807 2748
rect 9807 2692 9811 2748
rect 9747 2688 9811 2692
rect 9827 2748 9891 2752
rect 9827 2692 9831 2748
rect 9831 2692 9887 2748
rect 9887 2692 9891 2748
rect 9827 2688 9891 2692
rect 9907 2748 9971 2752
rect 9907 2692 9911 2748
rect 9911 2692 9967 2748
rect 9967 2692 9971 2748
rect 9907 2688 9971 2692
rect 9987 2748 10051 2752
rect 9987 2692 9991 2748
rect 9991 2692 10047 2748
rect 10047 2692 10051 2748
rect 9987 2688 10051 2692
rect 2351 2204 2415 2208
rect 2351 2148 2355 2204
rect 2355 2148 2411 2204
rect 2411 2148 2415 2204
rect 2351 2144 2415 2148
rect 2431 2204 2495 2208
rect 2431 2148 2435 2204
rect 2435 2148 2491 2204
rect 2491 2148 2495 2204
rect 2431 2144 2495 2148
rect 2511 2204 2575 2208
rect 2511 2148 2515 2204
rect 2515 2148 2571 2204
rect 2571 2148 2575 2204
rect 2511 2144 2575 2148
rect 2591 2204 2655 2208
rect 2591 2148 2595 2204
rect 2595 2148 2651 2204
rect 2651 2148 2655 2204
rect 2591 2144 2655 2148
rect 7282 2204 7346 2208
rect 7282 2148 7286 2204
rect 7286 2148 7342 2204
rect 7342 2148 7346 2204
rect 7282 2144 7346 2148
rect 7362 2204 7426 2208
rect 7362 2148 7366 2204
rect 7366 2148 7422 2204
rect 7422 2148 7426 2204
rect 7362 2144 7426 2148
rect 7442 2204 7506 2208
rect 7442 2148 7446 2204
rect 7446 2148 7502 2204
rect 7502 2148 7506 2204
rect 7442 2144 7506 2148
rect 7522 2204 7586 2208
rect 7522 2148 7526 2204
rect 7526 2148 7582 2204
rect 7582 2148 7586 2204
rect 7522 2144 7586 2148
rect 12212 2204 12276 2208
rect 12212 2148 12216 2204
rect 12216 2148 12272 2204
rect 12272 2148 12276 2204
rect 12212 2144 12276 2148
rect 12292 2204 12356 2208
rect 12292 2148 12296 2204
rect 12296 2148 12352 2204
rect 12352 2148 12356 2204
rect 12292 2144 12356 2148
rect 12372 2204 12436 2208
rect 12372 2148 12376 2204
rect 12376 2148 12432 2204
rect 12432 2148 12436 2204
rect 12372 2144 12436 2148
rect 12452 2204 12516 2208
rect 12452 2148 12456 2204
rect 12456 2148 12512 2204
rect 12512 2148 12516 2204
rect 12452 2144 12516 2148
<< metal4 >>
rect 2343 6560 2663 6576
rect 2343 6496 2351 6560
rect 2415 6496 2431 6560
rect 2495 6496 2511 6560
rect 2575 6496 2591 6560
rect 2655 6496 2663 6560
rect 2343 5472 2663 6496
rect 2343 5408 2351 5472
rect 2415 5408 2431 5472
rect 2495 5408 2511 5472
rect 2575 5408 2591 5472
rect 2655 5408 2663 5472
rect 2343 4384 2663 5408
rect 2343 4320 2351 4384
rect 2415 4320 2431 4384
rect 2495 4320 2511 4384
rect 2575 4320 2591 4384
rect 2655 4320 2663 4384
rect 2343 3296 2663 4320
rect 2343 3232 2351 3296
rect 2415 3232 2431 3296
rect 2495 3232 2511 3296
rect 2575 3232 2591 3296
rect 2655 3232 2663 3296
rect 2343 2208 2663 3232
rect 2343 2144 2351 2208
rect 2415 2144 2431 2208
rect 2495 2144 2511 2208
rect 2575 2144 2591 2208
rect 2655 2144 2663 2208
rect 2343 2128 2663 2144
rect 4808 6016 5129 6576
rect 4808 5952 4816 6016
rect 4880 5952 4896 6016
rect 4960 5952 4976 6016
rect 5040 5952 5056 6016
rect 5120 5952 5129 6016
rect 4808 4928 5129 5952
rect 4808 4864 4816 4928
rect 4880 4864 4896 4928
rect 4960 4864 4976 4928
rect 5040 4864 5056 4928
rect 5120 4864 5129 4928
rect 4808 3840 5129 4864
rect 4808 3776 4816 3840
rect 4880 3776 4896 3840
rect 4960 3776 4976 3840
rect 5040 3776 5056 3840
rect 5120 3776 5129 3840
rect 4808 2752 5129 3776
rect 4808 2688 4816 2752
rect 4880 2688 4896 2752
rect 4960 2688 4976 2752
rect 5040 2688 5056 2752
rect 5120 2688 5129 2752
rect 4808 2128 5129 2688
rect 7274 6560 7594 6576
rect 7274 6496 7282 6560
rect 7346 6496 7362 6560
rect 7426 6496 7442 6560
rect 7506 6496 7522 6560
rect 7586 6496 7594 6560
rect 7274 5472 7594 6496
rect 7274 5408 7282 5472
rect 7346 5408 7362 5472
rect 7426 5408 7442 5472
rect 7506 5408 7522 5472
rect 7586 5408 7594 5472
rect 7274 4384 7594 5408
rect 7274 4320 7282 4384
rect 7346 4320 7362 4384
rect 7426 4320 7442 4384
rect 7506 4320 7522 4384
rect 7586 4320 7594 4384
rect 7274 3296 7594 4320
rect 7274 3232 7282 3296
rect 7346 3232 7362 3296
rect 7426 3232 7442 3296
rect 7506 3232 7522 3296
rect 7586 3232 7594 3296
rect 7274 2208 7594 3232
rect 7274 2144 7282 2208
rect 7346 2144 7362 2208
rect 7426 2144 7442 2208
rect 7506 2144 7522 2208
rect 7586 2144 7594 2208
rect 7274 2128 7594 2144
rect 9739 6016 10059 6576
rect 9739 5952 9747 6016
rect 9811 5952 9827 6016
rect 9891 5952 9907 6016
rect 9971 5952 9987 6016
rect 10051 5952 10059 6016
rect 9739 4928 10059 5952
rect 9739 4864 9747 4928
rect 9811 4864 9827 4928
rect 9891 4864 9907 4928
rect 9971 4864 9987 4928
rect 10051 4864 10059 4928
rect 9739 3840 10059 4864
rect 9739 3776 9747 3840
rect 9811 3776 9827 3840
rect 9891 3776 9907 3840
rect 9971 3776 9987 3840
rect 10051 3776 10059 3840
rect 9739 2752 10059 3776
rect 9739 2688 9747 2752
rect 9811 2688 9827 2752
rect 9891 2688 9907 2752
rect 9971 2688 9987 2752
rect 10051 2688 10059 2752
rect 9739 2128 10059 2688
rect 12204 6560 12524 6576
rect 12204 6496 12212 6560
rect 12276 6496 12292 6560
rect 12356 6496 12372 6560
rect 12436 6496 12452 6560
rect 12516 6496 12524 6560
rect 12204 5472 12524 6496
rect 12204 5408 12212 5472
rect 12276 5408 12292 5472
rect 12356 5408 12372 5472
rect 12436 5408 12452 5472
rect 12516 5408 12524 5472
rect 12204 4384 12524 5408
rect 12204 4320 12212 4384
rect 12276 4320 12292 4384
rect 12356 4320 12372 4384
rect 12436 4320 12452 4384
rect 12516 4320 12524 4384
rect 12204 3296 12524 4320
rect 12204 3232 12212 3296
rect 12276 3232 12292 3296
rect 12356 3232 12372 3296
rect 12436 3232 12452 3296
rect 12516 3232 12524 3296
rect 12204 2208 12524 3232
rect 12204 2144 12212 2208
rect 12276 2144 12292 2208
rect 12356 2144 12372 2208
rect 12436 2144 12452 2208
rect 12516 2144 12524 2208
rect 12204 2128 12524 2144
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 38 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1605641404
transform 1 0 38 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 314 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1605641404
transform 1 0 1418 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1605641404
transform 1 0 314 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1605641404
transform 1 0 1418 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_16 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 2890 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 2522 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1605641404
transform 1 0 2982 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1605641404
transform 1 0 2522 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1605641404
transform 1 0 4086 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1605641404
transform 1 0 3626 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_17
timestamp 1605641404
transform 1 0 5742 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_21
timestamp 1605641404
transform 1 0 5650 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 5190 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63
timestamp 1605641404
transform 1 0 5834 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 4730 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 5466 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_62
timestamp 1605641404
transform 1 0 5742 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6386 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 7674 0 1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1605641404
transform 1 0 6478 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6386 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_83
timestamp 1605641404
transform 1 0 7674 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_68
timestamp 1605641404
transform 1 0 6294 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_73
timestamp 1605641404
transform 1 0 6754 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_81
timestamp 1605641404
transform 1 0 7490 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_18
timestamp 1605641404
transform 1 0 8594 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1605641404
transform 1 0 8410 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1605641404
transform 1 0 8686 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_96
timestamp 1605641404
transform 1 0 8870 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1605641404
transform 1 0 9790 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_108
timestamp 1605641404
transform 1 0 9974 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_19
timestamp 1605641404
transform 1 0 11446 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_22
timestamp 1605641404
transform 1 0 11262 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1605641404
transform 1 0 10894 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1605641404
transform 1 0 11538 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1605641404
transform 1 0 11078 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1605641404
transform 1 0 11354 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1605641404
transform 1 0 12642 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1605641404
transform 1 0 13746 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1605641404
transform 1 0 12458 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_147
timestamp 1605641404
transform 1 0 13562 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1605641404
transform -1 0 14758 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1605641404
transform -1 0 14758 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_20
timestamp 1605641404
transform 1 0 14298 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156
timestamp 1605641404
transform 1 0 14390 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_155
timestamp 1605641404
transform 1 0 14298 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1605641404
transform 1 0 38 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1605641404
transform 1 0 314 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1605641404
transform 1 0 1418 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_23
timestamp 1605641404
transform 1 0 2890 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1605641404
transform 1 0 2522 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1605641404
transform 1 0 2982 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1605641404
transform 1 0 4086 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1605641404
transform 1 0 5190 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1605641404
transform 1 0 6294 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1605641404
transform 1 0 7398 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 8594 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_24
timestamp 1605641404
transform 1 0 8502 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_96
timestamp 1605641404
transform 1 0 8870 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_108
timestamp 1605641404
transform 1 0 9974 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 11354 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_2_120
timestamp 1605641404
transform 1 0 11078 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_139
timestamp 1605641404
transform 1 0 12826 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1605641404
transform 1 0 13930 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1605641404
transform -1 0 14758 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_25
timestamp 1605641404
transform 1 0 14114 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_154
timestamp 1605641404
transform 1 0 14206 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1605641404
transform 1 0 38 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1605641404
transform 1 0 314 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1605641404
transform 1 0 1418 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1605641404
transform 1 0 2522 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1605641404
transform 1 0 3626 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_26
timestamp 1605641404
transform 1 0 5650 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1605641404
transform 1 0 4730 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1605641404
transform 1 0 5466 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1605641404
transform 1 0 5742 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1605641404
transform 1 0 6846 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1605641404
transform 1 0 7950 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1605641404
transform 1 0 9054 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1605641404
transform 1 0 10158 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_27
timestamp 1605641404
transform 1 0 11262 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1605641404
transform 1 0 11354 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1605641404
transform 1 0 12458 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_147
timestamp 1605641404
transform 1 0 13562 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1605641404
transform -1 0 14758 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_155
timestamp 1605641404
transform 1 0 14298 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1605641404
transform 1 0 38 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1605641404
transform 1 0 314 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1605641404
transform 1 0 1418 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_28
timestamp 1605641404
transform 1 0 2890 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1605641404
transform 1 0 2522 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1605641404
transform 1 0 2982 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1605641404
transform 1 0 4086 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1605641404
transform 1 0 5190 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1605641404
transform 1 0 6294 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1605641404
transform 1 0 7398 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_29
timestamp 1605641404
transform 1 0 8502 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1605641404
transform 1 0 8594 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1605641404
transform 1 0 9698 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_117
timestamp 1605641404
transform 1 0 10802 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 11722 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_125
timestamp 1605641404
transform 1 0 11538 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_136
timestamp 1605641404
transform 1 0 12550 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_148
timestamp 1605641404
transform 1 0 13654 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1605641404
transform -1 0 14758 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_30
timestamp 1605641404
transform 1 0 14114 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1605641404
transform 1 0 14022 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_154
timestamp 1605641404
transform 1 0 14206 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1605641404
transform 1 0 38 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1605641404
transform 1 0 314 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1605641404
transform 1 0 1418 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1605641404
transform 1 0 2522 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1605641404
transform 1 0 3626 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_31
timestamp 1605641404
transform 1 0 5650 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1605641404
transform 1 0 4730 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1605641404
transform 1 0 5466 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1605641404
transform 1 0 5742 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1605641404
transform 1 0 6846 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1605641404
transform 1 0 7950 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1605641404
transform 1 0 9054 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1605641404
transform 1 0 10158 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_32
timestamp 1605641404
transform 1 0 11262 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1605641404
transform 1 0 11354 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1605641404
transform 1 0 12458 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_147
timestamp 1605641404
transform 1 0 13562 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1605641404
transform -1 0 14758 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_155
timestamp 1605641404
transform 1 0 14298 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1605641404
transform 1 0 38 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1605641404
transform 1 0 38 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1605641404
transform 1 0 314 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1605641404
transform 1 0 1418 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1605641404
transform 1 0 314 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1605641404
transform 1 0 1418 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_33
timestamp 1605641404
transform 1 0 2890 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_36
timestamp 1605641404
transform 1 0 2890 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1605641404
transform 1 0 2522 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1605641404
transform 1 0 2982 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1605641404
transform 1 0 2522 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_32
timestamp 1605641404
transform 1 0 2982 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1605641404
transform 1 0 4086 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_44
timestamp 1605641404
transform 1 0 4086 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_37
timestamp 1605641404
transform 1 0 5742 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1605641404
transform 1 0 5190 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_56
timestamp 1605641404
transform 1 0 5190 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_63
timestamp 1605641404
transform 1 0 5834 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1605641404
transform 1 0 6294 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1605641404
transform 1 0 7398 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_75
timestamp 1605641404
transform 1 0 6938 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_34
timestamp 1605641404
transform 1 0 8502 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_38
timestamp 1605641404
transform 1 0 8594 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1605641404
transform 1 0 8594 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_87
timestamp 1605641404
transform 1 0 8042 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_94
timestamp 1605641404
transform 1 0 8686 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1605641404
transform 1 0 9698 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1605641404
transform 1 0 10802 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_106
timestamp 1605641404
transform 1 0 9790 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_39
timestamp 1605641404
transform 1 0 11446 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1605641404
transform 1 0 11906 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_118
timestamp 1605641404
transform 1 0 10894 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1605641404
transform 1 0 11538 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1605641404
transform 1 0 13010 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1605641404
transform 1 0 12642 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_149
timestamp 1605641404
transform 1 0 13746 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1605641404
transform -1 0 14758 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1605641404
transform -1 0 14758 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_35
timestamp 1605641404
transform 1 0 14114 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_40
timestamp 1605641404
transform 1 0 14298 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_154
timestamp 1605641404
transform 1 0 14206 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_156
timestamp 1605641404
transform 1 0 14390 0 1 5984
box -38 -48 130 592
<< labels >>
rlabel metal3 s 15454 7760 15934 7880 6 IO_ISOL_N
port 0 nsew default input
rlabel metal2 s 4012 0 4068 480 6 bottom_width_0_height_0__pin_0_
port 1 nsew default input
rlabel metal2 s 7416 0 7472 480 6 bottom_width_0_height_0__pin_1_lower
port 2 nsew default tristate
rlabel metal2 s 608 0 664 480 6 bottom_width_0_height_0__pin_1_upper
port 3 nsew default tristate
rlabel metal3 s 15454 3272 15934 3392 6 ccff_head
port 4 nsew default input
rlabel metal3 s 15454 5584 15934 5704 6 ccff_tail
port 5 nsew default tristate
rlabel metal2 s 10820 0 10876 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 6 nsew default tristate
rlabel metal2 s 14224 0 14280 480 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 7 nsew default input
rlabel metal2 s 7416 8520 7472 9000 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 8 nsew default tristate
rlabel metal3 s 15454 1096 15934 1216 6 prog_clk
port 9 nsew default input
rlabel metal4 s 2343 2128 2663 6576 6 VPWR
port 10 nsew default input
rlabel metal4 s 4809 2128 5129 6576 6 VGND
port 11 nsew default input
<< properties >>
string FIXED_BBOX 0 0 15934 9000
<< end >>
