VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga_top
  CLASS BLOCK ;
  FOREIGN fpga_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 1188.700 BY 1276.880 ;
  PIN Test_en
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1070.960 51.880 1071.560 ;
    END
  END Test_en
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1137.080 1055.320 1139.480 1055.920 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 97.880 51.880 98.480 ;
    END
  END ccff_tail
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1179.080 51.880 1179.680 ;
    END
  END clk
  PIN gfpga_pad_GPIO_A[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 117.650 1231.720 117.930 1234.120 ;
    END
  END gfpga_pad_GPIO_A[0]
  PIN gfpga_pad_GPIO_A[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 253.810 1231.720 254.090 1234.120 ;
    END
  END gfpga_pad_GPIO_A[1]
  PIN gfpga_pad_GPIO_A[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1137.080 103.320 1139.480 103.920 ;
    END
  END gfpga_pad_GPIO_A[2]
  PIN gfpga_pad_GPIO_A[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1137.080 222.320 1139.480 222.920 ;
    END
  END gfpga_pad_GPIO_A[3]
  PIN gfpga_pad_GPIO_A[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 117.650 44.120 117.930 46.520 ;
    END
  END gfpga_pad_GPIO_A[4]
  PIN gfpga_pad_GPIO_A[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 253.810 44.120 254.090 46.520 ;
    END
  END gfpga_pad_GPIO_A[5]
  PIN gfpga_pad_GPIO_A[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 206.000 51.880 206.600 ;
    END
  END gfpga_pad_GPIO_A[6]
  PIN gfpga_pad_GPIO_A[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 314.120 51.880 314.720 ;
    END
  END gfpga_pad_GPIO_A[7]
  PIN gfpga_pad_GPIO_IE[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 389.970 1231.720 390.250 1234.120 ;
    END
  END gfpga_pad_GPIO_IE[0]
  PIN gfpga_pad_GPIO_IE[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 526.130 1231.720 526.410 1234.120 ;
    END
  END gfpga_pad_GPIO_IE[1]
  PIN gfpga_pad_GPIO_IE[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1137.080 341.320 1139.480 341.920 ;
    END
  END gfpga_pad_GPIO_IE[2]
  PIN gfpga_pad_GPIO_IE[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1137.080 460.320 1139.480 460.920 ;
    END
  END gfpga_pad_GPIO_IE[3]
  PIN gfpga_pad_GPIO_IE[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 389.970 44.120 390.250 46.520 ;
    END
  END gfpga_pad_GPIO_IE[4]
  PIN gfpga_pad_GPIO_IE[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 526.130 44.120 526.410 46.520 ;
    END
  END gfpga_pad_GPIO_IE[5]
  PIN gfpga_pad_GPIO_IE[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 422.240 51.880 422.840 ;
    END
  END gfpga_pad_GPIO_IE[6]
  PIN gfpga_pad_GPIO_IE[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 530.360 51.880 530.960 ;
    END
  END gfpga_pad_GPIO_IE[7]
  PIN gfpga_pad_GPIO_OE[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 662.750 1231.720 663.030 1234.120 ;
    END
  END gfpga_pad_GPIO_OE[0]
  PIN gfpga_pad_GPIO_OE[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 798.910 1231.720 799.190 1234.120 ;
    END
  END gfpga_pad_GPIO_OE[1]
  PIN gfpga_pad_GPIO_OE[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1137.080 579.320 1139.480 579.920 ;
    END
  END gfpga_pad_GPIO_OE[2]
  PIN gfpga_pad_GPIO_OE[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1137.080 698.320 1139.480 698.920 ;
    END
  END gfpga_pad_GPIO_OE[3]
  PIN gfpga_pad_GPIO_OE[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 662.750 44.120 663.030 46.520 ;
    END
  END gfpga_pad_GPIO_OE[4]
  PIN gfpga_pad_GPIO_OE[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 798.910 44.120 799.190 46.520 ;
    END
  END gfpga_pad_GPIO_OE[5]
  PIN gfpga_pad_GPIO_OE[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 638.480 51.880 639.080 ;
    END
  END gfpga_pad_GPIO_OE[6]
  PIN gfpga_pad_GPIO_OE[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 746.600 51.880 747.200 ;
    END
  END gfpga_pad_GPIO_OE[7]
  PIN gfpga_pad_GPIO_Y[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 935.070 1231.720 935.350 1234.120 ;
    END
  END gfpga_pad_GPIO_Y[0]
  PIN gfpga_pad_GPIO_Y[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1071.230 1231.720 1071.510 1234.120 ;
    END
  END gfpga_pad_GPIO_Y[1]
  PIN gfpga_pad_GPIO_Y[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 1137.080 817.320 1139.480 817.920 ;
    END
  END gfpga_pad_GPIO_Y[2]
  PIN gfpga_pad_GPIO_Y[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 1137.080 936.320 1139.480 936.920 ;
    END
  END gfpga_pad_GPIO_Y[3]
  PIN gfpga_pad_GPIO_Y[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 935.070 44.120 935.350 46.520 ;
    END
  END gfpga_pad_GPIO_Y[4]
  PIN gfpga_pad_GPIO_Y[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1071.230 44.120 1071.510 46.520 ;
    END
  END gfpga_pad_GPIO_Y[5]
  PIN gfpga_pad_GPIO_Y[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 854.720 51.880 855.320 ;
    END
  END gfpga_pad_GPIO_Y[6]
  PIN gfpga_pad_GPIO_Y[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 962.840 51.880 963.440 ;
    END
  END gfpga_pad_GPIO_Y[7]
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1137.080 1174.320 1139.480 1174.920 ;
    END
  END prog_clk
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 25.000 25.000 1163.700 45.000 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.000 1188.700 20.000 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 75.000 74.915 1114.235 1203.005 ;
      LAYER met1 ;
        RECT 66.570 51.980 1117.990 1224.560 ;
      LAYER met2 ;
        RECT 52.330 1231.440 117.370 1231.720 ;
        RECT 118.210 1231.440 253.530 1231.720 ;
        RECT 254.370 1231.440 389.690 1231.720 ;
        RECT 390.530 1231.440 525.850 1231.720 ;
        RECT 526.690 1231.440 662.470 1231.720 ;
        RECT 663.310 1231.440 798.630 1231.720 ;
        RECT 799.470 1231.440 934.790 1231.720 ;
        RECT 935.630 1231.440 1070.950 1231.720 ;
        RECT 1071.790 1231.440 1126.250 1231.720 ;
        RECT 52.330 46.800 1126.250 1231.440 ;
        RECT 52.330 46.520 117.370 46.800 ;
        RECT 118.210 46.520 253.530 46.800 ;
        RECT 254.370 46.520 389.690 46.800 ;
        RECT 390.530 46.520 525.850 46.800 ;
        RECT 526.690 46.520 662.470 46.800 ;
        RECT 663.310 46.520 798.630 46.800 ;
        RECT 799.470 46.520 934.790 46.800 ;
        RECT 935.630 46.520 1070.950 46.800 ;
        RECT 1071.790 46.520 1126.250 46.800 ;
      LAYER met3 ;
        RECT 51.880 1180.080 1137.080 1203.085 ;
        RECT 52.280 1178.680 1137.080 1180.080 ;
        RECT 51.880 1175.320 1137.080 1178.680 ;
        RECT 51.880 1173.920 1136.680 1175.320 ;
        RECT 51.880 1071.960 1137.080 1173.920 ;
        RECT 52.280 1070.560 1137.080 1071.960 ;
        RECT 51.880 1056.320 1137.080 1070.560 ;
        RECT 51.880 1054.920 1136.680 1056.320 ;
        RECT 51.880 963.840 1137.080 1054.920 ;
        RECT 52.280 962.440 1137.080 963.840 ;
        RECT 51.880 937.320 1137.080 962.440 ;
        RECT 51.880 935.920 1136.680 937.320 ;
        RECT 51.880 855.720 1137.080 935.920 ;
        RECT 52.280 854.320 1137.080 855.720 ;
        RECT 51.880 818.320 1137.080 854.320 ;
        RECT 51.880 816.920 1136.680 818.320 ;
        RECT 51.880 747.600 1137.080 816.920 ;
        RECT 52.280 746.200 1137.080 747.600 ;
        RECT 51.880 699.320 1137.080 746.200 ;
        RECT 51.880 697.920 1136.680 699.320 ;
        RECT 51.880 639.480 1137.080 697.920 ;
        RECT 52.280 638.080 1137.080 639.480 ;
        RECT 51.880 580.320 1137.080 638.080 ;
        RECT 51.880 578.920 1136.680 580.320 ;
        RECT 51.880 531.360 1137.080 578.920 ;
        RECT 52.280 529.960 1137.080 531.360 ;
        RECT 51.880 461.320 1137.080 529.960 ;
        RECT 51.880 459.920 1136.680 461.320 ;
        RECT 51.880 423.240 1137.080 459.920 ;
        RECT 52.280 421.840 1137.080 423.240 ;
        RECT 51.880 342.320 1137.080 421.840 ;
        RECT 51.880 340.920 1136.680 342.320 ;
        RECT 51.880 315.120 1137.080 340.920 ;
        RECT 52.280 313.720 1137.080 315.120 ;
        RECT 51.880 223.320 1137.080 313.720 ;
        RECT 51.880 221.920 1136.680 223.320 ;
        RECT 51.880 207.000 1137.080 221.920 ;
        RECT 52.280 205.600 1137.080 207.000 ;
        RECT 51.880 104.320 1137.080 205.600 ;
        RECT 51.880 102.920 1136.680 104.320 ;
        RECT 51.880 98.880 1137.080 102.920 ;
        RECT 52.280 97.480 1137.080 98.880 ;
        RECT 51.880 71.095 1137.080 97.480 ;
      LAYER met4 ;
        RECT 0.000 0.000 1188.700 1276.880 ;
      LAYER met5 ;
        RECT 0.000 79.200 1188.700 1276.880 ;
  END
END fpga_top
END LIBRARY

