magic
tech sky130A
magscale 1 2
timestamp 1605003818
<< locali >>
rect 11069 25143 11103 25381
rect 14473 21879 14507 21981
rect 15853 20247 15887 20349
rect 23489 20247 23523 20485
rect 3341 19703 3375 19873
rect 11897 18615 11931 18853
rect 18889 18071 18923 18309
rect 11989 15895 12023 16065
rect 16129 13787 16163 13957
rect 4629 12699 4663 12869
rect 6837 12631 6871 12937
rect 9229 11611 9263 11849
rect 10425 11679 10459 11849
rect 3709 9979 3743 10149
rect 19901 7191 19935 7293
rect 13277 5015 13311 5253
rect 18153 3927 18187 4097
rect 2237 2839 2271 2941
<< viali >>
rect 8769 25449 8803 25483
rect 10517 25449 10551 25483
rect 20177 25449 20211 25483
rect 21465 25449 21499 25483
rect 11069 25381 11103 25415
rect 14381 25381 14415 25415
rect 15853 25381 15887 25415
rect 1409 25313 1443 25347
rect 8585 25313 8619 25347
rect 10333 25313 10367 25347
rect 10977 25313 11011 25347
rect 8493 25245 8527 25279
rect 7849 25177 7883 25211
rect 9229 25177 9263 25211
rect 9597 25177 9631 25211
rect 9965 25177 9999 25211
rect 11437 25313 11471 25347
rect 12173 25313 12207 25347
rect 13001 25313 13035 25347
rect 14105 25313 14139 25347
rect 17141 25313 17175 25347
rect 17693 25313 17727 25347
rect 18521 25313 18555 25347
rect 18889 25313 18923 25347
rect 19993 25313 20027 25347
rect 21281 25313 21315 25347
rect 22753 25313 22787 25347
rect 22845 25313 22879 25347
rect 24409 25313 24443 25347
rect 12817 25245 12851 25279
rect 15945 25245 15979 25279
rect 16129 25245 16163 25279
rect 16865 25245 16899 25279
rect 23029 25245 23063 25279
rect 24501 25245 24535 25279
rect 24593 25245 24627 25279
rect 11253 25177 11287 25211
rect 17325 25177 17359 25211
rect 19073 25177 19107 25211
rect 22109 25177 22143 25211
rect 25053 25177 25087 25211
rect 1593 25109 1627 25143
rect 11069 25109 11103 25143
rect 11621 25109 11655 25143
rect 13185 25109 13219 25143
rect 13553 25109 13587 25143
rect 13921 25109 13955 25143
rect 14841 25109 14875 25143
rect 15301 25109 15335 25143
rect 15485 25109 15519 25143
rect 16589 25109 16623 25143
rect 18061 25109 18095 25143
rect 21005 25109 21039 25143
rect 22385 25109 22419 25143
rect 24041 25109 24075 25143
rect 1593 24905 1627 24939
rect 7113 24905 7147 24939
rect 7665 24905 7699 24939
rect 8769 24905 8803 24939
rect 23029 24905 23063 24939
rect 8493 24837 8527 24871
rect 9873 24837 9907 24871
rect 9597 24769 9631 24803
rect 11437 24769 11471 24803
rect 11805 24769 11839 24803
rect 13645 24769 13679 24803
rect 14289 24769 14323 24803
rect 15209 24769 15243 24803
rect 15393 24769 15427 24803
rect 16865 24769 16899 24803
rect 18245 24769 18279 24803
rect 21557 24769 21591 24803
rect 22477 24769 22511 24803
rect 22661 24769 22695 24803
rect 25053 24769 25087 24803
rect 25513 24769 25547 24803
rect 1409 24701 1443 24735
rect 2513 24701 2547 24735
rect 7481 24701 7515 24735
rect 8033 24701 8067 24735
rect 8585 24701 8619 24735
rect 9137 24701 9171 24735
rect 9689 24701 9723 24735
rect 10333 24701 10367 24735
rect 11161 24701 11195 24735
rect 13461 24701 13495 24735
rect 15117 24701 15151 24735
rect 16129 24701 16163 24735
rect 17325 24701 17359 24735
rect 18061 24701 18095 24735
rect 19809 24701 19843 24735
rect 20913 24701 20947 24735
rect 24317 24701 24351 24735
rect 24961 24701 24995 24735
rect 10701 24633 10735 24667
rect 12725 24633 12759 24667
rect 14657 24633 14691 24667
rect 21833 24633 21867 24667
rect 22385 24633 22419 24667
rect 24869 24633 24903 24667
rect 2053 24565 2087 24599
rect 2421 24565 2455 24599
rect 2697 24565 2731 24599
rect 3065 24565 3099 24599
rect 10793 24565 10827 24599
rect 11253 24565 11287 24599
rect 12173 24565 12207 24599
rect 13001 24565 13035 24599
rect 14749 24565 14783 24599
rect 15853 24565 15887 24599
rect 16313 24565 16347 24599
rect 16681 24565 16715 24599
rect 16773 24565 16807 24599
rect 17785 24565 17819 24599
rect 18889 24565 18923 24599
rect 19349 24565 19383 24599
rect 19993 24565 20027 24599
rect 20453 24565 20487 24599
rect 20729 24565 20763 24599
rect 21097 24565 21131 24599
rect 22017 24565 22051 24599
rect 23489 24565 23523 24599
rect 23949 24565 23983 24599
rect 24501 24565 24535 24599
rect 1593 24361 1627 24395
rect 2697 24361 2731 24395
rect 6377 24361 6411 24395
rect 7573 24361 7607 24395
rect 8309 24361 8343 24395
rect 8677 24361 8711 24395
rect 12081 24361 12115 24395
rect 19901 24361 19935 24395
rect 21465 24361 21499 24395
rect 22109 24361 22143 24395
rect 6101 24293 6135 24327
rect 13737 24293 13771 24327
rect 14841 24293 14875 24327
rect 16405 24293 16439 24327
rect 23305 24293 23339 24327
rect 1409 24225 1443 24259
rect 2513 24225 2547 24259
rect 6193 24225 6227 24259
rect 7389 24225 7423 24259
rect 8493 24225 8527 24259
rect 10517 24225 10551 24259
rect 10609 24225 10643 24259
rect 11621 24225 11655 24259
rect 12173 24225 12207 24259
rect 13645 24225 13679 24259
rect 15669 24225 15703 24259
rect 17233 24225 17267 24259
rect 18429 24225 18463 24259
rect 19165 24225 19199 24259
rect 19717 24225 19751 24259
rect 21373 24225 21407 24259
rect 22477 24225 22511 24259
rect 23765 24225 23799 24259
rect 23857 24225 23891 24259
rect 24501 24225 24535 24259
rect 24961 24225 24995 24259
rect 10793 24157 10827 24191
rect 12265 24157 12299 24191
rect 13185 24157 13219 24191
rect 13829 24157 13863 24191
rect 15761 24157 15795 24191
rect 15945 24157 15979 24191
rect 17325 24157 17359 24191
rect 17417 24157 17451 24191
rect 18705 24157 18739 24191
rect 19625 24157 19659 24191
rect 21557 24157 21591 24191
rect 23949 24157 23983 24191
rect 3157 24089 3191 24123
rect 4353 24089 4387 24123
rect 4905 24089 4939 24123
rect 10149 24089 10183 24123
rect 11253 24089 11287 24123
rect 14473 24089 14507 24123
rect 16773 24089 16807 24123
rect 22753 24089 22787 24123
rect 23397 24089 23431 24123
rect 25145 24089 25179 24123
rect 2053 24021 2087 24055
rect 2329 24021 2363 24055
rect 5273 24021 5307 24055
rect 6745 24021 6779 24055
rect 7205 24021 7239 24055
rect 9413 24021 9447 24055
rect 9873 24021 9907 24055
rect 11713 24021 11747 24055
rect 12817 24021 12851 24055
rect 13277 24021 13311 24055
rect 15301 24021 15335 24055
rect 16865 24021 16899 24055
rect 18153 24021 18187 24055
rect 20361 24021 20395 24055
rect 20729 24021 20763 24055
rect 21005 24021 21039 24055
rect 1593 23817 1627 23851
rect 2697 23817 2731 23851
rect 3525 23817 3559 23851
rect 6653 23817 6687 23851
rect 8401 23817 8435 23851
rect 9321 23817 9355 23851
rect 11437 23817 11471 23851
rect 15577 23817 15611 23851
rect 16037 23817 16071 23851
rect 18061 23817 18095 23851
rect 21281 23817 21315 23851
rect 24961 23817 24995 23851
rect 5181 23749 5215 23783
rect 7297 23749 7331 23783
rect 12449 23749 12483 23783
rect 13461 23749 13495 23783
rect 13829 23749 13863 23783
rect 17141 23749 17175 23783
rect 20177 23749 20211 23783
rect 21741 23749 21775 23783
rect 3065 23681 3099 23715
rect 4721 23681 4755 23715
rect 5825 23681 5859 23715
rect 8769 23681 8803 23715
rect 9781 23681 9815 23715
rect 9965 23681 9999 23715
rect 12909 23681 12943 23715
rect 13093 23681 13127 23715
rect 15209 23681 15243 23715
rect 16589 23681 16623 23715
rect 16681 23681 16715 23715
rect 18613 23681 18647 23715
rect 19073 23681 19107 23715
rect 20729 23681 20763 23715
rect 22293 23681 22327 23715
rect 23489 23681 23523 23715
rect 24317 23681 24351 23715
rect 1409 23613 1443 23647
rect 2513 23613 2547 23647
rect 3617 23613 3651 23647
rect 4169 23613 4203 23647
rect 6193 23613 6227 23647
rect 7113 23613 7147 23647
rect 8217 23613 8251 23647
rect 9229 23613 9263 23647
rect 10701 23613 10735 23647
rect 11253 23613 11287 23647
rect 11805 23613 11839 23647
rect 14933 23613 14967 23647
rect 24133 23613 24167 23647
rect 25237 23613 25271 23647
rect 25789 23613 25823 23647
rect 10425 23545 10459 23579
rect 12173 23545 12207 23579
rect 15025 23545 15059 23579
rect 16497 23545 16531 23579
rect 18521 23545 18555 23579
rect 19717 23545 19751 23579
rect 20637 23545 20671 23579
rect 21557 23545 21591 23579
rect 22201 23545 22235 23579
rect 24041 23545 24075 23579
rect 26249 23545 26283 23579
rect 2053 23477 2087 23511
rect 2329 23477 2363 23511
rect 3801 23477 3835 23511
rect 4997 23477 5031 23511
rect 5549 23477 5583 23511
rect 5641 23477 5675 23511
rect 7849 23477 7883 23511
rect 9689 23477 9723 23511
rect 11069 23477 11103 23511
rect 12817 23477 12851 23511
rect 14381 23477 14415 23511
rect 14565 23477 14599 23511
rect 16129 23477 16163 23511
rect 17509 23477 17543 23511
rect 18429 23477 18463 23511
rect 19993 23477 20027 23511
rect 20545 23477 20579 23511
rect 22109 23477 22143 23511
rect 22753 23477 22787 23511
rect 23673 23477 23707 23511
rect 25421 23477 25455 23511
rect 3709 23273 3743 23307
rect 6561 23273 6595 23307
rect 11069 23273 11103 23307
rect 12265 23273 12299 23307
rect 13645 23273 13679 23307
rect 16865 23273 16899 23307
rect 17233 23273 17267 23307
rect 18061 23273 18095 23307
rect 18429 23273 18463 23307
rect 21097 23273 21131 23307
rect 23305 23273 23339 23307
rect 23489 23273 23523 23307
rect 24869 23273 24903 23307
rect 1685 23205 1719 23239
rect 2513 23205 2547 23239
rect 5181 23205 5215 23239
rect 6653 23205 6687 23239
rect 13369 23205 13403 23239
rect 14105 23205 14139 23239
rect 18889 23205 18923 23239
rect 23857 23205 23891 23239
rect 25329 23205 25363 23239
rect 2237 23137 2271 23171
rect 4905 23137 4939 23171
rect 8125 23137 8159 23171
rect 10609 23137 10643 23171
rect 12633 23137 12667 23171
rect 13829 23137 13863 23171
rect 15669 23137 15703 23171
rect 18797 23137 18831 23171
rect 21465 23137 21499 23171
rect 25053 23137 25087 23171
rect 6837 23069 6871 23103
rect 8217 23069 8251 23103
rect 8309 23069 8343 23103
rect 11161 23069 11195 23103
rect 11345 23069 11379 23103
rect 12725 23069 12759 23103
rect 12909 23069 12943 23103
rect 15761 23069 15795 23103
rect 15945 23069 15979 23103
rect 17325 23069 17359 23103
rect 17417 23069 17451 23103
rect 18981 23069 19015 23103
rect 19441 23069 19475 23103
rect 19809 23069 19843 23103
rect 21557 23069 21591 23103
rect 21741 23069 21775 23103
rect 22201 23069 22235 23103
rect 23949 23069 23983 23103
rect 24041 23069 24075 23103
rect 5733 23001 5767 23035
rect 6193 23001 6227 23035
rect 7757 23001 7791 23035
rect 9321 23001 9355 23035
rect 10241 23001 10275 23035
rect 15301 23001 15335 23035
rect 22477 23001 22511 23035
rect 2053 22933 2087 22967
rect 2973 22933 3007 22967
rect 4353 22933 4387 22967
rect 4813 22933 4847 22967
rect 6101 22933 6135 22967
rect 7481 22933 7515 22967
rect 9045 22933 9079 22967
rect 10701 22933 10735 22967
rect 11805 22933 11839 22967
rect 12173 22933 12207 22967
rect 14565 22933 14599 22967
rect 15025 22933 15059 22967
rect 16313 22933 16347 22967
rect 16773 22933 16807 22967
rect 20177 22933 20211 22967
rect 20729 22933 20763 22967
rect 23029 22933 23063 22967
rect 24593 22933 24627 22967
rect 2697 22729 2731 22763
rect 3801 22729 3835 22763
rect 4997 22729 5031 22763
rect 6561 22729 6595 22763
rect 8769 22729 8803 22763
rect 9229 22729 9263 22763
rect 10793 22729 10827 22763
rect 11805 22729 11839 22763
rect 12265 22729 12299 22763
rect 14289 22729 14323 22763
rect 15117 22729 15151 22763
rect 16313 22729 16347 22763
rect 16681 22729 16715 22763
rect 17417 22729 17451 22763
rect 19073 22729 19107 22763
rect 19625 22729 19659 22763
rect 21465 22729 21499 22763
rect 23857 22729 23891 22763
rect 14749 22661 14783 22695
rect 18061 22661 18095 22695
rect 20729 22661 20763 22695
rect 25053 22661 25087 22695
rect 5641 22593 5675 22627
rect 5825 22593 5859 22627
rect 6193 22593 6227 22627
rect 7205 22593 7239 22627
rect 7941 22593 7975 22627
rect 9781 22593 9815 22627
rect 10333 22593 10367 22627
rect 11345 22593 11379 22627
rect 12909 22593 12943 22627
rect 13093 22593 13127 22627
rect 15669 22593 15703 22627
rect 15761 22593 15795 22627
rect 18521 22593 18555 22627
rect 18613 22593 18647 22627
rect 20177 22593 20211 22627
rect 22109 22593 22143 22627
rect 22569 22593 22603 22627
rect 24501 22593 24535 22627
rect 24685 22593 24719 22627
rect 1409 22525 1443 22559
rect 2513 22525 2547 22559
rect 3157 22525 3191 22559
rect 3617 22525 3651 22559
rect 4721 22525 4755 22559
rect 7757 22525 7791 22559
rect 9689 22525 9723 22559
rect 14105 22525 14139 22559
rect 15577 22525 15611 22559
rect 16865 22525 16899 22559
rect 19441 22525 19475 22559
rect 19993 22525 20027 22559
rect 21833 22525 21867 22559
rect 2053 22457 2087 22491
rect 5549 22457 5583 22491
rect 7849 22457 7883 22491
rect 8401 22457 8435 22491
rect 10609 22457 10643 22491
rect 11253 22457 11287 22491
rect 12817 22457 12851 22491
rect 13829 22457 13863 22491
rect 20085 22457 20119 22491
rect 23489 22457 23523 22491
rect 24409 22457 24443 22491
rect 1593 22389 1627 22423
rect 2421 22389 2455 22423
rect 3433 22389 3467 22423
rect 4261 22389 4295 22423
rect 5181 22389 5215 22423
rect 7389 22389 7423 22423
rect 9597 22389 9631 22423
rect 11161 22389 11195 22423
rect 12449 22389 12483 22423
rect 13553 22389 13587 22423
rect 15209 22389 15243 22423
rect 17049 22389 17083 22423
rect 17785 22389 17819 22423
rect 18429 22389 18463 22423
rect 21097 22389 21131 22423
rect 21925 22389 21959 22423
rect 23121 22389 23155 22423
rect 24041 22389 24075 22423
rect 2789 22185 2823 22219
rect 6929 22185 6963 22219
rect 12909 22185 12943 22219
rect 15301 22185 15335 22219
rect 16865 22185 16899 22219
rect 20729 22185 20763 22219
rect 21925 22185 21959 22219
rect 23397 22185 23431 22219
rect 23949 22185 23983 22219
rect 14105 22117 14139 22151
rect 18797 22117 18831 22151
rect 20913 22117 20947 22151
rect 21833 22117 21867 22151
rect 1961 22049 1995 22083
rect 2237 22049 2271 22083
rect 3893 22049 3927 22083
rect 5089 22049 5123 22083
rect 7288 22049 7322 22083
rect 9873 22049 9907 22083
rect 10517 22049 10551 22083
rect 11244 22049 11278 22083
rect 14013 22049 14047 22083
rect 15669 22049 15703 22083
rect 17233 22049 17267 22083
rect 19625 22049 19659 22083
rect 22293 22049 22327 22083
rect 23029 22049 23063 22083
rect 24317 22049 24351 22083
rect 5181 21981 5215 22015
rect 5365 21981 5399 22015
rect 7021 21981 7055 22015
rect 10977 21981 11011 22015
rect 14289 21981 14323 22015
rect 14473 21981 14507 22015
rect 15761 21981 15795 22015
rect 15945 21981 15979 22015
rect 16405 21981 16439 22015
rect 17325 21981 17359 22015
rect 17509 21981 17543 22015
rect 18889 21981 18923 22015
rect 19073 21981 19107 22015
rect 22385 21981 22419 22015
rect 22477 21981 22511 22015
rect 24409 21981 24443 22015
rect 24593 21981 24627 22015
rect 3157 21913 3191 21947
rect 4721 21913 4755 21947
rect 5733 21913 5767 21947
rect 10057 21913 10091 21947
rect 13553 21913 13587 21947
rect 14749 21913 14783 21947
rect 16773 21913 16807 21947
rect 21465 21913 21499 21947
rect 1593 21845 1627 21879
rect 3525 21845 3559 21879
rect 4261 21845 4295 21879
rect 6285 21845 6319 21879
rect 8401 21845 8435 21879
rect 9229 21845 9263 21879
rect 10885 21845 10919 21879
rect 12357 21845 12391 21879
rect 13645 21845 13679 21879
rect 14473 21845 14507 21879
rect 15117 21845 15151 21879
rect 18153 21845 18187 21879
rect 18429 21845 18463 21879
rect 20085 21845 20119 21879
rect 23765 21845 23799 21879
rect 2697 21641 2731 21675
rect 4261 21641 4295 21675
rect 5641 21641 5675 21675
rect 8217 21641 8251 21675
rect 10701 21641 10735 21675
rect 12265 21641 12299 21675
rect 12449 21641 12483 21675
rect 14013 21641 14047 21675
rect 17233 21641 17267 21675
rect 21189 21641 21223 21675
rect 22201 21641 22235 21675
rect 23397 21641 23431 21675
rect 25421 21641 25455 21675
rect 17785 21573 17819 21607
rect 19625 21573 19659 21607
rect 2237 21505 2271 21539
rect 3249 21505 3283 21539
rect 4721 21505 4755 21539
rect 4813 21505 4847 21539
rect 6837 21505 6871 21539
rect 9321 21505 9355 21539
rect 12909 21505 12943 21539
rect 13001 21505 13035 21539
rect 14933 21505 14967 21539
rect 18613 21505 18647 21539
rect 19533 21505 19567 21539
rect 20085 21505 20119 21539
rect 20269 21505 20303 21539
rect 20729 21505 20763 21539
rect 21833 21505 21867 21539
rect 24225 21505 24259 21539
rect 1409 21437 1443 21471
rect 3709 21437 3743 21471
rect 4169 21437 4203 21471
rect 6009 21437 6043 21471
rect 7104 21437 7138 21471
rect 9577 21437 9611 21471
rect 21557 21437 21591 21471
rect 23121 21437 23155 21471
rect 24133 21437 24167 21471
rect 25237 21437 25271 21471
rect 25789 21437 25823 21471
rect 1685 21369 1719 21403
rect 2605 21369 2639 21403
rect 3157 21369 3191 21403
rect 6653 21369 6687 21403
rect 9137 21369 9171 21403
rect 13737 21369 13771 21403
rect 14841 21369 14875 21403
rect 15200 21369 15234 21403
rect 18521 21369 18555 21403
rect 24041 21369 24075 21403
rect 25053 21369 25087 21403
rect 3065 21301 3099 21335
rect 4629 21301 4663 21335
rect 5365 21301 5399 21335
rect 8861 21301 8895 21335
rect 11345 21301 11379 21335
rect 11805 21301 11839 21335
rect 12817 21301 12851 21335
rect 14473 21301 14507 21335
rect 16313 21301 16347 21335
rect 16957 21301 16991 21335
rect 18061 21301 18095 21335
rect 18429 21301 18463 21335
rect 19073 21301 19107 21335
rect 19993 21301 20027 21335
rect 21097 21301 21131 21335
rect 21649 21301 21683 21335
rect 22569 21301 22603 21335
rect 23673 21301 23707 21335
rect 24777 21301 24811 21335
rect 2421 21097 2455 21131
rect 6929 21097 6963 21131
rect 8033 21097 8067 21131
rect 14105 21097 14139 21131
rect 14749 21097 14783 21131
rect 17233 21097 17267 21131
rect 18797 21097 18831 21131
rect 19993 21097 20027 21131
rect 23305 21097 23339 21131
rect 24317 21097 24351 21131
rect 25237 21097 25271 21131
rect 2881 21029 2915 21063
rect 5080 21029 5114 21063
rect 15577 21029 15611 21063
rect 16120 21029 16154 21063
rect 21373 21029 21407 21063
rect 24685 21029 24719 21063
rect 2789 20961 2823 20995
rect 4813 20961 4847 20995
rect 7573 20961 7607 20995
rect 8401 20961 8435 20995
rect 8493 20961 8527 20995
rect 9689 20961 9723 20995
rect 9956 20961 9990 20995
rect 11805 20961 11839 20995
rect 12725 20961 12759 20995
rect 12992 20961 13026 20995
rect 18705 20961 18739 20995
rect 21281 20961 21315 20995
rect 22017 20961 22051 20995
rect 23213 20961 23247 20995
rect 23673 20961 23707 20995
rect 2053 20893 2087 20927
rect 3065 20893 3099 20927
rect 7941 20893 7975 20927
rect 8677 20893 8711 20927
rect 9321 20893 9355 20927
rect 12173 20893 12207 20927
rect 15853 20893 15887 20927
rect 18981 20893 19015 20927
rect 21465 20893 21499 20927
rect 23765 20893 23799 20927
rect 23949 20893 23983 20927
rect 25329 20893 25363 20927
rect 25421 20893 25455 20927
rect 11069 20825 11103 20859
rect 18337 20825 18371 20859
rect 20913 20825 20947 20859
rect 22385 20825 22419 20859
rect 1593 20757 1627 20791
rect 3709 20757 3743 20791
rect 4261 20757 4295 20791
rect 4629 20757 4663 20791
rect 6193 20757 6227 20791
rect 12541 20757 12575 20791
rect 15117 20757 15151 20791
rect 18153 20757 18187 20791
rect 19625 20757 19659 20791
rect 20453 20757 20487 20791
rect 22845 20757 22879 20791
rect 24869 20757 24903 20791
rect 2697 20553 2731 20587
rect 2973 20553 3007 20587
rect 3157 20553 3191 20587
rect 4721 20553 4755 20587
rect 8309 20553 8343 20587
rect 9873 20553 9907 20587
rect 12449 20553 12483 20587
rect 13553 20553 13587 20587
rect 14657 20553 14691 20587
rect 16221 20553 16255 20587
rect 18061 20553 18095 20587
rect 19073 20553 19107 20587
rect 19625 20553 19659 20587
rect 21005 20553 21039 20587
rect 21189 20553 21223 20587
rect 22661 20553 22695 20587
rect 23673 20553 23707 20587
rect 1593 20485 1627 20519
rect 4261 20485 4295 20519
rect 7021 20485 7055 20519
rect 19441 20485 19475 20519
rect 23489 20485 23523 20519
rect 24961 20485 24995 20519
rect 25973 20485 26007 20519
rect 2237 20417 2271 20451
rect 3617 20417 3651 20451
rect 3801 20417 3835 20451
rect 5181 20417 5215 20451
rect 5273 20417 5307 20451
rect 7481 20417 7515 20451
rect 8861 20417 8895 20451
rect 9321 20417 9355 20451
rect 10425 20417 10459 20451
rect 10885 20417 10919 20451
rect 12173 20417 12207 20451
rect 13001 20417 13035 20451
rect 14565 20417 14599 20451
rect 15301 20417 15335 20451
rect 16773 20417 16807 20451
rect 17233 20417 17267 20451
rect 18705 20417 18739 20451
rect 20085 20417 20119 20451
rect 20177 20417 20211 20451
rect 21741 20417 21775 20451
rect 22201 20417 22235 20451
rect 6837 20349 6871 20383
rect 12817 20349 12851 20383
rect 13829 20349 13863 20383
rect 15025 20349 15059 20383
rect 15853 20349 15887 20383
rect 16589 20349 16623 20383
rect 18429 20349 18463 20383
rect 21557 20349 21591 20383
rect 23029 20349 23063 20383
rect 1961 20281 1995 20315
rect 3525 20281 3559 20315
rect 5089 20281 5123 20315
rect 6561 20281 6595 20315
rect 7849 20281 7883 20315
rect 8677 20281 8711 20315
rect 10333 20281 10367 20315
rect 11253 20281 11287 20315
rect 11897 20281 11931 20315
rect 12909 20281 12943 20315
rect 15117 20281 15151 20315
rect 16037 20281 16071 20315
rect 16681 20281 16715 20315
rect 18521 20281 18555 20315
rect 24133 20417 24167 20451
rect 24225 20417 24259 20451
rect 24041 20349 24075 20383
rect 25237 20349 25271 20383
rect 25513 20281 25547 20315
rect 2053 20213 2087 20247
rect 4537 20213 4571 20247
rect 5733 20213 5767 20247
rect 6193 20213 6227 20247
rect 8125 20213 8159 20247
rect 8769 20213 8803 20247
rect 9781 20213 9815 20247
rect 10241 20213 10275 20247
rect 15669 20213 15703 20247
rect 15853 20213 15887 20247
rect 17785 20213 17819 20247
rect 19993 20213 20027 20247
rect 21649 20213 21683 20247
rect 23397 20213 23431 20247
rect 23489 20213 23523 20247
rect 2421 20009 2455 20043
rect 6101 20009 6135 20043
rect 8217 20009 8251 20043
rect 8769 20009 8803 20043
rect 9965 20009 9999 20043
rect 11529 20009 11563 20043
rect 13093 20009 13127 20043
rect 14657 20009 14691 20043
rect 15025 20009 15059 20043
rect 17785 20009 17819 20043
rect 20361 20009 20395 20043
rect 20913 20009 20947 20043
rect 22477 20009 22511 20043
rect 24041 20009 24075 20043
rect 24501 20009 24535 20043
rect 25421 20009 25455 20043
rect 2789 19941 2823 19975
rect 10333 19941 10367 19975
rect 11897 19941 11931 19975
rect 13001 19941 13035 19975
rect 15660 19941 15694 19975
rect 18122 19941 18156 19975
rect 20729 19941 20763 19975
rect 21281 19941 21315 19975
rect 25789 19941 25823 19975
rect 2881 19873 2915 19907
rect 3341 19873 3375 19907
rect 3525 19873 3559 19907
rect 4333 19873 4367 19907
rect 7093 19873 7127 19907
rect 12633 19873 12667 19907
rect 13461 19873 13495 19907
rect 13553 19873 13587 19907
rect 14105 19873 14139 19907
rect 15393 19873 15427 19907
rect 17877 19873 17911 19907
rect 22845 19873 22879 19907
rect 24409 19873 24443 19907
rect 2145 19805 2179 19839
rect 3065 19805 3099 19839
rect 4077 19805 4111 19839
rect 6837 19805 6871 19839
rect 10425 19805 10459 19839
rect 10609 19805 10643 19839
rect 11989 19805 12023 19839
rect 12081 19805 12115 19839
rect 13645 19805 13679 19839
rect 21373 19805 21407 19839
rect 21465 19805 21499 19839
rect 22937 19805 22971 19839
rect 23121 19805 23155 19839
rect 24593 19805 24627 19839
rect 9505 19737 9539 19771
rect 1685 19669 1719 19703
rect 3341 19669 3375 19703
rect 3801 19669 3835 19703
rect 5457 19669 5491 19703
rect 6377 19669 6411 19703
rect 11069 19669 11103 19703
rect 11345 19669 11379 19703
rect 16773 19669 16807 19703
rect 17417 19669 17451 19703
rect 19257 19669 19291 19703
rect 19809 19669 19843 19703
rect 21925 19669 21959 19703
rect 22385 19669 22419 19703
rect 23673 19669 23707 19703
rect 25053 19669 25087 19703
rect 26249 19669 26283 19703
rect 3433 19465 3467 19499
rect 9321 19465 9355 19499
rect 9781 19465 9815 19499
rect 12817 19465 12851 19499
rect 15393 19465 15427 19499
rect 16497 19465 16531 19499
rect 21005 19465 21039 19499
rect 22569 19465 22603 19499
rect 23489 19465 23523 19499
rect 24685 19397 24719 19431
rect 2697 19329 2731 19363
rect 4169 19329 4203 19363
rect 5825 19329 5859 19363
rect 7941 19329 7975 19363
rect 8861 19329 8895 19363
rect 15945 19329 15979 19363
rect 16773 19329 16807 19363
rect 21741 19329 21775 19363
rect 24317 19329 24351 19363
rect 2421 19261 2455 19295
rect 4077 19261 4111 19295
rect 4721 19261 4755 19295
rect 5549 19261 5583 19295
rect 7205 19261 7239 19295
rect 7757 19261 7791 19295
rect 8677 19261 8711 19295
rect 9873 19261 9907 19295
rect 10140 19261 10174 19295
rect 12909 19261 12943 19295
rect 13165 19261 13199 19295
rect 16957 19261 16991 19295
rect 17509 19261 17543 19295
rect 18705 19261 18739 19295
rect 22845 19261 22879 19295
rect 24041 19261 24075 19295
rect 24133 19261 24167 19295
rect 25053 19261 25087 19295
rect 25237 19261 25271 19295
rect 25789 19261 25823 19295
rect 26249 19261 26283 19295
rect 2513 19193 2547 19227
rect 5641 19193 5675 19227
rect 7665 19193 7699 19227
rect 14933 19193 14967 19227
rect 15853 19193 15887 19227
rect 17877 19193 17911 19227
rect 18950 19193 18984 19227
rect 21649 19193 21683 19227
rect 1869 19125 1903 19159
rect 2053 19125 2087 19159
rect 3065 19125 3099 19159
rect 3617 19125 3651 19159
rect 3985 19125 4019 19159
rect 4997 19125 5031 19159
rect 5181 19125 5215 19159
rect 6193 19125 6227 19159
rect 6653 19125 6687 19159
rect 7297 19125 7331 19159
rect 8401 19125 8435 19159
rect 11253 19125 11287 19159
rect 11897 19125 11931 19159
rect 12173 19125 12207 19159
rect 14289 19125 14323 19159
rect 15301 19125 15335 19159
rect 15761 19125 15795 19159
rect 18337 19125 18371 19159
rect 20085 19125 20119 19159
rect 21189 19125 21223 19159
rect 21557 19125 21591 19159
rect 23673 19125 23707 19159
rect 25421 19125 25455 19159
rect 2421 18921 2455 18955
rect 2881 18921 2915 18955
rect 4261 18921 4295 18955
rect 6745 18921 6779 18955
rect 8585 18921 8619 18955
rect 9505 18921 9539 18955
rect 11069 18921 11103 18955
rect 13553 18921 13587 18955
rect 15117 18921 15151 18955
rect 16313 18921 16347 18955
rect 16865 18921 16899 18955
rect 18153 18921 18187 18955
rect 18429 18921 18463 18955
rect 18889 18921 18923 18955
rect 19625 18921 19659 18955
rect 20729 18921 20763 18955
rect 21925 18921 21959 18955
rect 22477 18921 22511 18955
rect 25053 18921 25087 18955
rect 2789 18853 2823 18887
rect 7297 18853 7331 18887
rect 11897 18853 11931 18887
rect 11989 18853 12023 18887
rect 18797 18853 18831 18887
rect 22937 18853 22971 18887
rect 23765 18853 23799 18887
rect 25421 18853 25455 18887
rect 4077 18785 4111 18819
rect 5641 18785 5675 18819
rect 5733 18785 5767 18819
rect 7205 18785 7239 18819
rect 8401 18785 8435 18819
rect 9945 18785 9979 18819
rect 3065 18717 3099 18751
rect 5181 18717 5215 18751
rect 5825 18717 5859 18751
rect 7389 18717 7423 18751
rect 9689 18717 9723 18751
rect 1777 18649 1811 18683
rect 3709 18649 3743 18683
rect 4721 18649 4755 18683
rect 12440 18785 12474 18819
rect 15669 18785 15703 18819
rect 17233 18785 17267 18819
rect 21281 18785 21315 18819
rect 22845 18785 22879 18819
rect 24409 18785 24443 18819
rect 12173 18717 12207 18751
rect 15761 18717 15795 18751
rect 15945 18717 15979 18751
rect 17325 18717 17359 18751
rect 17417 18717 17451 18751
rect 19073 18717 19107 18751
rect 21373 18717 21407 18751
rect 21557 18717 21591 18751
rect 23029 18717 23063 18751
rect 24501 18717 24535 18751
rect 24593 18717 24627 18751
rect 14473 18649 14507 18683
rect 2145 18581 2179 18615
rect 5273 18581 5307 18615
rect 6285 18581 6319 18615
rect 6837 18581 6871 18615
rect 7941 18581 7975 18615
rect 8309 18581 8343 18615
rect 9137 18581 9171 18615
rect 11621 18581 11655 18615
rect 11897 18581 11931 18615
rect 14197 18581 14231 18615
rect 15301 18581 15335 18615
rect 16681 18581 16715 18615
rect 20269 18581 20303 18615
rect 20913 18581 20947 18615
rect 22385 18581 22419 18615
rect 24041 18581 24075 18615
rect 25881 18581 25915 18615
rect 26157 18581 26191 18615
rect 2053 18377 2087 18411
rect 3157 18377 3191 18411
rect 3617 18377 3651 18411
rect 6285 18377 6319 18411
rect 10517 18377 10551 18411
rect 11529 18377 11563 18411
rect 12633 18377 12667 18411
rect 13369 18377 13403 18411
rect 18061 18377 18095 18411
rect 21649 18377 21683 18411
rect 22109 18377 22143 18411
rect 25053 18377 25087 18411
rect 25421 18377 25455 18411
rect 5181 18309 5215 18343
rect 12265 18309 12299 18343
rect 16865 18309 16899 18343
rect 18889 18309 18923 18343
rect 22937 18309 22971 18343
rect 2513 18241 2547 18275
rect 2697 18241 2731 18275
rect 4077 18241 4111 18275
rect 4169 18241 4203 18275
rect 5825 18241 5859 18275
rect 11069 18241 11103 18275
rect 14013 18241 14047 18275
rect 14197 18241 14231 18275
rect 15485 18241 15519 18275
rect 18613 18241 18647 18275
rect 2421 18173 2455 18207
rect 3525 18173 3559 18207
rect 4721 18173 4755 18207
rect 5549 18173 5583 18207
rect 6653 18173 6687 18207
rect 7757 18173 7791 18207
rect 10425 18173 10459 18207
rect 10885 18173 10919 18207
rect 12437 18173 12471 18207
rect 13921 18173 13955 18207
rect 14565 18173 14599 18207
rect 18429 18173 18463 18207
rect 5641 18105 5675 18139
rect 8024 18105 8058 18139
rect 15752 18105 15786 18139
rect 17509 18105 17543 18139
rect 19073 18241 19107 18275
rect 19625 18241 19659 18275
rect 24133 18241 24167 18275
rect 24225 18241 24259 18275
rect 19717 18173 19751 18207
rect 19984 18173 20018 18207
rect 22201 18173 22235 18207
rect 25237 18173 25271 18207
rect 25789 18173 25823 18207
rect 22477 18105 22511 18139
rect 24041 18105 24075 18139
rect 1685 18037 1719 18071
rect 3985 18037 4019 18071
rect 5089 18037 5123 18071
rect 7113 18037 7147 18071
rect 7665 18037 7699 18071
rect 9137 18037 9171 18071
rect 10057 18037 10091 18071
rect 10977 18037 11011 18071
rect 13001 18037 13035 18071
rect 13553 18037 13587 18071
rect 14933 18037 14967 18071
rect 15393 18037 15427 18071
rect 17877 18037 17911 18071
rect 18521 18037 18555 18071
rect 18889 18037 18923 18071
rect 21097 18037 21131 18071
rect 23489 18037 23523 18071
rect 23673 18037 23707 18071
rect 24685 18037 24719 18071
rect 26249 18037 26283 18071
rect 2421 17833 2455 17867
rect 3433 17833 3467 17867
rect 5549 17833 5583 17867
rect 6561 17833 6595 17867
rect 7113 17833 7147 17867
rect 10701 17833 10735 17867
rect 11253 17833 11287 17867
rect 14105 17833 14139 17867
rect 15025 17833 15059 17867
rect 15301 17833 15335 17867
rect 18337 17833 18371 17867
rect 20269 17833 20303 17867
rect 22109 17833 22143 17867
rect 22477 17833 22511 17867
rect 24593 17833 24627 17867
rect 26341 17833 26375 17867
rect 6193 17765 6227 17799
rect 8493 17765 8527 17799
rect 11069 17765 11103 17799
rect 11621 17765 11655 17799
rect 11713 17765 11747 17799
rect 12909 17765 12943 17799
rect 13277 17765 13311 17799
rect 14013 17765 14047 17799
rect 17202 17765 17236 17799
rect 23673 17765 23707 17799
rect 2789 17697 2823 17731
rect 4436 17697 4470 17731
rect 7021 17697 7055 17731
rect 8217 17697 8251 17731
rect 10057 17697 10091 17731
rect 10149 17697 10183 17731
rect 15669 17697 15703 17731
rect 16957 17697 16991 17731
rect 19533 17697 19567 17731
rect 20729 17697 20763 17731
rect 21373 17697 21407 17731
rect 22937 17697 22971 17731
rect 24501 17697 24535 17731
rect 1409 17629 1443 17663
rect 2881 17629 2915 17663
rect 3065 17629 3099 17663
rect 4169 17629 4203 17663
rect 7205 17629 7239 17663
rect 10241 17629 10275 17663
rect 11805 17629 11839 17663
rect 14289 17629 14323 17663
rect 15761 17629 15795 17663
rect 15945 17629 15979 17663
rect 19717 17629 19751 17663
rect 21465 17629 21499 17663
rect 21649 17629 21683 17663
rect 23029 17629 23063 17663
rect 23121 17629 23155 17663
rect 24685 17629 24719 17663
rect 7757 17561 7791 17595
rect 9321 17561 9355 17595
rect 13645 17561 13679 17595
rect 14749 17561 14783 17595
rect 19349 17561 19383 17595
rect 22569 17561 22603 17595
rect 24133 17561 24167 17595
rect 1961 17493 1995 17527
rect 2329 17493 2363 17527
rect 3801 17493 3835 17527
rect 6653 17493 6687 17527
rect 8125 17493 8159 17527
rect 8953 17493 8987 17527
rect 9689 17493 9723 17527
rect 12541 17493 12575 17527
rect 16313 17493 16347 17527
rect 16773 17493 16807 17527
rect 18981 17493 19015 17527
rect 21005 17493 21039 17527
rect 25145 17493 25179 17527
rect 25605 17493 25639 17527
rect 25881 17493 25915 17527
rect 2789 17289 2823 17323
rect 5733 17289 5767 17323
rect 6653 17289 6687 17323
rect 8217 17289 8251 17323
rect 11437 17289 11471 17323
rect 14565 17289 14599 17323
rect 16129 17289 16163 17323
rect 16957 17289 16991 17323
rect 18061 17289 18095 17323
rect 19717 17289 19751 17323
rect 19993 17289 20027 17323
rect 23673 17289 23707 17323
rect 24685 17289 24719 17323
rect 25053 17289 25087 17323
rect 4629 17221 4663 17255
rect 10425 17221 10459 17255
rect 17233 17221 17267 17255
rect 23489 17221 23523 17255
rect 2053 17153 2087 17187
rect 3709 17153 3743 17187
rect 5181 17153 5215 17187
rect 5273 17153 5307 17187
rect 6193 17153 6227 17187
rect 8861 17153 8895 17187
rect 9873 17153 9907 17187
rect 10701 17153 10735 17187
rect 12265 17153 12299 17187
rect 13001 17153 13035 17187
rect 14749 17153 14783 17187
rect 18705 17153 18739 17187
rect 24225 17153 24259 17187
rect 1777 17085 1811 17119
rect 6837 17085 6871 17119
rect 7104 17085 7138 17119
rect 9689 17085 9723 17119
rect 10885 17085 10919 17119
rect 12909 17085 12943 17119
rect 17417 17085 17451 17119
rect 18429 17085 18463 17119
rect 19809 17085 19843 17119
rect 20913 17085 20947 17119
rect 24133 17085 24167 17119
rect 25237 17085 25271 17119
rect 2513 17017 2547 17051
rect 5089 17017 5123 17051
rect 9781 17017 9815 17051
rect 11897 17017 11931 17051
rect 12817 17017 12851 17051
rect 13737 17017 13771 17051
rect 14289 17017 14323 17051
rect 15016 17017 15050 17051
rect 17877 17017 17911 17051
rect 20821 17017 20855 17051
rect 21158 17017 21192 17051
rect 24041 17017 24075 17051
rect 1409 16949 1443 16983
rect 1869 16949 1903 16983
rect 3157 16949 3191 16983
rect 3525 16949 3559 16983
rect 3617 16949 3651 16983
rect 4261 16949 4295 16983
rect 4721 16949 4755 16983
rect 9137 16949 9171 16983
rect 9321 16949 9355 16983
rect 11069 16949 11103 16983
rect 12449 16949 12483 16983
rect 18521 16949 18555 16983
rect 19073 16949 19107 16983
rect 20453 16949 20487 16983
rect 22293 16949 22327 16983
rect 22937 16949 22971 16983
rect 25421 16949 25455 16983
rect 25789 16949 25823 16983
rect 26157 16949 26191 16983
rect 2513 16745 2547 16779
rect 2973 16745 3007 16779
rect 3525 16745 3559 16779
rect 4537 16745 4571 16779
rect 5641 16745 5675 16779
rect 7665 16745 7699 16779
rect 9689 16745 9723 16779
rect 10057 16745 10091 16779
rect 11529 16745 11563 16779
rect 13093 16745 13127 16779
rect 13645 16745 13679 16779
rect 14013 16745 14047 16779
rect 14197 16745 14231 16779
rect 14749 16745 14783 16779
rect 15485 16745 15519 16779
rect 16589 16745 16623 16779
rect 17233 16745 17267 16779
rect 18061 16745 18095 16779
rect 20085 16745 20119 16779
rect 22293 16745 22327 16779
rect 22937 16745 22971 16779
rect 23213 16745 23247 16779
rect 23397 16745 23431 16779
rect 23857 16745 23891 16779
rect 24409 16745 24443 16779
rect 1777 16677 1811 16711
rect 5549 16677 5583 16711
rect 9321 16677 9355 16711
rect 15117 16677 15151 16711
rect 21180 16677 21214 16711
rect 25237 16677 25271 16711
rect 1869 16609 1903 16643
rect 2789 16609 2823 16643
rect 3801 16609 3835 16643
rect 4445 16609 4479 16643
rect 6009 16609 6043 16643
rect 6101 16609 6135 16643
rect 7573 16609 7607 16643
rect 8309 16609 8343 16643
rect 10149 16609 10183 16643
rect 11980 16609 12014 16643
rect 15853 16609 15887 16643
rect 17049 16609 17083 16643
rect 18420 16609 18454 16643
rect 20729 16609 20763 16643
rect 23765 16609 23799 16643
rect 24961 16609 24995 16643
rect 25697 16609 25731 16643
rect 2053 16541 2087 16575
rect 4629 16541 4663 16575
rect 6285 16541 6319 16575
rect 7757 16541 7791 16575
rect 10333 16541 10367 16575
rect 11713 16541 11747 16575
rect 15945 16541 15979 16575
rect 16037 16541 16071 16575
rect 18153 16541 18187 16575
rect 20913 16541 20947 16575
rect 24041 16541 24075 16575
rect 5089 16473 5123 16507
rect 11069 16473 11103 16507
rect 16957 16473 16991 16507
rect 1409 16405 1443 16439
rect 4077 16405 4111 16439
rect 6745 16405 6779 16439
rect 7021 16405 7055 16439
rect 7205 16405 7239 16439
rect 8769 16405 8803 16439
rect 10701 16405 10735 16439
rect 17693 16405 17727 16439
rect 19533 16405 19567 16439
rect 24777 16405 24811 16439
rect 26065 16405 26099 16439
rect 8677 16201 8711 16235
rect 9781 16201 9815 16235
rect 10241 16201 10275 16235
rect 11253 16201 11287 16235
rect 12449 16201 12483 16235
rect 13553 16201 13587 16235
rect 14473 16201 14507 16235
rect 15945 16201 15979 16235
rect 16497 16201 16531 16235
rect 17049 16201 17083 16235
rect 17509 16201 17543 16235
rect 20729 16201 20763 16235
rect 23121 16201 23155 16235
rect 24685 16201 24719 16235
rect 25053 16201 25087 16235
rect 2697 16133 2731 16167
rect 4721 16133 4755 16167
rect 6193 16133 6227 16167
rect 11805 16133 11839 16167
rect 23673 16133 23707 16167
rect 2053 16065 2087 16099
rect 3709 16065 3743 16099
rect 5273 16065 5307 16099
rect 7665 16065 7699 16099
rect 9137 16065 9171 16099
rect 9321 16065 9355 16099
rect 10793 16065 10827 16099
rect 11989 16065 12023 16099
rect 12265 16065 12299 16099
rect 13001 16065 13035 16099
rect 14565 16065 14599 16099
rect 20637 16065 20671 16099
rect 21373 16065 21407 16099
rect 24225 16065 24259 16099
rect 4169 15997 4203 16031
rect 4537 15997 4571 16031
rect 5181 15997 5215 16031
rect 6469 15997 6503 16031
rect 10609 15997 10643 16031
rect 1777 15929 1811 15963
rect 3065 15929 3099 15963
rect 5825 15929 5859 15963
rect 7481 15929 7515 15963
rect 8217 15929 8251 15963
rect 10057 15929 10091 15963
rect 13829 15997 13863 16031
rect 17785 15997 17819 16031
rect 18061 15997 18095 16031
rect 21097 15997 21131 16031
rect 21833 15997 21867 16031
rect 22477 15997 22511 16031
rect 25237 15997 25271 16031
rect 25973 15997 26007 16031
rect 14810 15929 14844 15963
rect 18328 15929 18362 15963
rect 20269 15929 20303 15963
rect 21189 15929 21223 15963
rect 24041 15929 24075 15963
rect 25513 15929 25547 15963
rect 1409 15861 1443 15895
rect 1869 15861 1903 15895
rect 3157 15861 3191 15895
rect 3525 15861 3559 15895
rect 3617 15861 3651 15895
rect 5089 15861 5123 15895
rect 6285 15861 6319 15895
rect 7113 15861 7147 15895
rect 7573 15861 7607 15895
rect 8585 15861 8619 15895
rect 9045 15861 9079 15895
rect 10701 15861 10735 15895
rect 11989 15861 12023 15895
rect 12817 15861 12851 15895
rect 12909 15861 12943 15895
rect 17601 15861 17635 15895
rect 19441 15861 19475 15895
rect 22293 15861 22327 15895
rect 22661 15861 22695 15895
rect 23489 15861 23523 15895
rect 24133 15861 24167 15895
rect 26341 15861 26375 15895
rect 2697 15657 2731 15691
rect 4537 15657 4571 15691
rect 5181 15657 5215 15691
rect 5733 15657 5767 15691
rect 6101 15657 6135 15691
rect 8585 15657 8619 15691
rect 9229 15657 9263 15691
rect 9689 15657 9723 15691
rect 10333 15657 10367 15691
rect 12081 15657 12115 15691
rect 13185 15657 13219 15691
rect 14289 15657 14323 15691
rect 16589 15657 16623 15691
rect 19625 15657 19659 15691
rect 20361 15657 20395 15691
rect 21925 15657 21959 15691
rect 22477 15657 22511 15691
rect 22845 15657 22879 15691
rect 24041 15657 24075 15691
rect 25053 15657 25087 15691
rect 26249 15657 26283 15691
rect 2605 15589 2639 15623
rect 3709 15589 3743 15623
rect 6530 15589 6564 15623
rect 8309 15589 8343 15623
rect 10968 15589 11002 15623
rect 13553 15589 13587 15623
rect 15853 15589 15887 15623
rect 21373 15589 21407 15623
rect 22385 15589 22419 15623
rect 24409 15589 24443 15623
rect 5089 15521 5123 15555
rect 8953 15521 8987 15555
rect 10701 15521 10735 15555
rect 16497 15521 16531 15555
rect 18061 15521 18095 15555
rect 21281 15521 21315 15555
rect 22937 15521 22971 15555
rect 2789 15453 2823 15487
rect 3249 15453 3283 15487
rect 5273 15453 5307 15487
rect 6285 15453 6319 15487
rect 13645 15453 13679 15487
rect 13737 15453 13771 15487
rect 16681 15453 16715 15487
rect 17601 15453 17635 15487
rect 18153 15453 18187 15487
rect 18337 15453 18371 15487
rect 19717 15453 19751 15487
rect 19809 15453 19843 15487
rect 21465 15453 21499 15487
rect 23029 15453 23063 15487
rect 23765 15453 23799 15487
rect 24501 15453 24535 15487
rect 24685 15453 24719 15487
rect 2237 15385 2271 15419
rect 4721 15385 4755 15419
rect 8769 15385 8803 15419
rect 16129 15385 16163 15419
rect 17141 15385 17175 15419
rect 19257 15385 19291 15419
rect 20729 15385 20763 15419
rect 25421 15385 25455 15419
rect 1685 15317 1719 15351
rect 2053 15317 2087 15351
rect 7665 15317 7699 15351
rect 12725 15317 12759 15351
rect 13001 15317 13035 15351
rect 14657 15317 14691 15351
rect 14933 15317 14967 15351
rect 15485 15317 15519 15351
rect 17693 15317 17727 15351
rect 18797 15317 18831 15351
rect 19165 15317 19199 15351
rect 20913 15317 20947 15351
rect 25789 15317 25823 15351
rect 4813 15113 4847 15147
rect 11253 15113 11287 15147
rect 12449 15113 12483 15147
rect 16221 15113 16255 15147
rect 19441 15113 19475 15147
rect 20453 15113 20487 15147
rect 22385 15113 22419 15147
rect 23029 15113 23063 15147
rect 24685 15113 24719 15147
rect 26341 15113 26375 15147
rect 2329 15045 2363 15079
rect 9137 15045 9171 15079
rect 23397 15045 23431 15079
rect 13001 14977 13035 15011
rect 18061 14977 18095 15011
rect 19993 14977 20027 15011
rect 24133 14977 24167 15011
rect 24225 14977 24259 15011
rect 1501 14909 1535 14943
rect 2789 14909 2823 14943
rect 5273 14909 5307 14943
rect 6837 14909 6871 14943
rect 7093 14909 7127 14943
rect 9321 14909 9355 14943
rect 9577 14909 9611 14943
rect 12173 14909 12207 14943
rect 14013 14909 14047 14943
rect 16865 14909 16899 14943
rect 17509 14909 17543 14943
rect 17877 14909 17911 14943
rect 18328 14909 18362 14943
rect 20729 14909 20763 14943
rect 21005 14909 21039 14943
rect 25053 14909 25087 14943
rect 25237 14909 25271 14943
rect 25973 14909 26007 14943
rect 1777 14841 1811 14875
rect 2697 14841 2731 14875
rect 3034 14841 3068 14875
rect 5549 14841 5583 14875
rect 8769 14841 8803 14875
rect 12909 14841 12943 14875
rect 14280 14841 14314 14875
rect 21250 14841 21284 14875
rect 25513 14841 25547 14875
rect 4169 14773 4203 14807
rect 5089 14773 5123 14807
rect 6285 14773 6319 14807
rect 6561 14773 6595 14807
rect 8217 14773 8251 14807
rect 10701 14773 10735 14807
rect 11805 14773 11839 14807
rect 12817 14773 12851 14807
rect 13553 14773 13587 14807
rect 13921 14773 13955 14807
rect 15393 14773 15427 14807
rect 16497 14773 16531 14807
rect 17049 14773 17083 14807
rect 20545 14773 20579 14807
rect 23673 14773 23707 14807
rect 24041 14773 24075 14807
rect 1409 14569 1443 14603
rect 2513 14569 2547 14603
rect 3433 14569 3467 14603
rect 6009 14569 6043 14603
rect 6929 14569 6963 14603
rect 9045 14569 9079 14603
rect 9229 14569 9263 14603
rect 10057 14569 10091 14603
rect 11805 14569 11839 14603
rect 13369 14569 13403 14603
rect 15393 14569 15427 14603
rect 16865 14569 16899 14603
rect 17969 14569 18003 14603
rect 19349 14569 19383 14603
rect 19901 14569 19935 14603
rect 20361 14569 20395 14603
rect 20729 14569 20763 14603
rect 21741 14569 21775 14603
rect 22569 14569 22603 14603
rect 23397 14569 23431 14603
rect 25881 14569 25915 14603
rect 26249 14569 26283 14603
rect 1777 14501 1811 14535
rect 7021 14501 7055 14535
rect 7573 14501 7607 14535
rect 8033 14501 8067 14535
rect 10692 14501 10726 14535
rect 17785 14501 17819 14535
rect 22845 14501 22879 14535
rect 23673 14501 23707 14535
rect 24124 14501 24158 14535
rect 4077 14433 4111 14467
rect 4344 14433 4378 14467
rect 8125 14433 8159 14467
rect 9413 14433 9447 14467
rect 13277 14433 13311 14467
rect 16773 14433 16807 14467
rect 18337 14433 18371 14467
rect 19717 14433 19751 14467
rect 21649 14433 21683 14467
rect 1869 14365 1903 14399
rect 2053 14365 2087 14399
rect 2973 14365 3007 14399
rect 6469 14365 6503 14399
rect 7205 14365 7239 14399
rect 10425 14365 10459 14399
rect 12449 14365 12483 14399
rect 13461 14365 13495 14399
rect 16221 14365 16255 14399
rect 17049 14365 17083 14399
rect 18429 14365 18463 14399
rect 18613 14365 18647 14399
rect 21833 14365 21867 14399
rect 23857 14365 23891 14399
rect 3801 14297 3835 14331
rect 6561 14297 6595 14331
rect 12817 14297 12851 14331
rect 16405 14297 16439 14331
rect 21281 14297 21315 14331
rect 2881 14229 2915 14263
rect 5457 14229 5491 14263
rect 8309 14229 8343 14263
rect 8769 14229 8803 14263
rect 12909 14229 12943 14263
rect 14013 14229 14047 14263
rect 14289 14229 14323 14263
rect 14657 14229 14691 14263
rect 15117 14229 15151 14263
rect 21189 14229 21223 14263
rect 25237 14229 25271 14263
rect 2973 14025 3007 14059
rect 3525 14025 3559 14059
rect 4261 14025 4295 14059
rect 5181 14025 5215 14059
rect 8493 14025 8527 14059
rect 10057 14025 10091 14059
rect 11069 14025 11103 14059
rect 13001 14025 13035 14059
rect 14473 14025 14507 14059
rect 15209 14025 15243 14059
rect 17417 14025 17451 14059
rect 20821 14025 20855 14059
rect 22661 14025 22695 14059
rect 23489 14025 23523 14059
rect 25053 14025 25087 14059
rect 25697 14025 25731 14059
rect 26065 14025 26099 14059
rect 26341 14025 26375 14059
rect 4721 13957 4755 13991
rect 6837 13957 6871 13991
rect 8401 13957 8435 13991
rect 16129 13957 16163 13991
rect 16221 13957 16255 13991
rect 20361 13957 20395 13991
rect 22293 13957 22327 13991
rect 1593 13889 1627 13923
rect 5641 13889 5675 13923
rect 5825 13889 5859 13923
rect 6653 13889 6687 13923
rect 7297 13889 7331 13923
rect 7389 13889 7423 13923
rect 7849 13889 7883 13923
rect 8953 13889 8987 13923
rect 9137 13889 9171 13923
rect 10609 13889 10643 13923
rect 11805 13889 11839 13923
rect 15577 13889 15611 13923
rect 15945 13889 15979 13923
rect 1860 13821 1894 13855
rect 4077 13821 4111 13855
rect 5089 13821 5123 13855
rect 6193 13821 6227 13855
rect 9597 13821 9631 13855
rect 10517 13821 10551 13855
rect 11437 13821 11471 13855
rect 13093 13821 13127 13855
rect 13360 13821 13394 13855
rect 16957 13889 16991 13923
rect 20729 13889 20763 13923
rect 21373 13889 21407 13923
rect 16865 13821 16899 13855
rect 17785 13821 17819 13855
rect 18061 13821 18095 13855
rect 18317 13821 18351 13855
rect 21189 13821 21223 13855
rect 21281 13821 21315 13855
rect 21925 13821 21959 13855
rect 22477 13821 22511 13855
rect 23673 13821 23707 13855
rect 23940 13821 23974 13855
rect 3893 13753 3927 13787
rect 12173 13753 12207 13787
rect 16129 13753 16163 13787
rect 5549 13685 5583 13719
rect 7205 13685 7239 13719
rect 8861 13685 8895 13719
rect 9965 13685 9999 13719
rect 10425 13685 10459 13719
rect 16405 13685 16439 13719
rect 16773 13685 16807 13719
rect 19441 13685 19475 13719
rect 23121 13685 23155 13719
rect 4721 13481 4755 13515
rect 5733 13481 5767 13515
rect 6193 13481 6227 13515
rect 7665 13481 7699 13515
rect 8585 13481 8619 13515
rect 9229 13481 9263 13515
rect 12173 13481 12207 13515
rect 12633 13481 12667 13515
rect 13369 13481 13403 13515
rect 17325 13481 17359 13515
rect 17785 13481 17819 13515
rect 18153 13481 18187 13515
rect 19533 13481 19567 13515
rect 19901 13481 19935 13515
rect 21189 13481 21223 13515
rect 21649 13481 21683 13515
rect 23489 13481 23523 13515
rect 24041 13481 24075 13515
rect 24961 13481 24995 13515
rect 26065 13481 26099 13515
rect 5089 13413 5123 13447
rect 6552 13413 6586 13447
rect 8861 13413 8895 13447
rect 9956 13413 9990 13447
rect 11989 13413 12023 13447
rect 13645 13413 13679 13447
rect 14933 13413 14967 13447
rect 17693 13413 17727 13447
rect 18797 13413 18831 13447
rect 20269 13413 20303 13447
rect 21925 13413 21959 13447
rect 22354 13413 22388 13447
rect 1409 13345 1443 13379
rect 1676 13345 1710 13379
rect 4629 13345 4663 13379
rect 6285 13345 6319 13379
rect 9689 13345 9723 13379
rect 12541 13345 12575 13379
rect 14013 13345 14047 13379
rect 15301 13345 15335 13379
rect 15568 13345 15602 13379
rect 18245 13345 18279 13379
rect 19165 13345 19199 13379
rect 19717 13345 19751 13379
rect 21005 13345 21039 13379
rect 22109 13345 22143 13379
rect 5181 13277 5215 13311
rect 5273 13277 5307 13311
rect 12817 13277 12851 13311
rect 14197 13277 14231 13311
rect 18429 13277 18463 13311
rect 20729 13277 20763 13311
rect 25053 13277 25087 13311
rect 25145 13277 25179 13311
rect 11621 13209 11655 13243
rect 2789 13141 2823 13175
rect 3341 13141 3375 13175
rect 3709 13141 3743 13175
rect 11069 13141 11103 13175
rect 16681 13141 16715 13175
rect 24501 13141 24535 13175
rect 24593 13141 24627 13175
rect 25605 13141 25639 13175
rect 3985 12937 4019 12971
rect 4905 12937 4939 12971
rect 6653 12937 6687 12971
rect 6837 12937 6871 12971
rect 6929 12937 6963 12971
rect 9873 12937 9907 12971
rect 10425 12937 10459 12971
rect 11805 12937 11839 12971
rect 12265 12937 12299 12971
rect 14841 12937 14875 12971
rect 16405 12937 16439 12971
rect 17509 12937 17543 12971
rect 17877 12937 17911 12971
rect 18429 12937 18463 12971
rect 21005 12937 21039 12971
rect 24777 12937 24811 12971
rect 25973 12937 26007 12971
rect 26341 12937 26375 12971
rect 4353 12869 4387 12903
rect 4629 12869 4663 12903
rect 1593 12801 1627 12835
rect 5457 12801 5491 12835
rect 6285 12733 6319 12767
rect 1860 12665 1894 12699
rect 4629 12665 4663 12699
rect 5365 12665 5399 12699
rect 7941 12869 7975 12903
rect 14657 12869 14691 12903
rect 20453 12869 20487 12903
rect 23673 12869 23707 12903
rect 7573 12801 7607 12835
rect 11345 12801 11379 12835
rect 12909 12801 12943 12835
rect 13001 12801 13035 12835
rect 13737 12801 13771 12835
rect 13829 12801 13863 12835
rect 14289 12801 14323 12835
rect 15393 12801 15427 12835
rect 16221 12801 16255 12835
rect 17049 12801 17083 12835
rect 21465 12801 21499 12835
rect 21649 12801 21683 12835
rect 22385 12801 22419 12835
rect 22569 12801 22603 12835
rect 24225 12801 24259 12835
rect 25053 12801 25087 12835
rect 25513 12801 25547 12835
rect 7297 12733 7331 12767
rect 8309 12733 8343 12767
rect 8493 12733 8527 12767
rect 12817 12733 12851 12767
rect 13645 12733 13679 12767
rect 15301 12733 15335 12767
rect 16773 12733 16807 12767
rect 18521 12733 18555 12767
rect 18777 12733 18811 12767
rect 24041 12733 24075 12767
rect 25237 12733 25271 12767
rect 8738 12665 8772 12699
rect 11161 12665 11195 12699
rect 15945 12665 15979 12699
rect 16865 12665 16899 12699
rect 23489 12665 23523 12699
rect 2973 12597 3007 12631
rect 3525 12597 3559 12631
rect 4721 12597 4755 12631
rect 5273 12597 5307 12631
rect 6837 12597 6871 12631
rect 7389 12597 7423 12631
rect 10793 12597 10827 12631
rect 12449 12597 12483 12631
rect 13277 12597 13311 12631
rect 15209 12597 15243 12631
rect 19901 12597 19935 12631
rect 20821 12597 20855 12631
rect 21373 12597 21407 12631
rect 22017 12597 22051 12631
rect 23121 12597 23155 12631
rect 24133 12597 24167 12631
rect 1409 12393 1443 12427
rect 2881 12393 2915 12427
rect 3433 12393 3467 12427
rect 4261 12393 4295 12427
rect 6837 12393 6871 12427
rect 7757 12393 7791 12427
rect 9137 12393 9171 12427
rect 10885 12393 10919 12427
rect 12081 12393 12115 12427
rect 12541 12393 12575 12427
rect 15117 12393 15151 12427
rect 15577 12393 15611 12427
rect 22201 12393 22235 12427
rect 22845 12393 22879 12427
rect 25145 12393 25179 12427
rect 26157 12393 26191 12427
rect 2329 12325 2363 12359
rect 5724 12325 5758 12359
rect 9873 12325 9907 12359
rect 10425 12325 10459 12359
rect 16304 12325 16338 12359
rect 2789 12257 2823 12291
rect 3801 12257 3835 12291
rect 4077 12257 4111 12291
rect 5457 12257 5491 12291
rect 8401 12257 8435 12291
rect 9505 12257 9539 12291
rect 11253 12257 11287 12291
rect 11345 12257 11379 12291
rect 12633 12257 12667 12291
rect 14473 12257 14507 12291
rect 16037 12257 16071 12291
rect 18061 12257 18095 12291
rect 18705 12257 18739 12291
rect 19533 12257 19567 12291
rect 21281 12257 21315 12291
rect 22661 12257 22695 12291
rect 23765 12257 23799 12291
rect 24032 12257 24066 12291
rect 3065 12189 3099 12223
rect 8493 12189 8527 12223
rect 8677 12189 8711 12223
rect 11437 12189 11471 12223
rect 19625 12189 19659 12223
rect 19809 12189 19843 12223
rect 20729 12189 20763 12223
rect 21373 12189 21407 12223
rect 21557 12189 21591 12223
rect 22569 12189 22603 12223
rect 23213 12189 23247 12223
rect 1869 12121 1903 12155
rect 2421 12121 2455 12155
rect 10793 12121 10827 12155
rect 13921 12121 13955 12155
rect 4997 12053 5031 12087
rect 5365 12053 5399 12087
rect 7389 12053 7423 12087
rect 8033 12053 8067 12087
rect 14657 12053 14691 12087
rect 15945 12053 15979 12087
rect 17417 12053 17451 12087
rect 18981 12053 19015 12087
rect 19165 12053 19199 12087
rect 20177 12053 20211 12087
rect 20913 12053 20947 12087
rect 23673 12053 23707 12087
rect 25697 12053 25731 12087
rect 1593 11849 1627 11883
rect 5549 11849 5583 11883
rect 9229 11849 9263 11883
rect 10333 11849 10367 11883
rect 10425 11849 10459 11883
rect 11897 11849 11931 11883
rect 16405 11849 16439 11883
rect 17509 11849 17543 11883
rect 22569 11849 22603 11883
rect 23673 11849 23707 11883
rect 25421 11849 25455 11883
rect 2513 11781 2547 11815
rect 3065 11713 3099 11747
rect 3157 11713 3191 11747
rect 6653 11713 6687 11747
rect 7297 11713 7331 11747
rect 7389 11713 7423 11747
rect 8953 11713 8987 11747
rect 1409 11645 1443 11679
rect 1961 11645 1995 11679
rect 4169 11645 4203 11679
rect 13921 11781 13955 11815
rect 23489 11781 23523 11815
rect 10701 11713 10735 11747
rect 11345 11713 11379 11747
rect 16957 11713 16991 11747
rect 18613 11713 18647 11747
rect 20453 11713 20487 11747
rect 20545 11713 20579 11747
rect 21465 11713 21499 11747
rect 22017 11713 22051 11747
rect 22109 11713 22143 11747
rect 24225 11713 24259 11747
rect 9413 11645 9447 11679
rect 10425 11645 10459 11679
rect 11161 11645 11195 11679
rect 12541 11645 12575 11679
rect 15301 11645 15335 11679
rect 17785 11645 17819 11679
rect 18521 11645 18555 11679
rect 19901 11645 19935 11679
rect 21925 11645 21959 11679
rect 23121 11645 23155 11679
rect 25237 11645 25271 11679
rect 25789 11645 25823 11679
rect 4436 11577 4470 11611
rect 7205 11577 7239 11611
rect 8769 11577 8803 11611
rect 8861 11577 8895 11611
rect 9229 11577 9263 11611
rect 9965 11577 9999 11611
rect 11253 11577 11287 11611
rect 12173 11577 12207 11611
rect 12808 11577 12842 11611
rect 15209 11577 15243 11611
rect 15945 11577 15979 11611
rect 16865 11577 16899 11611
rect 18429 11577 18463 11611
rect 19257 11577 19291 11611
rect 20361 11577 20395 11611
rect 24133 11577 24167 11611
rect 24685 11577 24719 11611
rect 2605 11509 2639 11543
rect 2973 11509 3007 11543
rect 3617 11509 3651 11543
rect 4077 11509 4111 11543
rect 6193 11509 6227 11543
rect 6837 11509 6871 11543
rect 7849 11509 7883 11543
rect 8217 11509 8251 11543
rect 8401 11509 8435 11543
rect 10793 11509 10827 11543
rect 14565 11509 14599 11543
rect 15485 11509 15519 11543
rect 16313 11509 16347 11543
rect 16773 11509 16807 11543
rect 18061 11509 18095 11543
rect 19993 11509 20027 11543
rect 21097 11509 21131 11543
rect 21557 11509 21591 11543
rect 24041 11509 24075 11543
rect 25053 11509 25087 11543
rect 26157 11509 26191 11543
rect 2421 11305 2455 11339
rect 2881 11305 2915 11339
rect 3893 11305 3927 11339
rect 6009 11305 6043 11339
rect 6561 11305 6595 11339
rect 7757 11305 7791 11339
rect 8585 11305 8619 11339
rect 9413 11305 9447 11339
rect 10701 11305 10735 11339
rect 13185 11305 13219 11339
rect 17049 11305 17083 11339
rect 20361 11305 20395 11339
rect 21925 11305 21959 11339
rect 22293 11305 22327 11339
rect 22661 11305 22695 11339
rect 23121 11305 23155 11339
rect 25053 11305 25087 11339
rect 25697 11305 25731 11339
rect 26065 11305 26099 11339
rect 2329 11237 2363 11271
rect 3525 11237 3559 11271
rect 6929 11237 6963 11271
rect 8493 11237 8527 11271
rect 14013 11237 14047 11271
rect 18604 11237 18638 11271
rect 23940 11237 23974 11271
rect 2789 11169 2823 11203
rect 4077 11169 4111 11203
rect 4344 11169 4378 11203
rect 9045 11169 9079 11203
rect 10609 11169 10643 11203
rect 11805 11169 11839 11203
rect 12072 11169 12106 11203
rect 15936 11169 15970 11203
rect 17693 11169 17727 11203
rect 21281 11169 21315 11203
rect 21373 11169 21407 11203
rect 22477 11169 22511 11203
rect 23673 11169 23707 11203
rect 1409 11101 1443 11135
rect 3065 11101 3099 11135
rect 7021 11101 7055 11135
rect 7113 11101 7147 11135
rect 10885 11101 10919 11135
rect 15669 11101 15703 11135
rect 18337 11101 18371 11135
rect 21557 11101 21591 11135
rect 1961 11033 1995 11067
rect 5457 11033 5491 11067
rect 8125 11033 8159 11067
rect 9873 11033 9907 11067
rect 10241 11033 10275 11067
rect 11253 11033 11287 11067
rect 15485 11033 15519 11067
rect 18061 11033 18095 11067
rect 19717 11033 19751 11067
rect 20913 11033 20947 11067
rect 6377 10965 6411 10999
rect 11713 10965 11747 10999
rect 14381 10965 14415 10999
rect 14749 10965 14783 10999
rect 20729 10965 20763 10999
rect 23397 10965 23431 10999
rect 1409 10761 1443 10795
rect 2513 10761 2547 10795
rect 5365 10761 5399 10795
rect 6285 10761 6319 10795
rect 7941 10761 7975 10795
rect 10425 10761 10459 10795
rect 11069 10761 11103 10795
rect 11345 10761 11379 10795
rect 12173 10761 12207 10795
rect 13461 10761 13495 10795
rect 15577 10761 15611 10795
rect 16405 10761 16439 10795
rect 19533 10761 19567 10795
rect 21005 10761 21039 10795
rect 22477 10761 22511 10795
rect 23029 10761 23063 10795
rect 23489 10761 23523 10795
rect 25053 10761 25087 10795
rect 5733 10693 5767 10727
rect 8217 10693 8251 10727
rect 11897 10693 11931 10727
rect 13829 10693 13863 10727
rect 14013 10693 14047 10727
rect 15025 10693 15059 10727
rect 19349 10693 19383 10727
rect 20545 10693 20579 10727
rect 21097 10693 21131 10727
rect 2053 10625 2087 10659
rect 7297 10625 7331 10659
rect 7389 10625 7423 10659
rect 8953 10625 8987 10659
rect 13093 10625 13127 10659
rect 14473 10625 14507 10659
rect 14565 10625 14599 10659
rect 16957 10625 16991 10659
rect 17417 10625 17451 10659
rect 18245 10625 18279 10659
rect 20085 10625 20119 10659
rect 21557 10625 21591 10659
rect 21741 10625 21775 10659
rect 22109 10625 22143 10659
rect 1777 10557 1811 10591
rect 1869 10557 1903 10591
rect 3065 10557 3099 10591
rect 5549 10557 5583 10591
rect 6653 10557 6687 10591
rect 9045 10557 9079 10591
rect 9312 10557 9346 10591
rect 12817 10557 12851 10591
rect 15945 10557 15979 10591
rect 17877 10557 17911 10591
rect 18429 10557 18463 10591
rect 19993 10557 20027 10591
rect 21465 10557 21499 10591
rect 23673 10557 23707 10591
rect 23929 10557 23963 10591
rect 2973 10489 3007 10523
rect 3332 10489 3366 10523
rect 5089 10489 5123 10523
rect 7205 10489 7239 10523
rect 14381 10489 14415 10523
rect 16773 10489 16807 10523
rect 19073 10489 19107 10523
rect 19901 10489 19935 10523
rect 4445 10421 4479 10455
rect 6837 10421 6871 10455
rect 12449 10421 12483 10455
rect 12909 10421 12943 10455
rect 16221 10421 16255 10455
rect 16865 10421 16899 10455
rect 18613 10421 18647 10455
rect 25605 10421 25639 10455
rect 25973 10421 26007 10455
rect 26341 10421 26375 10455
rect 1961 10217 1995 10251
rect 2421 10217 2455 10251
rect 4077 10217 4111 10251
rect 6101 10217 6135 10251
rect 7573 10217 7607 10251
rect 8217 10217 8251 10251
rect 8585 10217 8619 10251
rect 9689 10217 9723 10251
rect 10701 10217 10735 10251
rect 13829 10217 13863 10251
rect 14289 10217 14323 10251
rect 17693 10217 17727 10251
rect 19073 10217 19107 10251
rect 19257 10217 19291 10251
rect 19625 10217 19659 10251
rect 22845 10217 22879 10251
rect 23213 10217 23247 10251
rect 23857 10217 23891 10251
rect 24501 10217 24535 10251
rect 24777 10217 24811 10251
rect 25513 10217 25547 10251
rect 25881 10217 25915 10251
rect 26249 10217 26283 10251
rect 2881 10149 2915 10183
rect 3709 10149 3743 10183
rect 4445 10149 4479 10183
rect 6009 10149 6043 10183
rect 9229 10149 9263 10183
rect 10149 10149 10183 10183
rect 11774 10149 11808 10183
rect 15568 10149 15602 10183
rect 20269 10149 20303 10183
rect 20729 10149 20763 10183
rect 21180 10149 21214 10183
rect 2789 10081 2823 10115
rect 1409 10013 1443 10047
rect 3065 10013 3099 10047
rect 4537 10081 4571 10115
rect 8953 10081 8987 10115
rect 10057 10081 10091 10115
rect 11529 10081 11563 10115
rect 14105 10081 14139 10115
rect 18061 10081 18095 10115
rect 18153 10081 18187 10115
rect 23765 10081 23799 10115
rect 24961 10081 24995 10115
rect 4721 10013 4755 10047
rect 6285 10013 6319 10047
rect 6745 10013 6779 10047
rect 7665 10013 7699 10047
rect 7757 10013 7791 10047
rect 10241 10013 10275 10047
rect 15025 10013 15059 10047
rect 15301 10013 15335 10047
rect 18797 10013 18831 10047
rect 19717 10013 19751 10047
rect 19901 10013 19935 10047
rect 20913 10013 20947 10047
rect 23949 10013 23983 10047
rect 3709 9945 3743 9979
rect 3893 9945 3927 9979
rect 5641 9945 5675 9979
rect 7205 9945 7239 9979
rect 12909 9945 12943 9979
rect 23397 9945 23431 9979
rect 2237 9877 2271 9911
rect 3525 9877 3559 9911
rect 5181 9877 5215 9911
rect 7113 9877 7147 9911
rect 8769 9877 8803 9911
rect 11069 9877 11103 9911
rect 13461 9877 13495 9911
rect 14657 9877 14691 9911
rect 16681 9877 16715 9911
rect 17233 9877 17267 9911
rect 17877 9877 17911 9911
rect 18337 9877 18371 9911
rect 22293 9877 22327 9911
rect 25145 9877 25179 9911
rect 4445 9673 4479 9707
rect 11529 9673 11563 9707
rect 12173 9673 12207 9707
rect 13461 9673 13495 9707
rect 13829 9673 13863 9707
rect 14013 9673 14047 9707
rect 19165 9673 19199 9707
rect 22109 9673 22143 9707
rect 25605 9673 25639 9707
rect 1961 9605 1995 9639
rect 5181 9605 5215 9639
rect 6285 9605 6319 9639
rect 12449 9605 12483 9639
rect 15577 9605 15611 9639
rect 17877 9605 17911 9639
rect 18981 9605 19015 9639
rect 20269 9605 20303 9639
rect 20637 9605 20671 9639
rect 23121 9605 23155 9639
rect 25053 9605 25087 9639
rect 26433 9605 26467 9639
rect 1685 9537 1719 9571
rect 5733 9537 5767 9571
rect 8125 9537 8159 9571
rect 13093 9537 13127 9571
rect 14473 9537 14507 9571
rect 14565 9537 14599 9571
rect 15393 9537 15427 9571
rect 16129 9537 16163 9571
rect 16589 9537 16623 9571
rect 19625 9537 19659 9571
rect 19809 9537 19843 9571
rect 2145 9469 2179 9503
rect 5641 9469 5675 9503
rect 7389 9469 7423 9503
rect 7849 9469 7883 9503
rect 8953 9469 8987 9503
rect 9045 9469 9079 9503
rect 9312 9469 9346 9503
rect 12817 9469 12851 9503
rect 16037 9469 16071 9503
rect 16957 9469 16991 9503
rect 17333 9469 17367 9503
rect 18061 9469 18095 9503
rect 18613 9469 18647 9503
rect 19533 9469 19567 9503
rect 20729 9469 20763 9503
rect 22753 9469 22787 9503
rect 23673 9469 23707 9503
rect 23940 9469 23974 9503
rect 2390 9401 2424 9435
rect 6653 9401 6687 9435
rect 20974 9401 21008 9435
rect 23489 9401 23523 9435
rect 3525 9333 3559 9367
rect 4169 9333 4203 9367
rect 5089 9333 5123 9367
rect 5549 9333 5583 9367
rect 7481 9333 7515 9367
rect 7941 9333 7975 9367
rect 8493 9333 8527 9367
rect 10425 9333 10459 9367
rect 11069 9333 11103 9367
rect 12909 9333 12943 9367
rect 14381 9333 14415 9367
rect 15945 9333 15979 9367
rect 17141 9333 17175 9367
rect 18245 9333 18279 9367
rect 25973 9333 26007 9367
rect 1409 9129 1443 9163
rect 2237 9129 2271 9163
rect 2881 9129 2915 9163
rect 4077 9129 4111 9163
rect 5273 9129 5307 9163
rect 9137 9129 9171 9163
rect 10057 9129 10091 9163
rect 10885 9129 10919 9163
rect 14657 9129 14691 9163
rect 19993 9129 20027 9163
rect 20269 9129 20303 9163
rect 21373 9129 21407 9163
rect 22937 9129 22971 9163
rect 23489 9129 23523 9163
rect 24501 9129 24535 9163
rect 25421 9129 25455 9163
rect 25789 9129 25823 9163
rect 26249 9129 26283 9163
rect 4445 9061 4479 9095
rect 6368 9061 6402 9095
rect 9505 9061 9539 9095
rect 11161 9061 11195 9095
rect 17325 9061 17359 9095
rect 18236 9061 18270 9095
rect 22293 9061 22327 9095
rect 23857 9061 23891 9095
rect 2789 8993 2823 9027
rect 3893 8993 3927 9027
rect 6009 8993 6043 9027
rect 8125 8993 8159 9027
rect 11785 8993 11819 9027
rect 14105 8993 14139 9027
rect 15568 8993 15602 9027
rect 17969 8993 18003 9027
rect 20637 8993 20671 9027
rect 21281 8993 21315 9027
rect 22845 8993 22879 9027
rect 24409 8993 24443 9027
rect 2973 8925 3007 8959
rect 4537 8925 4571 8959
rect 4629 8925 4663 8959
rect 6101 8925 6135 8959
rect 8585 8925 8619 8959
rect 10149 8925 10183 8959
rect 10241 8925 10275 8959
rect 11529 8925 11563 8959
rect 13461 8925 13495 8959
rect 15025 8925 15059 8959
rect 15301 8925 15335 8959
rect 17877 8925 17911 8959
rect 21465 8925 21499 8959
rect 21925 8925 21959 8959
rect 23029 8925 23063 8959
rect 24593 8925 24627 8959
rect 2421 8857 2455 8891
rect 5641 8857 5675 8891
rect 9689 8857 9723 8891
rect 13921 8857 13955 8891
rect 20453 8857 20487 8891
rect 3433 8789 3467 8823
rect 5825 8789 5859 8823
rect 7481 8789 7515 8823
rect 8401 8789 8435 8823
rect 12909 8789 12943 8823
rect 14289 8789 14323 8823
rect 16681 8789 16715 8823
rect 19349 8789 19383 8823
rect 20913 8789 20947 8823
rect 22477 8789 22511 8823
rect 24041 8789 24075 8823
rect 25053 8789 25087 8823
rect 2697 8585 2731 8619
rect 5641 8585 5675 8619
rect 6285 8585 6319 8619
rect 9321 8585 9355 8619
rect 11805 8585 11839 8619
rect 12449 8585 12483 8619
rect 13921 8585 13955 8619
rect 15393 8585 15427 8619
rect 17877 8585 17911 8619
rect 19993 8585 20027 8619
rect 20453 8585 20487 8619
rect 21557 8585 21591 8619
rect 22385 8585 22419 8619
rect 23673 8585 23707 8619
rect 24777 8585 24811 8619
rect 25053 8585 25087 8619
rect 26157 8585 26191 8619
rect 2237 8517 2271 8551
rect 7021 8517 7055 8551
rect 12265 8517 12299 8551
rect 20545 8517 20579 8551
rect 1685 8449 1719 8483
rect 3249 8449 3283 8483
rect 8493 8449 8527 8483
rect 10333 8449 10367 8483
rect 11345 8449 11379 8483
rect 12909 8449 12943 8483
rect 13093 8449 13127 8483
rect 16037 8449 16071 8483
rect 18061 8449 18095 8483
rect 21189 8449 21223 8483
rect 24133 8449 24167 8483
rect 24225 8449 24259 8483
rect 1409 8381 1443 8415
rect 3065 8381 3099 8415
rect 4261 8381 4295 8415
rect 6837 8381 6871 8415
rect 7389 8381 7423 8415
rect 7849 8381 7883 8415
rect 8401 8381 8435 8415
rect 9045 8381 9079 8415
rect 9505 8381 9539 8415
rect 11253 8381 11287 8415
rect 14013 8381 14047 8415
rect 14280 8381 14314 8415
rect 16405 8381 16439 8415
rect 16528 8381 16562 8415
rect 21925 8381 21959 8415
rect 22477 8381 22511 8415
rect 25237 8381 25271 8415
rect 25789 8381 25823 8415
rect 4169 8313 4203 8347
rect 4506 8313 4540 8347
rect 6653 8313 6687 8347
rect 8309 8313 8343 8347
rect 9781 8313 9815 8347
rect 10609 8313 10643 8347
rect 11161 8313 11195 8347
rect 12817 8313 12851 8347
rect 13553 8313 13587 8347
rect 16773 8313 16807 8347
rect 17509 8313 17543 8347
rect 18306 8313 18340 8347
rect 20913 8313 20947 8347
rect 23029 8313 23063 8347
rect 2605 8245 2639 8279
rect 3157 8245 3191 8279
rect 3709 8245 3743 8279
rect 7941 8245 7975 8279
rect 10793 8245 10827 8279
rect 19441 8245 19475 8279
rect 21005 8245 21039 8279
rect 22661 8245 22695 8279
rect 23397 8245 23431 8279
rect 24041 8245 24075 8279
rect 25421 8245 25455 8279
rect 2789 8041 2823 8075
rect 3801 8041 3835 8075
rect 4353 8041 4387 8075
rect 5089 8041 5123 8075
rect 5825 8041 5859 8075
rect 8401 8041 8435 8075
rect 9413 8041 9447 8075
rect 10517 8041 10551 8075
rect 11345 8041 11379 8075
rect 11713 8041 11747 8075
rect 11897 8041 11931 8075
rect 13277 8041 13311 8075
rect 13461 8041 13495 8075
rect 15301 8041 15335 8075
rect 17693 8041 17727 8075
rect 18797 8041 18831 8075
rect 20269 8041 20303 8075
rect 22937 8041 22971 8075
rect 23305 8041 23339 8075
rect 24041 8041 24075 8075
rect 24501 8041 24535 8075
rect 25973 8041 26007 8075
rect 26341 8041 26375 8075
rect 13001 7973 13035 8007
rect 14933 7973 14967 8007
rect 15853 7973 15887 8007
rect 16221 7973 16255 8007
rect 18337 7973 18371 8007
rect 21180 7973 21214 8007
rect 1676 7905 1710 7939
rect 5181 7905 5215 7939
rect 6745 7905 6779 7939
rect 8309 7905 8343 7939
rect 12265 7905 12299 7939
rect 13829 7905 13863 7939
rect 13921 7905 13955 7939
rect 16569 7905 16603 7939
rect 19165 7905 19199 7939
rect 19809 7905 19843 7939
rect 23397 7905 23431 7939
rect 24869 7905 24903 7939
rect 1409 7837 1443 7871
rect 5365 7837 5399 7871
rect 6837 7837 6871 7871
rect 7021 7837 7055 7871
rect 8493 7837 8527 7871
rect 10609 7837 10643 7871
rect 10793 7837 10827 7871
rect 12357 7837 12391 7871
rect 12449 7837 12483 7871
rect 14105 7837 14139 7871
rect 16313 7837 16347 7871
rect 19257 7837 19291 7871
rect 19349 7837 19383 7871
rect 20913 7837 20947 7871
rect 24961 7837 24995 7871
rect 25053 7837 25087 7871
rect 7665 7769 7699 7803
rect 3341 7701 3375 7735
rect 4721 7701 4755 7735
rect 6101 7701 6135 7735
rect 6377 7701 6411 7735
rect 7941 7701 7975 7735
rect 8953 7701 8987 7735
rect 9965 7701 9999 7735
rect 10149 7701 10183 7735
rect 14473 7701 14507 7735
rect 18613 7701 18647 7735
rect 20545 7701 20579 7735
rect 22293 7701 22327 7735
rect 23581 7701 23615 7735
rect 25513 7701 25547 7735
rect 1501 7497 1535 7531
rect 2513 7497 2547 7531
rect 3985 7497 4019 7531
rect 5457 7497 5491 7531
rect 8585 7497 8619 7531
rect 9781 7497 9815 7531
rect 11253 7497 11287 7531
rect 11897 7497 11931 7531
rect 13553 7497 13587 7531
rect 15025 7497 15059 7531
rect 15577 7497 15611 7531
rect 15853 7497 15887 7531
rect 17509 7497 17543 7531
rect 19349 7497 19383 7531
rect 20085 7497 20119 7531
rect 23397 7497 23431 7531
rect 23949 7497 23983 7531
rect 26433 7497 26467 7531
rect 7573 7429 7607 7463
rect 12173 7429 12207 7463
rect 18245 7429 18279 7463
rect 21649 7429 21683 7463
rect 24961 7429 24995 7463
rect 2145 7361 2179 7395
rect 4445 7361 4479 7395
rect 4537 7361 4571 7395
rect 8033 7361 8067 7395
rect 8125 7361 8159 7395
rect 13093 7361 13127 7395
rect 14473 7361 14507 7395
rect 14565 7361 14599 7395
rect 17049 7361 17083 7395
rect 17877 7361 17911 7395
rect 18889 7361 18923 7395
rect 20729 7361 20763 7395
rect 22201 7361 22235 7395
rect 22293 7361 22327 7395
rect 24593 7361 24627 7395
rect 26065 7361 26099 7395
rect 3525 7293 3559 7327
rect 5641 7293 5675 7327
rect 7941 7293 7975 7327
rect 9321 7293 9355 7327
rect 9873 7293 9907 7327
rect 10129 7293 10163 7327
rect 12817 7293 12851 7327
rect 16773 7293 16807 7327
rect 19901 7293 19935 7327
rect 20637 7293 20671 7327
rect 21281 7293 21315 7327
rect 24317 7293 24351 7327
rect 25513 7293 25547 7327
rect 1961 7225 1995 7259
rect 3893 7225 3927 7259
rect 7113 7225 7147 7259
rect 9045 7225 9079 7259
rect 13921 7225 13955 7259
rect 16221 7225 16255 7259
rect 16865 7225 16899 7259
rect 18613 7225 18647 7259
rect 25329 7225 25363 7259
rect 1869 7157 1903 7191
rect 2973 7157 3007 7191
rect 4353 7157 4387 7191
rect 4997 7157 5031 7191
rect 5825 7157 5859 7191
rect 6469 7157 6503 7191
rect 7389 7157 7423 7191
rect 9137 7157 9171 7191
rect 12449 7157 12483 7191
rect 12909 7157 12943 7191
rect 14013 7157 14047 7191
rect 14381 7157 14415 7191
rect 16405 7157 16439 7191
rect 18705 7157 18739 7191
rect 19625 7157 19659 7191
rect 19901 7157 19935 7191
rect 20177 7157 20211 7191
rect 20545 7157 20579 7191
rect 21741 7157 21775 7191
rect 22109 7157 22143 7191
rect 23121 7157 23155 7191
rect 24409 7157 24443 7191
rect 25697 7157 25731 7191
rect 4353 6953 4387 6987
rect 7205 6953 7239 6987
rect 7665 6953 7699 6987
rect 10057 6953 10091 6987
rect 12173 6953 12207 6987
rect 12449 6953 12483 6987
rect 13093 6953 13127 6987
rect 13645 6953 13679 6987
rect 16589 6953 16623 6987
rect 17877 6953 17911 6987
rect 18981 6953 19015 6987
rect 20269 6953 20303 6987
rect 21925 6953 21959 6987
rect 25697 6953 25731 6987
rect 13001 6885 13035 6919
rect 14013 6885 14047 6919
rect 17417 6885 17451 6919
rect 18245 6885 18279 6919
rect 23572 6885 23606 6919
rect 1501 6817 1535 6851
rect 1768 6817 1802 6851
rect 5069 6817 5103 6851
rect 6745 6817 6779 6851
rect 7757 6817 7791 6851
rect 8677 6817 8711 6851
rect 10405 6817 10439 6851
rect 16129 6817 16163 6851
rect 17693 6817 17727 6851
rect 19441 6817 19475 6851
rect 21281 6817 21315 6851
rect 23029 6817 23063 6851
rect 4813 6749 4847 6783
rect 7849 6749 7883 6783
rect 10149 6749 10183 6783
rect 13185 6749 13219 6783
rect 14197 6749 14231 6783
rect 15485 6749 15519 6783
rect 16681 6749 16715 6783
rect 16773 6749 16807 6783
rect 18337 6749 18371 6783
rect 18521 6749 18555 6783
rect 19625 6749 19659 6783
rect 21373 6749 21407 6783
rect 21557 6749 21591 6783
rect 23305 6749 23339 6783
rect 7297 6681 7331 6715
rect 9045 6681 9079 6715
rect 16221 6681 16255 6715
rect 19349 6681 19383 6715
rect 20913 6681 20947 6715
rect 22661 6681 22695 6715
rect 24685 6681 24719 6715
rect 25329 6681 25363 6715
rect 2881 6613 2915 6647
rect 3433 6613 3467 6647
rect 3893 6613 3927 6647
rect 4629 6613 4663 6647
rect 6193 6613 6227 6647
rect 8401 6613 8435 6647
rect 9413 6613 9447 6647
rect 11529 6613 11563 6647
rect 12633 6613 12667 6647
rect 14657 6613 14691 6647
rect 15025 6613 15059 6647
rect 20637 6613 20671 6647
rect 22293 6613 22327 6647
rect 25973 6613 26007 6647
rect 3801 6409 3835 6443
rect 4905 6409 4939 6443
rect 9781 6409 9815 6443
rect 14749 6409 14783 6443
rect 17417 6409 17451 6443
rect 17785 6409 17819 6443
rect 19441 6409 19475 6443
rect 20361 6409 20395 6443
rect 21833 6409 21867 6443
rect 23121 6409 23155 6443
rect 23397 6409 23431 6443
rect 25053 6409 25087 6443
rect 26065 6409 26099 6443
rect 26341 6409 26375 6443
rect 4813 6273 4847 6307
rect 5457 6273 5491 6307
rect 15209 6273 15243 6307
rect 18521 6273 18555 6307
rect 18705 6273 18739 6307
rect 19809 6273 19843 6307
rect 2421 6205 2455 6239
rect 4445 6205 4479 6239
rect 5273 6205 5307 6239
rect 7389 6205 7423 6239
rect 9873 6205 9907 6239
rect 12449 6205 12483 6239
rect 12716 6205 12750 6239
rect 15301 6205 15335 6239
rect 15568 6205 15602 6239
rect 19073 6205 19107 6239
rect 20453 6205 20487 6239
rect 23673 6205 23707 6239
rect 2329 6137 2363 6171
rect 2666 6137 2700 6171
rect 6285 6137 6319 6171
rect 7634 6137 7668 6171
rect 9413 6137 9447 6171
rect 10118 6137 10152 6171
rect 20698 6137 20732 6171
rect 23918 6137 23952 6171
rect 25605 6137 25639 6171
rect 1409 6069 1443 6103
rect 1869 6069 1903 6103
rect 5365 6069 5399 6103
rect 6653 6069 6687 6103
rect 7297 6069 7331 6103
rect 8769 6069 8803 6103
rect 11253 6069 11287 6103
rect 11897 6069 11931 6103
rect 12173 6069 12207 6103
rect 13829 6069 13863 6103
rect 14381 6069 14415 6103
rect 16681 6069 16715 6103
rect 18061 6069 18095 6103
rect 18429 6069 18463 6103
rect 22385 6069 22419 6103
rect 1409 5865 1443 5899
rect 3433 5865 3467 5899
rect 4261 5865 4295 5899
rect 4721 5865 4755 5899
rect 5273 5865 5307 5899
rect 7205 5865 7239 5899
rect 7849 5865 7883 5899
rect 9689 5865 9723 5899
rect 11529 5865 11563 5899
rect 11897 5865 11931 5899
rect 14105 5865 14139 5899
rect 15669 5865 15703 5899
rect 15761 5865 15795 5899
rect 16681 5865 16715 5899
rect 16865 5865 16899 5899
rect 17693 5865 17727 5899
rect 18245 5865 18279 5899
rect 21189 5865 21223 5899
rect 22937 5865 22971 5899
rect 23673 5865 23707 5899
rect 24041 5865 24075 5899
rect 25053 5865 25087 5899
rect 25421 5865 25455 5899
rect 25881 5865 25915 5899
rect 26157 5865 26191 5899
rect 2881 5797 2915 5831
rect 6193 5797 6227 5831
rect 21824 5797 21858 5831
rect 1777 5729 1811 5763
rect 1869 5729 1903 5763
rect 4629 5729 4663 5763
rect 6285 5729 6319 5763
rect 7757 5729 7791 5763
rect 10057 5729 10091 5763
rect 12245 5729 12279 5763
rect 18337 5729 18371 5763
rect 19441 5729 19475 5763
rect 21557 5729 21591 5763
rect 24409 5729 24443 5763
rect 24501 5729 24535 5763
rect 2053 5661 2087 5695
rect 2973 5661 3007 5695
rect 4905 5661 4939 5695
rect 5733 5661 5767 5695
rect 6469 5661 6503 5695
rect 8033 5661 8067 5695
rect 8861 5661 8895 5695
rect 10149 5661 10183 5695
rect 10241 5661 10275 5695
rect 11989 5661 12023 5695
rect 15853 5661 15887 5695
rect 17417 5661 17451 5695
rect 18429 5661 18463 5695
rect 19625 5661 19659 5695
rect 24593 5661 24627 5695
rect 3893 5593 3927 5627
rect 5825 5593 5859 5627
rect 7389 5593 7423 5627
rect 15301 5593 15335 5627
rect 17877 5593 17911 5627
rect 19349 5593 19383 5627
rect 2513 5525 2547 5559
rect 6929 5525 6963 5559
rect 8493 5525 8527 5559
rect 9229 5525 9263 5559
rect 10701 5525 10735 5559
rect 11161 5525 11195 5559
rect 13369 5525 13403 5559
rect 14473 5525 14507 5559
rect 15117 5525 15151 5559
rect 16405 5525 16439 5559
rect 18981 5525 19015 5559
rect 20453 5525 20487 5559
rect 2973 5321 3007 5355
rect 4353 5321 4387 5355
rect 4721 5321 4755 5355
rect 5181 5321 5215 5355
rect 7573 5321 7607 5355
rect 10149 5321 10183 5355
rect 11897 5321 11931 5355
rect 13461 5321 13495 5355
rect 13829 5321 13863 5355
rect 14013 5321 14047 5355
rect 15393 5321 15427 5355
rect 16589 5321 16623 5355
rect 18245 5321 18279 5355
rect 18613 5321 18647 5355
rect 21281 5321 21315 5355
rect 22293 5321 22327 5355
rect 23121 5321 23155 5355
rect 23673 5321 23707 5355
rect 24685 5321 24719 5355
rect 26341 5321 26375 5355
rect 6285 5253 6319 5287
rect 7113 5253 7147 5287
rect 10701 5253 10735 5287
rect 13277 5253 13311 5287
rect 15577 5253 15611 5287
rect 16957 5253 16991 5287
rect 17325 5253 17359 5287
rect 23489 5253 23523 5287
rect 2053 5185 2087 5219
rect 3617 5185 3651 5219
rect 5089 5185 5123 5219
rect 5641 5185 5675 5219
rect 5733 5185 5767 5219
rect 7481 5185 7515 5219
rect 8217 5185 8251 5219
rect 9689 5185 9723 5219
rect 11253 5185 11287 5219
rect 12173 5185 12207 5219
rect 13001 5185 13035 5219
rect 1777 5117 1811 5151
rect 2881 5117 2915 5151
rect 3433 5117 3467 5151
rect 5549 5117 5583 5151
rect 7941 5117 7975 5151
rect 9597 5117 9631 5151
rect 3341 5049 3375 5083
rect 6653 5049 6687 5083
rect 9505 5049 9539 5083
rect 10609 5049 10643 5083
rect 11161 5049 11195 5083
rect 14473 5185 14507 5219
rect 14565 5185 14599 5219
rect 16037 5185 16071 5219
rect 16129 5185 16163 5219
rect 21833 5185 21867 5219
rect 24225 5185 24259 5219
rect 25513 5185 25547 5219
rect 14381 5117 14415 5151
rect 15945 5117 15979 5151
rect 18797 5117 18831 5151
rect 21649 5117 21683 5151
rect 24133 5117 24167 5151
rect 25237 5117 25271 5151
rect 25973 5117 26007 5151
rect 17877 5049 17911 5083
rect 19064 5049 19098 5083
rect 21097 5049 21131 5083
rect 22661 5049 22695 5083
rect 24041 5049 24075 5083
rect 1409 4981 1443 5015
rect 1869 4981 1903 5015
rect 2421 4981 2455 5015
rect 8033 4981 8067 5015
rect 8677 4981 8711 5015
rect 8953 4981 8987 5015
rect 9137 4981 9171 5015
rect 11069 4981 11103 5015
rect 12449 4981 12483 5015
rect 12817 4981 12851 5015
rect 12909 4981 12943 5015
rect 13277 4981 13311 5015
rect 20177 4981 20211 5015
rect 20729 4981 20763 5015
rect 21741 4981 21775 5015
rect 25053 4981 25087 5015
rect 1501 4777 1535 4811
rect 1961 4777 1995 4811
rect 2513 4777 2547 4811
rect 4077 4777 4111 4811
rect 4445 4777 4479 4811
rect 5549 4777 5583 4811
rect 5733 4777 5767 4811
rect 7297 4777 7331 4811
rect 7757 4777 7791 4811
rect 9229 4777 9263 4811
rect 9689 4777 9723 4811
rect 10149 4777 10183 4811
rect 12357 4777 12391 4811
rect 13277 4777 13311 4811
rect 13461 4777 13495 4811
rect 13921 4777 13955 4811
rect 15117 4777 15151 4811
rect 19441 4777 19475 4811
rect 20637 4777 20671 4811
rect 20913 4777 20947 4811
rect 23765 4777 23799 4811
rect 24501 4777 24535 4811
rect 26249 4777 26283 4811
rect 1869 4709 1903 4743
rect 3065 4709 3099 4743
rect 5273 4709 5307 4743
rect 6193 4709 6227 4743
rect 6837 4709 6871 4743
rect 8401 4709 8435 4743
rect 10057 4709 10091 4743
rect 12909 4709 12943 4743
rect 22845 4709 22879 4743
rect 25421 4709 25455 4743
rect 3433 4641 3467 4675
rect 3893 4641 3927 4675
rect 6101 4641 6135 4675
rect 7665 4641 7699 4675
rect 11345 4641 11379 4675
rect 12265 4641 12299 4675
rect 13829 4641 13863 4675
rect 15568 4641 15602 4675
rect 18061 4641 18095 4675
rect 18328 4641 18362 4675
rect 21281 4641 21315 4675
rect 24409 4641 24443 4675
rect 25789 4641 25823 4675
rect 2145 4573 2179 4607
rect 4537 4573 4571 4607
rect 4721 4573 4755 4607
rect 6285 4573 6319 4607
rect 7205 4573 7239 4607
rect 7941 4573 7975 4607
rect 8861 4573 8895 4607
rect 10241 4573 10275 4607
rect 12449 4573 12483 4607
rect 14013 4573 14047 4607
rect 15301 4573 15335 4607
rect 17601 4573 17635 4607
rect 21373 4573 21407 4607
rect 21465 4573 21499 4607
rect 22937 4573 22971 4607
rect 23121 4573 23155 4607
rect 24593 4573 24627 4607
rect 10793 4505 10827 4539
rect 11805 4505 11839 4539
rect 21925 4505 21959 4539
rect 24041 4505 24075 4539
rect 11897 4437 11931 4471
rect 14565 4437 14599 4471
rect 16681 4437 16715 4471
rect 17969 4437 18003 4471
rect 19993 4437 20027 4471
rect 22385 4437 22419 4471
rect 22477 4437 22511 4471
rect 25053 4437 25087 4471
rect 2513 4233 2547 4267
rect 5917 4233 5951 4267
rect 9689 4233 9723 4267
rect 11897 4233 11931 4267
rect 13921 4233 13955 4267
rect 15577 4233 15611 4267
rect 18429 4233 18463 4267
rect 19441 4233 19475 4267
rect 21097 4233 21131 4267
rect 22661 4233 22695 4267
rect 26157 4233 26191 4267
rect 10793 4165 10827 4199
rect 17877 4165 17911 4199
rect 19901 4165 19935 4199
rect 2053 4097 2087 4131
rect 3985 4097 4019 4131
rect 7021 4097 7055 4131
rect 10241 4097 10275 4131
rect 11161 4097 11195 4131
rect 13001 4097 13035 4131
rect 14565 4097 14599 4131
rect 15117 4097 15151 4131
rect 16221 4097 16255 4131
rect 18153 4097 18187 4131
rect 18245 4097 18279 4131
rect 18889 4097 18923 4131
rect 19073 4097 19107 4131
rect 20453 4097 20487 4131
rect 20545 4097 20579 4131
rect 22201 4097 22235 4131
rect 22937 4097 22971 4131
rect 24133 4097 24167 4131
rect 24317 4097 24351 4131
rect 25053 4097 25087 4131
rect 3893 4029 3927 4063
rect 7205 4029 7239 4063
rect 7461 4029 7495 4063
rect 10057 4029 10091 4063
rect 11253 4029 11287 4063
rect 12909 4029 12943 4063
rect 14381 4029 14415 4063
rect 15485 4029 15519 4063
rect 16037 4029 16071 4063
rect 16681 4029 16715 4063
rect 1869 3961 1903 3995
rect 2881 3961 2915 3995
rect 3525 3961 3559 3995
rect 4230 3961 4264 3995
rect 9505 3961 9539 3995
rect 10149 3961 10183 3995
rect 12265 3961 12299 3995
rect 12817 3961 12851 3995
rect 15945 3961 15979 3995
rect 17509 3961 17543 3995
rect 25237 4029 25271 4063
rect 25789 4029 25823 4063
rect 21925 3961 21959 3995
rect 22017 3961 22051 3995
rect 23489 3961 23523 3995
rect 24777 3961 24811 3995
rect 1409 3893 1443 3927
rect 1777 3893 1811 3927
rect 2973 3893 3007 3927
rect 5365 3893 5399 3927
rect 6377 3893 6411 3927
rect 8585 3893 8619 3927
rect 9137 3893 9171 3927
rect 11437 3893 11471 3927
rect 12449 3893 12483 3927
rect 13461 3893 13495 3927
rect 14013 3893 14047 3927
rect 14473 3893 14507 3927
rect 16957 3893 16991 3927
rect 18153 3893 18187 3927
rect 18797 3893 18831 3927
rect 19993 3893 20027 3927
rect 20361 3893 20395 3927
rect 21373 3893 21407 3927
rect 21557 3893 21591 3927
rect 23673 3893 23707 3927
rect 24041 3893 24075 3927
rect 25421 3893 25455 3927
rect 1409 3689 1443 3723
rect 1777 3689 1811 3723
rect 1869 3689 1903 3723
rect 2421 3689 2455 3723
rect 6101 3689 6135 3723
rect 6469 3689 6503 3723
rect 7665 3689 7699 3723
rect 7849 3689 7883 3723
rect 8217 3689 8251 3723
rect 9689 3689 9723 3723
rect 10057 3689 10091 3723
rect 11253 3689 11287 3723
rect 12541 3689 12575 3723
rect 12817 3689 12851 3723
rect 13277 3689 13311 3723
rect 15301 3689 15335 3723
rect 15761 3689 15795 3723
rect 16865 3689 16899 3723
rect 17325 3689 17359 3723
rect 18889 3689 18923 3723
rect 19901 3689 19935 3723
rect 21373 3689 21407 3723
rect 22385 3689 22419 3723
rect 22845 3689 22879 3723
rect 22937 3689 22971 3723
rect 24041 3689 24075 3723
rect 24409 3689 24443 3723
rect 24501 3689 24535 3723
rect 25421 3689 25455 3723
rect 26249 3689 26283 3723
rect 2789 3621 2823 3655
rect 3433 3621 3467 3655
rect 3893 3621 3927 3655
rect 4344 3621 4378 3655
rect 6837 3621 6871 3655
rect 11621 3621 11655 3655
rect 16313 3621 16347 3655
rect 16773 3621 16807 3655
rect 17233 3621 17267 3655
rect 18797 3621 18831 3655
rect 21281 3621 21315 3655
rect 21925 3621 21959 3655
rect 4077 3553 4111 3587
rect 6561 3553 6595 3587
rect 10701 3553 10735 3587
rect 11069 3553 11103 3587
rect 13185 3553 13219 3587
rect 15117 3553 15151 3587
rect 15669 3553 15703 3587
rect 23765 3553 23799 3587
rect 25789 3553 25823 3587
rect 2053 3485 2087 3519
rect 2973 3485 3007 3519
rect 8309 3485 8343 3519
rect 8401 3485 8435 3519
rect 9045 3485 9079 3519
rect 10149 3485 10183 3519
rect 10241 3485 10275 3519
rect 11713 3485 11747 3519
rect 11805 3485 11839 3519
rect 13369 3485 13403 3519
rect 14013 3485 14047 3519
rect 14381 3485 14415 3519
rect 15853 3485 15887 3519
rect 17417 3485 17451 3519
rect 18981 3485 19015 3519
rect 21465 3485 21499 3519
rect 23121 3485 23155 3519
rect 24593 3485 24627 3519
rect 18429 3417 18463 3451
rect 19625 3417 19659 3451
rect 20913 3417 20947 3451
rect 25053 3417 25087 3451
rect 5457 3349 5491 3383
rect 7389 3349 7423 3383
rect 9505 3349 9539 3383
rect 18061 3349 18095 3383
rect 20269 3349 20303 3383
rect 20729 3349 20763 3383
rect 22477 3349 22511 3383
rect 1409 3145 1443 3179
rect 3617 3145 3651 3179
rect 5181 3145 5215 3179
rect 6561 3145 6595 3179
rect 7113 3145 7147 3179
rect 8585 3145 8619 3179
rect 9597 3145 9631 3179
rect 11069 3145 11103 3179
rect 11989 3145 12023 3179
rect 17049 3145 17083 3179
rect 18061 3145 18095 3179
rect 19073 3145 19107 3179
rect 19625 3145 19659 3179
rect 20729 3145 20763 3179
rect 21189 3145 21223 3179
rect 22569 3145 22603 3179
rect 22937 3145 22971 3179
rect 23489 3145 23523 3179
rect 24777 3145 24811 3179
rect 25053 3145 25087 3179
rect 26065 3145 26099 3179
rect 26341 3145 26375 3179
rect 2789 3077 2823 3111
rect 9229 3077 9263 3111
rect 11713 3077 11747 3111
rect 13829 3077 13863 3111
rect 23673 3077 23707 3111
rect 2053 3009 2087 3043
rect 3525 3009 3559 3043
rect 4169 3009 4203 3043
rect 5825 3009 5859 3043
rect 7205 3009 7239 3043
rect 17417 3009 17451 3043
rect 18613 3009 18647 3043
rect 19441 3009 19475 3043
rect 20085 3009 20119 3043
rect 20177 3009 20211 3043
rect 21833 3009 21867 3043
rect 24317 3009 24351 3043
rect 2237 2941 2271 2975
rect 4721 2941 4755 2975
rect 5641 2941 5675 2975
rect 6285 2941 6319 2975
rect 9689 2941 9723 2975
rect 12449 2941 12483 2975
rect 15117 2941 15151 2975
rect 17785 2941 17819 2975
rect 18429 2941 18463 2975
rect 18521 2941 18555 2975
rect 21557 2941 21591 2975
rect 24133 2941 24167 2975
rect 25237 2941 25271 2975
rect 1777 2873 1811 2907
rect 2513 2873 2547 2907
rect 3985 2873 4019 2907
rect 5089 2873 5123 2907
rect 5549 2873 5583 2907
rect 7472 2873 7506 2907
rect 9934 2873 9968 2907
rect 12716 2873 12750 2907
rect 14657 2873 14691 2907
rect 15362 2873 15396 2907
rect 19993 2873 20027 2907
rect 21097 2873 21131 2907
rect 21649 2873 21683 2907
rect 24041 2873 24075 2907
rect 25513 2873 25547 2907
rect 1869 2805 1903 2839
rect 2237 2805 2271 2839
rect 4077 2805 4111 2839
rect 14933 2805 14967 2839
rect 16497 2805 16531 2839
rect 1961 2601 1995 2635
rect 2789 2601 2823 2635
rect 3525 2601 3559 2635
rect 6285 2601 6319 2635
rect 8585 2601 8619 2635
rect 9597 2601 9631 2635
rect 11437 2601 11471 2635
rect 14841 2601 14875 2635
rect 15485 2601 15519 2635
rect 15945 2601 15979 2635
rect 18337 2601 18371 2635
rect 18797 2601 18831 2635
rect 21189 2601 21223 2635
rect 23029 2601 23063 2635
rect 24041 2601 24075 2635
rect 25053 2601 25087 2635
rect 26433 2601 26467 2635
rect 1685 2533 1719 2567
rect 6745 2533 6779 2567
rect 7472 2533 7506 2567
rect 9229 2533 9263 2567
rect 10324 2533 10358 2567
rect 12449 2533 12483 2567
rect 13154 2533 13188 2567
rect 18153 2533 18187 2567
rect 21649 2533 21683 2567
rect 23857 2533 23891 2567
rect 24501 2533 24535 2567
rect 25421 2533 25455 2567
rect 25605 2533 25639 2567
rect 4353 2465 4387 2499
rect 4620 2465 4654 2499
rect 7205 2465 7239 2499
rect 10057 2465 10091 2499
rect 12909 2465 12943 2499
rect 15853 2465 15887 2499
rect 17049 2465 17083 2499
rect 18705 2465 18739 2499
rect 19993 2465 20027 2499
rect 21557 2465 21591 2499
rect 22845 2465 22879 2499
rect 23397 2465 23431 2499
rect 24409 2465 24443 2499
rect 26065 2465 26099 2499
rect 2881 2397 2915 2431
rect 3065 2397 3099 2431
rect 3893 2397 3927 2431
rect 12081 2397 12115 2431
rect 16129 2397 16163 2431
rect 18889 2397 18923 2431
rect 19349 2397 19383 2431
rect 20545 2397 20579 2431
rect 21741 2397 21775 2431
rect 22201 2397 22235 2431
rect 22569 2397 22603 2431
rect 24685 2397 24719 2431
rect 2421 2329 2455 2363
rect 14289 2329 14323 2363
rect 15301 2329 15335 2363
rect 5733 2261 5767 2295
rect 16589 2261 16623 2295
rect 16957 2261 16991 2295
rect 17233 2261 17267 2295
rect 17693 2261 17727 2295
rect 19809 2261 19843 2295
rect 20177 2261 20211 2295
rect 20913 2261 20947 2295
<< metal1 >>
rect 2866 27412 2872 27464
rect 2924 27452 2930 27464
rect 3786 27452 3792 27464
rect 2924 27424 3792 27452
rect 2924 27412 2930 27424
rect 3786 27412 3792 27424
rect 3844 27412 3850 27464
rect 21082 26800 21088 26852
rect 21140 26840 21146 26852
rect 24670 26840 24676 26852
rect 21140 26812 24676 26840
rect 21140 26800 21146 26812
rect 24670 26800 24676 26812
rect 24728 26800 24734 26852
rect 20070 26392 20076 26444
rect 20128 26432 20134 26444
rect 24762 26432 24768 26444
rect 20128 26404 24768 26432
rect 20128 26392 20134 26404
rect 24762 26392 24768 26404
rect 24820 26392 24826 26444
rect 11882 26324 11888 26376
rect 11940 26364 11946 26376
rect 17954 26364 17960 26376
rect 11940 26336 17960 26364
rect 11940 26324 11946 26336
rect 17954 26324 17960 26336
rect 18012 26324 18018 26376
rect 8294 26188 8300 26240
rect 8352 26228 8358 26240
rect 18230 26228 18236 26240
rect 8352 26200 18236 26228
rect 8352 26188 8358 26200
rect 18230 26188 18236 26200
rect 18288 26188 18294 26240
rect 7742 26120 7748 26172
rect 7800 26160 7806 26172
rect 17126 26160 17132 26172
rect 7800 26132 17132 26160
rect 7800 26120 7806 26132
rect 17126 26120 17132 26132
rect 17184 26120 17190 26172
rect 8754 26052 8760 26104
rect 8812 26092 8818 26104
rect 18322 26092 18328 26104
rect 8812 26064 18328 26092
rect 8812 26052 8818 26064
rect 18322 26052 18328 26064
rect 18380 26052 18386 26104
rect 7834 25984 7840 26036
rect 7892 26024 7898 26036
rect 13078 26024 13084 26036
rect 7892 25996 13084 26024
rect 7892 25984 7898 25996
rect 13078 25984 13084 25996
rect 13136 25984 13142 26036
rect 13170 25984 13176 26036
rect 13228 26024 13234 26036
rect 24670 26024 24676 26036
rect 13228 25996 24676 26024
rect 13228 25984 13234 25996
rect 24670 25984 24676 25996
rect 24728 25984 24734 26036
rect 8938 25916 8944 25968
rect 8996 25956 9002 25968
rect 16574 25956 16580 25968
rect 8996 25928 16580 25956
rect 8996 25916 9002 25928
rect 16574 25916 16580 25928
rect 16632 25916 16638 25968
rect 17218 25916 17224 25968
rect 17276 25956 17282 25968
rect 22370 25956 22376 25968
rect 17276 25928 22376 25956
rect 17276 25916 17282 25928
rect 22370 25916 22376 25928
rect 22428 25916 22434 25968
rect 6362 25848 6368 25900
rect 6420 25888 6426 25900
rect 17770 25888 17776 25900
rect 6420 25860 17776 25888
rect 6420 25848 6426 25860
rect 17770 25848 17776 25860
rect 17828 25848 17834 25900
rect 8846 25780 8852 25832
rect 8904 25820 8910 25832
rect 19518 25820 19524 25832
rect 8904 25792 19524 25820
rect 8904 25780 8910 25792
rect 19518 25780 19524 25792
rect 19576 25780 19582 25832
rect 22462 25780 22468 25832
rect 22520 25820 22526 25832
rect 26510 25820 26516 25832
rect 22520 25792 26516 25820
rect 22520 25780 22526 25792
rect 26510 25780 26516 25792
rect 26568 25780 26574 25832
rect 7466 25712 7472 25764
rect 7524 25752 7530 25764
rect 18874 25752 18880 25764
rect 7524 25724 18880 25752
rect 7524 25712 7530 25724
rect 18874 25712 18880 25724
rect 18932 25712 18938 25764
rect 18966 25712 18972 25764
rect 19024 25752 19030 25764
rect 25866 25752 25872 25764
rect 19024 25724 25872 25752
rect 19024 25712 19030 25724
rect 25866 25712 25872 25724
rect 25924 25712 25930 25764
rect 9122 25644 9128 25696
rect 9180 25684 9186 25696
rect 21266 25684 21272 25696
rect 9180 25656 21272 25684
rect 9180 25644 9186 25656
rect 21266 25644 21272 25656
rect 21324 25644 21330 25696
rect 22186 25644 22192 25696
rect 22244 25684 22250 25696
rect 24762 25684 24768 25696
rect 22244 25656 24768 25684
rect 22244 25644 22250 25656
rect 24762 25644 24768 25656
rect 24820 25644 24826 25696
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 8757 25483 8815 25489
rect 8757 25449 8769 25483
rect 8803 25480 8815 25483
rect 8938 25480 8944 25492
rect 8803 25452 8944 25480
rect 8803 25449 8815 25452
rect 8757 25443 8815 25449
rect 8938 25440 8944 25452
rect 8996 25440 9002 25492
rect 10505 25483 10563 25489
rect 10505 25449 10517 25483
rect 10551 25480 10563 25483
rect 17218 25480 17224 25492
rect 10551 25452 17224 25480
rect 10551 25449 10563 25452
rect 10505 25443 10563 25449
rect 17218 25440 17224 25452
rect 17276 25440 17282 25492
rect 19978 25440 19984 25492
rect 20036 25440 20042 25492
rect 20165 25483 20223 25489
rect 20165 25449 20177 25483
rect 20211 25449 20223 25483
rect 20165 25443 20223 25449
rect 21453 25483 21511 25489
rect 21453 25449 21465 25483
rect 21499 25480 21511 25483
rect 24762 25480 24768 25492
rect 21499 25452 24768 25480
rect 21499 25449 21511 25452
rect 21453 25443 21511 25449
rect 11057 25415 11115 25421
rect 11057 25381 11069 25415
rect 11103 25412 11115 25415
rect 14369 25415 14427 25421
rect 14369 25412 14381 25415
rect 11103 25384 14381 25412
rect 11103 25381 11115 25384
rect 11057 25375 11115 25381
rect 14369 25381 14381 25384
rect 14415 25381 14427 25415
rect 14369 25375 14427 25381
rect 14642 25372 14648 25424
rect 14700 25412 14706 25424
rect 15654 25412 15660 25424
rect 14700 25384 15660 25412
rect 14700 25372 14706 25384
rect 15654 25372 15660 25384
rect 15712 25372 15718 25424
rect 15841 25415 15899 25421
rect 15841 25412 15853 25415
rect 15764 25384 15853 25412
rect 15764 25356 15792 25384
rect 15841 25381 15853 25384
rect 15887 25381 15899 25415
rect 15841 25375 15899 25381
rect 15930 25372 15936 25424
rect 15988 25412 15994 25424
rect 19996 25412 20024 25440
rect 15988 25384 20024 25412
rect 20180 25412 20208 25443
rect 24762 25440 24768 25452
rect 24820 25440 24826 25492
rect 24578 25412 24584 25424
rect 20180 25384 24584 25412
rect 15988 25372 15994 25384
rect 24578 25372 24584 25384
rect 24636 25372 24642 25424
rect 1394 25344 1400 25356
rect 1355 25316 1400 25344
rect 1394 25304 1400 25316
rect 1452 25304 1458 25356
rect 8573 25347 8631 25353
rect 8573 25313 8585 25347
rect 8619 25344 8631 25347
rect 8662 25344 8668 25356
rect 8619 25316 8668 25344
rect 8619 25313 8631 25316
rect 8573 25307 8631 25313
rect 8662 25304 8668 25316
rect 8720 25304 8726 25356
rect 9306 25304 9312 25356
rect 9364 25344 9370 25356
rect 9582 25344 9588 25356
rect 9364 25316 9588 25344
rect 9364 25304 9370 25316
rect 9582 25304 9588 25316
rect 9640 25304 9646 25356
rect 10321 25347 10379 25353
rect 10321 25313 10333 25347
rect 10367 25344 10379 25347
rect 10962 25344 10968 25356
rect 10367 25316 10968 25344
rect 10367 25313 10379 25316
rect 10321 25307 10379 25313
rect 10962 25304 10968 25316
rect 11020 25304 11026 25356
rect 11425 25347 11483 25353
rect 11425 25313 11437 25347
rect 11471 25344 11483 25347
rect 11606 25344 11612 25356
rect 11471 25316 11612 25344
rect 11471 25313 11483 25316
rect 11425 25307 11483 25313
rect 11606 25304 11612 25316
rect 11664 25304 11670 25356
rect 11790 25304 11796 25356
rect 11848 25344 11854 25356
rect 12161 25347 12219 25353
rect 12161 25344 12173 25347
rect 11848 25316 12173 25344
rect 11848 25304 11854 25316
rect 12161 25313 12173 25316
rect 12207 25313 12219 25347
rect 12986 25344 12992 25356
rect 12947 25316 12992 25344
rect 12161 25307 12219 25313
rect 12986 25304 12992 25316
rect 13044 25304 13050 25356
rect 13906 25304 13912 25356
rect 13964 25344 13970 25356
rect 14093 25347 14151 25353
rect 14093 25344 14105 25347
rect 13964 25316 14105 25344
rect 13964 25304 13970 25316
rect 14093 25313 14105 25316
rect 14139 25313 14151 25347
rect 14093 25307 14151 25313
rect 15746 25304 15752 25356
rect 15804 25304 15810 25356
rect 17126 25344 17132 25356
rect 15856 25316 16988 25344
rect 17087 25316 17132 25344
rect 8481 25279 8539 25285
rect 8481 25245 8493 25279
rect 8527 25276 8539 25279
rect 12805 25279 12863 25285
rect 12805 25276 12817 25279
rect 8527 25248 12817 25276
rect 8527 25245 8539 25248
rect 8481 25239 8539 25245
rect 12805 25245 12817 25248
rect 12851 25276 12863 25279
rect 13814 25276 13820 25288
rect 12851 25248 13820 25276
rect 12851 25245 12863 25248
rect 12805 25239 12863 25245
rect 13814 25236 13820 25248
rect 13872 25276 13878 25288
rect 15856 25276 15884 25316
rect 13872 25248 15884 25276
rect 13872 25236 13878 25248
rect 15930 25236 15936 25288
rect 15988 25276 15994 25288
rect 16114 25276 16120 25288
rect 15988 25248 16033 25276
rect 16075 25248 16120 25276
rect 15988 25236 15994 25248
rect 16114 25236 16120 25248
rect 16172 25236 16178 25288
rect 16482 25236 16488 25288
rect 16540 25276 16546 25288
rect 16853 25279 16911 25285
rect 16853 25276 16865 25279
rect 16540 25248 16865 25276
rect 16540 25236 16546 25248
rect 16853 25245 16865 25248
rect 16899 25245 16911 25279
rect 16960 25276 16988 25316
rect 17126 25304 17132 25316
rect 17184 25304 17190 25356
rect 17681 25347 17739 25353
rect 17681 25344 17693 25347
rect 17236 25316 17693 25344
rect 17236 25276 17264 25316
rect 17681 25313 17693 25316
rect 17727 25344 17739 25347
rect 18509 25347 18567 25353
rect 18509 25344 18521 25347
rect 17727 25316 18521 25344
rect 17727 25313 17739 25316
rect 17681 25307 17739 25313
rect 18509 25313 18521 25316
rect 18555 25313 18567 25347
rect 18874 25344 18880 25356
rect 18835 25316 18880 25344
rect 18509 25307 18567 25313
rect 18874 25304 18880 25316
rect 18932 25304 18938 25356
rect 19981 25347 20039 25353
rect 19981 25313 19993 25347
rect 20027 25344 20039 25347
rect 20622 25344 20628 25356
rect 20027 25316 20628 25344
rect 20027 25313 20039 25316
rect 19981 25307 20039 25313
rect 20622 25304 20628 25316
rect 20680 25304 20686 25356
rect 21174 25304 21180 25356
rect 21232 25344 21238 25356
rect 21269 25347 21327 25353
rect 21269 25344 21281 25347
rect 21232 25316 21281 25344
rect 21232 25304 21238 25316
rect 21269 25313 21281 25316
rect 21315 25313 21327 25347
rect 22738 25344 22744 25356
rect 22699 25316 22744 25344
rect 21269 25307 21327 25313
rect 22738 25304 22744 25316
rect 22796 25304 22802 25356
rect 22833 25347 22891 25353
rect 22833 25313 22845 25347
rect 22879 25344 22891 25347
rect 22922 25344 22928 25356
rect 22879 25316 22928 25344
rect 22879 25313 22891 25316
rect 22833 25307 22891 25313
rect 22922 25304 22928 25316
rect 22980 25304 22986 25356
rect 24026 25304 24032 25356
rect 24084 25344 24090 25356
rect 24397 25347 24455 25353
rect 24397 25344 24409 25347
rect 24084 25316 24409 25344
rect 24084 25304 24090 25316
rect 24397 25313 24409 25316
rect 24443 25313 24455 25347
rect 24397 25307 24455 25313
rect 22462 25276 22468 25288
rect 16960 25248 17264 25276
rect 17328 25248 22468 25276
rect 16853 25239 16911 25245
rect 7098 25168 7104 25220
rect 7156 25208 7162 25220
rect 7837 25211 7895 25217
rect 7837 25208 7849 25211
rect 7156 25180 7849 25208
rect 7156 25168 7162 25180
rect 7837 25177 7849 25180
rect 7883 25208 7895 25211
rect 9217 25211 9275 25217
rect 9217 25208 9229 25211
rect 7883 25180 9229 25208
rect 7883 25177 7895 25180
rect 7837 25171 7895 25177
rect 9217 25177 9229 25180
rect 9263 25208 9275 25211
rect 9585 25211 9643 25217
rect 9585 25208 9597 25211
rect 9263 25180 9597 25208
rect 9263 25177 9275 25180
rect 9217 25171 9275 25177
rect 9585 25177 9597 25180
rect 9631 25208 9643 25211
rect 9766 25208 9772 25220
rect 9631 25180 9772 25208
rect 9631 25177 9643 25180
rect 9585 25171 9643 25177
rect 9766 25168 9772 25180
rect 9824 25208 9830 25220
rect 9953 25211 10011 25217
rect 9953 25208 9965 25211
rect 9824 25180 9965 25208
rect 9824 25168 9830 25180
rect 9953 25177 9965 25180
rect 9999 25208 10011 25211
rect 11241 25211 11299 25217
rect 11241 25208 11253 25211
rect 9999 25180 11253 25208
rect 9999 25177 10011 25180
rect 9953 25171 10011 25177
rect 11241 25177 11253 25180
rect 11287 25208 11299 25211
rect 11790 25208 11796 25220
rect 11287 25180 11796 25208
rect 11287 25177 11299 25180
rect 11241 25171 11299 25177
rect 11790 25168 11796 25180
rect 11848 25168 11854 25220
rect 17218 25208 17224 25220
rect 11900 25180 15884 25208
rect 1581 25143 1639 25149
rect 1581 25109 1593 25143
rect 1627 25140 1639 25143
rect 2774 25140 2780 25152
rect 1627 25112 2780 25140
rect 1627 25109 1639 25112
rect 1581 25103 1639 25109
rect 2774 25100 2780 25112
rect 2832 25100 2838 25152
rect 7374 25100 7380 25152
rect 7432 25140 7438 25152
rect 11057 25143 11115 25149
rect 11057 25140 11069 25143
rect 7432 25112 11069 25140
rect 7432 25100 7438 25112
rect 11057 25109 11069 25112
rect 11103 25109 11115 25143
rect 11057 25103 11115 25109
rect 11609 25143 11667 25149
rect 11609 25109 11621 25143
rect 11655 25140 11667 25143
rect 11900 25140 11928 25180
rect 11655 25112 11928 25140
rect 11655 25109 11667 25112
rect 11609 25103 11667 25109
rect 13170 25100 13176 25152
rect 13228 25140 13234 25152
rect 13538 25140 13544 25152
rect 13228 25112 13273 25140
rect 13499 25112 13544 25140
rect 13228 25100 13234 25112
rect 13538 25100 13544 25112
rect 13596 25100 13602 25152
rect 13906 25140 13912 25152
rect 13867 25112 13912 25140
rect 13906 25100 13912 25112
rect 13964 25100 13970 25152
rect 14734 25100 14740 25152
rect 14792 25140 14798 25152
rect 14829 25143 14887 25149
rect 14829 25140 14841 25143
rect 14792 25112 14841 25140
rect 14792 25100 14798 25112
rect 14829 25109 14841 25112
rect 14875 25109 14887 25143
rect 15286 25140 15292 25152
rect 15247 25112 15292 25140
rect 14829 25103 14887 25109
rect 15286 25100 15292 25112
rect 15344 25100 15350 25152
rect 15470 25140 15476 25152
rect 15431 25112 15476 25140
rect 15470 25100 15476 25112
rect 15528 25100 15534 25152
rect 15856 25140 15884 25180
rect 16040 25180 17224 25208
rect 16040 25140 16068 25180
rect 17218 25168 17224 25180
rect 17276 25168 17282 25220
rect 17328 25217 17356 25248
rect 22462 25236 22468 25248
rect 22520 25236 22526 25288
rect 23014 25276 23020 25288
rect 22975 25248 23020 25276
rect 23014 25236 23020 25248
rect 23072 25236 23078 25288
rect 23566 25236 23572 25288
rect 23624 25276 23630 25288
rect 24489 25279 24547 25285
rect 24489 25276 24501 25279
rect 23624 25248 24501 25276
rect 23624 25236 23630 25248
rect 24489 25245 24501 25248
rect 24535 25245 24547 25279
rect 24489 25239 24547 25245
rect 24581 25279 24639 25285
rect 24581 25245 24593 25279
rect 24627 25245 24639 25279
rect 24581 25239 24639 25245
rect 17313 25211 17371 25217
rect 17313 25177 17325 25211
rect 17359 25177 17371 25211
rect 18966 25208 18972 25220
rect 17313 25171 17371 25177
rect 17420 25180 18972 25208
rect 15856 25112 16068 25140
rect 16577 25143 16635 25149
rect 16577 25109 16589 25143
rect 16623 25140 16635 25143
rect 16758 25140 16764 25152
rect 16623 25112 16764 25140
rect 16623 25109 16635 25112
rect 16577 25103 16635 25109
rect 16758 25100 16764 25112
rect 16816 25100 16822 25152
rect 16850 25100 16856 25152
rect 16908 25140 16914 25152
rect 17420 25140 17448 25180
rect 18966 25168 18972 25180
rect 19024 25168 19030 25220
rect 19061 25211 19119 25217
rect 19061 25177 19073 25211
rect 19107 25208 19119 25211
rect 21818 25208 21824 25220
rect 19107 25180 21824 25208
rect 19107 25177 19119 25180
rect 19061 25171 19119 25177
rect 21818 25168 21824 25180
rect 21876 25168 21882 25220
rect 22097 25211 22155 25217
rect 22097 25177 22109 25211
rect 22143 25208 22155 25211
rect 23032 25208 23060 25236
rect 24596 25208 24624 25239
rect 25038 25208 25044 25220
rect 22143 25180 25044 25208
rect 22143 25177 22155 25180
rect 22097 25171 22155 25177
rect 25038 25168 25044 25180
rect 25096 25168 25102 25220
rect 18046 25140 18052 25152
rect 16908 25112 17448 25140
rect 18007 25112 18052 25140
rect 16908 25100 16914 25112
rect 18046 25100 18052 25112
rect 18104 25100 18110 25152
rect 20990 25140 20996 25152
rect 20951 25112 20996 25140
rect 20990 25100 20996 25112
rect 21048 25100 21054 25152
rect 22373 25143 22431 25149
rect 22373 25109 22385 25143
rect 22419 25140 22431 25143
rect 23474 25140 23480 25152
rect 22419 25112 23480 25140
rect 22419 25109 22431 25112
rect 22373 25103 22431 25109
rect 23474 25100 23480 25112
rect 23532 25100 23538 25152
rect 24029 25143 24087 25149
rect 24029 25109 24041 25143
rect 24075 25140 24087 25143
rect 24118 25140 24124 25152
rect 24075 25112 24124 25140
rect 24075 25109 24087 25112
rect 24029 25103 24087 25109
rect 24118 25100 24124 25112
rect 24176 25100 24182 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1578 24936 1584 24948
rect 1539 24908 1584 24936
rect 1578 24896 1584 24908
rect 1636 24896 1642 24948
rect 7098 24936 7104 24948
rect 7059 24908 7104 24936
rect 7098 24896 7104 24908
rect 7156 24896 7162 24948
rect 7650 24936 7656 24948
rect 7611 24908 7656 24936
rect 7650 24896 7656 24908
rect 7708 24896 7714 24948
rect 8754 24936 8760 24948
rect 8715 24908 8760 24936
rect 8754 24896 8760 24908
rect 8812 24896 8818 24948
rect 9306 24896 9312 24948
rect 9364 24936 9370 24948
rect 13906 24936 13912 24948
rect 9364 24908 13912 24936
rect 9364 24896 9370 24908
rect 13906 24896 13912 24908
rect 13964 24896 13970 24948
rect 14642 24896 14648 24948
rect 14700 24896 14706 24948
rect 16850 24936 16856 24948
rect 15120 24908 16856 24936
rect 8481 24871 8539 24877
rect 8481 24837 8493 24871
rect 8527 24868 8539 24871
rect 8662 24868 8668 24880
rect 8527 24840 8668 24868
rect 8527 24837 8539 24840
rect 8481 24831 8539 24837
rect 8662 24828 8668 24840
rect 8720 24828 8726 24880
rect 9861 24871 9919 24877
rect 9861 24837 9873 24871
rect 9907 24868 9919 24871
rect 9950 24868 9956 24880
rect 9907 24840 9956 24868
rect 9907 24837 9919 24840
rect 9861 24831 9919 24837
rect 9950 24828 9956 24840
rect 10008 24828 10014 24880
rect 10686 24828 10692 24880
rect 10744 24868 10750 24880
rect 14660 24868 14688 24896
rect 10744 24840 14688 24868
rect 10744 24828 10750 24840
rect 14918 24828 14924 24880
rect 14976 24868 14982 24880
rect 15120 24868 15148 24908
rect 16850 24896 16856 24908
rect 16908 24896 16914 24948
rect 17218 24896 17224 24948
rect 17276 24936 17282 24948
rect 22646 24936 22652 24948
rect 17276 24908 22652 24936
rect 17276 24896 17282 24908
rect 22646 24896 22652 24908
rect 22704 24896 22710 24948
rect 22922 24896 22928 24948
rect 22980 24936 22986 24948
rect 23017 24939 23075 24945
rect 23017 24936 23029 24939
rect 22980 24908 23029 24936
rect 22980 24896 22986 24908
rect 23017 24905 23029 24908
rect 23063 24905 23075 24939
rect 23017 24899 23075 24905
rect 15470 24868 15476 24880
rect 14976 24840 15148 24868
rect 15212 24840 15476 24868
rect 14976 24828 14982 24840
rect 9490 24760 9496 24812
rect 9548 24800 9554 24812
rect 9585 24803 9643 24809
rect 9585 24800 9597 24803
rect 9548 24772 9597 24800
rect 9548 24760 9554 24772
rect 9585 24769 9597 24772
rect 9631 24800 9643 24803
rect 11422 24800 11428 24812
rect 9631 24772 11284 24800
rect 11383 24772 11428 24800
rect 9631 24769 9643 24772
rect 9585 24763 9643 24769
rect 1397 24735 1455 24741
rect 1397 24701 1409 24735
rect 1443 24732 1455 24735
rect 2501 24735 2559 24741
rect 1443 24704 2452 24732
rect 1443 24701 1455 24704
rect 1397 24695 1455 24701
rect 2424 24608 2452 24704
rect 2501 24701 2513 24735
rect 2547 24732 2559 24735
rect 7469 24735 7527 24741
rect 2547 24704 3096 24732
rect 2547 24701 2559 24704
rect 2501 24695 2559 24701
rect 3068 24608 3096 24704
rect 7469 24701 7481 24735
rect 7515 24732 7527 24735
rect 7558 24732 7564 24744
rect 7515 24704 7564 24732
rect 7515 24701 7527 24704
rect 7469 24695 7527 24701
rect 7558 24692 7564 24704
rect 7616 24732 7622 24744
rect 8021 24735 8079 24741
rect 8021 24732 8033 24735
rect 7616 24704 8033 24732
rect 7616 24692 7622 24704
rect 8021 24701 8033 24704
rect 8067 24701 8079 24735
rect 8021 24695 8079 24701
rect 8573 24735 8631 24741
rect 8573 24701 8585 24735
rect 8619 24732 8631 24735
rect 8754 24732 8760 24744
rect 8619 24704 8760 24732
rect 8619 24701 8631 24704
rect 8573 24695 8631 24701
rect 8754 24692 8760 24704
rect 8812 24732 8818 24744
rect 9692 24741 9720 24772
rect 9125 24735 9183 24741
rect 9125 24732 9137 24735
rect 8812 24704 9137 24732
rect 8812 24692 8818 24704
rect 9125 24701 9137 24704
rect 9171 24701 9183 24735
rect 9125 24695 9183 24701
rect 9677 24735 9735 24741
rect 9677 24701 9689 24735
rect 9723 24732 9735 24735
rect 10321 24735 10379 24741
rect 9723 24704 9757 24732
rect 9723 24701 9735 24704
rect 9677 24695 9735 24701
rect 10321 24701 10333 24735
rect 10367 24732 10379 24735
rect 11146 24732 11152 24744
rect 10367 24704 11152 24732
rect 10367 24701 10379 24704
rect 10321 24695 10379 24701
rect 11146 24692 11152 24704
rect 11204 24692 11210 24744
rect 11256 24732 11284 24772
rect 11422 24760 11428 24772
rect 11480 24760 11486 24812
rect 11606 24760 11612 24812
rect 11664 24800 11670 24812
rect 11793 24803 11851 24809
rect 11793 24800 11805 24803
rect 11664 24772 11805 24800
rect 11664 24760 11670 24772
rect 11793 24769 11805 24772
rect 11839 24800 11851 24803
rect 11974 24800 11980 24812
rect 11839 24772 11980 24800
rect 11839 24769 11851 24772
rect 11793 24763 11851 24769
rect 11974 24760 11980 24772
rect 12032 24760 12038 24812
rect 13630 24800 13636 24812
rect 13591 24772 13636 24800
rect 13630 24760 13636 24772
rect 13688 24760 13694 24812
rect 15212 24809 15240 24840
rect 15470 24828 15476 24840
rect 15528 24828 15534 24880
rect 16298 24828 16304 24880
rect 16356 24868 16362 24880
rect 18046 24868 18052 24880
rect 16356 24840 18052 24868
rect 16356 24828 16362 24840
rect 18046 24828 18052 24840
rect 18104 24828 18110 24880
rect 19978 24828 19984 24880
rect 20036 24868 20042 24880
rect 22186 24868 22192 24880
rect 20036 24840 22192 24868
rect 20036 24828 20042 24840
rect 22186 24828 22192 24840
rect 22244 24828 22250 24880
rect 22940 24868 22968 24896
rect 22296 24840 22968 24868
rect 14277 24803 14335 24809
rect 14277 24769 14289 24803
rect 14323 24800 14335 24803
rect 15197 24803 15255 24809
rect 15197 24800 15209 24803
rect 14323 24772 15209 24800
rect 14323 24769 14335 24772
rect 14277 24763 14335 24769
rect 15197 24769 15209 24772
rect 15243 24769 15255 24803
rect 15197 24763 15255 24769
rect 15381 24803 15439 24809
rect 15381 24769 15393 24803
rect 15427 24800 15439 24803
rect 16850 24800 16856 24812
rect 15427 24772 16856 24800
rect 15427 24769 15439 24772
rect 15381 24763 15439 24769
rect 16850 24760 16856 24772
rect 16908 24760 16914 24812
rect 17126 24760 17132 24812
rect 17184 24760 17190 24812
rect 12250 24732 12256 24744
rect 11256 24704 12256 24732
rect 12250 24692 12256 24704
rect 12308 24692 12314 24744
rect 13078 24692 13084 24744
rect 13136 24732 13142 24744
rect 13449 24735 13507 24741
rect 13449 24732 13461 24735
rect 13136 24704 13461 24732
rect 13136 24692 13142 24704
rect 13449 24701 13461 24704
rect 13495 24732 13507 24735
rect 13538 24732 13544 24744
rect 13495 24704 13544 24732
rect 13495 24701 13507 24704
rect 13449 24695 13507 24701
rect 13538 24692 13544 24704
rect 13596 24692 13602 24744
rect 15102 24732 15108 24744
rect 15063 24704 15108 24732
rect 15102 24692 15108 24704
rect 15160 24692 15166 24744
rect 15746 24692 15752 24744
rect 15804 24732 15810 24744
rect 15930 24732 15936 24744
rect 15804 24704 15936 24732
rect 15804 24692 15810 24704
rect 15930 24692 15936 24704
rect 15988 24732 15994 24744
rect 16117 24735 16175 24741
rect 16117 24732 16129 24735
rect 15988 24704 16129 24732
rect 15988 24692 15994 24704
rect 16117 24701 16129 24704
rect 16163 24701 16175 24735
rect 17144 24732 17172 24760
rect 18064 24741 18092 24828
rect 18230 24800 18236 24812
rect 18191 24772 18236 24800
rect 18230 24760 18236 24772
rect 18288 24760 18294 24812
rect 21174 24760 21180 24812
rect 21232 24800 21238 24812
rect 21545 24803 21603 24809
rect 21545 24800 21557 24803
rect 21232 24772 21557 24800
rect 21232 24760 21238 24772
rect 21545 24769 21557 24772
rect 21591 24800 21603 24803
rect 22296 24800 22324 24840
rect 22462 24800 22468 24812
rect 21591 24772 22324 24800
rect 22423 24772 22468 24800
rect 21591 24769 21603 24772
rect 21545 24763 21603 24769
rect 22462 24760 22468 24772
rect 22520 24760 22526 24812
rect 22646 24800 22652 24812
rect 22607 24772 22652 24800
rect 22646 24760 22652 24772
rect 22704 24800 22710 24812
rect 23014 24800 23020 24812
rect 22704 24772 23020 24800
rect 22704 24760 22710 24772
rect 23014 24760 23020 24772
rect 23072 24760 23078 24812
rect 25038 24800 25044 24812
rect 24999 24772 25044 24800
rect 25038 24760 25044 24772
rect 25096 24800 25102 24812
rect 25501 24803 25559 24809
rect 25501 24800 25513 24803
rect 25096 24772 25513 24800
rect 25096 24760 25102 24772
rect 25501 24769 25513 24772
rect 25547 24769 25559 24803
rect 25501 24763 25559 24769
rect 17313 24735 17371 24741
rect 17313 24732 17325 24735
rect 16117 24695 16175 24701
rect 16224 24704 17325 24732
rect 10689 24667 10747 24673
rect 10689 24633 10701 24667
rect 10735 24664 10747 24667
rect 12713 24667 12771 24673
rect 10735 24636 11284 24664
rect 10735 24633 10747 24636
rect 10689 24627 10747 24633
rect 11256 24608 11284 24636
rect 12713 24633 12725 24667
rect 12759 24664 12771 24667
rect 13262 24664 13268 24676
rect 12759 24636 13268 24664
rect 12759 24633 12771 24636
rect 12713 24627 12771 24633
rect 13262 24624 13268 24636
rect 13320 24624 13326 24676
rect 14645 24667 14703 24673
rect 14645 24633 14657 24667
rect 14691 24664 14703 24667
rect 16022 24664 16028 24676
rect 14691 24636 16028 24664
rect 14691 24633 14703 24636
rect 14645 24627 14703 24633
rect 16022 24624 16028 24636
rect 16080 24624 16086 24676
rect 1394 24556 1400 24608
rect 1452 24596 1458 24608
rect 2038 24596 2044 24608
rect 1452 24568 2044 24596
rect 1452 24556 1458 24568
rect 2038 24556 2044 24568
rect 2096 24556 2102 24608
rect 2406 24596 2412 24608
rect 2367 24568 2412 24596
rect 2406 24556 2412 24568
rect 2464 24556 2470 24608
rect 2498 24556 2504 24608
rect 2556 24596 2562 24608
rect 2685 24599 2743 24605
rect 2685 24596 2697 24599
rect 2556 24568 2697 24596
rect 2556 24556 2562 24568
rect 2685 24565 2697 24568
rect 2731 24565 2743 24599
rect 3050 24596 3056 24608
rect 3011 24568 3056 24596
rect 2685 24559 2743 24565
rect 3050 24556 3056 24568
rect 3108 24556 3114 24608
rect 10781 24599 10839 24605
rect 10781 24565 10793 24599
rect 10827 24596 10839 24599
rect 10962 24596 10968 24608
rect 10827 24568 10968 24596
rect 10827 24565 10839 24568
rect 10781 24559 10839 24565
rect 10962 24556 10968 24568
rect 11020 24556 11026 24608
rect 11238 24596 11244 24608
rect 11199 24568 11244 24596
rect 11238 24556 11244 24568
rect 11296 24556 11302 24608
rect 12158 24596 12164 24608
rect 12119 24568 12164 24596
rect 12158 24556 12164 24568
rect 12216 24556 12222 24608
rect 12986 24596 12992 24608
rect 12947 24568 12992 24596
rect 12986 24556 12992 24568
rect 13044 24556 13050 24608
rect 14734 24596 14740 24608
rect 14695 24568 14740 24596
rect 14734 24556 14740 24568
rect 14792 24556 14798 24608
rect 15838 24596 15844 24608
rect 15799 24568 15844 24596
rect 15838 24556 15844 24568
rect 15896 24556 15902 24608
rect 15930 24556 15936 24608
rect 15988 24596 15994 24608
rect 16224 24596 16252 24704
rect 17313 24701 17325 24704
rect 17359 24701 17371 24735
rect 17313 24695 17371 24701
rect 18049 24735 18107 24741
rect 18049 24701 18061 24735
rect 18095 24701 18107 24735
rect 19794 24732 19800 24744
rect 19707 24704 19800 24732
rect 18049 24695 18107 24701
rect 17126 24664 17132 24676
rect 16316 24636 17132 24664
rect 16316 24605 16344 24636
rect 17126 24624 17132 24636
rect 17184 24624 17190 24676
rect 17328 24664 17356 24695
rect 19794 24692 19800 24704
rect 19852 24732 19858 24744
rect 20901 24735 20959 24741
rect 19852 24704 20484 24732
rect 19852 24692 19858 24704
rect 19242 24664 19248 24676
rect 17328 24636 19248 24664
rect 19242 24624 19248 24636
rect 19300 24624 19306 24676
rect 15988 24568 16252 24596
rect 16301 24599 16359 24605
rect 15988 24556 15994 24568
rect 16301 24565 16313 24599
rect 16347 24565 16359 24599
rect 16666 24596 16672 24608
rect 16627 24568 16672 24596
rect 16301 24559 16359 24565
rect 16666 24556 16672 24568
rect 16724 24556 16730 24608
rect 16758 24556 16764 24608
rect 16816 24596 16822 24608
rect 17770 24596 17776 24608
rect 16816 24568 16861 24596
rect 17731 24568 17776 24596
rect 16816 24556 16822 24568
rect 17770 24556 17776 24568
rect 17828 24556 17834 24608
rect 18874 24596 18880 24608
rect 18835 24568 18880 24596
rect 18874 24556 18880 24568
rect 18932 24556 18938 24608
rect 19334 24596 19340 24608
rect 19295 24568 19340 24596
rect 19334 24556 19340 24568
rect 19392 24556 19398 24608
rect 19981 24599 20039 24605
rect 19981 24565 19993 24599
rect 20027 24596 20039 24599
rect 20070 24596 20076 24608
rect 20027 24568 20076 24596
rect 20027 24565 20039 24568
rect 19981 24559 20039 24565
rect 20070 24556 20076 24568
rect 20128 24556 20134 24608
rect 20456 24605 20484 24704
rect 20901 24701 20913 24735
rect 20947 24732 20959 24735
rect 20990 24732 20996 24744
rect 20947 24704 20996 24732
rect 20947 24701 20959 24704
rect 20901 24695 20959 24701
rect 20990 24692 20996 24704
rect 21048 24732 21054 24744
rect 21450 24732 21456 24744
rect 21048 24704 21456 24732
rect 21048 24692 21054 24704
rect 21450 24692 21456 24704
rect 21508 24692 21514 24744
rect 22922 24692 22928 24744
rect 22980 24732 22986 24744
rect 24305 24735 24363 24741
rect 24305 24732 24317 24735
rect 22980 24704 24317 24732
rect 22980 24692 22986 24704
rect 24305 24701 24317 24704
rect 24351 24732 24363 24735
rect 24949 24735 25007 24741
rect 24949 24732 24961 24735
rect 24351 24704 24961 24732
rect 24351 24701 24363 24704
rect 24305 24695 24363 24701
rect 24949 24701 24961 24704
rect 24995 24701 25007 24735
rect 24949 24695 25007 24701
rect 21818 24664 21824 24676
rect 21731 24636 21824 24664
rect 21818 24624 21824 24636
rect 21876 24664 21882 24676
rect 22373 24667 22431 24673
rect 22373 24664 22385 24667
rect 21876 24636 22385 24664
rect 21876 24624 21882 24636
rect 22373 24633 22385 24636
rect 22419 24633 22431 24667
rect 24026 24664 24032 24676
rect 22373 24627 22431 24633
rect 23492 24636 24032 24664
rect 20441 24599 20499 24605
rect 20441 24565 20453 24599
rect 20487 24596 20499 24599
rect 20530 24596 20536 24608
rect 20487 24568 20536 24596
rect 20487 24565 20499 24568
rect 20441 24559 20499 24565
rect 20530 24556 20536 24568
rect 20588 24556 20594 24608
rect 20714 24596 20720 24608
rect 20675 24568 20720 24596
rect 20714 24556 20720 24568
rect 20772 24556 20778 24608
rect 21082 24596 21088 24608
rect 21043 24568 21088 24596
rect 21082 24556 21088 24568
rect 21140 24556 21146 24608
rect 21910 24556 21916 24608
rect 21968 24596 21974 24608
rect 22005 24599 22063 24605
rect 22005 24596 22017 24599
rect 21968 24568 22017 24596
rect 21968 24556 21974 24568
rect 22005 24565 22017 24568
rect 22051 24565 22063 24599
rect 22005 24559 22063 24565
rect 22554 24556 22560 24608
rect 22612 24596 22618 24608
rect 23492 24605 23520 24636
rect 24026 24624 24032 24636
rect 24084 24624 24090 24676
rect 24578 24624 24584 24676
rect 24636 24664 24642 24676
rect 24857 24667 24915 24673
rect 24857 24664 24869 24667
rect 24636 24636 24869 24664
rect 24636 24624 24642 24636
rect 24857 24633 24869 24636
rect 24903 24633 24915 24667
rect 24857 24627 24915 24633
rect 23477 24599 23535 24605
rect 23477 24596 23489 24599
rect 22612 24568 23489 24596
rect 22612 24556 22618 24568
rect 23477 24565 23489 24568
rect 23523 24565 23535 24599
rect 23477 24559 23535 24565
rect 23566 24556 23572 24608
rect 23624 24596 23630 24608
rect 23937 24599 23995 24605
rect 23937 24596 23949 24599
rect 23624 24568 23949 24596
rect 23624 24556 23630 24568
rect 23937 24565 23949 24568
rect 23983 24565 23995 24599
rect 23937 24559 23995 24565
rect 24489 24599 24547 24605
rect 24489 24565 24501 24599
rect 24535 24596 24547 24599
rect 24670 24596 24676 24608
rect 24535 24568 24676 24596
rect 24535 24565 24547 24568
rect 24489 24559 24547 24565
rect 24670 24556 24676 24568
rect 24728 24556 24734 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1486 24352 1492 24404
rect 1544 24392 1550 24404
rect 1581 24395 1639 24401
rect 1581 24392 1593 24395
rect 1544 24364 1593 24392
rect 1544 24352 1550 24364
rect 1581 24361 1593 24364
rect 1627 24361 1639 24395
rect 2682 24392 2688 24404
rect 2643 24364 2688 24392
rect 1581 24355 1639 24361
rect 2682 24352 2688 24364
rect 2740 24352 2746 24404
rect 6362 24392 6368 24404
rect 6323 24364 6368 24392
rect 6362 24352 6368 24364
rect 6420 24352 6426 24404
rect 7561 24395 7619 24401
rect 7561 24361 7573 24395
rect 7607 24392 7619 24395
rect 7742 24392 7748 24404
rect 7607 24364 7748 24392
rect 7607 24361 7619 24364
rect 7561 24355 7619 24361
rect 7742 24352 7748 24364
rect 7800 24352 7806 24404
rect 8294 24392 8300 24404
rect 8255 24364 8300 24392
rect 8294 24352 8300 24364
rect 8352 24352 8358 24404
rect 8665 24395 8723 24401
rect 8665 24361 8677 24395
rect 8711 24392 8723 24395
rect 8846 24392 8852 24404
rect 8711 24364 8852 24392
rect 8711 24361 8723 24364
rect 8665 24355 8723 24361
rect 8846 24352 8852 24364
rect 8904 24352 8910 24404
rect 11054 24352 11060 24404
rect 11112 24392 11118 24404
rect 11606 24392 11612 24404
rect 11112 24364 11612 24392
rect 11112 24352 11118 24364
rect 11606 24352 11612 24364
rect 11664 24352 11670 24404
rect 12069 24395 12127 24401
rect 12069 24361 12081 24395
rect 12115 24392 12127 24395
rect 12158 24392 12164 24404
rect 12115 24364 12164 24392
rect 12115 24361 12127 24364
rect 12069 24355 12127 24361
rect 12158 24352 12164 24364
rect 12216 24352 12222 24404
rect 12434 24352 12440 24404
rect 12492 24392 12498 24404
rect 18230 24392 18236 24404
rect 12492 24364 18236 24392
rect 12492 24352 12498 24364
rect 18230 24352 18236 24364
rect 18288 24352 18294 24404
rect 19889 24395 19947 24401
rect 19889 24361 19901 24395
rect 19935 24392 19947 24395
rect 19978 24392 19984 24404
rect 19935 24364 19984 24392
rect 19935 24361 19947 24364
rect 19889 24355 19947 24361
rect 19978 24352 19984 24364
rect 20036 24352 20042 24404
rect 21358 24352 21364 24404
rect 21416 24392 21422 24404
rect 21453 24395 21511 24401
rect 21453 24392 21465 24395
rect 21416 24364 21465 24392
rect 21416 24352 21422 24364
rect 21453 24361 21465 24364
rect 21499 24361 21511 24395
rect 21453 24355 21511 24361
rect 22097 24395 22155 24401
rect 22097 24361 22109 24395
rect 22143 24392 22155 24395
rect 22462 24392 22468 24404
rect 22143 24364 22468 24392
rect 22143 24361 22155 24364
rect 22097 24355 22155 24361
rect 22462 24352 22468 24364
rect 22520 24352 22526 24404
rect 6089 24327 6147 24333
rect 6089 24293 6101 24327
rect 6135 24324 6147 24327
rect 7098 24324 7104 24336
rect 6135 24296 7104 24324
rect 6135 24293 6147 24296
rect 6089 24287 6147 24293
rect 7098 24284 7104 24296
rect 7156 24284 7162 24336
rect 13538 24284 13544 24336
rect 13596 24324 13602 24336
rect 13725 24327 13783 24333
rect 13725 24324 13737 24327
rect 13596 24296 13737 24324
rect 13596 24284 13602 24296
rect 13725 24293 13737 24296
rect 13771 24293 13783 24327
rect 13725 24287 13783 24293
rect 14829 24327 14887 24333
rect 14829 24293 14841 24327
rect 14875 24324 14887 24327
rect 16393 24327 16451 24333
rect 16393 24324 16405 24327
rect 14875 24296 16405 24324
rect 14875 24293 14887 24296
rect 14829 24287 14887 24293
rect 16393 24293 16405 24296
rect 16439 24324 16451 24327
rect 16850 24324 16856 24336
rect 16439 24296 16856 24324
rect 16439 24293 16451 24296
rect 16393 24287 16451 24293
rect 16850 24284 16856 24296
rect 16908 24324 16914 24336
rect 17402 24324 17408 24336
rect 16908 24296 17408 24324
rect 16908 24284 16914 24296
rect 17402 24284 17408 24296
rect 17460 24284 17466 24336
rect 23293 24327 23351 24333
rect 23293 24293 23305 24327
rect 23339 24324 23351 24327
rect 23339 24296 23888 24324
rect 23339 24293 23351 24296
rect 23293 24287 23351 24293
rect 23860 24268 23888 24296
rect 23934 24284 23940 24336
rect 23992 24324 23998 24336
rect 23992 24296 24992 24324
rect 23992 24284 23998 24296
rect 24964 24268 24992 24296
rect 1397 24259 1455 24265
rect 1397 24225 1409 24259
rect 1443 24256 1455 24259
rect 2130 24256 2136 24268
rect 1443 24228 2136 24256
rect 1443 24225 1455 24228
rect 1397 24219 1455 24225
rect 2130 24216 2136 24228
rect 2188 24216 2194 24268
rect 2501 24259 2559 24265
rect 2501 24225 2513 24259
rect 2547 24256 2559 24259
rect 2590 24256 2596 24268
rect 2547 24228 2596 24256
rect 2547 24225 2559 24228
rect 2501 24219 2559 24225
rect 2590 24216 2596 24228
rect 2648 24216 2654 24268
rect 6178 24256 6184 24268
rect 6139 24228 6184 24256
rect 6178 24216 6184 24228
rect 6236 24216 6242 24268
rect 7374 24256 7380 24268
rect 7335 24228 7380 24256
rect 7374 24216 7380 24228
rect 7432 24216 7438 24268
rect 8478 24256 8484 24268
rect 8439 24228 8484 24256
rect 8478 24216 8484 24228
rect 8536 24216 8542 24268
rect 10502 24256 10508 24268
rect 10463 24228 10508 24256
rect 10502 24216 10508 24228
rect 10560 24216 10566 24268
rect 10597 24259 10655 24265
rect 10597 24225 10609 24259
rect 10643 24256 10655 24259
rect 10870 24256 10876 24268
rect 10643 24228 10876 24256
rect 10643 24225 10655 24228
rect 10597 24219 10655 24225
rect 10870 24216 10876 24228
rect 10928 24216 10934 24268
rect 11609 24259 11667 24265
rect 11609 24225 11621 24259
rect 11655 24256 11667 24259
rect 12161 24259 12219 24265
rect 12161 24256 12173 24259
rect 11655 24228 12173 24256
rect 11655 24225 11667 24228
rect 11609 24219 11667 24225
rect 12161 24225 12173 24228
rect 12207 24256 12219 24259
rect 12342 24256 12348 24268
rect 12207 24228 12348 24256
rect 12207 24225 12219 24228
rect 12161 24219 12219 24225
rect 12342 24216 12348 24228
rect 12400 24216 12406 24268
rect 13446 24216 13452 24268
rect 13504 24256 13510 24268
rect 13633 24259 13691 24265
rect 13633 24256 13645 24259
rect 13504 24228 13645 24256
rect 13504 24216 13510 24228
rect 13633 24225 13645 24228
rect 13679 24225 13691 24259
rect 13633 24219 13691 24225
rect 15470 24216 15476 24268
rect 15528 24256 15534 24268
rect 15657 24259 15715 24265
rect 15657 24256 15669 24259
rect 15528 24228 15669 24256
rect 15528 24216 15534 24228
rect 15657 24225 15669 24228
rect 15703 24225 15715 24259
rect 15657 24219 15715 24225
rect 16022 24216 16028 24268
rect 16080 24256 16086 24268
rect 17221 24259 17279 24265
rect 16080 24228 17172 24256
rect 16080 24216 16086 24228
rect 10778 24188 10784 24200
rect 10739 24160 10784 24188
rect 10778 24148 10784 24160
rect 10836 24148 10842 24200
rect 12066 24148 12072 24200
rect 12124 24188 12130 24200
rect 12253 24191 12311 24197
rect 12253 24188 12265 24191
rect 12124 24160 12265 24188
rect 12124 24148 12130 24160
rect 12253 24157 12265 24160
rect 12299 24157 12311 24191
rect 12253 24151 12311 24157
rect 13173 24191 13231 24197
rect 13173 24157 13185 24191
rect 13219 24188 13231 24191
rect 13354 24188 13360 24200
rect 13219 24160 13360 24188
rect 13219 24157 13231 24160
rect 13173 24151 13231 24157
rect 13354 24148 13360 24160
rect 13412 24148 13418 24200
rect 13817 24191 13875 24197
rect 13817 24157 13829 24191
rect 13863 24157 13875 24191
rect 13817 24151 13875 24157
rect 3145 24123 3203 24129
rect 3145 24120 3157 24123
rect 2332 24092 3157 24120
rect 2332 24061 2360 24092
rect 3145 24089 3157 24092
rect 3191 24120 3203 24123
rect 3510 24120 3516 24132
rect 3191 24092 3516 24120
rect 3191 24089 3203 24092
rect 3145 24083 3203 24089
rect 3510 24080 3516 24092
rect 3568 24120 3574 24132
rect 4341 24123 4399 24129
rect 4341 24120 4353 24123
rect 3568 24092 4353 24120
rect 3568 24080 3574 24092
rect 4341 24089 4353 24092
rect 4387 24120 4399 24123
rect 4893 24123 4951 24129
rect 4893 24120 4905 24123
rect 4387 24092 4905 24120
rect 4387 24089 4399 24092
rect 4341 24083 4399 24089
rect 4893 24089 4905 24092
rect 4939 24120 4951 24123
rect 4939 24092 6316 24120
rect 4939 24089 4951 24092
rect 4893 24083 4951 24089
rect 6288 24064 6316 24092
rect 9674 24080 9680 24132
rect 9732 24120 9738 24132
rect 10137 24123 10195 24129
rect 10137 24120 10149 24123
rect 9732 24092 10149 24120
rect 9732 24080 9738 24092
rect 10137 24089 10149 24092
rect 10183 24089 10195 24123
rect 10137 24083 10195 24089
rect 11241 24123 11299 24129
rect 11241 24089 11253 24123
rect 11287 24120 11299 24123
rect 11422 24120 11428 24132
rect 11287 24092 11428 24120
rect 11287 24089 11299 24092
rect 11241 24083 11299 24089
rect 11422 24080 11428 24092
rect 11480 24120 11486 24132
rect 13538 24120 13544 24132
rect 11480 24092 13544 24120
rect 11480 24080 11486 24092
rect 13538 24080 13544 24092
rect 13596 24120 13602 24132
rect 13832 24120 13860 24151
rect 15562 24148 15568 24200
rect 15620 24188 15626 24200
rect 15749 24191 15807 24197
rect 15749 24188 15761 24191
rect 15620 24160 15761 24188
rect 15620 24148 15626 24160
rect 15749 24157 15761 24160
rect 15795 24157 15807 24191
rect 15749 24151 15807 24157
rect 15933 24191 15991 24197
rect 15933 24157 15945 24191
rect 15979 24188 15991 24191
rect 16206 24188 16212 24200
rect 15979 24160 16212 24188
rect 15979 24157 15991 24160
rect 15933 24151 15991 24157
rect 13596 24092 13860 24120
rect 14461 24123 14519 24129
rect 13596 24080 13602 24092
rect 14461 24089 14473 24123
rect 14507 24120 14519 24123
rect 15948 24120 15976 24151
rect 16206 24148 16212 24160
rect 16264 24148 16270 24200
rect 14507 24092 15976 24120
rect 14507 24089 14519 24092
rect 14461 24083 14519 24089
rect 16666 24080 16672 24132
rect 16724 24120 16730 24132
rect 16761 24123 16819 24129
rect 16761 24120 16773 24123
rect 16724 24092 16773 24120
rect 16724 24080 16730 24092
rect 16761 24089 16773 24092
rect 16807 24120 16819 24123
rect 17034 24120 17040 24132
rect 16807 24092 17040 24120
rect 16807 24089 16819 24092
rect 16761 24083 16819 24089
rect 17034 24080 17040 24092
rect 17092 24080 17098 24132
rect 17144 24120 17172 24228
rect 17221 24225 17233 24259
rect 17267 24256 17279 24259
rect 17494 24256 17500 24268
rect 17267 24228 17500 24256
rect 17267 24225 17279 24228
rect 17221 24219 17279 24225
rect 17494 24216 17500 24228
rect 17552 24216 17558 24268
rect 17954 24216 17960 24268
rect 18012 24256 18018 24268
rect 18417 24259 18475 24265
rect 18417 24256 18429 24259
rect 18012 24228 18429 24256
rect 18012 24216 18018 24228
rect 18417 24225 18429 24228
rect 18463 24256 18475 24259
rect 19153 24259 19211 24265
rect 19153 24256 19165 24259
rect 18463 24228 19165 24256
rect 18463 24225 18475 24228
rect 18417 24219 18475 24225
rect 19153 24225 19165 24228
rect 19199 24225 19211 24259
rect 19153 24219 19211 24225
rect 19705 24259 19763 24265
rect 19705 24225 19717 24259
rect 19751 24256 19763 24259
rect 20346 24256 20352 24268
rect 19751 24228 20352 24256
rect 19751 24225 19763 24228
rect 19705 24219 19763 24225
rect 20346 24216 20352 24228
rect 20404 24216 20410 24268
rect 21266 24216 21272 24268
rect 21324 24256 21330 24268
rect 21361 24259 21419 24265
rect 21361 24256 21373 24259
rect 21324 24228 21373 24256
rect 21324 24216 21330 24228
rect 21361 24225 21373 24228
rect 21407 24225 21419 24259
rect 21361 24219 21419 24225
rect 22465 24259 22523 24265
rect 22465 24225 22477 24259
rect 22511 24256 22523 24259
rect 22738 24256 22744 24268
rect 22511 24228 22744 24256
rect 22511 24225 22523 24228
rect 22465 24219 22523 24225
rect 22738 24216 22744 24228
rect 22796 24216 22802 24268
rect 23750 24256 23756 24268
rect 23711 24228 23756 24256
rect 23750 24216 23756 24228
rect 23808 24216 23814 24268
rect 23842 24216 23848 24268
rect 23900 24256 23906 24268
rect 24486 24256 24492 24268
rect 23900 24228 23945 24256
rect 24447 24228 24492 24256
rect 23900 24216 23906 24228
rect 24486 24216 24492 24228
rect 24544 24216 24550 24268
rect 24946 24256 24952 24268
rect 24859 24228 24952 24256
rect 24946 24216 24952 24228
rect 25004 24216 25010 24268
rect 17310 24188 17316 24200
rect 17271 24160 17316 24188
rect 17310 24148 17316 24160
rect 17368 24148 17374 24200
rect 17405 24191 17463 24197
rect 17405 24157 17417 24191
rect 17451 24157 17463 24191
rect 18690 24188 18696 24200
rect 18651 24160 18696 24188
rect 17405 24151 17463 24157
rect 17420 24120 17448 24151
rect 18690 24148 18696 24160
rect 18748 24148 18754 24200
rect 19613 24191 19671 24197
rect 19613 24157 19625 24191
rect 19659 24188 19671 24191
rect 20714 24188 20720 24200
rect 19659 24160 20720 24188
rect 19659 24157 19671 24160
rect 19613 24151 19671 24157
rect 20714 24148 20720 24160
rect 20772 24148 20778 24200
rect 21545 24191 21603 24197
rect 21545 24157 21557 24191
rect 21591 24157 21603 24191
rect 21545 24151 21603 24157
rect 18598 24120 18604 24132
rect 17144 24092 18604 24120
rect 18598 24080 18604 24092
rect 18656 24080 18662 24132
rect 21560 24120 21588 24151
rect 23290 24148 23296 24200
rect 23348 24188 23354 24200
rect 23937 24191 23995 24197
rect 23937 24188 23949 24191
rect 23348 24160 23949 24188
rect 23348 24148 23354 24160
rect 23937 24157 23949 24160
rect 23983 24157 23995 24191
rect 23937 24151 23995 24157
rect 22646 24120 22652 24132
rect 21560 24092 22652 24120
rect 22646 24080 22652 24092
rect 22704 24120 22710 24132
rect 22741 24123 22799 24129
rect 22741 24120 22753 24123
rect 22704 24092 22753 24120
rect 22704 24080 22710 24092
rect 22741 24089 22753 24092
rect 22787 24089 22799 24123
rect 22741 24083 22799 24089
rect 22830 24080 22836 24132
rect 22888 24120 22894 24132
rect 23385 24123 23443 24129
rect 23385 24120 23397 24123
rect 22888 24092 23397 24120
rect 22888 24080 22894 24092
rect 23385 24089 23397 24092
rect 23431 24089 23443 24123
rect 25130 24120 25136 24132
rect 25091 24092 25136 24120
rect 23385 24083 23443 24089
rect 25130 24080 25136 24092
rect 25188 24080 25194 24132
rect 2041 24055 2099 24061
rect 2041 24021 2053 24055
rect 2087 24052 2099 24055
rect 2317 24055 2375 24061
rect 2317 24052 2329 24055
rect 2087 24024 2329 24052
rect 2087 24021 2099 24024
rect 2041 24015 2099 24021
rect 2317 24021 2329 24024
rect 2363 24021 2375 24055
rect 5258 24052 5264 24064
rect 5219 24024 5264 24052
rect 2317 24015 2375 24021
rect 5258 24012 5264 24024
rect 5316 24012 5322 24064
rect 6270 24012 6276 24064
rect 6328 24052 6334 24064
rect 6733 24055 6791 24061
rect 6733 24052 6745 24055
rect 6328 24024 6745 24052
rect 6328 24012 6334 24024
rect 6733 24021 6745 24024
rect 6779 24021 6791 24055
rect 7190 24052 7196 24064
rect 7151 24024 7196 24052
rect 6733 24015 6791 24021
rect 7190 24012 7196 24024
rect 7248 24012 7254 24064
rect 9398 24052 9404 24064
rect 9359 24024 9404 24052
rect 9398 24012 9404 24024
rect 9456 24012 9462 24064
rect 9766 24012 9772 24064
rect 9824 24052 9830 24064
rect 9861 24055 9919 24061
rect 9861 24052 9873 24055
rect 9824 24024 9873 24052
rect 9824 24012 9830 24024
rect 9861 24021 9873 24024
rect 9907 24021 9919 24055
rect 11698 24052 11704 24064
rect 11659 24024 11704 24052
rect 9861 24015 9919 24021
rect 11698 24012 11704 24024
rect 11756 24012 11762 24064
rect 12802 24052 12808 24064
rect 12763 24024 12808 24052
rect 12802 24012 12808 24024
rect 12860 24012 12866 24064
rect 13170 24012 13176 24064
rect 13228 24052 13234 24064
rect 13265 24055 13323 24061
rect 13265 24052 13277 24055
rect 13228 24024 13277 24052
rect 13228 24012 13234 24024
rect 13265 24021 13277 24024
rect 13311 24021 13323 24055
rect 15286 24052 15292 24064
rect 15247 24024 15292 24052
rect 13265 24015 13323 24021
rect 15286 24012 15292 24024
rect 15344 24012 15350 24064
rect 16850 24052 16856 24064
rect 16811 24024 16856 24052
rect 16850 24012 16856 24024
rect 16908 24012 16914 24064
rect 18138 24052 18144 24064
rect 18099 24024 18144 24052
rect 18138 24012 18144 24024
rect 18196 24012 18202 24064
rect 20346 24052 20352 24064
rect 20307 24024 20352 24052
rect 20346 24012 20352 24024
rect 20404 24012 20410 24064
rect 20717 24055 20775 24061
rect 20717 24021 20729 24055
rect 20763 24052 20775 24055
rect 20898 24052 20904 24064
rect 20763 24024 20904 24052
rect 20763 24021 20775 24024
rect 20717 24015 20775 24021
rect 20898 24012 20904 24024
rect 20956 24012 20962 24064
rect 20993 24055 21051 24061
rect 20993 24021 21005 24055
rect 21039 24052 21051 24055
rect 21818 24052 21824 24064
rect 21039 24024 21824 24052
rect 21039 24021 21051 24024
rect 20993 24015 21051 24021
rect 21818 24012 21824 24024
rect 21876 24012 21882 24064
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1581 23851 1639 23857
rect 1581 23817 1593 23851
rect 1627 23848 1639 23851
rect 1670 23848 1676 23860
rect 1627 23820 1676 23848
rect 1627 23817 1639 23820
rect 1581 23811 1639 23817
rect 1670 23808 1676 23820
rect 1728 23808 1734 23860
rect 2314 23808 2320 23860
rect 2372 23848 2378 23860
rect 2685 23851 2743 23857
rect 2685 23848 2697 23851
rect 2372 23820 2697 23848
rect 2372 23808 2378 23820
rect 2685 23817 2697 23820
rect 2731 23817 2743 23851
rect 3510 23848 3516 23860
rect 3471 23820 3516 23848
rect 2685 23811 2743 23817
rect 3510 23808 3516 23820
rect 3568 23808 3574 23860
rect 6641 23851 6699 23857
rect 6641 23817 6653 23851
rect 6687 23848 6699 23851
rect 7374 23848 7380 23860
rect 6687 23820 7380 23848
rect 6687 23817 6699 23820
rect 6641 23811 6699 23817
rect 7374 23808 7380 23820
rect 7432 23808 7438 23860
rect 8389 23851 8447 23857
rect 8389 23817 8401 23851
rect 8435 23848 8447 23851
rect 9122 23848 9128 23860
rect 8435 23820 9128 23848
rect 8435 23817 8447 23820
rect 8389 23811 8447 23817
rect 9122 23808 9128 23820
rect 9180 23808 9186 23860
rect 9306 23848 9312 23860
rect 9267 23820 9312 23848
rect 9306 23808 9312 23820
rect 9364 23808 9370 23860
rect 9858 23808 9864 23860
rect 9916 23848 9922 23860
rect 11238 23848 11244 23860
rect 9916 23820 11244 23848
rect 9916 23808 9922 23820
rect 11238 23808 11244 23820
rect 11296 23808 11302 23860
rect 11425 23851 11483 23857
rect 11425 23817 11437 23851
rect 11471 23848 11483 23851
rect 11514 23848 11520 23860
rect 11471 23820 11520 23848
rect 11471 23817 11483 23820
rect 11425 23811 11483 23817
rect 11514 23808 11520 23820
rect 11572 23808 11578 23860
rect 15470 23848 15476 23860
rect 11900 23820 15476 23848
rect 4062 23740 4068 23792
rect 4120 23780 4126 23792
rect 5169 23783 5227 23789
rect 5169 23780 5181 23783
rect 4120 23752 5181 23780
rect 4120 23740 4126 23752
rect 5169 23749 5181 23752
rect 5215 23749 5227 23783
rect 5169 23743 5227 23749
rect 7285 23783 7343 23789
rect 7285 23749 7297 23783
rect 7331 23780 7343 23783
rect 7466 23780 7472 23792
rect 7331 23752 7472 23780
rect 7331 23749 7343 23752
rect 7285 23743 7343 23749
rect 7466 23740 7472 23752
rect 7524 23740 7530 23792
rect 8662 23740 8668 23792
rect 8720 23780 8726 23792
rect 11900 23780 11928 23820
rect 15470 23808 15476 23820
rect 15528 23848 15534 23860
rect 15565 23851 15623 23857
rect 15565 23848 15577 23851
rect 15528 23820 15577 23848
rect 15528 23808 15534 23820
rect 15565 23817 15577 23820
rect 15611 23817 15623 23851
rect 16022 23848 16028 23860
rect 15983 23820 16028 23848
rect 15565 23811 15623 23817
rect 8720 23752 11928 23780
rect 12437 23783 12495 23789
rect 8720 23740 8726 23752
rect 12437 23749 12449 23783
rect 12483 23780 12495 23783
rect 12710 23780 12716 23792
rect 12483 23752 12716 23780
rect 12483 23749 12495 23752
rect 12437 23743 12495 23749
rect 12710 23740 12716 23752
rect 12768 23740 12774 23792
rect 13446 23780 13452 23792
rect 13407 23752 13452 23780
rect 13446 23740 13452 23752
rect 13504 23740 13510 23792
rect 13630 23740 13636 23792
rect 13688 23780 13694 23792
rect 13817 23783 13875 23789
rect 13817 23780 13829 23783
rect 13688 23752 13829 23780
rect 13688 23740 13694 23752
rect 13817 23749 13829 23752
rect 13863 23780 13875 23783
rect 14274 23780 14280 23792
rect 13863 23752 14280 23780
rect 13863 23749 13875 23752
rect 13817 23743 13875 23749
rect 14274 23740 14280 23752
rect 14332 23740 14338 23792
rect 15580 23780 15608 23811
rect 16022 23808 16028 23820
rect 16080 23808 16086 23860
rect 16758 23808 16764 23860
rect 16816 23848 16822 23860
rect 18049 23851 18107 23857
rect 18049 23848 18061 23851
rect 16816 23820 18061 23848
rect 16816 23808 16822 23820
rect 18049 23817 18061 23820
rect 18095 23817 18107 23851
rect 18049 23811 18107 23817
rect 21269 23851 21327 23857
rect 21269 23817 21281 23851
rect 21315 23848 21327 23851
rect 21358 23848 21364 23860
rect 21315 23820 21364 23848
rect 21315 23817 21327 23820
rect 21269 23811 21327 23817
rect 21358 23808 21364 23820
rect 21416 23808 21422 23860
rect 24946 23848 24952 23860
rect 24907 23820 24952 23848
rect 24946 23808 24952 23820
rect 25004 23848 25010 23860
rect 26050 23848 26056 23860
rect 25004 23820 26056 23848
rect 25004 23808 25010 23820
rect 26050 23808 26056 23820
rect 26108 23808 26114 23860
rect 17129 23783 17187 23789
rect 17129 23780 17141 23783
rect 15580 23752 17141 23780
rect 17129 23749 17141 23752
rect 17175 23780 17187 23783
rect 17310 23780 17316 23792
rect 17175 23752 17316 23780
rect 17175 23749 17187 23752
rect 17129 23743 17187 23749
rect 17310 23740 17316 23752
rect 17368 23740 17374 23792
rect 20162 23780 20168 23792
rect 20123 23752 20168 23780
rect 20162 23740 20168 23752
rect 20220 23740 20226 23792
rect 21729 23783 21787 23789
rect 21729 23749 21741 23783
rect 21775 23780 21787 23783
rect 21775 23752 22416 23780
rect 21775 23749 21787 23752
rect 21729 23743 21787 23749
rect 1946 23672 1952 23724
rect 2004 23712 2010 23724
rect 2590 23712 2596 23724
rect 2004 23684 2596 23712
rect 2004 23672 2010 23684
rect 2590 23672 2596 23684
rect 2648 23712 2654 23724
rect 3053 23715 3111 23721
rect 3053 23712 3065 23715
rect 2648 23684 3065 23712
rect 2648 23672 2654 23684
rect 3053 23681 3065 23684
rect 3099 23681 3111 23715
rect 3053 23675 3111 23681
rect 4709 23715 4767 23721
rect 4709 23681 4721 23715
rect 4755 23712 4767 23715
rect 5813 23715 5871 23721
rect 5813 23712 5825 23715
rect 4755 23684 5825 23712
rect 4755 23681 4767 23684
rect 4709 23675 4767 23681
rect 5813 23681 5825 23684
rect 5859 23712 5871 23715
rect 6086 23712 6092 23724
rect 5859 23684 6092 23712
rect 5859 23681 5871 23684
rect 5813 23675 5871 23681
rect 6086 23672 6092 23684
rect 6144 23672 6150 23724
rect 8478 23672 8484 23724
rect 8536 23712 8542 23724
rect 8757 23715 8815 23721
rect 8757 23712 8769 23715
rect 8536 23684 8769 23712
rect 8536 23672 8542 23684
rect 8757 23681 8769 23684
rect 8803 23712 8815 23715
rect 8938 23712 8944 23724
rect 8803 23684 8944 23712
rect 8803 23681 8815 23684
rect 8757 23675 8815 23681
rect 8938 23672 8944 23684
rect 8996 23672 9002 23724
rect 9398 23672 9404 23724
rect 9456 23712 9462 23724
rect 9769 23715 9827 23721
rect 9769 23712 9781 23715
rect 9456 23684 9781 23712
rect 9456 23672 9462 23684
rect 9769 23681 9781 23684
rect 9815 23681 9827 23715
rect 9950 23712 9956 23724
rect 9911 23684 9956 23712
rect 9769 23675 9827 23681
rect 9950 23672 9956 23684
rect 10008 23672 10014 23724
rect 12894 23712 12900 23724
rect 12855 23684 12900 23712
rect 12894 23672 12900 23684
rect 12952 23672 12958 23724
rect 13081 23715 13139 23721
rect 13081 23681 13093 23715
rect 13127 23712 13139 23715
rect 13354 23712 13360 23724
rect 13127 23684 13360 23712
rect 13127 23681 13139 23684
rect 13081 23675 13139 23681
rect 13354 23672 13360 23684
rect 13412 23672 13418 23724
rect 15197 23715 15255 23721
rect 15197 23681 15209 23715
rect 15243 23681 15255 23715
rect 15197 23675 15255 23681
rect 1397 23647 1455 23653
rect 1397 23613 1409 23647
rect 1443 23644 1455 23647
rect 1670 23644 1676 23656
rect 1443 23616 1676 23644
rect 1443 23613 1455 23616
rect 1397 23607 1455 23613
rect 1670 23604 1676 23616
rect 1728 23604 1734 23656
rect 2501 23647 2559 23653
rect 2501 23644 2513 23647
rect 2332 23616 2513 23644
rect 2041 23511 2099 23517
rect 2041 23477 2053 23511
rect 2087 23508 2099 23511
rect 2130 23508 2136 23520
rect 2087 23480 2136 23508
rect 2087 23477 2099 23480
rect 2041 23471 2099 23477
rect 2130 23468 2136 23480
rect 2188 23468 2194 23520
rect 2222 23468 2228 23520
rect 2280 23508 2286 23520
rect 2332 23517 2360 23616
rect 2501 23613 2513 23616
rect 2547 23613 2559 23647
rect 2501 23607 2559 23613
rect 2682 23604 2688 23656
rect 2740 23644 2746 23656
rect 3605 23647 3663 23653
rect 3605 23644 3617 23647
rect 2740 23616 3617 23644
rect 2740 23604 2746 23616
rect 3605 23613 3617 23616
rect 3651 23644 3663 23647
rect 4157 23647 4215 23653
rect 4157 23644 4169 23647
rect 3651 23616 4169 23644
rect 3651 23613 3663 23616
rect 3605 23607 3663 23613
rect 4157 23613 4169 23616
rect 4203 23613 4215 23647
rect 4157 23607 4215 23613
rect 5534 23604 5540 23656
rect 5592 23644 5598 23656
rect 6178 23644 6184 23656
rect 5592 23616 6184 23644
rect 5592 23604 5598 23616
rect 6178 23604 6184 23616
rect 6236 23604 6242 23656
rect 7101 23647 7159 23653
rect 7101 23613 7113 23647
rect 7147 23644 7159 23647
rect 7190 23644 7196 23656
rect 7147 23616 7196 23644
rect 7147 23613 7159 23616
rect 7101 23607 7159 23613
rect 7190 23604 7196 23616
rect 7248 23604 7254 23656
rect 8205 23647 8263 23653
rect 8205 23613 8217 23647
rect 8251 23644 8263 23647
rect 8294 23644 8300 23656
rect 8251 23616 8300 23644
rect 8251 23613 8263 23616
rect 8205 23607 8263 23613
rect 8294 23604 8300 23616
rect 8352 23604 8358 23656
rect 9217 23647 9275 23653
rect 9217 23613 9229 23647
rect 9263 23644 9275 23647
rect 9968 23644 9996 23672
rect 9263 23616 9996 23644
rect 9263 23613 9275 23616
rect 9217 23607 9275 23613
rect 10502 23604 10508 23656
rect 10560 23644 10566 23656
rect 10689 23647 10747 23653
rect 10689 23644 10701 23647
rect 10560 23616 10701 23644
rect 10560 23604 10566 23616
rect 10689 23613 10701 23616
rect 10735 23644 10747 23647
rect 11054 23644 11060 23656
rect 10735 23616 11060 23644
rect 10735 23613 10747 23616
rect 10689 23607 10747 23613
rect 11054 23604 11060 23616
rect 11112 23604 11118 23656
rect 11238 23644 11244 23656
rect 11199 23616 11244 23644
rect 11238 23604 11244 23616
rect 11296 23644 11302 23656
rect 11793 23647 11851 23653
rect 11793 23644 11805 23647
rect 11296 23616 11805 23644
rect 11296 23604 11302 23616
rect 11793 23613 11805 23616
rect 11839 23644 11851 23647
rect 12434 23644 12440 23656
rect 11839 23616 12440 23644
rect 11839 23613 11851 23616
rect 11793 23607 11851 23613
rect 12434 23604 12440 23616
rect 12492 23604 12498 23656
rect 5258 23536 5264 23588
rect 5316 23576 5322 23588
rect 10413 23579 10471 23585
rect 5316 23548 5672 23576
rect 5316 23536 5322 23548
rect 2317 23511 2375 23517
rect 2317 23508 2329 23511
rect 2280 23480 2329 23508
rect 2280 23468 2286 23480
rect 2317 23477 2329 23480
rect 2363 23477 2375 23511
rect 2317 23471 2375 23477
rect 3510 23468 3516 23520
rect 3568 23508 3574 23520
rect 3789 23511 3847 23517
rect 3789 23508 3801 23511
rect 3568 23480 3801 23508
rect 3568 23468 3574 23480
rect 3789 23477 3801 23480
rect 3835 23477 3847 23511
rect 3789 23471 3847 23477
rect 4614 23468 4620 23520
rect 4672 23508 4678 23520
rect 4985 23511 5043 23517
rect 4985 23508 4997 23511
rect 4672 23480 4997 23508
rect 4672 23468 4678 23480
rect 4985 23477 4997 23480
rect 5031 23508 5043 23511
rect 5442 23508 5448 23520
rect 5031 23480 5448 23508
rect 5031 23477 5043 23480
rect 4985 23471 5043 23477
rect 5442 23468 5448 23480
rect 5500 23508 5506 23520
rect 5644 23517 5672 23548
rect 10413 23545 10425 23579
rect 10459 23576 10471 23579
rect 10778 23576 10784 23588
rect 10459 23548 10784 23576
rect 10459 23545 10471 23548
rect 10413 23539 10471 23545
rect 10778 23536 10784 23548
rect 10836 23536 10842 23588
rect 11514 23536 11520 23588
rect 11572 23576 11578 23588
rect 12161 23579 12219 23585
rect 12161 23576 12173 23579
rect 11572 23548 12173 23576
rect 11572 23536 11578 23548
rect 12161 23545 12173 23548
rect 12207 23576 12219 23579
rect 12912 23576 12940 23672
rect 14550 23604 14556 23656
rect 14608 23644 14614 23656
rect 14921 23647 14979 23653
rect 14921 23644 14933 23647
rect 14608 23616 14933 23644
rect 14608 23604 14614 23616
rect 14921 23613 14933 23616
rect 14967 23613 14979 23647
rect 15212 23644 15240 23675
rect 16114 23672 16120 23724
rect 16172 23712 16178 23724
rect 16482 23712 16488 23724
rect 16172 23684 16488 23712
rect 16172 23672 16178 23684
rect 16482 23672 16488 23684
rect 16540 23712 16546 23724
rect 16577 23715 16635 23721
rect 16577 23712 16589 23715
rect 16540 23684 16589 23712
rect 16540 23672 16546 23684
rect 16577 23681 16589 23684
rect 16623 23681 16635 23715
rect 16577 23675 16635 23681
rect 16669 23715 16727 23721
rect 16669 23681 16681 23715
rect 16715 23681 16727 23715
rect 18598 23712 18604 23724
rect 18559 23684 18604 23712
rect 16669 23675 16727 23681
rect 16206 23644 16212 23656
rect 15212 23616 16212 23644
rect 14921 23607 14979 23613
rect 16206 23604 16212 23616
rect 16264 23644 16270 23656
rect 16684 23644 16712 23675
rect 18598 23672 18604 23684
rect 18656 23712 18662 23724
rect 18966 23712 18972 23724
rect 18656 23684 18972 23712
rect 18656 23672 18662 23684
rect 18966 23672 18972 23684
rect 19024 23712 19030 23724
rect 19061 23715 19119 23721
rect 19061 23712 19073 23715
rect 19024 23684 19073 23712
rect 19024 23672 19030 23684
rect 19061 23681 19073 23684
rect 19107 23681 19119 23715
rect 20717 23715 20775 23721
rect 20717 23712 20729 23715
rect 19061 23675 19119 23681
rect 20088 23684 20729 23712
rect 16264 23616 16712 23644
rect 16264 23604 16270 23616
rect 20088 23588 20116 23684
rect 20717 23681 20729 23684
rect 20763 23681 20775 23715
rect 22278 23712 22284 23724
rect 22239 23684 22284 23712
rect 20717 23675 20775 23681
rect 22278 23672 22284 23684
rect 22336 23672 22342 23724
rect 20898 23604 20904 23656
rect 20956 23644 20962 23656
rect 22388 23644 22416 23752
rect 23477 23715 23535 23721
rect 23477 23681 23489 23715
rect 23523 23712 23535 23715
rect 24302 23712 24308 23724
rect 23523 23684 24308 23712
rect 23523 23681 23535 23684
rect 23477 23675 23535 23681
rect 24302 23672 24308 23684
rect 24360 23672 24366 23724
rect 24121 23647 24179 23653
rect 24121 23644 24133 23647
rect 20956 23616 21680 23644
rect 22388 23616 24133 23644
rect 20956 23604 20962 23616
rect 15013 23579 15071 23585
rect 15013 23576 15025 23579
rect 12207 23548 12940 23576
rect 14384 23548 15025 23576
rect 12207 23545 12219 23548
rect 12161 23539 12219 23545
rect 5537 23511 5595 23517
rect 5537 23508 5549 23511
rect 5500 23480 5549 23508
rect 5500 23468 5506 23480
rect 5537 23477 5549 23480
rect 5583 23477 5595 23511
rect 5537 23471 5595 23477
rect 5629 23511 5687 23517
rect 5629 23477 5641 23511
rect 5675 23508 5687 23511
rect 6362 23508 6368 23520
rect 5675 23480 6368 23508
rect 5675 23477 5687 23480
rect 5629 23471 5687 23477
rect 6362 23468 6368 23480
rect 6420 23468 6426 23520
rect 7837 23511 7895 23517
rect 7837 23477 7849 23511
rect 7883 23508 7895 23511
rect 8294 23508 8300 23520
rect 7883 23480 8300 23508
rect 7883 23477 7895 23480
rect 7837 23471 7895 23477
rect 8294 23468 8300 23480
rect 8352 23468 8358 23520
rect 9674 23508 9680 23520
rect 9635 23480 9680 23508
rect 9674 23468 9680 23480
rect 9732 23468 9738 23520
rect 11054 23508 11060 23520
rect 11015 23480 11060 23508
rect 11054 23468 11060 23480
rect 11112 23468 11118 23520
rect 12802 23508 12808 23520
rect 12763 23480 12808 23508
rect 12802 23468 12808 23480
rect 12860 23468 12866 23520
rect 13906 23468 13912 23520
rect 13964 23508 13970 23520
rect 14384 23517 14412 23548
rect 15013 23545 15025 23548
rect 15059 23545 15071 23579
rect 15013 23539 15071 23545
rect 16485 23579 16543 23585
rect 16485 23545 16497 23579
rect 16531 23576 16543 23579
rect 17770 23576 17776 23588
rect 16531 23548 17776 23576
rect 16531 23545 16543 23548
rect 16485 23539 16543 23545
rect 17770 23536 17776 23548
rect 17828 23536 17834 23588
rect 18138 23536 18144 23588
rect 18196 23576 18202 23588
rect 18509 23579 18567 23585
rect 18509 23576 18521 23579
rect 18196 23548 18521 23576
rect 18196 23536 18202 23548
rect 18509 23545 18521 23548
rect 18555 23576 18567 23579
rect 19150 23576 19156 23588
rect 18555 23548 19156 23576
rect 18555 23545 18567 23548
rect 18509 23539 18567 23545
rect 19150 23536 19156 23548
rect 19208 23536 19214 23588
rect 19705 23579 19763 23585
rect 19705 23545 19717 23579
rect 19751 23576 19763 23579
rect 20070 23576 20076 23588
rect 19751 23548 20076 23576
rect 19751 23545 19763 23548
rect 19705 23539 19763 23545
rect 20070 23536 20076 23548
rect 20128 23536 20134 23588
rect 20625 23579 20683 23585
rect 20625 23576 20637 23579
rect 20180 23548 20637 23576
rect 14369 23511 14427 23517
rect 14369 23508 14381 23511
rect 13964 23480 14381 23508
rect 13964 23468 13970 23480
rect 14369 23477 14381 23480
rect 14415 23477 14427 23511
rect 14369 23471 14427 23477
rect 14553 23511 14611 23517
rect 14553 23477 14565 23511
rect 14599 23508 14611 23511
rect 15102 23508 15108 23520
rect 14599 23480 15108 23508
rect 14599 23477 14611 23480
rect 14553 23471 14611 23477
rect 15102 23468 15108 23480
rect 15160 23468 15166 23520
rect 16117 23511 16175 23517
rect 16117 23477 16129 23511
rect 16163 23508 16175 23511
rect 16390 23508 16396 23520
rect 16163 23480 16396 23508
rect 16163 23477 16175 23480
rect 16117 23471 16175 23477
rect 16390 23468 16396 23480
rect 16448 23468 16454 23520
rect 17494 23508 17500 23520
rect 17455 23480 17500 23508
rect 17494 23468 17500 23480
rect 17552 23468 17558 23520
rect 18046 23468 18052 23520
rect 18104 23508 18110 23520
rect 18417 23511 18475 23517
rect 18417 23508 18429 23511
rect 18104 23480 18429 23508
rect 18104 23468 18110 23480
rect 18417 23477 18429 23480
rect 18463 23508 18475 23511
rect 18782 23508 18788 23520
rect 18463 23480 18788 23508
rect 18463 23477 18475 23480
rect 18417 23471 18475 23477
rect 18782 23468 18788 23480
rect 18840 23468 18846 23520
rect 19426 23468 19432 23520
rect 19484 23508 19490 23520
rect 19981 23511 20039 23517
rect 19981 23508 19993 23511
rect 19484 23480 19993 23508
rect 19484 23468 19490 23480
rect 19981 23477 19993 23480
rect 20027 23508 20039 23511
rect 20180 23508 20208 23548
rect 20625 23545 20637 23548
rect 20671 23545 20683 23579
rect 20625 23539 20683 23545
rect 21266 23536 21272 23588
rect 21324 23576 21330 23588
rect 21545 23579 21603 23585
rect 21545 23576 21557 23579
rect 21324 23548 21557 23576
rect 21324 23536 21330 23548
rect 21545 23545 21557 23548
rect 21591 23545 21603 23579
rect 21652 23576 21680 23616
rect 24121 23613 24133 23616
rect 24167 23644 24179 23647
rect 24854 23644 24860 23656
rect 24167 23616 24860 23644
rect 24167 23613 24179 23616
rect 24121 23607 24179 23613
rect 24854 23604 24860 23616
rect 24912 23604 24918 23656
rect 25222 23644 25228 23656
rect 25183 23616 25228 23644
rect 25222 23604 25228 23616
rect 25280 23644 25286 23656
rect 25777 23647 25835 23653
rect 25777 23644 25789 23647
rect 25280 23616 25789 23644
rect 25280 23604 25286 23616
rect 25777 23613 25789 23616
rect 25823 23613 25835 23647
rect 25777 23607 25835 23613
rect 22189 23579 22247 23585
rect 22189 23576 22201 23579
rect 21652 23548 22201 23576
rect 21545 23539 21603 23545
rect 22189 23545 22201 23548
rect 22235 23545 22247 23579
rect 22189 23539 22247 23545
rect 23474 23536 23480 23588
rect 23532 23576 23538 23588
rect 24029 23579 24087 23585
rect 24029 23576 24041 23579
rect 23532 23548 24041 23576
rect 23532 23536 23538 23548
rect 24029 23545 24041 23548
rect 24075 23576 24087 23579
rect 26237 23579 26295 23585
rect 26237 23576 26249 23579
rect 24075 23548 26249 23576
rect 24075 23545 24087 23548
rect 24029 23539 24087 23545
rect 26237 23545 26249 23548
rect 26283 23545 26295 23579
rect 26237 23539 26295 23545
rect 20027 23480 20208 23508
rect 20027 23477 20039 23480
rect 19981 23471 20039 23477
rect 20254 23468 20260 23520
rect 20312 23508 20318 23520
rect 20533 23511 20591 23517
rect 20533 23508 20545 23511
rect 20312 23480 20545 23508
rect 20312 23468 20318 23480
rect 20533 23477 20545 23480
rect 20579 23477 20591 23511
rect 20533 23471 20591 23477
rect 22094 23468 22100 23520
rect 22152 23508 22158 23520
rect 22738 23508 22744 23520
rect 22152 23480 22197 23508
rect 22699 23480 22744 23508
rect 22152 23468 22158 23480
rect 22738 23468 22744 23480
rect 22796 23468 22802 23520
rect 23658 23508 23664 23520
rect 23619 23480 23664 23508
rect 23658 23468 23664 23480
rect 23716 23468 23722 23520
rect 25406 23508 25412 23520
rect 25367 23480 25412 23508
rect 25406 23468 25412 23480
rect 25464 23468 25470 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 3697 23307 3755 23313
rect 3697 23273 3709 23307
rect 3743 23304 3755 23307
rect 4062 23304 4068 23316
rect 3743 23276 4068 23304
rect 3743 23273 3755 23276
rect 3697 23267 3755 23273
rect 4062 23264 4068 23276
rect 4120 23264 4126 23316
rect 5902 23264 5908 23316
rect 5960 23304 5966 23316
rect 6546 23304 6552 23316
rect 5960 23276 6552 23304
rect 5960 23264 5966 23276
rect 6546 23264 6552 23276
rect 6604 23264 6610 23316
rect 11054 23304 11060 23316
rect 11015 23276 11060 23304
rect 11054 23264 11060 23276
rect 11112 23264 11118 23316
rect 12158 23264 12164 23316
rect 12216 23304 12222 23316
rect 12253 23307 12311 23313
rect 12253 23304 12265 23307
rect 12216 23276 12265 23304
rect 12216 23264 12222 23276
rect 12253 23273 12265 23276
rect 12299 23273 12311 23307
rect 13630 23304 13636 23316
rect 13591 23276 13636 23304
rect 12253 23267 12311 23273
rect 13630 23264 13636 23276
rect 13688 23264 13694 23316
rect 16758 23264 16764 23316
rect 16816 23304 16822 23316
rect 16853 23307 16911 23313
rect 16853 23304 16865 23307
rect 16816 23276 16865 23304
rect 16816 23264 16822 23276
rect 16853 23273 16865 23276
rect 16899 23273 16911 23307
rect 16853 23267 16911 23273
rect 16942 23264 16948 23316
rect 17000 23304 17006 23316
rect 17218 23304 17224 23316
rect 17000 23276 17224 23304
rect 17000 23264 17006 23276
rect 17218 23264 17224 23276
rect 17276 23264 17282 23316
rect 18046 23304 18052 23316
rect 18007 23276 18052 23304
rect 18046 23264 18052 23276
rect 18104 23264 18110 23316
rect 18414 23304 18420 23316
rect 18375 23276 18420 23304
rect 18414 23264 18420 23276
rect 18472 23264 18478 23316
rect 20714 23264 20720 23316
rect 20772 23304 20778 23316
rect 21085 23307 21143 23313
rect 21085 23304 21097 23307
rect 20772 23276 21097 23304
rect 20772 23264 20778 23276
rect 21085 23273 21097 23276
rect 21131 23304 21143 23307
rect 22002 23304 22008 23316
rect 21131 23276 22008 23304
rect 21131 23273 21143 23276
rect 21085 23267 21143 23273
rect 22002 23264 22008 23276
rect 22060 23264 22066 23316
rect 23290 23304 23296 23316
rect 23251 23276 23296 23304
rect 23290 23264 23296 23276
rect 23348 23264 23354 23316
rect 23474 23304 23480 23316
rect 23435 23276 23480 23304
rect 23474 23264 23480 23276
rect 23532 23264 23538 23316
rect 24854 23304 24860 23316
rect 24815 23276 24860 23304
rect 24854 23264 24860 23276
rect 24912 23264 24918 23316
rect 1670 23236 1676 23248
rect 1631 23208 1676 23236
rect 1670 23196 1676 23208
rect 1728 23196 1734 23248
rect 2406 23196 2412 23248
rect 2464 23236 2470 23248
rect 2501 23239 2559 23245
rect 2501 23236 2513 23239
rect 2464 23208 2513 23236
rect 2464 23196 2470 23208
rect 2501 23205 2513 23208
rect 2547 23205 2559 23239
rect 2501 23199 2559 23205
rect 5169 23239 5227 23245
rect 5169 23205 5181 23239
rect 5215 23236 5227 23239
rect 5534 23236 5540 23248
rect 5215 23208 5540 23236
rect 5215 23205 5227 23208
rect 5169 23199 5227 23205
rect 5534 23196 5540 23208
rect 5592 23196 5598 23248
rect 6178 23196 6184 23248
rect 6236 23236 6242 23248
rect 6641 23239 6699 23245
rect 6641 23236 6653 23239
rect 6236 23208 6653 23236
rect 6236 23196 6242 23208
rect 6641 23205 6653 23208
rect 6687 23205 6699 23239
rect 6641 23199 6699 23205
rect 11790 23196 11796 23248
rect 11848 23236 11854 23248
rect 12066 23236 12072 23248
rect 11848 23208 12072 23236
rect 11848 23196 11854 23208
rect 12066 23196 12072 23208
rect 12124 23196 12130 23248
rect 13357 23239 13415 23245
rect 13357 23205 13369 23239
rect 13403 23236 13415 23239
rect 13538 23236 13544 23248
rect 13403 23208 13544 23236
rect 13403 23205 13415 23208
rect 13357 23199 13415 23205
rect 13538 23196 13544 23208
rect 13596 23196 13602 23248
rect 14090 23236 14096 23248
rect 14051 23208 14096 23236
rect 14090 23196 14096 23208
rect 14148 23196 14154 23248
rect 15930 23236 15936 23248
rect 15396 23208 15936 23236
rect 2225 23171 2283 23177
rect 2225 23137 2237 23171
rect 2271 23137 2283 23171
rect 4890 23168 4896 23180
rect 4851 23140 4896 23168
rect 2225 23131 2283 23137
rect 2240 23100 2268 23131
rect 4890 23128 4896 23140
rect 4948 23128 4954 23180
rect 7098 23128 7104 23180
rect 7156 23168 7162 23180
rect 8110 23168 8116 23180
rect 7156 23140 8116 23168
rect 7156 23128 7162 23140
rect 8110 23128 8116 23140
rect 8168 23128 8174 23180
rect 10597 23171 10655 23177
rect 10597 23137 10609 23171
rect 10643 23168 10655 23171
rect 10643 23140 11376 23168
rect 10643 23137 10655 23140
rect 10597 23131 10655 23137
rect 2406 23100 2412 23112
rect 2240 23072 2412 23100
rect 2406 23060 2412 23072
rect 2464 23060 2470 23112
rect 6825 23103 6883 23109
rect 6825 23069 6837 23103
rect 6871 23100 6883 23103
rect 7006 23100 7012 23112
rect 6871 23072 7012 23100
rect 6871 23069 6883 23072
rect 6825 23063 6883 23069
rect 7006 23060 7012 23072
rect 7064 23060 7070 23112
rect 8018 23060 8024 23112
rect 8076 23100 8082 23112
rect 8205 23103 8263 23109
rect 8205 23100 8217 23103
rect 8076 23072 8217 23100
rect 8076 23060 8082 23072
rect 8205 23069 8217 23072
rect 8251 23069 8263 23103
rect 8205 23063 8263 23069
rect 8294 23060 8300 23112
rect 8352 23100 8358 23112
rect 11146 23100 11152 23112
rect 8352 23072 8397 23100
rect 11107 23072 11152 23100
rect 8352 23060 8358 23072
rect 11146 23060 11152 23072
rect 11204 23060 11210 23112
rect 11348 23109 11376 23140
rect 12434 23128 12440 23180
rect 12492 23168 12498 23180
rect 12621 23171 12679 23177
rect 12621 23168 12633 23171
rect 12492 23140 12633 23168
rect 12492 23128 12498 23140
rect 12621 23137 12633 23140
rect 12667 23137 12679 23171
rect 12621 23131 12679 23137
rect 13817 23171 13875 23177
rect 13817 23137 13829 23171
rect 13863 23168 13875 23171
rect 14182 23168 14188 23180
rect 13863 23140 14188 23168
rect 13863 23137 13875 23140
rect 13817 23131 13875 23137
rect 14182 23128 14188 23140
rect 14240 23128 14246 23180
rect 11333 23103 11391 23109
rect 11333 23069 11345 23103
rect 11379 23100 11391 23103
rect 12066 23100 12072 23112
rect 11379 23072 12072 23100
rect 11379 23069 11391 23072
rect 11333 23063 11391 23069
rect 12066 23060 12072 23072
rect 12124 23060 12130 23112
rect 12710 23100 12716 23112
rect 12671 23072 12716 23100
rect 12710 23060 12716 23072
rect 12768 23060 12774 23112
rect 12897 23103 12955 23109
rect 12897 23069 12909 23103
rect 12943 23100 12955 23103
rect 13354 23100 13360 23112
rect 12943 23072 13360 23100
rect 12943 23069 12955 23072
rect 12897 23063 12955 23069
rect 13354 23060 13360 23072
rect 13412 23060 13418 23112
rect 13630 23060 13636 23112
rect 13688 23100 13694 23112
rect 15396 23100 15424 23208
rect 15930 23196 15936 23208
rect 15988 23196 15994 23248
rect 17236 23236 17264 23264
rect 18877 23239 18935 23245
rect 18877 23236 18889 23239
rect 17236 23208 18889 23236
rect 18877 23205 18889 23208
rect 18923 23236 18935 23239
rect 19058 23236 19064 23248
rect 18923 23208 19064 23236
rect 18923 23205 18935 23208
rect 18877 23199 18935 23205
rect 19058 23196 19064 23208
rect 19116 23196 19122 23248
rect 15562 23128 15568 23180
rect 15620 23168 15626 23180
rect 15657 23171 15715 23177
rect 15657 23168 15669 23171
rect 15620 23140 15669 23168
rect 15620 23128 15626 23140
rect 15657 23137 15669 23140
rect 15703 23137 15715 23171
rect 15657 23131 15715 23137
rect 17770 23128 17776 23180
rect 17828 23168 17834 23180
rect 18785 23171 18843 23177
rect 18785 23168 18797 23171
rect 17828 23140 18797 23168
rect 17828 23128 17834 23140
rect 18785 23137 18797 23140
rect 18831 23137 18843 23171
rect 18785 23131 18843 23137
rect 21358 23128 21364 23180
rect 21416 23168 21422 23180
rect 21453 23171 21511 23177
rect 21453 23168 21465 23171
rect 21416 23140 21465 23168
rect 21416 23128 21422 23140
rect 21453 23137 21465 23140
rect 21499 23137 21511 23171
rect 23308 23168 23336 23264
rect 23845 23239 23903 23245
rect 23845 23205 23857 23239
rect 23891 23236 23903 23239
rect 24026 23236 24032 23248
rect 23891 23208 24032 23236
rect 23891 23205 23903 23208
rect 23845 23199 23903 23205
rect 24026 23196 24032 23208
rect 24084 23196 24090 23248
rect 25314 23236 25320 23248
rect 25275 23208 25320 23236
rect 25314 23196 25320 23208
rect 25372 23196 25378 23248
rect 25038 23168 25044 23180
rect 23308 23140 24808 23168
rect 24999 23140 25044 23168
rect 21453 23131 21511 23137
rect 13688 23072 15424 23100
rect 13688 23060 13694 23072
rect 15470 23060 15476 23112
rect 15528 23100 15534 23112
rect 15749 23103 15807 23109
rect 15749 23100 15761 23103
rect 15528 23072 15761 23100
rect 15528 23060 15534 23072
rect 15749 23069 15761 23072
rect 15795 23069 15807 23103
rect 15930 23100 15936 23112
rect 15891 23072 15936 23100
rect 15749 23063 15807 23069
rect 15930 23060 15936 23072
rect 15988 23060 15994 23112
rect 16574 23060 16580 23112
rect 16632 23100 16638 23112
rect 17313 23103 17371 23109
rect 17313 23100 17325 23103
rect 16632 23072 17325 23100
rect 16632 23060 16638 23072
rect 17313 23069 17325 23072
rect 17359 23069 17371 23103
rect 17313 23063 17371 23069
rect 17405 23103 17463 23109
rect 17405 23069 17417 23103
rect 17451 23069 17463 23103
rect 17405 23063 17463 23069
rect 5534 22992 5540 23044
rect 5592 23032 5598 23044
rect 5721 23035 5779 23041
rect 5721 23032 5733 23035
rect 5592 23004 5733 23032
rect 5592 22992 5598 23004
rect 5721 23001 5733 23004
rect 5767 23032 5779 23035
rect 6181 23035 6239 23041
rect 6181 23032 6193 23035
rect 5767 23004 6193 23032
rect 5767 23001 5779 23004
rect 5721 22995 5779 23001
rect 6181 23001 6193 23004
rect 6227 23001 6239 23035
rect 6181 22995 6239 23001
rect 6730 22992 6736 23044
rect 6788 23032 6794 23044
rect 7745 23035 7803 23041
rect 7745 23032 7757 23035
rect 6788 23004 7757 23032
rect 6788 22992 6794 23004
rect 7745 23001 7757 23004
rect 7791 23001 7803 23035
rect 9309 23035 9367 23041
rect 9309 23032 9321 23035
rect 7745 22995 7803 23001
rect 8956 23004 9321 23032
rect 2038 22964 2044 22976
rect 1999 22936 2044 22964
rect 2038 22924 2044 22936
rect 2096 22924 2102 22976
rect 2590 22924 2596 22976
rect 2648 22964 2654 22976
rect 2961 22967 3019 22973
rect 2961 22964 2973 22967
rect 2648 22936 2973 22964
rect 2648 22924 2654 22936
rect 2961 22933 2973 22936
rect 3007 22933 3019 22967
rect 4338 22964 4344 22976
rect 4299 22936 4344 22964
rect 2961 22927 3019 22933
rect 4338 22924 4344 22936
rect 4396 22924 4402 22976
rect 4798 22964 4804 22976
rect 4759 22936 4804 22964
rect 4798 22924 4804 22936
rect 4856 22924 4862 22976
rect 6089 22967 6147 22973
rect 6089 22933 6101 22967
rect 6135 22964 6147 22967
rect 6270 22964 6276 22976
rect 6135 22936 6276 22964
rect 6135 22933 6147 22936
rect 6089 22927 6147 22933
rect 6270 22924 6276 22936
rect 6328 22924 6334 22976
rect 7466 22964 7472 22976
rect 7427 22936 7472 22964
rect 7466 22924 7472 22936
rect 7524 22924 7530 22976
rect 8294 22924 8300 22976
rect 8352 22964 8358 22976
rect 8956 22964 8984 23004
rect 9309 23001 9321 23004
rect 9355 23032 9367 23035
rect 9674 23032 9680 23044
rect 9355 23004 9680 23032
rect 9355 23001 9367 23004
rect 9309 22995 9367 23001
rect 9674 22992 9680 23004
rect 9732 22992 9738 23044
rect 10229 23035 10287 23041
rect 10229 23001 10241 23035
rect 10275 23032 10287 23035
rect 10870 23032 10876 23044
rect 10275 23004 10876 23032
rect 10275 23001 10287 23004
rect 10229 22995 10287 23001
rect 10870 22992 10876 23004
rect 10928 22992 10934 23044
rect 14734 22992 14740 23044
rect 14792 23032 14798 23044
rect 15289 23035 15347 23041
rect 15289 23032 15301 23035
rect 14792 23004 15301 23032
rect 14792 22992 14798 23004
rect 15289 23001 15301 23004
rect 15335 23001 15347 23035
rect 15289 22995 15347 23001
rect 16942 22992 16948 23044
rect 17000 23032 17006 23044
rect 17420 23032 17448 23063
rect 18966 23060 18972 23112
rect 19024 23100 19030 23112
rect 19429 23103 19487 23109
rect 19429 23100 19441 23103
rect 19024 23072 19441 23100
rect 19024 23060 19030 23072
rect 19429 23069 19441 23072
rect 19475 23100 19487 23103
rect 19794 23100 19800 23112
rect 19475 23072 19800 23100
rect 19475 23069 19487 23072
rect 19429 23063 19487 23069
rect 19794 23060 19800 23072
rect 19852 23060 19858 23112
rect 21545 23103 21603 23109
rect 21545 23069 21557 23103
rect 21591 23069 21603 23103
rect 21545 23063 21603 23069
rect 21729 23103 21787 23109
rect 21729 23069 21741 23103
rect 21775 23100 21787 23103
rect 22094 23100 22100 23112
rect 21775 23072 22100 23100
rect 21775 23069 21787 23072
rect 21729 23063 21787 23069
rect 17000 23004 17448 23032
rect 17000 22992 17006 23004
rect 17678 22992 17684 23044
rect 17736 23032 17742 23044
rect 18984 23032 19012 23060
rect 17736 23004 19012 23032
rect 21560 23032 21588 23063
rect 22094 23060 22100 23072
rect 22152 23060 22158 23112
rect 22189 23103 22247 23109
rect 22189 23069 22201 23103
rect 22235 23100 22247 23103
rect 22278 23100 22284 23112
rect 22235 23072 22284 23100
rect 22235 23069 22247 23072
rect 22189 23063 22247 23069
rect 22278 23060 22284 23072
rect 22336 23100 22342 23112
rect 23934 23100 23940 23112
rect 22336 23072 23244 23100
rect 23895 23072 23940 23100
rect 22336 23060 22342 23072
rect 23216 23044 23244 23072
rect 23934 23060 23940 23072
rect 23992 23060 23998 23112
rect 24029 23103 24087 23109
rect 24029 23069 24041 23103
rect 24075 23069 24087 23103
rect 24780 23100 24808 23140
rect 25038 23128 25044 23140
rect 25096 23128 25102 23180
rect 25314 23100 25320 23112
rect 24780 23072 25320 23100
rect 24029 23063 24087 23069
rect 22462 23032 22468 23044
rect 21560 23004 22468 23032
rect 17736 22992 17742 23004
rect 22462 22992 22468 23004
rect 22520 22992 22526 23044
rect 23198 22992 23204 23044
rect 23256 23032 23262 23044
rect 24044 23032 24072 23063
rect 25314 23060 25320 23072
rect 25372 23060 25378 23112
rect 23256 23004 24072 23032
rect 23256 22992 23262 23004
rect 8352 22936 8984 22964
rect 9033 22967 9091 22973
rect 8352 22924 8358 22936
rect 9033 22933 9045 22967
rect 9079 22964 9091 22967
rect 9122 22964 9128 22976
rect 9079 22936 9128 22964
rect 9079 22933 9091 22936
rect 9033 22927 9091 22933
rect 9122 22924 9128 22936
rect 9180 22924 9186 22976
rect 10686 22964 10692 22976
rect 10647 22936 10692 22964
rect 10686 22924 10692 22936
rect 10744 22924 10750 22976
rect 11790 22964 11796 22976
rect 11751 22936 11796 22964
rect 11790 22924 11796 22936
rect 11848 22924 11854 22976
rect 12158 22964 12164 22976
rect 12119 22936 12164 22964
rect 12158 22924 12164 22936
rect 12216 22924 12222 22976
rect 14550 22964 14556 22976
rect 14511 22936 14556 22964
rect 14550 22924 14556 22936
rect 14608 22924 14614 22976
rect 15013 22967 15071 22973
rect 15013 22933 15025 22967
rect 15059 22964 15071 22967
rect 16206 22964 16212 22976
rect 15059 22936 16212 22964
rect 15059 22933 15071 22936
rect 15013 22927 15071 22933
rect 16206 22924 16212 22936
rect 16264 22964 16270 22976
rect 16301 22967 16359 22973
rect 16301 22964 16313 22967
rect 16264 22936 16313 22964
rect 16264 22924 16270 22936
rect 16301 22933 16313 22936
rect 16347 22933 16359 22967
rect 16758 22964 16764 22976
rect 16719 22936 16764 22964
rect 16301 22927 16359 22933
rect 16758 22924 16764 22936
rect 16816 22924 16822 22976
rect 20162 22964 20168 22976
rect 20123 22936 20168 22964
rect 20162 22924 20168 22936
rect 20220 22924 20226 22976
rect 20714 22964 20720 22976
rect 20675 22936 20720 22964
rect 20714 22924 20720 22936
rect 20772 22924 20778 22976
rect 23014 22964 23020 22976
rect 22975 22936 23020 22964
rect 23014 22924 23020 22936
rect 23072 22924 23078 22976
rect 24581 22967 24639 22973
rect 24581 22933 24593 22967
rect 24627 22964 24639 22967
rect 24854 22964 24860 22976
rect 24627 22936 24860 22964
rect 24627 22933 24639 22936
rect 24581 22927 24639 22933
rect 24854 22924 24860 22936
rect 24912 22924 24918 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 1578 22720 1584 22772
rect 1636 22760 1642 22772
rect 2685 22763 2743 22769
rect 2685 22760 2697 22763
rect 1636 22732 2697 22760
rect 1636 22720 1642 22732
rect 2685 22729 2697 22732
rect 2731 22729 2743 22763
rect 2685 22723 2743 22729
rect 3234 22720 3240 22772
rect 3292 22760 3298 22772
rect 3789 22763 3847 22769
rect 3789 22760 3801 22763
rect 3292 22732 3801 22760
rect 3292 22720 3298 22732
rect 3789 22729 3801 22732
rect 3835 22729 3847 22763
rect 4982 22760 4988 22772
rect 4943 22732 4988 22760
rect 3789 22723 3847 22729
rect 4982 22720 4988 22732
rect 5040 22720 5046 22772
rect 6546 22760 6552 22772
rect 6507 22732 6552 22760
rect 6546 22720 6552 22732
rect 6604 22720 6610 22772
rect 8110 22720 8116 22772
rect 8168 22760 8174 22772
rect 8757 22763 8815 22769
rect 8757 22760 8769 22763
rect 8168 22732 8769 22760
rect 8168 22720 8174 22732
rect 8757 22729 8769 22732
rect 8803 22729 8815 22763
rect 8757 22723 8815 22729
rect 9217 22763 9275 22769
rect 9217 22729 9229 22763
rect 9263 22760 9275 22763
rect 9398 22760 9404 22772
rect 9263 22732 9404 22760
rect 9263 22729 9275 22732
rect 9217 22723 9275 22729
rect 6086 22692 6092 22704
rect 6012 22664 6092 22692
rect 5534 22584 5540 22636
rect 5592 22624 5598 22636
rect 5629 22627 5687 22633
rect 5629 22624 5641 22627
rect 5592 22596 5641 22624
rect 5592 22584 5598 22596
rect 5629 22593 5641 22596
rect 5675 22593 5687 22627
rect 5629 22587 5687 22593
rect 5813 22627 5871 22633
rect 5813 22593 5825 22627
rect 5859 22624 5871 22627
rect 6012 22624 6040 22664
rect 6086 22652 6092 22664
rect 6144 22652 6150 22704
rect 6178 22624 6184 22636
rect 5859 22596 6040 22624
rect 6139 22596 6184 22624
rect 5859 22593 5871 22596
rect 5813 22587 5871 22593
rect 1397 22559 1455 22565
rect 1397 22525 1409 22559
rect 1443 22556 1455 22559
rect 2501 22559 2559 22565
rect 1443 22528 2084 22556
rect 1443 22525 1455 22528
rect 1397 22519 1455 22525
rect 2056 22497 2084 22528
rect 2501 22525 2513 22559
rect 2547 22556 2559 22559
rect 3142 22556 3148 22568
rect 2547 22528 3148 22556
rect 2547 22525 2559 22528
rect 2501 22519 2559 22525
rect 3142 22516 3148 22528
rect 3200 22516 3206 22568
rect 3605 22559 3663 22565
rect 3605 22525 3617 22559
rect 3651 22556 3663 22559
rect 4709 22559 4767 22565
rect 3651 22528 4292 22556
rect 3651 22525 3663 22528
rect 3605 22519 3663 22525
rect 2041 22491 2099 22497
rect 2041 22457 2053 22491
rect 2087 22488 2099 22491
rect 2314 22488 2320 22500
rect 2087 22460 2320 22488
rect 2087 22457 2099 22460
rect 2041 22451 2099 22457
rect 2314 22448 2320 22460
rect 2372 22448 2378 22500
rect 1578 22420 1584 22432
rect 1539 22392 1584 22420
rect 1578 22380 1584 22392
rect 1636 22380 1642 22432
rect 2406 22420 2412 22432
rect 2367 22392 2412 22420
rect 2406 22380 2412 22392
rect 2464 22380 2470 22432
rect 3326 22380 3332 22432
rect 3384 22420 3390 22432
rect 4264 22429 4292 22528
rect 4709 22525 4721 22559
rect 4755 22556 4767 22559
rect 5828 22556 5856 22587
rect 6178 22584 6184 22596
rect 6236 22624 6242 22636
rect 7193 22627 7251 22633
rect 7193 22624 7205 22627
rect 6236 22596 7205 22624
rect 6236 22584 6242 22596
rect 7193 22593 7205 22596
rect 7239 22593 7251 22627
rect 7193 22587 7251 22593
rect 6546 22556 6552 22568
rect 4755 22528 6552 22556
rect 4755 22525 4767 22528
rect 4709 22519 4767 22525
rect 6546 22516 6552 22528
rect 6604 22516 6610 22568
rect 4982 22448 4988 22500
rect 5040 22488 5046 22500
rect 5537 22491 5595 22497
rect 5537 22488 5549 22491
rect 5040 22460 5549 22488
rect 5040 22448 5046 22460
rect 5537 22457 5549 22460
rect 5583 22488 5595 22491
rect 7098 22488 7104 22500
rect 5583 22460 7104 22488
rect 5583 22457 5595 22460
rect 5537 22451 5595 22457
rect 7098 22448 7104 22460
rect 7156 22448 7162 22500
rect 7208 22488 7236 22587
rect 7282 22584 7288 22636
rect 7340 22624 7346 22636
rect 7926 22624 7932 22636
rect 7340 22596 7932 22624
rect 7340 22584 7346 22596
rect 7926 22584 7932 22596
rect 7984 22584 7990 22636
rect 7466 22516 7472 22568
rect 7524 22556 7530 22568
rect 7745 22559 7803 22565
rect 7745 22556 7757 22559
rect 7524 22528 7757 22556
rect 7524 22516 7530 22528
rect 7745 22525 7757 22528
rect 7791 22525 7803 22559
rect 7745 22519 7803 22525
rect 7837 22491 7895 22497
rect 7837 22488 7849 22491
rect 7208 22460 7849 22488
rect 7837 22457 7849 22460
rect 7883 22488 7895 22491
rect 8018 22488 8024 22500
rect 7883 22460 8024 22488
rect 7883 22457 7895 22460
rect 7837 22451 7895 22457
rect 8018 22448 8024 22460
rect 8076 22488 8082 22500
rect 8389 22491 8447 22497
rect 8389 22488 8401 22491
rect 8076 22460 8401 22488
rect 8076 22448 8082 22460
rect 8389 22457 8401 22460
rect 8435 22457 8447 22491
rect 8772 22488 8800 22723
rect 9398 22720 9404 22732
rect 9456 22720 9462 22772
rect 10781 22763 10839 22769
rect 10781 22729 10793 22763
rect 10827 22760 10839 22763
rect 11054 22760 11060 22772
rect 10827 22732 11060 22760
rect 10827 22729 10839 22732
rect 10781 22723 10839 22729
rect 11054 22720 11060 22732
rect 11112 22720 11118 22772
rect 11422 22720 11428 22772
rect 11480 22760 11486 22772
rect 11793 22763 11851 22769
rect 11793 22760 11805 22763
rect 11480 22732 11805 22760
rect 11480 22720 11486 22732
rect 11793 22729 11805 22732
rect 11839 22729 11851 22763
rect 11793 22723 11851 22729
rect 12253 22763 12311 22769
rect 12253 22729 12265 22763
rect 12299 22760 12311 22763
rect 12434 22760 12440 22772
rect 12299 22732 12440 22760
rect 12299 22729 12311 22732
rect 12253 22723 12311 22729
rect 9214 22584 9220 22636
rect 9272 22624 9278 22636
rect 9769 22627 9827 22633
rect 9769 22624 9781 22627
rect 9272 22596 9781 22624
rect 9272 22584 9278 22596
rect 9769 22593 9781 22596
rect 9815 22593 9827 22627
rect 9769 22587 9827 22593
rect 10321 22627 10379 22633
rect 10321 22593 10333 22627
rect 10367 22624 10379 22627
rect 11238 22624 11244 22636
rect 10367 22596 11244 22624
rect 10367 22593 10379 22596
rect 10321 22587 10379 22593
rect 11238 22584 11244 22596
rect 11296 22624 11302 22636
rect 11333 22627 11391 22633
rect 11333 22624 11345 22627
rect 11296 22596 11345 22624
rect 11296 22584 11302 22596
rect 11333 22593 11345 22596
rect 11379 22593 11391 22627
rect 11808 22624 11836 22723
rect 12434 22720 12440 22732
rect 12492 22760 12498 22772
rect 13630 22760 13636 22772
rect 12492 22732 13636 22760
rect 12492 22720 12498 22732
rect 13630 22720 13636 22732
rect 13688 22720 13694 22772
rect 14277 22763 14335 22769
rect 14277 22729 14289 22763
rect 14323 22760 14335 22763
rect 14826 22760 14832 22772
rect 14323 22732 14832 22760
rect 14323 22729 14335 22732
rect 14277 22723 14335 22729
rect 14826 22720 14832 22732
rect 14884 22720 14890 22772
rect 15105 22763 15163 22769
rect 15105 22729 15117 22763
rect 15151 22760 15163 22763
rect 15562 22760 15568 22772
rect 15151 22732 15568 22760
rect 15151 22729 15163 22732
rect 15105 22723 15163 22729
rect 15562 22720 15568 22732
rect 15620 22760 15626 22772
rect 16022 22760 16028 22772
rect 15620 22732 16028 22760
rect 15620 22720 15626 22732
rect 16022 22720 16028 22732
rect 16080 22760 16086 22772
rect 16301 22763 16359 22769
rect 16301 22760 16313 22763
rect 16080 22732 16313 22760
rect 16080 22720 16086 22732
rect 16301 22729 16313 22732
rect 16347 22729 16359 22763
rect 16301 22723 16359 22729
rect 12342 22652 12348 22704
rect 12400 22692 12406 22704
rect 14737 22695 14795 22701
rect 12400 22664 14596 22692
rect 12400 22652 12406 22664
rect 12250 22624 12256 22636
rect 11808 22596 12256 22624
rect 11333 22587 11391 22593
rect 12250 22584 12256 22596
rect 12308 22624 12314 22636
rect 12897 22627 12955 22633
rect 12897 22624 12909 22627
rect 12308 22596 12909 22624
rect 12308 22584 12314 22596
rect 12897 22593 12909 22596
rect 12943 22593 12955 22627
rect 12897 22587 12955 22593
rect 13081 22627 13139 22633
rect 13081 22593 13093 22627
rect 13127 22624 13139 22627
rect 13538 22624 13544 22636
rect 13127 22596 13544 22624
rect 13127 22593 13139 22596
rect 13081 22587 13139 22593
rect 13538 22584 13544 22596
rect 13596 22584 13602 22636
rect 9122 22516 9128 22568
rect 9180 22556 9186 22568
rect 9677 22559 9735 22565
rect 9677 22556 9689 22559
rect 9180 22528 9689 22556
rect 9180 22516 9186 22528
rect 9677 22525 9689 22528
rect 9723 22556 9735 22559
rect 10686 22556 10692 22568
rect 9723 22528 10692 22556
rect 9723 22525 9735 22528
rect 9677 22519 9735 22525
rect 10686 22516 10692 22528
rect 10744 22516 10750 22568
rect 13262 22516 13268 22568
rect 13320 22556 13326 22568
rect 14093 22559 14151 22565
rect 14093 22556 14105 22559
rect 13320 22528 14105 22556
rect 13320 22516 13326 22528
rect 14093 22525 14105 22528
rect 14139 22556 14151 22559
rect 14458 22556 14464 22568
rect 14139 22528 14464 22556
rect 14139 22525 14151 22528
rect 14093 22519 14151 22525
rect 14458 22516 14464 22528
rect 14516 22516 14522 22568
rect 9306 22488 9312 22500
rect 8772 22460 9312 22488
rect 8389 22451 8447 22457
rect 9306 22448 9312 22460
rect 9364 22448 9370 22500
rect 10502 22448 10508 22500
rect 10560 22488 10566 22500
rect 10597 22491 10655 22497
rect 10597 22488 10609 22491
rect 10560 22460 10609 22488
rect 10560 22448 10566 22460
rect 10597 22457 10609 22460
rect 10643 22488 10655 22491
rect 11241 22491 11299 22497
rect 11241 22488 11253 22491
rect 10643 22460 11253 22488
rect 10643 22457 10655 22460
rect 10597 22451 10655 22457
rect 11241 22457 11253 22460
rect 11287 22488 11299 22491
rect 12805 22491 12863 22497
rect 12805 22488 12817 22491
rect 11287 22460 12817 22488
rect 11287 22457 11299 22460
rect 11241 22451 11299 22457
rect 12805 22457 12817 22460
rect 12851 22488 12863 22491
rect 12894 22488 12900 22500
rect 12851 22460 12900 22488
rect 12851 22457 12863 22460
rect 12805 22451 12863 22457
rect 12894 22448 12900 22460
rect 12952 22448 12958 22500
rect 13354 22448 13360 22500
rect 13412 22488 13418 22500
rect 13817 22491 13875 22497
rect 13817 22488 13829 22491
rect 13412 22460 13829 22488
rect 13412 22448 13418 22460
rect 13817 22457 13829 22460
rect 13863 22457 13875 22491
rect 14568 22488 14596 22664
rect 14737 22661 14749 22695
rect 14783 22692 14795 22695
rect 16316 22692 16344 22723
rect 16574 22720 16580 22772
rect 16632 22760 16638 22772
rect 16669 22763 16727 22769
rect 16669 22760 16681 22763
rect 16632 22732 16681 22760
rect 16632 22720 16638 22732
rect 16669 22729 16681 22732
rect 16715 22729 16727 22763
rect 16669 22723 16727 22729
rect 17218 22720 17224 22772
rect 17276 22760 17282 22772
rect 17405 22763 17463 22769
rect 17405 22760 17417 22763
rect 17276 22732 17417 22760
rect 17276 22720 17282 22732
rect 17405 22729 17417 22732
rect 17451 22729 17463 22763
rect 19058 22760 19064 22772
rect 19019 22732 19064 22760
rect 17405 22723 17463 22729
rect 19058 22720 19064 22732
rect 19116 22720 19122 22772
rect 19610 22760 19616 22772
rect 19571 22732 19616 22760
rect 19610 22720 19616 22732
rect 19668 22720 19674 22772
rect 20898 22720 20904 22772
rect 20956 22760 20962 22772
rect 21453 22763 21511 22769
rect 21453 22760 21465 22763
rect 20956 22732 21465 22760
rect 20956 22720 20962 22732
rect 21453 22729 21465 22732
rect 21499 22729 21511 22763
rect 23842 22760 23848 22772
rect 23803 22732 23848 22760
rect 21453 22723 21511 22729
rect 23842 22720 23848 22732
rect 23900 22760 23906 22772
rect 23900 22732 24532 22760
rect 23900 22720 23906 22732
rect 18049 22695 18107 22701
rect 14783 22664 15792 22692
rect 16316 22664 16620 22692
rect 14783 22661 14795 22664
rect 14737 22655 14795 22661
rect 14642 22584 14648 22636
rect 14700 22624 14706 22636
rect 14918 22624 14924 22636
rect 14700 22596 14924 22624
rect 14700 22584 14706 22596
rect 14918 22584 14924 22596
rect 14976 22584 14982 22636
rect 15378 22584 15384 22636
rect 15436 22624 15442 22636
rect 15764 22633 15792 22664
rect 15657 22627 15715 22633
rect 15657 22624 15669 22627
rect 15436 22596 15669 22624
rect 15436 22584 15442 22596
rect 15657 22593 15669 22596
rect 15703 22593 15715 22627
rect 15657 22587 15715 22593
rect 15749 22627 15807 22633
rect 15749 22593 15761 22627
rect 15795 22624 15807 22627
rect 16482 22624 16488 22636
rect 15795 22596 16488 22624
rect 15795 22593 15807 22596
rect 15749 22587 15807 22593
rect 16482 22584 16488 22596
rect 16540 22584 16546 22636
rect 15562 22556 15568 22568
rect 15523 22528 15568 22556
rect 15562 22516 15568 22528
rect 15620 22516 15626 22568
rect 16592 22556 16620 22664
rect 18049 22661 18061 22695
rect 18095 22692 18107 22695
rect 18690 22692 18696 22704
rect 18095 22664 18696 22692
rect 18095 22661 18107 22664
rect 18049 22655 18107 22661
rect 18690 22652 18696 22664
rect 18748 22652 18754 22704
rect 20717 22695 20775 22701
rect 20717 22692 20729 22695
rect 18800 22664 20729 22692
rect 16758 22584 16764 22636
rect 16816 22624 16822 22636
rect 18509 22627 18567 22633
rect 18509 22624 18521 22627
rect 16816 22596 18521 22624
rect 16816 22584 16822 22596
rect 18509 22593 18521 22596
rect 18555 22593 18567 22627
rect 18509 22587 18567 22593
rect 18601 22627 18659 22633
rect 18601 22593 18613 22627
rect 18647 22624 18659 22627
rect 18800 22624 18828 22664
rect 20717 22661 20729 22664
rect 20763 22661 20775 22695
rect 20717 22655 20775 22661
rect 23566 22652 23572 22704
rect 23624 22692 23630 22704
rect 23750 22692 23756 22704
rect 23624 22664 23756 22692
rect 23624 22652 23630 22664
rect 23750 22652 23756 22664
rect 23808 22652 23814 22704
rect 18647 22596 18828 22624
rect 18647 22593 18659 22596
rect 18601 22587 18659 22593
rect 16853 22559 16911 22565
rect 16853 22556 16865 22559
rect 16592 22528 16865 22556
rect 16853 22525 16865 22528
rect 16899 22525 16911 22559
rect 16853 22519 16911 22525
rect 17310 22516 17316 22568
rect 17368 22556 17374 22568
rect 18616 22556 18644 22587
rect 19794 22584 19800 22636
rect 19852 22624 19858 22636
rect 20165 22627 20223 22633
rect 20165 22624 20177 22627
rect 19852 22596 20177 22624
rect 19852 22584 19858 22596
rect 20165 22593 20177 22596
rect 20211 22593 20223 22627
rect 22094 22624 22100 22636
rect 22007 22596 22100 22624
rect 20165 22587 20223 22593
rect 22094 22584 22100 22596
rect 22152 22624 22158 22636
rect 24504 22633 24532 22732
rect 25038 22692 25044 22704
rect 24999 22664 25044 22692
rect 25038 22652 25044 22664
rect 25096 22652 25102 22704
rect 22557 22627 22615 22633
rect 22557 22624 22569 22627
rect 22152 22596 22569 22624
rect 22152 22584 22158 22596
rect 22557 22593 22569 22596
rect 22603 22624 22615 22627
rect 24489 22627 24547 22633
rect 22603 22596 23980 22624
rect 22603 22593 22615 22596
rect 22557 22587 22615 22593
rect 17368 22528 18644 22556
rect 19429 22559 19487 22565
rect 17368 22516 17374 22528
rect 19429 22525 19441 22559
rect 19475 22556 19487 22559
rect 19981 22559 20039 22565
rect 19981 22556 19993 22559
rect 19475 22528 19993 22556
rect 19475 22525 19487 22528
rect 19429 22519 19487 22525
rect 19981 22525 19993 22528
rect 20027 22556 20039 22559
rect 20346 22556 20352 22568
rect 20027 22528 20352 22556
rect 20027 22525 20039 22528
rect 19981 22519 20039 22525
rect 20346 22516 20352 22528
rect 20404 22516 20410 22568
rect 20714 22516 20720 22568
rect 20772 22556 20778 22568
rect 21726 22556 21732 22568
rect 20772 22528 21732 22556
rect 20772 22516 20778 22528
rect 21726 22516 21732 22528
rect 21784 22556 21790 22568
rect 21821 22559 21879 22565
rect 21821 22556 21833 22559
rect 21784 22528 21833 22556
rect 21784 22516 21790 22528
rect 21821 22525 21833 22528
rect 21867 22525 21879 22559
rect 21821 22519 21879 22525
rect 23382 22516 23388 22568
rect 23440 22556 23446 22568
rect 23566 22556 23572 22568
rect 23440 22528 23572 22556
rect 23440 22516 23446 22528
rect 23566 22516 23572 22528
rect 23624 22516 23630 22568
rect 23842 22516 23848 22568
rect 23900 22516 23906 22568
rect 23952 22556 23980 22596
rect 24489 22593 24501 22627
rect 24535 22593 24547 22627
rect 24489 22587 24547 22593
rect 24673 22627 24731 22633
rect 24673 22593 24685 22627
rect 24719 22624 24731 22627
rect 24854 22624 24860 22636
rect 24719 22596 24860 22624
rect 24719 22593 24731 22596
rect 24673 22587 24731 22593
rect 24688 22556 24716 22587
rect 24854 22584 24860 22596
rect 24912 22584 24918 22636
rect 23952 22528 24716 22556
rect 18322 22488 18328 22500
rect 14568 22460 18328 22488
rect 13817 22451 13875 22457
rect 18322 22448 18328 22460
rect 18380 22448 18386 22500
rect 19518 22448 19524 22500
rect 19576 22488 19582 22500
rect 20073 22491 20131 22497
rect 20073 22488 20085 22491
rect 19576 22460 20085 22488
rect 19576 22448 19582 22460
rect 20073 22457 20085 22460
rect 20119 22457 20131 22491
rect 20073 22451 20131 22457
rect 23477 22491 23535 22497
rect 23477 22457 23489 22491
rect 23523 22488 23535 22491
rect 23860 22488 23888 22516
rect 24397 22491 24455 22497
rect 24397 22488 24409 22491
rect 23523 22460 24409 22488
rect 23523 22457 23535 22460
rect 23477 22451 23535 22457
rect 24397 22457 24409 22460
rect 24443 22457 24455 22491
rect 24397 22451 24455 22457
rect 3421 22423 3479 22429
rect 3421 22420 3433 22423
rect 3384 22392 3433 22420
rect 3384 22380 3390 22392
rect 3421 22389 3433 22392
rect 3467 22389 3479 22423
rect 3421 22383 3479 22389
rect 4249 22423 4307 22429
rect 4249 22389 4261 22423
rect 4295 22420 4307 22423
rect 4522 22420 4528 22432
rect 4295 22392 4528 22420
rect 4295 22389 4307 22392
rect 4249 22383 4307 22389
rect 4522 22380 4528 22392
rect 4580 22380 4586 22432
rect 5074 22380 5080 22432
rect 5132 22420 5138 22432
rect 5169 22423 5227 22429
rect 5169 22420 5181 22423
rect 5132 22392 5181 22420
rect 5132 22380 5138 22392
rect 5169 22389 5181 22392
rect 5215 22389 5227 22423
rect 5169 22383 5227 22389
rect 6178 22380 6184 22432
rect 6236 22420 6242 22432
rect 6638 22420 6644 22432
rect 6236 22392 6644 22420
rect 6236 22380 6242 22392
rect 6638 22380 6644 22392
rect 6696 22380 6702 22432
rect 7374 22420 7380 22432
rect 7335 22392 7380 22420
rect 7374 22380 7380 22392
rect 7432 22380 7438 22432
rect 8846 22380 8852 22432
rect 8904 22420 8910 22432
rect 9585 22423 9643 22429
rect 9585 22420 9597 22423
rect 8904 22392 9597 22420
rect 8904 22380 8910 22392
rect 9585 22389 9597 22392
rect 9631 22389 9643 22423
rect 9585 22383 9643 22389
rect 11054 22380 11060 22432
rect 11112 22420 11118 22432
rect 11149 22423 11207 22429
rect 11149 22420 11161 22423
rect 11112 22392 11161 22420
rect 11112 22380 11118 22392
rect 11149 22389 11161 22392
rect 11195 22389 11207 22423
rect 12434 22420 12440 22432
rect 12395 22392 12440 22420
rect 11149 22383 11207 22389
rect 12434 22380 12440 22392
rect 12492 22380 12498 22432
rect 13538 22420 13544 22432
rect 13499 22392 13544 22420
rect 13538 22380 13544 22392
rect 13596 22380 13602 22432
rect 15197 22423 15255 22429
rect 15197 22389 15209 22423
rect 15243 22420 15255 22423
rect 16298 22420 16304 22432
rect 15243 22392 16304 22420
rect 15243 22389 15255 22392
rect 15197 22383 15255 22389
rect 16298 22380 16304 22392
rect 16356 22380 16362 22432
rect 17034 22420 17040 22432
rect 16995 22392 17040 22420
rect 17034 22380 17040 22392
rect 17092 22380 17098 22432
rect 17770 22420 17776 22432
rect 17731 22392 17776 22420
rect 17770 22380 17776 22392
rect 17828 22380 17834 22432
rect 18138 22380 18144 22432
rect 18196 22420 18202 22432
rect 18417 22423 18475 22429
rect 18417 22420 18429 22423
rect 18196 22392 18429 22420
rect 18196 22380 18202 22392
rect 18417 22389 18429 22392
rect 18463 22389 18475 22423
rect 18417 22383 18475 22389
rect 19242 22380 19248 22432
rect 19300 22420 19306 22432
rect 21085 22423 21143 22429
rect 21085 22420 21097 22423
rect 19300 22392 21097 22420
rect 19300 22380 19306 22392
rect 21085 22389 21097 22392
rect 21131 22420 21143 22423
rect 21358 22420 21364 22432
rect 21131 22392 21364 22420
rect 21131 22389 21143 22392
rect 21085 22383 21143 22389
rect 21358 22380 21364 22392
rect 21416 22380 21422 22432
rect 21542 22380 21548 22432
rect 21600 22420 21606 22432
rect 21913 22423 21971 22429
rect 21913 22420 21925 22423
rect 21600 22392 21925 22420
rect 21600 22380 21606 22392
rect 21913 22389 21925 22392
rect 21959 22389 21971 22423
rect 21913 22383 21971 22389
rect 23109 22423 23167 22429
rect 23109 22389 23121 22423
rect 23155 22420 23167 22423
rect 23198 22420 23204 22432
rect 23155 22392 23204 22420
rect 23155 22389 23167 22392
rect 23109 22383 23167 22389
rect 23198 22380 23204 22392
rect 23256 22420 23262 22432
rect 23382 22420 23388 22432
rect 23256 22392 23388 22420
rect 23256 22380 23262 22392
rect 23382 22380 23388 22392
rect 23440 22380 23446 22432
rect 24026 22420 24032 22432
rect 23987 22392 24032 22420
rect 24026 22380 24032 22392
rect 24084 22380 24090 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 2777 22219 2835 22225
rect 2777 22185 2789 22219
rect 2823 22216 2835 22219
rect 2866 22216 2872 22228
rect 2823 22188 2872 22216
rect 2823 22185 2835 22188
rect 2777 22179 2835 22185
rect 2866 22176 2872 22188
rect 2924 22176 2930 22228
rect 5074 22216 5080 22228
rect 4172 22188 5080 22216
rect 1578 22040 1584 22092
rect 1636 22080 1642 22092
rect 1949 22083 2007 22089
rect 1949 22080 1961 22083
rect 1636 22052 1961 22080
rect 1636 22040 1642 22052
rect 1949 22049 1961 22052
rect 1995 22049 2007 22083
rect 1949 22043 2007 22049
rect 2225 22083 2283 22089
rect 2225 22049 2237 22083
rect 2271 22080 2283 22083
rect 2682 22080 2688 22092
rect 2271 22052 2688 22080
rect 2271 22049 2283 22052
rect 2225 22043 2283 22049
rect 2682 22040 2688 22052
rect 2740 22040 2746 22092
rect 3881 22083 3939 22089
rect 3881 22049 3893 22083
rect 3927 22080 3939 22083
rect 4172 22080 4200 22188
rect 5074 22176 5080 22188
rect 5132 22176 5138 22228
rect 6917 22219 6975 22225
rect 6917 22185 6929 22219
rect 6963 22216 6975 22219
rect 7282 22216 7288 22228
rect 6963 22188 7288 22216
rect 6963 22185 6975 22188
rect 6917 22179 6975 22185
rect 7282 22176 7288 22188
rect 7340 22176 7346 22228
rect 7926 22176 7932 22228
rect 7984 22216 7990 22228
rect 8662 22216 8668 22228
rect 7984 22188 8668 22216
rect 7984 22176 7990 22188
rect 8662 22176 8668 22188
rect 8720 22176 8726 22228
rect 9122 22176 9128 22228
rect 9180 22216 9186 22228
rect 9490 22216 9496 22228
rect 9180 22188 9496 22216
rect 9180 22176 9186 22188
rect 9490 22176 9496 22188
rect 9548 22176 9554 22228
rect 12894 22216 12900 22228
rect 12855 22188 12900 22216
rect 12894 22176 12900 22188
rect 12952 22176 12958 22228
rect 13262 22176 13268 22228
rect 13320 22216 13326 22228
rect 13446 22216 13452 22228
rect 13320 22188 13452 22216
rect 13320 22176 13326 22188
rect 13446 22176 13452 22188
rect 13504 22176 13510 22228
rect 15289 22219 15347 22225
rect 15289 22185 15301 22219
rect 15335 22216 15347 22219
rect 15562 22216 15568 22228
rect 15335 22188 15568 22216
rect 15335 22185 15347 22188
rect 15289 22179 15347 22185
rect 15562 22176 15568 22188
rect 15620 22176 15626 22228
rect 16853 22219 16911 22225
rect 16853 22216 16865 22219
rect 16592 22188 16865 22216
rect 7190 22108 7196 22160
rect 7248 22148 7254 22160
rect 7650 22148 7656 22160
rect 7248 22120 7656 22148
rect 7248 22108 7254 22120
rect 7650 22108 7656 22120
rect 7708 22108 7714 22160
rect 11146 22148 11152 22160
rect 11072 22120 11152 22148
rect 3927 22052 4200 22080
rect 3927 22049 3939 22052
rect 3881 22043 3939 22049
rect 4982 22040 4988 22092
rect 5040 22080 5046 22092
rect 7282 22089 7288 22092
rect 5077 22083 5135 22089
rect 5077 22080 5089 22083
rect 5040 22052 5089 22080
rect 5040 22040 5046 22052
rect 5077 22049 5089 22052
rect 5123 22049 5135 22083
rect 7276 22080 7288 22089
rect 7243 22052 7288 22080
rect 5077 22043 5135 22049
rect 7276 22043 7288 22052
rect 7282 22040 7288 22043
rect 7340 22040 7346 22092
rect 8662 22040 8668 22092
rect 8720 22080 8726 22092
rect 9861 22083 9919 22089
rect 9861 22080 9873 22083
rect 8720 22052 9873 22080
rect 8720 22040 8726 22052
rect 9861 22049 9873 22052
rect 9907 22080 9919 22083
rect 10134 22080 10140 22092
rect 9907 22052 10140 22080
rect 9907 22049 9919 22052
rect 9861 22043 9919 22049
rect 10134 22040 10140 22052
rect 10192 22040 10198 22092
rect 10505 22083 10563 22089
rect 10505 22049 10517 22083
rect 10551 22080 10563 22083
rect 11072 22080 11100 22120
rect 11146 22108 11152 22120
rect 11204 22148 11210 22160
rect 12342 22148 12348 22160
rect 11204 22120 12348 22148
rect 11204 22108 11210 22120
rect 12342 22108 12348 22120
rect 12400 22108 12406 22160
rect 12434 22108 12440 22160
rect 12492 22148 12498 22160
rect 14093 22151 14151 22157
rect 14093 22148 14105 22151
rect 12492 22120 14105 22148
rect 12492 22108 12498 22120
rect 13740 22092 13768 22120
rect 14093 22117 14105 22120
rect 14139 22117 14151 22151
rect 14093 22111 14151 22117
rect 11238 22089 11244 22092
rect 11232 22080 11244 22089
rect 10551 22052 11100 22080
rect 11199 22052 11244 22080
rect 10551 22049 10563 22052
rect 10505 22043 10563 22049
rect 11232 22043 11244 22052
rect 11238 22040 11244 22043
rect 11296 22040 11302 22092
rect 11974 22040 11980 22092
rect 12032 22040 12038 22092
rect 13722 22040 13728 22092
rect 13780 22040 13786 22092
rect 14001 22083 14059 22089
rect 14001 22049 14013 22083
rect 14047 22080 14059 22083
rect 14642 22080 14648 22092
rect 14047 22052 14648 22080
rect 14047 22049 14059 22052
rect 14001 22043 14059 22049
rect 14642 22040 14648 22052
rect 14700 22040 14706 22092
rect 15657 22083 15715 22089
rect 15657 22080 15669 22083
rect 15304 22052 15669 22080
rect 5166 22012 5172 22024
rect 5127 21984 5172 22012
rect 5166 21972 5172 21984
rect 5224 21972 5230 22024
rect 5353 22015 5411 22021
rect 5353 21981 5365 22015
rect 5399 22012 5411 22015
rect 5442 22012 5448 22024
rect 5399 21984 5448 22012
rect 5399 21981 5411 21984
rect 5353 21975 5411 21981
rect 5442 21972 5448 21984
rect 5500 21972 5506 22024
rect 7009 22015 7067 22021
rect 7009 21981 7021 22015
rect 7055 21981 7067 22015
rect 7009 21975 7067 21981
rect 3145 21947 3203 21953
rect 3145 21913 3157 21947
rect 3191 21944 3203 21947
rect 3602 21944 3608 21956
rect 3191 21916 3608 21944
rect 3191 21913 3203 21916
rect 3145 21907 3203 21913
rect 3602 21904 3608 21916
rect 3660 21904 3666 21956
rect 4709 21947 4767 21953
rect 4709 21913 4721 21947
rect 4755 21944 4767 21947
rect 4890 21944 4896 21956
rect 4755 21916 4896 21944
rect 4755 21913 4767 21916
rect 4709 21907 4767 21913
rect 4890 21904 4896 21916
rect 4948 21944 4954 21956
rect 5721 21947 5779 21953
rect 5721 21944 5733 21947
rect 4948 21916 5733 21944
rect 4948 21904 4954 21916
rect 5721 21913 5733 21916
rect 5767 21913 5779 21947
rect 5721 21907 5779 21913
rect 6638 21904 6644 21956
rect 6696 21944 6702 21956
rect 7024 21944 7052 21975
rect 8110 21972 8116 22024
rect 8168 22012 8174 22024
rect 8386 22012 8392 22024
rect 8168 21984 8392 22012
rect 8168 21972 8174 21984
rect 8386 21972 8392 21984
rect 8444 21972 8450 22024
rect 9674 21972 9680 22024
rect 9732 22012 9738 22024
rect 10965 22015 11023 22021
rect 10965 22012 10977 22015
rect 9732 21984 10977 22012
rect 9732 21972 9738 21984
rect 10965 21981 10977 21984
rect 11011 21981 11023 22015
rect 11992 22012 12020 22040
rect 14090 22012 14096 22024
rect 11992 21984 14096 22012
rect 10965 21975 11023 21981
rect 14090 21972 14096 21984
rect 14148 21972 14154 22024
rect 14277 22015 14335 22021
rect 14277 21981 14289 22015
rect 14323 22012 14335 22015
rect 14461 22015 14519 22021
rect 14461 22012 14473 22015
rect 14323 21984 14473 22012
rect 14323 21981 14335 21984
rect 14277 21975 14335 21981
rect 14461 21981 14473 21984
rect 14507 21981 14519 22015
rect 15304 22012 15332 22052
rect 15657 22049 15669 22052
rect 15703 22080 15715 22083
rect 16592 22080 16620 22188
rect 16853 22185 16865 22188
rect 16899 22185 16911 22219
rect 16853 22179 16911 22185
rect 20717 22219 20775 22225
rect 20717 22185 20729 22219
rect 20763 22216 20775 22219
rect 21174 22216 21180 22228
rect 20763 22188 21180 22216
rect 20763 22185 20775 22188
rect 20717 22179 20775 22185
rect 21174 22176 21180 22188
rect 21232 22216 21238 22228
rect 21542 22216 21548 22228
rect 21232 22188 21548 22216
rect 21232 22176 21238 22188
rect 21542 22176 21548 22188
rect 21600 22176 21606 22228
rect 21726 22176 21732 22228
rect 21784 22216 21790 22228
rect 21913 22219 21971 22225
rect 21913 22216 21925 22219
rect 21784 22188 21925 22216
rect 21784 22176 21790 22188
rect 21913 22185 21925 22188
rect 21959 22185 21971 22219
rect 21913 22179 21971 22185
rect 23385 22219 23443 22225
rect 23385 22185 23397 22219
rect 23431 22216 23443 22219
rect 23934 22216 23940 22228
rect 23431 22188 23940 22216
rect 23431 22185 23443 22188
rect 23385 22179 23443 22185
rect 23934 22176 23940 22188
rect 23992 22176 23998 22228
rect 24854 22176 24860 22228
rect 24912 22176 24918 22228
rect 18785 22151 18843 22157
rect 18785 22117 18797 22151
rect 18831 22148 18843 22151
rect 19058 22148 19064 22160
rect 18831 22120 19064 22148
rect 18831 22117 18843 22120
rect 18785 22111 18843 22117
rect 19058 22108 19064 22120
rect 19116 22108 19122 22160
rect 20898 22148 20904 22160
rect 20859 22120 20904 22148
rect 20898 22108 20904 22120
rect 20956 22108 20962 22160
rect 21821 22151 21879 22157
rect 21821 22117 21833 22151
rect 21867 22148 21879 22151
rect 22094 22148 22100 22160
rect 21867 22120 22100 22148
rect 21867 22117 21879 22120
rect 21821 22111 21879 22117
rect 22094 22108 22100 22120
rect 22152 22108 22158 22160
rect 24026 22148 24032 22160
rect 23400 22120 24032 22148
rect 17218 22080 17224 22092
rect 15703 22052 16620 22080
rect 17179 22052 17224 22080
rect 15703 22049 15715 22052
rect 15657 22043 15715 22049
rect 17218 22040 17224 22052
rect 17276 22040 17282 22092
rect 19518 22040 19524 22092
rect 19576 22080 19582 22092
rect 19613 22083 19671 22089
rect 19613 22080 19625 22083
rect 19576 22052 19625 22080
rect 19576 22040 19582 22052
rect 19613 22049 19625 22052
rect 19659 22049 19671 22083
rect 22278 22080 22284 22092
rect 22239 22052 22284 22080
rect 19613 22043 19671 22049
rect 22278 22040 22284 22052
rect 22336 22040 22342 22092
rect 23017 22083 23075 22089
rect 23017 22049 23029 22083
rect 23063 22080 23075 22083
rect 23400 22080 23428 22120
rect 24026 22108 24032 22120
rect 24084 22108 24090 22160
rect 23063 22052 23428 22080
rect 24305 22083 24363 22089
rect 23063 22049 23075 22052
rect 23017 22043 23075 22049
rect 24305 22049 24317 22083
rect 24351 22080 24363 22083
rect 24762 22080 24768 22092
rect 24351 22052 24768 22080
rect 24351 22049 24363 22052
rect 24305 22043 24363 22049
rect 24762 22040 24768 22052
rect 24820 22040 24826 22092
rect 14461 21975 14519 21981
rect 14660 21984 15332 22012
rect 6696 21916 7052 21944
rect 10045 21947 10103 21953
rect 6696 21904 6702 21916
rect 10045 21913 10057 21947
rect 10091 21944 10103 21947
rect 10686 21944 10692 21956
rect 10091 21916 10692 21944
rect 10091 21913 10103 21916
rect 10045 21907 10103 21913
rect 10686 21904 10692 21916
rect 10744 21904 10750 21956
rect 13541 21947 13599 21953
rect 13541 21913 13553 21947
rect 13587 21944 13599 21947
rect 14660 21944 14688 21984
rect 15562 21972 15568 22024
rect 15620 22012 15626 22024
rect 15749 22015 15807 22021
rect 15749 22012 15761 22015
rect 15620 21984 15761 22012
rect 15620 21972 15626 21984
rect 15749 21981 15761 21984
rect 15795 21981 15807 22015
rect 15749 21975 15807 21981
rect 15933 22015 15991 22021
rect 15933 21981 15945 22015
rect 15979 22012 15991 22015
rect 16298 22012 16304 22024
rect 15979 21984 16304 22012
rect 15979 21981 15991 21984
rect 15933 21975 15991 21981
rect 16298 21972 16304 21984
rect 16356 21972 16362 22024
rect 16393 22015 16451 22021
rect 16393 21981 16405 22015
rect 16439 22012 16451 22015
rect 16439 21984 16528 22012
rect 16439 21981 16451 21984
rect 16393 21975 16451 21981
rect 13587 21916 14688 21944
rect 14737 21947 14795 21953
rect 13587 21913 13599 21916
rect 13541 21907 13599 21913
rect 14737 21913 14749 21947
rect 14783 21944 14795 21947
rect 15470 21944 15476 21956
rect 14783 21916 15476 21944
rect 14783 21913 14795 21916
rect 14737 21907 14795 21913
rect 15470 21904 15476 21916
rect 15528 21904 15534 21956
rect 15838 21944 15844 21956
rect 15580 21916 15844 21944
rect 1394 21836 1400 21888
rect 1452 21876 1458 21888
rect 1581 21879 1639 21885
rect 1581 21876 1593 21879
rect 1452 21848 1593 21876
rect 1452 21836 1458 21848
rect 1581 21845 1593 21848
rect 1627 21845 1639 21879
rect 3510 21876 3516 21888
rect 3471 21848 3516 21876
rect 1581 21839 1639 21845
rect 3510 21836 3516 21848
rect 3568 21836 3574 21888
rect 4154 21836 4160 21888
rect 4212 21876 4218 21888
rect 4249 21879 4307 21885
rect 4249 21876 4261 21879
rect 4212 21848 4261 21876
rect 4212 21836 4218 21848
rect 4249 21845 4261 21848
rect 4295 21845 4307 21879
rect 4249 21839 4307 21845
rect 6273 21879 6331 21885
rect 6273 21845 6285 21879
rect 6319 21876 6331 21879
rect 6914 21876 6920 21888
rect 6319 21848 6920 21876
rect 6319 21845 6331 21848
rect 6273 21839 6331 21845
rect 6914 21836 6920 21848
rect 6972 21836 6978 21888
rect 8386 21876 8392 21888
rect 8347 21848 8392 21876
rect 8386 21836 8392 21848
rect 8444 21836 8450 21888
rect 9214 21876 9220 21888
rect 9175 21848 9220 21876
rect 9214 21836 9220 21848
rect 9272 21836 9278 21888
rect 10873 21879 10931 21885
rect 10873 21845 10885 21879
rect 10919 21876 10931 21879
rect 10962 21876 10968 21888
rect 10919 21848 10968 21876
rect 10919 21845 10931 21848
rect 10873 21839 10931 21845
rect 10962 21836 10968 21848
rect 11020 21836 11026 21888
rect 11974 21836 11980 21888
rect 12032 21876 12038 21888
rect 12345 21879 12403 21885
rect 12345 21876 12357 21879
rect 12032 21848 12357 21876
rect 12032 21836 12038 21848
rect 12345 21845 12357 21848
rect 12391 21845 12403 21879
rect 13630 21876 13636 21888
rect 13591 21848 13636 21876
rect 12345 21839 12403 21845
rect 13630 21836 13636 21848
rect 13688 21836 13694 21888
rect 14461 21879 14519 21885
rect 14461 21845 14473 21879
rect 14507 21876 14519 21879
rect 15105 21879 15163 21885
rect 15105 21876 15117 21879
rect 14507 21848 15117 21876
rect 14507 21845 14519 21848
rect 14461 21839 14519 21845
rect 15105 21845 15117 21848
rect 15151 21876 15163 21879
rect 15378 21876 15384 21888
rect 15151 21848 15384 21876
rect 15151 21845 15163 21848
rect 15105 21839 15163 21845
rect 15378 21836 15384 21848
rect 15436 21876 15442 21888
rect 15580 21876 15608 21916
rect 15838 21904 15844 21916
rect 15896 21944 15902 21956
rect 16500 21944 16528 21984
rect 16942 21972 16948 22024
rect 17000 22012 17006 22024
rect 17313 22015 17371 22021
rect 17313 22012 17325 22015
rect 17000 21984 17325 22012
rect 17000 21972 17006 21984
rect 17313 21981 17325 21984
rect 17359 21981 17371 22015
rect 17313 21975 17371 21981
rect 17497 22015 17555 22021
rect 17497 21981 17509 22015
rect 17543 22012 17555 22015
rect 17862 22012 17868 22024
rect 17543 21984 17868 22012
rect 17543 21981 17555 21984
rect 17497 21975 17555 21981
rect 15896 21916 16528 21944
rect 15896 21904 15902 21916
rect 15436 21848 15608 21876
rect 15436 21836 15442 21848
rect 15930 21836 15936 21888
rect 15988 21876 15994 21888
rect 16390 21876 16396 21888
rect 15988 21848 16396 21876
rect 15988 21836 15994 21848
rect 16390 21836 16396 21848
rect 16448 21836 16454 21888
rect 16500 21876 16528 21916
rect 16761 21947 16819 21953
rect 16761 21913 16773 21947
rect 16807 21944 16819 21947
rect 16850 21944 16856 21956
rect 16807 21916 16856 21944
rect 16807 21913 16819 21916
rect 16761 21907 16819 21913
rect 16850 21904 16856 21916
rect 16908 21904 16914 21956
rect 17512 21876 17540 21975
rect 17862 21972 17868 21984
rect 17920 21972 17926 22024
rect 18322 21972 18328 22024
rect 18380 22012 18386 22024
rect 18877 22015 18935 22021
rect 18877 22012 18889 22015
rect 18380 21984 18889 22012
rect 18380 21972 18386 21984
rect 18877 21981 18889 21984
rect 18923 21981 18935 22015
rect 18877 21975 18935 21981
rect 19061 22015 19119 22021
rect 19061 21981 19073 22015
rect 19107 22012 19119 22015
rect 19107 21984 20116 22012
rect 19107 21981 19119 21984
rect 19061 21975 19119 21981
rect 18138 21876 18144 21888
rect 16500 21848 17540 21876
rect 18099 21848 18144 21876
rect 18138 21836 18144 21848
rect 18196 21836 18202 21888
rect 18417 21879 18475 21885
rect 18417 21845 18429 21879
rect 18463 21876 18475 21879
rect 19242 21876 19248 21888
rect 18463 21848 19248 21876
rect 18463 21845 18475 21848
rect 18417 21839 18475 21845
rect 19242 21836 19248 21848
rect 19300 21836 19306 21888
rect 20088 21885 20116 21984
rect 22186 21972 22192 22024
rect 22244 22012 22250 22024
rect 22373 22015 22431 22021
rect 22373 22012 22385 22015
rect 22244 21984 22385 22012
rect 22244 21972 22250 21984
rect 22373 21981 22385 21984
rect 22419 21981 22431 22015
rect 22373 21975 22431 21981
rect 22465 22015 22523 22021
rect 22465 21981 22477 22015
rect 22511 21981 22523 22015
rect 22465 21975 22523 21981
rect 21453 21947 21511 21953
rect 21453 21913 21465 21947
rect 21499 21944 21511 21947
rect 21818 21944 21824 21956
rect 21499 21916 21824 21944
rect 21499 21913 21511 21916
rect 21453 21907 21511 21913
rect 21818 21904 21824 21916
rect 21876 21944 21882 21956
rect 22480 21944 22508 21975
rect 23290 21972 23296 22024
rect 23348 22012 23354 22024
rect 24397 22015 24455 22021
rect 24397 22012 24409 22015
rect 23348 21984 24409 22012
rect 23348 21972 23354 21984
rect 24397 21981 24409 21984
rect 24443 21981 24455 22015
rect 24397 21975 24455 21981
rect 24581 22015 24639 22021
rect 24581 21981 24593 22015
rect 24627 22012 24639 22015
rect 24872 22012 24900 22176
rect 24946 22012 24952 22024
rect 24627 21984 24952 22012
rect 24627 21981 24639 21984
rect 24581 21975 24639 21981
rect 24946 21972 24952 21984
rect 25004 21972 25010 22024
rect 21876 21916 22508 21944
rect 21876 21904 21882 21916
rect 23566 21904 23572 21956
rect 23624 21944 23630 21956
rect 24026 21944 24032 21956
rect 23624 21916 24032 21944
rect 23624 21904 23630 21916
rect 24026 21904 24032 21916
rect 24084 21904 24090 21956
rect 20073 21879 20131 21885
rect 20073 21845 20085 21879
rect 20119 21876 20131 21879
rect 20530 21876 20536 21888
rect 20119 21848 20536 21876
rect 20119 21845 20131 21848
rect 20073 21839 20131 21845
rect 20530 21836 20536 21848
rect 20588 21836 20594 21888
rect 23753 21879 23811 21885
rect 23753 21845 23765 21879
rect 23799 21876 23811 21879
rect 23934 21876 23940 21888
rect 23799 21848 23940 21876
rect 23799 21845 23811 21848
rect 23753 21839 23811 21845
rect 23934 21836 23940 21848
rect 23992 21836 23998 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 2685 21675 2743 21681
rect 2685 21641 2697 21675
rect 2731 21672 2743 21675
rect 3510 21672 3516 21684
rect 2731 21644 3516 21672
rect 2731 21641 2743 21644
rect 2685 21635 2743 21641
rect 3510 21632 3516 21644
rect 3568 21632 3574 21684
rect 4249 21675 4307 21681
rect 4249 21641 4261 21675
rect 4295 21672 4307 21675
rect 5166 21672 5172 21684
rect 4295 21644 5172 21672
rect 4295 21641 4307 21644
rect 4249 21635 4307 21641
rect 5166 21632 5172 21644
rect 5224 21672 5230 21684
rect 5629 21675 5687 21681
rect 5629 21672 5641 21675
rect 5224 21644 5641 21672
rect 5224 21632 5230 21644
rect 5629 21641 5641 21644
rect 5675 21641 5687 21675
rect 5629 21635 5687 21641
rect 6546 21632 6552 21684
rect 6604 21672 6610 21684
rect 8205 21675 8263 21681
rect 8205 21672 8217 21675
rect 6604 21644 8217 21672
rect 6604 21632 6610 21644
rect 8205 21641 8217 21644
rect 8251 21641 8263 21675
rect 9674 21672 9680 21684
rect 8205 21635 8263 21641
rect 9324 21644 9680 21672
rect 2225 21539 2283 21545
rect 2225 21505 2237 21539
rect 2271 21536 2283 21539
rect 3050 21536 3056 21548
rect 2271 21508 3056 21536
rect 2271 21505 2283 21508
rect 2225 21499 2283 21505
rect 3050 21496 3056 21508
rect 3108 21536 3114 21548
rect 3237 21539 3295 21545
rect 3237 21536 3249 21539
rect 3108 21508 3249 21536
rect 3108 21496 3114 21508
rect 3237 21505 3249 21508
rect 3283 21505 3295 21539
rect 3237 21499 3295 21505
rect 4338 21496 4344 21548
rect 4396 21536 4402 21548
rect 4706 21536 4712 21548
rect 4396 21508 4712 21536
rect 4396 21496 4402 21508
rect 4706 21496 4712 21508
rect 4764 21496 4770 21548
rect 4801 21539 4859 21545
rect 4801 21505 4813 21539
rect 4847 21536 4859 21539
rect 5166 21536 5172 21548
rect 4847 21508 5172 21536
rect 4847 21505 4859 21508
rect 4801 21499 4859 21505
rect 1394 21468 1400 21480
rect 1355 21440 1400 21468
rect 1394 21428 1400 21440
rect 1452 21428 1458 21480
rect 1578 21428 1584 21480
rect 1636 21468 1642 21480
rect 3697 21471 3755 21477
rect 3697 21468 3709 21471
rect 1636 21440 3709 21468
rect 1636 21428 1642 21440
rect 3697 21437 3709 21440
rect 3743 21437 3755 21471
rect 3697 21431 3755 21437
rect 4157 21471 4215 21477
rect 4157 21437 4169 21471
rect 4203 21468 4215 21471
rect 4816 21468 4844 21499
rect 5166 21496 5172 21508
rect 5224 21496 5230 21548
rect 6086 21496 6092 21548
rect 6144 21536 6150 21548
rect 6638 21536 6644 21548
rect 6144 21508 6644 21536
rect 6144 21496 6150 21508
rect 6638 21496 6644 21508
rect 6696 21536 6702 21548
rect 9324 21545 9352 21644
rect 9674 21632 9680 21644
rect 9732 21632 9738 21684
rect 9950 21632 9956 21684
rect 10008 21672 10014 21684
rect 10689 21675 10747 21681
rect 10689 21672 10701 21675
rect 10008 21644 10701 21672
rect 10008 21632 10014 21644
rect 10689 21641 10701 21644
rect 10735 21641 10747 21675
rect 12250 21672 12256 21684
rect 12211 21644 12256 21672
rect 10689 21635 10747 21641
rect 12250 21632 12256 21644
rect 12308 21632 12314 21684
rect 12342 21632 12348 21684
rect 12400 21672 12406 21684
rect 12437 21675 12495 21681
rect 12437 21672 12449 21675
rect 12400 21644 12449 21672
rect 12400 21632 12406 21644
rect 12437 21641 12449 21644
rect 12483 21641 12495 21675
rect 12437 21635 12495 21641
rect 13722 21632 13728 21684
rect 13780 21672 13786 21684
rect 14001 21675 14059 21681
rect 14001 21672 14013 21675
rect 13780 21644 14013 21672
rect 13780 21632 13786 21644
rect 14001 21641 14013 21644
rect 14047 21641 14059 21675
rect 14001 21635 14059 21641
rect 14090 21632 14096 21684
rect 14148 21672 14154 21684
rect 17218 21672 17224 21684
rect 14148 21644 15884 21672
rect 17179 21644 17224 21672
rect 14148 21632 14154 21644
rect 6825 21539 6883 21545
rect 6825 21536 6837 21539
rect 6696 21508 6837 21536
rect 6696 21496 6702 21508
rect 6825 21505 6837 21508
rect 6871 21505 6883 21539
rect 6825 21499 6883 21505
rect 9309 21539 9367 21545
rect 9309 21505 9321 21539
rect 9355 21505 9367 21539
rect 12268 21536 12296 21632
rect 15856 21604 15884 21644
rect 17218 21632 17224 21644
rect 17276 21632 17282 21684
rect 21174 21672 21180 21684
rect 21135 21644 21180 21672
rect 21174 21632 21180 21644
rect 21232 21632 21238 21684
rect 22186 21672 22192 21684
rect 22147 21644 22192 21672
rect 22186 21632 22192 21644
rect 22244 21632 22250 21684
rect 23290 21632 23296 21684
rect 23348 21672 23354 21684
rect 23385 21675 23443 21681
rect 23385 21672 23397 21675
rect 23348 21644 23397 21672
rect 23348 21632 23354 21644
rect 23385 21641 23397 21644
rect 23431 21641 23443 21675
rect 23385 21635 23443 21641
rect 23750 21632 23756 21684
rect 23808 21672 23814 21684
rect 24210 21672 24216 21684
rect 23808 21644 24216 21672
rect 23808 21632 23814 21644
rect 24210 21632 24216 21644
rect 24268 21632 24274 21684
rect 25406 21672 25412 21684
rect 25367 21644 25412 21672
rect 25406 21632 25412 21644
rect 25464 21632 25470 21684
rect 17034 21604 17040 21616
rect 15856 21576 17040 21604
rect 17034 21564 17040 21576
rect 17092 21604 17098 21616
rect 17773 21607 17831 21613
rect 17773 21604 17785 21607
rect 17092 21576 17785 21604
rect 17092 21564 17098 21576
rect 17773 21573 17785 21576
rect 17819 21604 17831 21607
rect 18322 21604 18328 21616
rect 17819 21576 18328 21604
rect 17819 21573 17831 21576
rect 17773 21567 17831 21573
rect 18322 21564 18328 21576
rect 18380 21564 18386 21616
rect 19613 21607 19671 21613
rect 19613 21573 19625 21607
rect 19659 21604 19671 21607
rect 19978 21604 19984 21616
rect 19659 21576 19984 21604
rect 19659 21573 19671 21576
rect 19613 21567 19671 21573
rect 19978 21564 19984 21576
rect 20036 21564 20042 21616
rect 21450 21604 21456 21616
rect 20088 21576 21456 21604
rect 12897 21539 12955 21545
rect 12897 21536 12909 21539
rect 12268 21508 12909 21536
rect 9309 21499 9367 21505
rect 12897 21505 12909 21508
rect 12943 21505 12955 21539
rect 12897 21499 12955 21505
rect 12989 21539 13047 21545
rect 12989 21505 13001 21539
rect 13035 21505 13047 21539
rect 12989 21499 13047 21505
rect 4203 21440 4844 21468
rect 4203 21437 4215 21440
rect 4157 21431 4215 21437
rect 4982 21428 4988 21480
rect 5040 21468 5046 21480
rect 5997 21471 6055 21477
rect 5997 21468 6009 21471
rect 5040 21440 6009 21468
rect 5040 21428 5046 21440
rect 5997 21437 6009 21440
rect 6043 21437 6055 21471
rect 5997 21431 6055 21437
rect 6914 21428 6920 21480
rect 6972 21468 6978 21480
rect 7092 21471 7150 21477
rect 7092 21468 7104 21471
rect 6972 21440 7104 21468
rect 6972 21428 6978 21440
rect 7092 21437 7104 21440
rect 7138 21468 7150 21471
rect 8386 21468 8392 21480
rect 7138 21440 8392 21468
rect 7138 21437 7150 21440
rect 7092 21431 7150 21437
rect 8386 21428 8392 21440
rect 8444 21428 8450 21480
rect 9030 21428 9036 21480
rect 9088 21468 9094 21480
rect 9214 21468 9220 21480
rect 9088 21440 9220 21468
rect 9088 21428 9094 21440
rect 9214 21428 9220 21440
rect 9272 21468 9278 21480
rect 9565 21471 9623 21477
rect 9565 21468 9577 21471
rect 9272 21440 9577 21468
rect 9272 21428 9278 21440
rect 9565 21437 9577 21440
rect 9611 21437 9623 21471
rect 13004 21468 13032 21499
rect 13814 21496 13820 21548
rect 13872 21536 13878 21548
rect 14918 21536 14924 21548
rect 13872 21508 14924 21536
rect 13872 21496 13878 21508
rect 14918 21496 14924 21508
rect 14976 21496 14982 21548
rect 16114 21496 16120 21548
rect 16172 21496 16178 21548
rect 18598 21536 18604 21548
rect 18559 21508 18604 21536
rect 18598 21496 18604 21508
rect 18656 21536 18662 21548
rect 19426 21536 19432 21548
rect 18656 21508 19432 21536
rect 18656 21496 18662 21508
rect 19426 21496 19432 21508
rect 19484 21496 19490 21548
rect 20088 21545 20116 21576
rect 21450 21564 21456 21576
rect 21508 21604 21514 21616
rect 21508 21576 25268 21604
rect 21508 21564 21514 21576
rect 19521 21539 19579 21545
rect 19521 21505 19533 21539
rect 19567 21536 19579 21539
rect 20073 21539 20131 21545
rect 20073 21536 20085 21539
rect 19567 21508 20085 21536
rect 19567 21505 19579 21508
rect 19521 21499 19579 21505
rect 20073 21505 20085 21508
rect 20119 21505 20131 21539
rect 20073 21499 20131 21505
rect 20257 21539 20315 21545
rect 20257 21505 20269 21539
rect 20303 21536 20315 21539
rect 20530 21536 20536 21548
rect 20303 21508 20536 21536
rect 20303 21505 20315 21508
rect 20257 21499 20315 21505
rect 20530 21496 20536 21508
rect 20588 21496 20594 21548
rect 20714 21536 20720 21548
rect 20675 21508 20720 21536
rect 20714 21496 20720 21508
rect 20772 21496 20778 21548
rect 21818 21536 21824 21548
rect 21779 21508 21824 21536
rect 21818 21496 21824 21508
rect 21876 21496 21882 21548
rect 23934 21496 23940 21548
rect 23992 21536 23998 21548
rect 24213 21539 24271 21545
rect 24213 21536 24225 21539
rect 23992 21508 24225 21536
rect 23992 21496 23998 21508
rect 24213 21505 24225 21508
rect 24259 21505 24271 21539
rect 24213 21499 24271 21505
rect 9565 21431 9623 21437
rect 11808 21440 13032 21468
rect 1670 21400 1676 21412
rect 1631 21372 1676 21400
rect 1670 21360 1676 21372
rect 1728 21360 1734 21412
rect 2593 21403 2651 21409
rect 2593 21369 2605 21403
rect 2639 21400 2651 21403
rect 3145 21403 3203 21409
rect 3145 21400 3157 21403
rect 2639 21372 3157 21400
rect 2639 21369 2651 21372
rect 2593 21363 2651 21369
rect 3145 21369 3157 21372
rect 3191 21400 3203 21403
rect 3234 21400 3240 21412
rect 3191 21372 3240 21400
rect 3191 21369 3203 21372
rect 3145 21363 3203 21369
rect 3234 21360 3240 21372
rect 3292 21360 3298 21412
rect 6641 21403 6699 21409
rect 6641 21369 6653 21403
rect 6687 21400 6699 21403
rect 7282 21400 7288 21412
rect 6687 21372 7288 21400
rect 6687 21369 6699 21372
rect 6641 21363 6699 21369
rect 7282 21360 7288 21372
rect 7340 21360 7346 21412
rect 8662 21360 8668 21412
rect 8720 21400 8726 21412
rect 9125 21403 9183 21409
rect 9125 21400 9137 21403
rect 8720 21372 9137 21400
rect 8720 21360 8726 21372
rect 9125 21369 9137 21372
rect 9171 21369 9183 21403
rect 9125 21363 9183 21369
rect 10594 21360 10600 21412
rect 10652 21400 10658 21412
rect 10962 21400 10968 21412
rect 10652 21372 10968 21400
rect 10652 21360 10658 21372
rect 10962 21360 10968 21372
rect 11020 21360 11026 21412
rect 2866 21292 2872 21344
rect 2924 21332 2930 21344
rect 3053 21335 3111 21341
rect 3053 21332 3065 21335
rect 2924 21304 3065 21332
rect 2924 21292 2930 21304
rect 3053 21301 3065 21304
rect 3099 21301 3111 21335
rect 3053 21295 3111 21301
rect 4154 21292 4160 21344
rect 4212 21332 4218 21344
rect 4617 21335 4675 21341
rect 4617 21332 4629 21335
rect 4212 21304 4629 21332
rect 4212 21292 4218 21304
rect 4617 21301 4629 21304
rect 4663 21301 4675 21335
rect 4617 21295 4675 21301
rect 5353 21335 5411 21341
rect 5353 21301 5365 21335
rect 5399 21332 5411 21335
rect 5442 21332 5448 21344
rect 5399 21304 5448 21332
rect 5399 21301 5411 21304
rect 5353 21295 5411 21301
rect 5442 21292 5448 21304
rect 5500 21292 5506 21344
rect 8846 21332 8852 21344
rect 8807 21304 8852 21332
rect 8846 21292 8852 21304
rect 8904 21292 8910 21344
rect 11238 21292 11244 21344
rect 11296 21332 11302 21344
rect 11333 21335 11391 21341
rect 11333 21332 11345 21335
rect 11296 21304 11345 21332
rect 11296 21292 11302 21304
rect 11333 21301 11345 21304
rect 11379 21332 11391 21335
rect 11422 21332 11428 21344
rect 11379 21304 11428 21332
rect 11379 21301 11391 21304
rect 11333 21295 11391 21301
rect 11422 21292 11428 21304
rect 11480 21332 11486 21344
rect 11808 21341 11836 21440
rect 13725 21403 13783 21409
rect 13725 21369 13737 21403
rect 13771 21400 13783 21403
rect 14090 21400 14096 21412
rect 13771 21372 14096 21400
rect 13771 21369 13783 21372
rect 13725 21363 13783 21369
rect 14090 21360 14096 21372
rect 14148 21400 14154 21412
rect 14829 21403 14887 21409
rect 14829 21400 14841 21403
rect 14148 21372 14841 21400
rect 14148 21360 14154 21372
rect 14829 21369 14841 21372
rect 14875 21400 14887 21403
rect 15188 21403 15246 21409
rect 15188 21400 15200 21403
rect 14875 21372 15200 21400
rect 14875 21369 14887 21372
rect 14829 21363 14887 21369
rect 15188 21369 15200 21372
rect 15234 21400 15246 21403
rect 15378 21400 15384 21412
rect 15234 21372 15384 21400
rect 15234 21369 15246 21372
rect 15188 21363 15246 21369
rect 15378 21360 15384 21372
rect 15436 21360 15442 21412
rect 16132 21344 16160 21496
rect 20732 21468 20760 21496
rect 21545 21471 21603 21477
rect 21545 21468 21557 21471
rect 20732 21440 21557 21468
rect 21545 21437 21557 21440
rect 21591 21437 21603 21471
rect 21545 21431 21603 21437
rect 23109 21471 23167 21477
rect 23109 21437 23121 21471
rect 23155 21468 23167 21471
rect 23566 21468 23572 21480
rect 23155 21440 23572 21468
rect 23155 21437 23167 21440
rect 23109 21431 23167 21437
rect 23566 21428 23572 21440
rect 23624 21468 23630 21480
rect 25240 21477 25268 21576
rect 24121 21471 24179 21477
rect 24121 21468 24133 21471
rect 23624 21440 24133 21468
rect 23624 21428 23630 21440
rect 24121 21437 24133 21440
rect 24167 21437 24179 21471
rect 24121 21431 24179 21437
rect 25225 21471 25283 21477
rect 25225 21437 25237 21471
rect 25271 21468 25283 21471
rect 25777 21471 25835 21477
rect 25777 21468 25789 21471
rect 25271 21440 25789 21468
rect 25271 21437 25283 21440
rect 25225 21431 25283 21437
rect 25777 21437 25789 21440
rect 25823 21437 25835 21471
rect 25777 21431 25835 21437
rect 17954 21360 17960 21412
rect 18012 21400 18018 21412
rect 18509 21403 18567 21409
rect 18509 21400 18521 21403
rect 18012 21372 18521 21400
rect 18012 21360 18018 21372
rect 18509 21369 18521 21372
rect 18555 21369 18567 21403
rect 18509 21363 18567 21369
rect 23290 21360 23296 21412
rect 23348 21400 23354 21412
rect 24029 21403 24087 21409
rect 24029 21400 24041 21403
rect 23348 21372 24041 21400
rect 23348 21360 23354 21372
rect 24029 21369 24041 21372
rect 24075 21400 24087 21403
rect 25041 21403 25099 21409
rect 25041 21400 25053 21403
rect 24075 21372 25053 21400
rect 24075 21369 24087 21372
rect 24029 21363 24087 21369
rect 25041 21369 25053 21372
rect 25087 21369 25099 21403
rect 25041 21363 25099 21369
rect 11793 21335 11851 21341
rect 11793 21332 11805 21335
rect 11480 21304 11805 21332
rect 11480 21292 11486 21304
rect 11793 21301 11805 21304
rect 11839 21301 11851 21335
rect 11793 21295 11851 21301
rect 12434 21292 12440 21344
rect 12492 21332 12498 21344
rect 12805 21335 12863 21341
rect 12805 21332 12817 21335
rect 12492 21304 12817 21332
rect 12492 21292 12498 21304
rect 12805 21301 12817 21304
rect 12851 21301 12863 21335
rect 12805 21295 12863 21301
rect 13354 21292 13360 21344
rect 13412 21332 13418 21344
rect 13814 21332 13820 21344
rect 13412 21304 13820 21332
rect 13412 21292 13418 21304
rect 13814 21292 13820 21304
rect 13872 21292 13878 21344
rect 14461 21335 14519 21341
rect 14461 21301 14473 21335
rect 14507 21332 14519 21335
rect 14642 21332 14648 21344
rect 14507 21304 14648 21332
rect 14507 21301 14519 21304
rect 14461 21295 14519 21301
rect 14642 21292 14648 21304
rect 14700 21292 14706 21344
rect 16114 21292 16120 21344
rect 16172 21292 16178 21344
rect 16298 21332 16304 21344
rect 16259 21304 16304 21332
rect 16298 21292 16304 21304
rect 16356 21292 16362 21344
rect 16942 21332 16948 21344
rect 16903 21304 16948 21332
rect 16942 21292 16948 21304
rect 17000 21292 17006 21344
rect 18046 21332 18052 21344
rect 18007 21304 18052 21332
rect 18046 21292 18052 21304
rect 18104 21292 18110 21344
rect 18322 21292 18328 21344
rect 18380 21332 18386 21344
rect 18417 21335 18475 21341
rect 18417 21332 18429 21335
rect 18380 21304 18429 21332
rect 18380 21292 18386 21304
rect 18417 21301 18429 21304
rect 18463 21301 18475 21335
rect 19058 21332 19064 21344
rect 19019 21304 19064 21332
rect 18417 21295 18475 21301
rect 19058 21292 19064 21304
rect 19116 21292 19122 21344
rect 19518 21292 19524 21344
rect 19576 21332 19582 21344
rect 19981 21335 20039 21341
rect 19981 21332 19993 21335
rect 19576 21304 19993 21332
rect 19576 21292 19582 21304
rect 19981 21301 19993 21304
rect 20027 21301 20039 21335
rect 19981 21295 20039 21301
rect 20898 21292 20904 21344
rect 20956 21332 20962 21344
rect 21085 21335 21143 21341
rect 21085 21332 21097 21335
rect 20956 21304 21097 21332
rect 20956 21292 20962 21304
rect 21085 21301 21097 21304
rect 21131 21332 21143 21335
rect 21637 21335 21695 21341
rect 21637 21332 21649 21335
rect 21131 21304 21649 21332
rect 21131 21301 21143 21304
rect 21085 21295 21143 21301
rect 21637 21301 21649 21304
rect 21683 21301 21695 21335
rect 21637 21295 21695 21301
rect 22278 21292 22284 21344
rect 22336 21332 22342 21344
rect 22557 21335 22615 21341
rect 22557 21332 22569 21335
rect 22336 21304 22569 21332
rect 22336 21292 22342 21304
rect 22557 21301 22569 21304
rect 22603 21301 22615 21335
rect 23658 21332 23664 21344
rect 23619 21304 23664 21332
rect 22557 21295 22615 21301
rect 23658 21292 23664 21304
rect 23716 21292 23722 21344
rect 24762 21332 24768 21344
rect 24675 21304 24768 21332
rect 24762 21292 24768 21304
rect 24820 21332 24826 21344
rect 25866 21332 25872 21344
rect 24820 21304 25872 21332
rect 24820 21292 24826 21304
rect 25866 21292 25872 21304
rect 25924 21292 25930 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 2406 21128 2412 21140
rect 2367 21100 2412 21128
rect 2406 21088 2412 21100
rect 2464 21088 2470 21140
rect 6914 21128 6920 21140
rect 6875 21100 6920 21128
rect 6914 21088 6920 21100
rect 6972 21088 6978 21140
rect 8021 21131 8079 21137
rect 8021 21097 8033 21131
rect 8067 21128 8079 21131
rect 8202 21128 8208 21140
rect 8067 21100 8208 21128
rect 8067 21097 8079 21100
rect 8021 21091 8079 21097
rect 8202 21088 8208 21100
rect 8260 21088 8266 21140
rect 13722 21128 13728 21140
rect 12728 21100 13728 21128
rect 1762 21020 1768 21072
rect 1820 21060 1826 21072
rect 2682 21060 2688 21072
rect 1820 21032 2688 21060
rect 1820 21020 1826 21032
rect 2682 21020 2688 21032
rect 2740 21060 2746 21072
rect 2869 21063 2927 21069
rect 2869 21060 2881 21063
rect 2740 21032 2881 21060
rect 2740 21020 2746 21032
rect 2869 21029 2881 21032
rect 2915 21060 2927 21063
rect 4246 21060 4252 21072
rect 2915 21032 4252 21060
rect 2915 21029 2927 21032
rect 2869 21023 2927 21029
rect 4246 21020 4252 21032
rect 4304 21020 4310 21072
rect 5068 21063 5126 21069
rect 5068 21029 5080 21063
rect 5114 21060 5126 21063
rect 5166 21060 5172 21072
rect 5114 21032 5172 21060
rect 5114 21029 5126 21032
rect 5068 21023 5126 21029
rect 5166 21020 5172 21032
rect 5224 21020 5230 21072
rect 8754 21020 8760 21072
rect 8812 21060 8818 21072
rect 9214 21060 9220 21072
rect 8812 21032 9220 21060
rect 8812 21020 8818 21032
rect 9214 21020 9220 21032
rect 9272 21020 9278 21072
rect 2777 20995 2835 21001
rect 2777 20961 2789 20995
rect 2823 20992 2835 20995
rect 2958 20992 2964 21004
rect 2823 20964 2964 20992
rect 2823 20961 2835 20964
rect 2777 20955 2835 20961
rect 2958 20952 2964 20964
rect 3016 20952 3022 21004
rect 4801 20995 4859 21001
rect 4801 20961 4813 20995
rect 4847 20992 4859 20995
rect 4890 20992 4896 21004
rect 4847 20964 4896 20992
rect 4847 20961 4859 20964
rect 4801 20955 4859 20961
rect 4890 20952 4896 20964
rect 4948 20952 4954 21004
rect 7561 20995 7619 21001
rect 7561 20961 7573 20995
rect 7607 20992 7619 20995
rect 8294 20992 8300 21004
rect 7607 20964 8300 20992
rect 7607 20961 7619 20964
rect 7561 20955 7619 20961
rect 8294 20952 8300 20964
rect 8352 20992 8358 21004
rect 8389 20995 8447 21001
rect 8389 20992 8401 20995
rect 8352 20964 8401 20992
rect 8352 20952 8358 20964
rect 8389 20961 8401 20964
rect 8435 20961 8447 20995
rect 8389 20955 8447 20961
rect 8481 20995 8539 21001
rect 8481 20961 8493 20995
rect 8527 20992 8539 20995
rect 9582 20992 9588 21004
rect 8527 20964 9588 20992
rect 8527 20961 8539 20964
rect 8481 20955 8539 20961
rect 2041 20927 2099 20933
rect 2041 20893 2053 20927
rect 2087 20924 2099 20927
rect 3050 20924 3056 20936
rect 2087 20896 3056 20924
rect 2087 20893 2099 20896
rect 2041 20887 2099 20893
rect 3050 20884 3056 20896
rect 3108 20884 3114 20936
rect 7929 20927 7987 20933
rect 7929 20893 7941 20927
rect 7975 20924 7987 20927
rect 8496 20924 8524 20955
rect 9582 20952 9588 20964
rect 9640 20952 9646 21004
rect 9674 20952 9680 21004
rect 9732 20992 9738 21004
rect 9950 21001 9956 21004
rect 9944 20992 9956 21001
rect 9732 20964 9777 20992
rect 9911 20964 9956 20992
rect 9732 20952 9738 20964
rect 9944 20955 9956 20964
rect 9950 20952 9956 20955
rect 10008 20952 10014 21004
rect 12728 21001 12756 21100
rect 13722 21088 13728 21100
rect 13780 21088 13786 21140
rect 14090 21128 14096 21140
rect 14051 21100 14096 21128
rect 14090 21088 14096 21100
rect 14148 21088 14154 21140
rect 14734 21128 14740 21140
rect 14695 21100 14740 21128
rect 14734 21088 14740 21100
rect 14792 21088 14798 21140
rect 16574 21088 16580 21140
rect 16632 21128 16638 21140
rect 17221 21131 17279 21137
rect 17221 21128 17233 21131
rect 16632 21100 17233 21128
rect 16632 21088 16638 21100
rect 17221 21097 17233 21100
rect 17267 21097 17279 21131
rect 17221 21091 17279 21097
rect 18598 21088 18604 21140
rect 18656 21128 18662 21140
rect 18785 21131 18843 21137
rect 18785 21128 18797 21131
rect 18656 21100 18797 21128
rect 18656 21088 18662 21100
rect 18785 21097 18797 21100
rect 18831 21097 18843 21131
rect 18785 21091 18843 21097
rect 19426 21088 19432 21140
rect 19484 21128 19490 21140
rect 19981 21131 20039 21137
rect 19981 21128 19993 21131
rect 19484 21100 19993 21128
rect 19484 21088 19490 21100
rect 19981 21097 19993 21100
rect 20027 21128 20039 21131
rect 20806 21128 20812 21140
rect 20027 21100 20812 21128
rect 20027 21097 20039 21100
rect 19981 21091 20039 21097
rect 20806 21088 20812 21100
rect 20864 21088 20870 21140
rect 23290 21128 23296 21140
rect 23251 21100 23296 21128
rect 23290 21088 23296 21100
rect 23348 21088 23354 21140
rect 23382 21088 23388 21140
rect 23440 21128 23446 21140
rect 24305 21131 24363 21137
rect 24305 21128 24317 21131
rect 23440 21100 24317 21128
rect 23440 21088 23446 21100
rect 24305 21097 24317 21100
rect 24351 21128 24363 21131
rect 24351 21100 24808 21128
rect 24351 21097 24363 21100
rect 24305 21091 24363 21097
rect 14182 21060 14188 21072
rect 12820 21032 14188 21060
rect 11793 20995 11851 21001
rect 11793 20961 11805 20995
rect 11839 20992 11851 20995
rect 12713 20995 12771 21001
rect 11839 20964 12664 20992
rect 11839 20961 11851 20964
rect 11793 20955 11851 20961
rect 7975 20896 8524 20924
rect 8665 20927 8723 20933
rect 7975 20893 7987 20896
rect 7929 20887 7987 20893
rect 8665 20893 8677 20927
rect 8711 20924 8723 20927
rect 8754 20924 8760 20936
rect 8711 20896 8760 20924
rect 8711 20893 8723 20896
rect 8665 20887 8723 20893
rect 8754 20884 8760 20896
rect 8812 20924 8818 20936
rect 9030 20924 9036 20936
rect 8812 20896 9036 20924
rect 8812 20884 8818 20896
rect 9030 20884 9036 20896
rect 9088 20924 9094 20936
rect 9309 20927 9367 20933
rect 9309 20924 9321 20927
rect 9088 20896 9321 20924
rect 9088 20884 9094 20896
rect 9309 20893 9321 20896
rect 9355 20893 9367 20927
rect 12158 20924 12164 20936
rect 12119 20896 12164 20924
rect 9309 20887 9367 20893
rect 12158 20884 12164 20896
rect 12216 20884 12222 20936
rect 12636 20924 12664 20964
rect 12713 20961 12725 20995
rect 12759 20961 12771 20995
rect 12713 20955 12771 20961
rect 12820 20924 12848 21032
rect 14182 21020 14188 21032
rect 14240 21020 14246 21072
rect 15378 21020 15384 21072
rect 15436 21060 15442 21072
rect 15565 21063 15623 21069
rect 15565 21060 15577 21063
rect 15436 21032 15577 21060
rect 15436 21020 15442 21032
rect 15565 21029 15577 21032
rect 15611 21060 15623 21063
rect 16108 21063 16166 21069
rect 16108 21060 16120 21063
rect 15611 21032 16120 21060
rect 15611 21029 15623 21032
rect 15565 21023 15623 21029
rect 16108 21029 16120 21032
rect 16154 21060 16166 21063
rect 16298 21060 16304 21072
rect 16154 21032 16304 21060
rect 16154 21029 16166 21032
rect 16108 21023 16166 21029
rect 16298 21020 16304 21032
rect 16356 21020 16362 21072
rect 21174 21020 21180 21072
rect 21232 21060 21238 21072
rect 21361 21063 21419 21069
rect 21361 21060 21373 21063
rect 21232 21032 21373 21060
rect 21232 21020 21238 21032
rect 21361 21029 21373 21032
rect 21407 21060 21419 21063
rect 24673 21063 24731 21069
rect 24673 21060 24685 21063
rect 21407 21032 24685 21060
rect 21407 21029 21419 21032
rect 21361 21023 21419 21029
rect 24673 21029 24685 21032
rect 24719 21029 24731 21063
rect 24780 21060 24808 21100
rect 24854 21088 24860 21140
rect 24912 21128 24918 21140
rect 25225 21131 25283 21137
rect 25225 21128 25237 21131
rect 24912 21100 25237 21128
rect 24912 21088 24918 21100
rect 25225 21097 25237 21100
rect 25271 21128 25283 21131
rect 25406 21128 25412 21140
rect 25271 21100 25412 21128
rect 25271 21097 25283 21100
rect 25225 21091 25283 21097
rect 25406 21088 25412 21100
rect 25464 21088 25470 21140
rect 24946 21060 24952 21072
rect 24780 21032 24952 21060
rect 24673 21023 24731 21029
rect 24946 21020 24952 21032
rect 25004 21020 25010 21072
rect 25314 21020 25320 21072
rect 25372 21020 25378 21072
rect 12980 20995 13038 21001
rect 12980 20961 12992 20995
rect 13026 20992 13038 20995
rect 13538 20992 13544 21004
rect 13026 20964 13544 20992
rect 13026 20961 13038 20964
rect 12980 20955 13038 20961
rect 13538 20952 13544 20964
rect 13596 20952 13602 21004
rect 14090 20952 14096 21004
rect 14148 20992 14154 21004
rect 16942 20992 16948 21004
rect 14148 20964 16948 20992
rect 14148 20952 14154 20964
rect 16942 20952 16948 20964
rect 17000 20952 17006 21004
rect 18598 20952 18604 21004
rect 18656 20992 18662 21004
rect 18693 20995 18751 21001
rect 18693 20992 18705 20995
rect 18656 20964 18705 20992
rect 18656 20952 18662 20964
rect 18693 20961 18705 20964
rect 18739 20961 18751 20995
rect 18693 20955 18751 20961
rect 20714 20952 20720 21004
rect 20772 20992 20778 21004
rect 21269 20995 21327 21001
rect 21269 20992 21281 20995
rect 20772 20964 21281 20992
rect 20772 20952 20778 20964
rect 21269 20961 21281 20964
rect 21315 20961 21327 20995
rect 21269 20955 21327 20961
rect 21818 20952 21824 21004
rect 21876 20992 21882 21004
rect 22005 20995 22063 21001
rect 22005 20992 22017 20995
rect 21876 20964 22017 20992
rect 21876 20952 21882 20964
rect 22005 20961 22017 20964
rect 22051 20992 22063 20995
rect 23106 20992 23112 21004
rect 22051 20964 23112 20992
rect 22051 20961 22063 20964
rect 22005 20955 22063 20961
rect 23106 20952 23112 20964
rect 23164 20952 23170 21004
rect 23201 20995 23259 21001
rect 23201 20961 23213 20995
rect 23247 20992 23259 20995
rect 23658 20992 23664 21004
rect 23247 20964 23664 20992
rect 23247 20961 23259 20964
rect 23201 20955 23259 20961
rect 23658 20952 23664 20964
rect 23716 20952 23722 21004
rect 25332 20992 25360 21020
rect 25332 20964 25452 20992
rect 12636 20896 12848 20924
rect 14918 20884 14924 20936
rect 14976 20924 14982 20936
rect 15841 20927 15899 20933
rect 15841 20924 15853 20927
rect 14976 20896 15853 20924
rect 14976 20884 14982 20896
rect 15841 20893 15853 20896
rect 15887 20893 15899 20927
rect 18966 20924 18972 20936
rect 18927 20896 18972 20924
rect 15841 20887 15899 20893
rect 18966 20884 18972 20896
rect 19024 20884 19030 20936
rect 20990 20884 20996 20936
rect 21048 20924 21054 20936
rect 21453 20927 21511 20933
rect 21453 20924 21465 20927
rect 21048 20896 21465 20924
rect 21048 20884 21054 20896
rect 21453 20893 21465 20896
rect 21499 20893 21511 20927
rect 21453 20887 21511 20893
rect 23474 20884 23480 20936
rect 23532 20924 23538 20936
rect 23753 20927 23811 20933
rect 23753 20924 23765 20927
rect 23532 20896 23765 20924
rect 23532 20884 23538 20896
rect 23753 20893 23765 20896
rect 23799 20893 23811 20927
rect 23753 20887 23811 20893
rect 23937 20927 23995 20933
rect 23937 20893 23949 20927
rect 23983 20924 23995 20927
rect 24670 20924 24676 20936
rect 23983 20896 24676 20924
rect 23983 20893 23995 20896
rect 23937 20887 23995 20893
rect 24670 20884 24676 20896
rect 24728 20884 24734 20936
rect 25038 20884 25044 20936
rect 25096 20924 25102 20936
rect 25424 20933 25452 20964
rect 25317 20927 25375 20933
rect 25317 20924 25329 20927
rect 25096 20896 25329 20924
rect 25096 20884 25102 20896
rect 25317 20893 25329 20896
rect 25363 20893 25375 20927
rect 25317 20887 25375 20893
rect 25409 20927 25467 20933
rect 25409 20893 25421 20927
rect 25455 20893 25467 20927
rect 25409 20887 25467 20893
rect 11054 20856 11060 20868
rect 11015 20828 11060 20856
rect 11054 20816 11060 20828
rect 11112 20816 11118 20868
rect 14182 20816 14188 20868
rect 14240 20856 14246 20868
rect 18325 20859 18383 20865
rect 18325 20856 18337 20859
rect 14240 20828 15691 20856
rect 14240 20816 14246 20828
rect 1486 20748 1492 20800
rect 1544 20788 1550 20800
rect 1581 20791 1639 20797
rect 1581 20788 1593 20791
rect 1544 20760 1593 20788
rect 1544 20748 1550 20760
rect 1581 20757 1593 20760
rect 1627 20757 1639 20791
rect 3694 20788 3700 20800
rect 3655 20760 3700 20788
rect 1581 20751 1639 20757
rect 3694 20748 3700 20760
rect 3752 20748 3758 20800
rect 4246 20788 4252 20800
rect 4207 20760 4252 20788
rect 4246 20748 4252 20760
rect 4304 20748 4310 20800
rect 4338 20748 4344 20800
rect 4396 20788 4402 20800
rect 4617 20791 4675 20797
rect 4617 20788 4629 20791
rect 4396 20760 4629 20788
rect 4396 20748 4402 20760
rect 4617 20757 4629 20760
rect 4663 20757 4675 20791
rect 4617 20751 4675 20757
rect 5442 20748 5448 20800
rect 5500 20788 5506 20800
rect 6181 20791 6239 20797
rect 6181 20788 6193 20791
rect 5500 20760 6193 20788
rect 5500 20748 5506 20760
rect 6181 20757 6193 20760
rect 6227 20788 6239 20791
rect 6822 20788 6828 20800
rect 6227 20760 6828 20788
rect 6227 20757 6239 20760
rect 6181 20751 6239 20757
rect 6822 20748 6828 20760
rect 6880 20748 6886 20800
rect 12434 20748 12440 20800
rect 12492 20788 12498 20800
rect 12529 20791 12587 20797
rect 12529 20788 12541 20791
rect 12492 20760 12541 20788
rect 12492 20748 12498 20760
rect 12529 20757 12541 20760
rect 12575 20788 12587 20791
rect 13354 20788 13360 20800
rect 12575 20760 13360 20788
rect 12575 20757 12587 20760
rect 12529 20751 12587 20757
rect 13354 20748 13360 20760
rect 13412 20748 13418 20800
rect 15105 20791 15163 20797
rect 15105 20757 15117 20791
rect 15151 20788 15163 20791
rect 15562 20788 15568 20800
rect 15151 20760 15568 20788
rect 15151 20757 15163 20760
rect 15105 20751 15163 20757
rect 15562 20748 15568 20760
rect 15620 20748 15626 20800
rect 15663 20788 15691 20828
rect 16776 20828 18337 20856
rect 16776 20788 16804 20828
rect 18325 20825 18337 20828
rect 18371 20825 18383 20859
rect 20898 20856 20904 20868
rect 20859 20828 20904 20856
rect 18325 20819 18383 20825
rect 20898 20816 20904 20828
rect 20956 20816 20962 20868
rect 22373 20859 22431 20865
rect 22373 20825 22385 20859
rect 22419 20856 22431 20859
rect 22419 20828 23428 20856
rect 22419 20825 22431 20828
rect 22373 20819 22431 20825
rect 15663 20760 16804 20788
rect 18141 20791 18199 20797
rect 18141 20757 18153 20791
rect 18187 20788 18199 20791
rect 18506 20788 18512 20800
rect 18187 20760 18512 20788
rect 18187 20757 18199 20760
rect 18141 20751 18199 20757
rect 18506 20748 18512 20760
rect 18564 20748 18570 20800
rect 19610 20788 19616 20800
rect 19571 20760 19616 20788
rect 19610 20748 19616 20760
rect 19668 20748 19674 20800
rect 19702 20748 19708 20800
rect 19760 20788 19766 20800
rect 20346 20788 20352 20800
rect 19760 20760 20352 20788
rect 19760 20748 19766 20760
rect 20346 20748 20352 20760
rect 20404 20748 20410 20800
rect 20441 20791 20499 20797
rect 20441 20757 20453 20791
rect 20487 20788 20499 20791
rect 20530 20788 20536 20800
rect 20487 20760 20536 20788
rect 20487 20757 20499 20760
rect 20441 20751 20499 20757
rect 20530 20748 20536 20760
rect 20588 20748 20594 20800
rect 22094 20748 22100 20800
rect 22152 20788 22158 20800
rect 22388 20788 22416 20819
rect 22830 20788 22836 20800
rect 22152 20760 22416 20788
rect 22743 20760 22836 20788
rect 22152 20748 22158 20760
rect 22830 20748 22836 20760
rect 22888 20788 22894 20800
rect 23290 20788 23296 20800
rect 22888 20760 23296 20788
rect 22888 20748 22894 20760
rect 23290 20748 23296 20760
rect 23348 20748 23354 20800
rect 23400 20788 23428 20828
rect 23750 20788 23756 20800
rect 23400 20760 23756 20788
rect 23750 20748 23756 20760
rect 23808 20748 23814 20800
rect 24854 20788 24860 20800
rect 24815 20760 24860 20788
rect 24854 20748 24860 20760
rect 24912 20748 24918 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 2682 20584 2688 20596
rect 2643 20556 2688 20584
rect 2682 20544 2688 20556
rect 2740 20544 2746 20596
rect 2958 20584 2964 20596
rect 2919 20556 2964 20584
rect 2958 20544 2964 20556
rect 3016 20544 3022 20596
rect 3145 20587 3203 20593
rect 3145 20553 3157 20587
rect 3191 20584 3203 20587
rect 4154 20584 4160 20596
rect 3191 20556 4160 20584
rect 3191 20553 3203 20556
rect 3145 20547 3203 20553
rect 4154 20544 4160 20556
rect 4212 20544 4218 20596
rect 4706 20584 4712 20596
rect 4667 20556 4712 20584
rect 4706 20544 4712 20556
rect 4764 20544 4770 20596
rect 8294 20584 8300 20596
rect 8255 20556 8300 20584
rect 8294 20544 8300 20556
rect 8352 20544 8358 20596
rect 9674 20544 9680 20596
rect 9732 20584 9738 20596
rect 9861 20587 9919 20593
rect 9861 20584 9873 20587
rect 9732 20556 9873 20584
rect 9732 20544 9738 20556
rect 9861 20553 9873 20556
rect 9907 20553 9919 20587
rect 9861 20547 9919 20553
rect 10686 20544 10692 20596
rect 10744 20584 10750 20596
rect 10870 20584 10876 20596
rect 10744 20556 10876 20584
rect 10744 20544 10750 20556
rect 10870 20544 10876 20556
rect 10928 20544 10934 20596
rect 12434 20544 12440 20596
rect 12492 20584 12498 20596
rect 13538 20584 13544 20596
rect 12492 20556 12537 20584
rect 13499 20556 13544 20584
rect 12492 20544 12498 20556
rect 13538 20544 13544 20556
rect 13596 20544 13602 20596
rect 14645 20587 14703 20593
rect 14645 20553 14657 20587
rect 14691 20584 14703 20587
rect 15286 20584 15292 20596
rect 14691 20556 15292 20584
rect 14691 20553 14703 20556
rect 14645 20547 14703 20553
rect 15286 20544 15292 20556
rect 15344 20544 15350 20596
rect 15470 20544 15476 20596
rect 15528 20584 15534 20596
rect 16209 20587 16267 20593
rect 16209 20584 16221 20587
rect 15528 20556 16221 20584
rect 15528 20544 15534 20556
rect 16209 20553 16221 20556
rect 16255 20553 16267 20587
rect 18046 20584 18052 20596
rect 18007 20556 18052 20584
rect 16209 20547 16267 20553
rect 18046 20544 18052 20556
rect 18104 20544 18110 20596
rect 18966 20544 18972 20596
rect 19024 20584 19030 20596
rect 19061 20587 19119 20593
rect 19061 20584 19073 20587
rect 19024 20556 19073 20584
rect 19024 20544 19030 20556
rect 19061 20553 19073 20556
rect 19107 20553 19119 20587
rect 19061 20547 19119 20553
rect 19613 20587 19671 20593
rect 19613 20553 19625 20587
rect 19659 20584 19671 20587
rect 20714 20584 20720 20596
rect 19659 20556 20720 20584
rect 19659 20553 19671 20556
rect 19613 20547 19671 20553
rect 20714 20544 20720 20556
rect 20772 20544 20778 20596
rect 20990 20584 20996 20596
rect 20951 20556 20996 20584
rect 20990 20544 20996 20556
rect 21048 20544 21054 20596
rect 21174 20584 21180 20596
rect 21135 20556 21180 20584
rect 21174 20544 21180 20556
rect 21232 20544 21238 20596
rect 22649 20587 22707 20593
rect 22649 20553 22661 20587
rect 22695 20584 22707 20587
rect 22738 20584 22744 20596
rect 22695 20556 22744 20584
rect 22695 20553 22707 20556
rect 22649 20547 22707 20553
rect 22738 20544 22744 20556
rect 22796 20544 22802 20596
rect 23566 20544 23572 20596
rect 23624 20584 23630 20596
rect 23661 20587 23719 20593
rect 23661 20584 23673 20587
rect 23624 20556 23673 20584
rect 23624 20544 23630 20556
rect 23661 20553 23673 20556
rect 23707 20553 23719 20587
rect 23661 20547 23719 20553
rect 25130 20544 25136 20596
rect 25188 20584 25194 20596
rect 26234 20584 26240 20596
rect 25188 20556 26240 20584
rect 25188 20544 25194 20556
rect 26234 20544 26240 20556
rect 26292 20544 26298 20596
rect 1581 20519 1639 20525
rect 1581 20485 1593 20519
rect 1627 20516 1639 20519
rect 2774 20516 2780 20528
rect 1627 20488 2780 20516
rect 1627 20485 1639 20488
rect 1581 20479 1639 20485
rect 2774 20476 2780 20488
rect 2832 20476 2838 20528
rect 3050 20476 3056 20528
rect 3108 20516 3114 20528
rect 4249 20519 4307 20525
rect 4249 20516 4261 20519
rect 3108 20488 4261 20516
rect 3108 20476 3114 20488
rect 4249 20485 4261 20488
rect 4295 20516 4307 20519
rect 6546 20516 6552 20528
rect 4295 20488 6552 20516
rect 4295 20485 4307 20488
rect 4249 20479 4307 20485
rect 6546 20476 6552 20488
rect 6604 20476 6610 20528
rect 7006 20516 7012 20528
rect 6967 20488 7012 20516
rect 7006 20476 7012 20488
rect 7064 20476 7070 20528
rect 11514 20476 11520 20528
rect 11572 20516 11578 20528
rect 11698 20516 11704 20528
rect 11572 20488 11704 20516
rect 11572 20476 11578 20488
rect 11698 20476 11704 20488
rect 11756 20476 11762 20528
rect 17862 20476 17868 20528
rect 17920 20516 17926 20528
rect 19429 20519 19487 20525
rect 19429 20516 19441 20519
rect 17920 20488 19441 20516
rect 17920 20476 17926 20488
rect 2225 20451 2283 20457
rect 2225 20417 2237 20451
rect 2271 20448 2283 20451
rect 3068 20448 3096 20476
rect 2271 20420 3096 20448
rect 2271 20417 2283 20420
rect 2225 20411 2283 20417
rect 3510 20408 3516 20460
rect 3568 20448 3574 20460
rect 3605 20451 3663 20457
rect 3605 20448 3617 20451
rect 3568 20420 3617 20448
rect 3568 20408 3574 20420
rect 3605 20417 3617 20420
rect 3651 20417 3663 20451
rect 3605 20411 3663 20417
rect 3789 20451 3847 20457
rect 3789 20417 3801 20451
rect 3835 20448 3847 20451
rect 4154 20448 4160 20460
rect 3835 20420 4160 20448
rect 3835 20417 3847 20420
rect 3789 20411 3847 20417
rect 4154 20408 4160 20420
rect 4212 20408 4218 20460
rect 5074 20408 5080 20460
rect 5132 20448 5138 20460
rect 5169 20451 5227 20457
rect 5169 20448 5181 20451
rect 5132 20420 5181 20448
rect 5132 20408 5138 20420
rect 5169 20417 5181 20420
rect 5215 20417 5227 20451
rect 5169 20411 5227 20417
rect 5261 20451 5319 20457
rect 5261 20417 5273 20451
rect 5307 20417 5319 20451
rect 5261 20411 5319 20417
rect 7469 20451 7527 20457
rect 7469 20417 7481 20451
rect 7515 20448 7527 20451
rect 8849 20451 8907 20457
rect 8849 20448 8861 20451
rect 7515 20420 8861 20448
rect 7515 20417 7527 20420
rect 7469 20411 7527 20417
rect 8849 20417 8861 20420
rect 8895 20448 8907 20451
rect 9309 20451 9367 20457
rect 9309 20448 9321 20451
rect 8895 20420 9321 20448
rect 8895 20417 8907 20420
rect 8849 20411 8907 20417
rect 9309 20417 9321 20420
rect 9355 20448 9367 20451
rect 9950 20448 9956 20460
rect 9355 20420 9956 20448
rect 9355 20417 9367 20420
rect 9309 20411 9367 20417
rect 5276 20380 5304 20411
rect 9950 20408 9956 20420
rect 10008 20448 10014 20460
rect 10413 20451 10471 20457
rect 10413 20448 10425 20451
rect 10008 20420 10425 20448
rect 10008 20408 10014 20420
rect 10413 20417 10425 20420
rect 10459 20448 10471 20451
rect 10873 20451 10931 20457
rect 10873 20448 10885 20451
rect 10459 20420 10885 20448
rect 10459 20417 10471 20420
rect 10413 20411 10471 20417
rect 10873 20417 10885 20420
rect 10919 20448 10931 20451
rect 11974 20448 11980 20460
rect 10919 20420 11980 20448
rect 10919 20417 10931 20420
rect 10873 20411 10931 20417
rect 11974 20408 11980 20420
rect 12032 20448 12038 20460
rect 12161 20451 12219 20457
rect 12161 20448 12173 20451
rect 12032 20420 12173 20448
rect 12032 20408 12038 20420
rect 12161 20417 12173 20420
rect 12207 20448 12219 20451
rect 12989 20451 13047 20457
rect 12989 20448 13001 20451
rect 12207 20420 13001 20448
rect 12207 20417 12219 20420
rect 12161 20411 12219 20417
rect 12989 20417 13001 20420
rect 13035 20417 13047 20451
rect 12989 20411 13047 20417
rect 14553 20451 14611 20457
rect 14553 20417 14565 20451
rect 14599 20448 14611 20451
rect 14918 20448 14924 20460
rect 14599 20420 14924 20448
rect 14599 20417 14611 20420
rect 14553 20411 14611 20417
rect 14918 20408 14924 20420
rect 14976 20448 14982 20460
rect 15289 20451 15347 20457
rect 15289 20448 15301 20451
rect 14976 20420 15301 20448
rect 14976 20408 14982 20420
rect 15289 20417 15301 20420
rect 15335 20448 15347 20451
rect 15378 20448 15384 20460
rect 15335 20420 15384 20448
rect 15335 20417 15347 20420
rect 15289 20411 15347 20417
rect 15378 20408 15384 20420
rect 15436 20408 15442 20460
rect 16758 20448 16764 20460
rect 16719 20420 16764 20448
rect 16758 20408 16764 20420
rect 16816 20448 16822 20460
rect 17221 20451 17279 20457
rect 17221 20448 17233 20451
rect 16816 20420 17233 20448
rect 16816 20408 16822 20420
rect 17221 20417 17233 20420
rect 17267 20417 17279 20451
rect 18506 20448 18512 20460
rect 17221 20411 17279 20417
rect 18432 20420 18512 20448
rect 6825 20383 6883 20389
rect 6825 20380 6837 20383
rect 4540 20352 5304 20380
rect 6564 20352 6837 20380
rect 1762 20272 1768 20324
rect 1820 20312 1826 20324
rect 1946 20312 1952 20324
rect 1820 20284 1952 20312
rect 1820 20272 1826 20284
rect 1946 20272 1952 20284
rect 2004 20272 2010 20324
rect 3326 20272 3332 20324
rect 3384 20312 3390 20324
rect 3513 20315 3571 20321
rect 3513 20312 3525 20315
rect 3384 20284 3525 20312
rect 3384 20272 3390 20284
rect 3513 20281 3525 20284
rect 3559 20281 3571 20315
rect 3513 20275 3571 20281
rect 1486 20204 1492 20256
rect 1544 20244 1550 20256
rect 2041 20247 2099 20253
rect 2041 20244 2053 20247
rect 1544 20216 2053 20244
rect 1544 20204 1550 20216
rect 2041 20213 2053 20216
rect 2087 20213 2099 20247
rect 2041 20207 2099 20213
rect 4154 20204 4160 20256
rect 4212 20244 4218 20256
rect 4540 20253 4568 20352
rect 6564 20324 6592 20352
rect 6825 20349 6837 20352
rect 6871 20349 6883 20383
rect 6825 20343 6883 20349
rect 7098 20340 7104 20392
rect 7156 20380 7162 20392
rect 7558 20380 7564 20392
rect 7156 20352 7564 20380
rect 7156 20340 7162 20352
rect 7558 20340 7564 20352
rect 7616 20340 7622 20392
rect 10042 20340 10048 20392
rect 10100 20380 10106 20392
rect 10778 20380 10784 20392
rect 10100 20352 10784 20380
rect 10100 20340 10106 20352
rect 10778 20340 10784 20352
rect 10836 20340 10842 20392
rect 12802 20380 12808 20392
rect 12715 20352 12808 20380
rect 12802 20340 12808 20352
rect 12860 20380 12866 20392
rect 13817 20383 13875 20389
rect 13817 20380 13829 20383
rect 12860 20352 13829 20380
rect 12860 20340 12866 20352
rect 13817 20349 13829 20352
rect 13863 20349 13875 20383
rect 13817 20343 13875 20349
rect 14734 20340 14740 20392
rect 14792 20380 14798 20392
rect 15013 20383 15071 20389
rect 15013 20380 15025 20383
rect 14792 20352 15025 20380
rect 14792 20340 14798 20352
rect 15013 20349 15025 20352
rect 15059 20349 15071 20383
rect 15013 20343 15071 20349
rect 15841 20383 15899 20389
rect 15841 20349 15853 20383
rect 15887 20380 15899 20383
rect 16577 20383 16635 20389
rect 16577 20380 16589 20383
rect 15887 20352 16589 20380
rect 15887 20349 15899 20352
rect 15841 20343 15899 20349
rect 16577 20349 16589 20352
rect 16623 20380 16635 20383
rect 17402 20380 17408 20392
rect 16623 20352 17408 20380
rect 16623 20349 16635 20352
rect 16577 20343 16635 20349
rect 17402 20340 17408 20352
rect 17460 20340 17466 20392
rect 18432 20389 18460 20420
rect 18506 20408 18512 20420
rect 18564 20408 18570 20460
rect 18708 20457 18736 20488
rect 19429 20485 19441 20488
rect 19475 20485 19487 20519
rect 19429 20479 19487 20485
rect 23477 20519 23535 20525
rect 23477 20485 23489 20519
rect 23523 20516 23535 20519
rect 24670 20516 24676 20528
rect 23523 20488 24676 20516
rect 23523 20485 23535 20488
rect 23477 20479 23535 20485
rect 18693 20451 18751 20457
rect 18693 20417 18705 20451
rect 18739 20417 18751 20451
rect 18693 20411 18751 20417
rect 19334 20408 19340 20460
rect 19392 20448 19398 20460
rect 20073 20451 20131 20457
rect 20073 20448 20085 20451
rect 19392 20420 20085 20448
rect 19392 20408 19398 20420
rect 20073 20417 20085 20420
rect 20119 20417 20131 20451
rect 20073 20411 20131 20417
rect 20162 20408 20168 20460
rect 20220 20448 20226 20460
rect 21729 20451 21787 20457
rect 21729 20448 21741 20451
rect 20220 20420 21741 20448
rect 20220 20408 20226 20420
rect 21729 20417 21741 20420
rect 21775 20448 21787 20451
rect 22189 20451 22247 20457
rect 22189 20448 22201 20451
rect 21775 20420 22201 20448
rect 21775 20417 21787 20420
rect 21729 20411 21787 20417
rect 22189 20417 22201 20420
rect 22235 20417 22247 20451
rect 22189 20411 22247 20417
rect 23290 20408 23296 20460
rect 23348 20448 23354 20460
rect 24228 20457 24256 20488
rect 24670 20476 24676 20488
rect 24728 20476 24734 20528
rect 24949 20519 25007 20525
rect 24949 20485 24961 20519
rect 24995 20516 25007 20519
rect 25314 20516 25320 20528
rect 24995 20488 25320 20516
rect 24995 20485 25007 20488
rect 24949 20479 25007 20485
rect 24121 20451 24179 20457
rect 24121 20448 24133 20451
rect 23348 20420 24133 20448
rect 23348 20408 23354 20420
rect 24121 20417 24133 20420
rect 24167 20417 24179 20451
rect 24121 20411 24179 20417
rect 24213 20451 24271 20457
rect 24213 20417 24225 20451
rect 24259 20417 24271 20451
rect 24213 20411 24271 20417
rect 24578 20408 24584 20460
rect 24636 20448 24642 20460
rect 24964 20448 24992 20479
rect 25314 20476 25320 20488
rect 25372 20476 25378 20528
rect 25958 20516 25964 20528
rect 25919 20488 25964 20516
rect 25958 20476 25964 20488
rect 26016 20476 26022 20528
rect 24636 20420 24992 20448
rect 24636 20408 24642 20420
rect 18417 20383 18475 20389
rect 18417 20349 18429 20383
rect 18463 20349 18475 20383
rect 18417 20343 18475 20349
rect 21545 20383 21603 20389
rect 21545 20349 21557 20383
rect 21591 20380 21603 20383
rect 22002 20380 22008 20392
rect 21591 20352 22008 20380
rect 21591 20349 21603 20352
rect 21545 20343 21603 20349
rect 22002 20340 22008 20352
rect 22060 20340 22066 20392
rect 23017 20383 23075 20389
rect 23017 20349 23029 20383
rect 23063 20380 23075 20383
rect 24029 20383 24087 20389
rect 24029 20380 24041 20383
rect 23063 20352 24041 20380
rect 23063 20349 23075 20352
rect 23017 20343 23075 20349
rect 24029 20349 24041 20352
rect 24075 20380 24087 20383
rect 24762 20380 24768 20392
rect 24075 20352 24768 20380
rect 24075 20349 24087 20352
rect 24029 20343 24087 20349
rect 24762 20340 24768 20352
rect 24820 20340 24826 20392
rect 25222 20380 25228 20392
rect 25183 20352 25228 20380
rect 25222 20340 25228 20352
rect 25280 20340 25286 20392
rect 4798 20272 4804 20324
rect 4856 20312 4862 20324
rect 5077 20315 5135 20321
rect 5077 20312 5089 20315
rect 4856 20284 5089 20312
rect 4856 20272 4862 20284
rect 5077 20281 5089 20284
rect 5123 20281 5135 20315
rect 6546 20312 6552 20324
rect 6507 20284 6552 20312
rect 5077 20275 5135 20281
rect 6546 20272 6552 20284
rect 6604 20272 6610 20324
rect 7837 20315 7895 20321
rect 7837 20281 7849 20315
rect 7883 20312 7895 20315
rect 8665 20315 8723 20321
rect 8665 20312 8677 20315
rect 7883 20284 8677 20312
rect 7883 20281 7895 20284
rect 7837 20275 7895 20281
rect 8665 20281 8677 20284
rect 8711 20312 8723 20315
rect 8846 20312 8852 20324
rect 8711 20284 8852 20312
rect 8711 20281 8723 20284
rect 8665 20275 8723 20281
rect 8846 20272 8852 20284
rect 8904 20272 8910 20324
rect 10321 20315 10379 20321
rect 10321 20281 10333 20315
rect 10367 20312 10379 20315
rect 10686 20312 10692 20324
rect 10367 20284 10692 20312
rect 10367 20281 10379 20284
rect 10321 20275 10379 20281
rect 10686 20272 10692 20284
rect 10744 20312 10750 20324
rect 11241 20315 11299 20321
rect 11241 20312 11253 20315
rect 10744 20284 11253 20312
rect 10744 20272 10750 20284
rect 11241 20281 11253 20284
rect 11287 20281 11299 20315
rect 11241 20275 11299 20281
rect 11514 20272 11520 20324
rect 11572 20312 11578 20324
rect 11885 20315 11943 20321
rect 11885 20312 11897 20315
rect 11572 20284 11897 20312
rect 11572 20272 11578 20284
rect 11885 20281 11897 20284
rect 11931 20312 11943 20315
rect 12897 20315 12955 20321
rect 12897 20312 12909 20315
rect 11931 20284 12909 20312
rect 11931 20281 11943 20284
rect 11885 20275 11943 20281
rect 12897 20281 12909 20284
rect 12943 20281 12955 20315
rect 12897 20275 12955 20281
rect 14182 20272 14188 20324
rect 14240 20312 14246 20324
rect 15105 20315 15163 20321
rect 15105 20312 15117 20315
rect 14240 20284 15117 20312
rect 14240 20272 14246 20284
rect 15105 20281 15117 20284
rect 15151 20281 15163 20315
rect 15105 20275 15163 20281
rect 15286 20272 15292 20324
rect 15344 20312 15350 20324
rect 16025 20315 16083 20321
rect 16025 20312 16037 20315
rect 15344 20284 16037 20312
rect 15344 20272 15350 20284
rect 16025 20281 16037 20284
rect 16071 20312 16083 20315
rect 16669 20315 16727 20321
rect 16669 20312 16681 20315
rect 16071 20284 16681 20312
rect 16071 20281 16083 20284
rect 16025 20275 16083 20281
rect 16669 20281 16681 20284
rect 16715 20281 16727 20315
rect 18509 20315 18567 20321
rect 18509 20312 18521 20315
rect 16669 20275 16727 20281
rect 17788 20284 18521 20312
rect 17788 20256 17816 20284
rect 18509 20281 18521 20284
rect 18555 20281 18567 20315
rect 18509 20275 18567 20281
rect 24946 20272 24952 20324
rect 25004 20312 25010 20324
rect 25501 20315 25559 20321
rect 25501 20312 25513 20315
rect 25004 20284 25513 20312
rect 25004 20272 25010 20284
rect 25501 20281 25513 20284
rect 25547 20281 25559 20315
rect 25501 20275 25559 20281
rect 4525 20247 4583 20253
rect 4525 20244 4537 20247
rect 4212 20216 4537 20244
rect 4212 20204 4218 20216
rect 4525 20213 4537 20216
rect 4571 20213 4583 20247
rect 4525 20207 4583 20213
rect 5166 20204 5172 20256
rect 5224 20244 5230 20256
rect 5442 20244 5448 20256
rect 5224 20216 5448 20244
rect 5224 20204 5230 20216
rect 5442 20204 5448 20216
rect 5500 20244 5506 20256
rect 5721 20247 5779 20253
rect 5721 20244 5733 20247
rect 5500 20216 5733 20244
rect 5500 20204 5506 20216
rect 5721 20213 5733 20216
rect 5767 20213 5779 20247
rect 5721 20207 5779 20213
rect 6181 20247 6239 20253
rect 6181 20213 6193 20247
rect 6227 20244 6239 20247
rect 6270 20244 6276 20256
rect 6227 20216 6276 20244
rect 6227 20213 6239 20216
rect 6181 20207 6239 20213
rect 6270 20204 6276 20216
rect 6328 20204 6334 20256
rect 7558 20204 7564 20256
rect 7616 20244 7622 20256
rect 8113 20247 8171 20253
rect 8113 20244 8125 20247
rect 7616 20216 8125 20244
rect 7616 20204 7622 20216
rect 8113 20213 8125 20216
rect 8159 20244 8171 20247
rect 8757 20247 8815 20253
rect 8757 20244 8769 20247
rect 8159 20216 8769 20244
rect 8159 20213 8171 20216
rect 8113 20207 8171 20213
rect 8757 20213 8769 20216
rect 8803 20244 8815 20247
rect 9030 20244 9036 20256
rect 8803 20216 9036 20244
rect 8803 20213 8815 20216
rect 8757 20207 8815 20213
rect 9030 20204 9036 20216
rect 9088 20204 9094 20256
rect 9769 20247 9827 20253
rect 9769 20213 9781 20247
rect 9815 20244 9827 20247
rect 9950 20244 9956 20256
rect 9815 20216 9956 20244
rect 9815 20213 9827 20216
rect 9769 20207 9827 20213
rect 9950 20204 9956 20216
rect 10008 20244 10014 20256
rect 10229 20247 10287 20253
rect 10229 20244 10241 20247
rect 10008 20216 10241 20244
rect 10008 20204 10014 20216
rect 10229 20213 10241 20216
rect 10275 20213 10287 20247
rect 10229 20207 10287 20213
rect 13722 20204 13728 20256
rect 13780 20244 13786 20256
rect 15194 20244 15200 20256
rect 13780 20216 15200 20244
rect 13780 20204 13786 20216
rect 15194 20204 15200 20216
rect 15252 20204 15258 20256
rect 15378 20204 15384 20256
rect 15436 20244 15442 20256
rect 15657 20247 15715 20253
rect 15657 20244 15669 20247
rect 15436 20216 15669 20244
rect 15436 20204 15442 20216
rect 15657 20213 15669 20216
rect 15703 20244 15715 20247
rect 15841 20247 15899 20253
rect 15841 20244 15853 20247
rect 15703 20216 15853 20244
rect 15703 20213 15715 20216
rect 15657 20207 15715 20213
rect 15841 20213 15853 20216
rect 15887 20213 15899 20247
rect 17770 20244 17776 20256
rect 17731 20216 17776 20244
rect 15841 20207 15899 20213
rect 17770 20204 17776 20216
rect 17828 20204 17834 20256
rect 19978 20244 19984 20256
rect 19939 20216 19984 20244
rect 19978 20204 19984 20216
rect 20036 20204 20042 20256
rect 21634 20244 21640 20256
rect 21595 20216 21640 20244
rect 21634 20204 21640 20216
rect 21692 20204 21698 20256
rect 23382 20244 23388 20256
rect 23343 20216 23388 20244
rect 23382 20204 23388 20216
rect 23440 20244 23446 20256
rect 23477 20247 23535 20253
rect 23477 20244 23489 20247
rect 23440 20216 23489 20244
rect 23440 20204 23446 20216
rect 23477 20213 23489 20216
rect 23523 20213 23535 20247
rect 23477 20207 23535 20213
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 2409 20043 2467 20049
rect 2409 20009 2421 20043
rect 2455 20040 2467 20043
rect 3326 20040 3332 20052
rect 2455 20012 3332 20040
rect 2455 20009 2467 20012
rect 2409 20003 2467 20009
rect 3326 20000 3332 20012
rect 3384 20000 3390 20052
rect 6086 20040 6092 20052
rect 5999 20012 6092 20040
rect 6086 20000 6092 20012
rect 6144 20040 6150 20052
rect 6730 20040 6736 20052
rect 6144 20012 6736 20040
rect 6144 20000 6150 20012
rect 6730 20000 6736 20012
rect 6788 20000 6794 20052
rect 7834 20000 7840 20052
rect 7892 20040 7898 20052
rect 8018 20040 8024 20052
rect 7892 20012 8024 20040
rect 7892 20000 7898 20012
rect 8018 20000 8024 20012
rect 8076 20040 8082 20052
rect 8205 20043 8263 20049
rect 8205 20040 8217 20043
rect 8076 20012 8217 20040
rect 8076 20000 8082 20012
rect 8205 20009 8217 20012
rect 8251 20009 8263 20043
rect 8754 20040 8760 20052
rect 8715 20012 8760 20040
rect 8205 20003 8263 20009
rect 8754 20000 8760 20012
rect 8812 20000 8818 20052
rect 9953 20043 10011 20049
rect 9953 20009 9965 20043
rect 9999 20040 10011 20043
rect 10778 20040 10784 20052
rect 9999 20012 10784 20040
rect 9999 20009 10011 20012
rect 9953 20003 10011 20009
rect 10778 20000 10784 20012
rect 10836 20000 10842 20052
rect 11514 20040 11520 20052
rect 11475 20012 11520 20040
rect 11514 20000 11520 20012
rect 11572 20000 11578 20052
rect 12342 20040 12348 20052
rect 11624 20012 12348 20040
rect 2777 19975 2835 19981
rect 2777 19941 2789 19975
rect 2823 19972 2835 19975
rect 3142 19972 3148 19984
rect 2823 19944 3148 19972
rect 2823 19941 2835 19944
rect 2777 19935 2835 19941
rect 3142 19932 3148 19944
rect 3200 19972 3206 19984
rect 3200 19944 3372 19972
rect 3200 19932 3206 19944
rect 2869 19907 2927 19913
rect 2869 19873 2881 19907
rect 2915 19904 2927 19907
rect 3234 19904 3240 19916
rect 2915 19876 3240 19904
rect 2915 19873 2927 19876
rect 2869 19867 2927 19873
rect 3234 19864 3240 19876
rect 3292 19864 3298 19916
rect 3344 19913 3372 19944
rect 8938 19932 8944 19984
rect 8996 19972 9002 19984
rect 10321 19975 10379 19981
rect 10321 19972 10333 19975
rect 8996 19944 10333 19972
rect 8996 19932 9002 19944
rect 10321 19941 10333 19944
rect 10367 19941 10379 19975
rect 10321 19935 10379 19941
rect 10410 19932 10416 19984
rect 10468 19972 10474 19984
rect 11624 19972 11652 20012
rect 12342 20000 12348 20012
rect 12400 20000 12406 20052
rect 13078 20040 13084 20052
rect 13039 20012 13084 20040
rect 13078 20000 13084 20012
rect 13136 20000 13142 20052
rect 14182 20000 14188 20052
rect 14240 20040 14246 20052
rect 14645 20043 14703 20049
rect 14645 20040 14657 20043
rect 14240 20012 14657 20040
rect 14240 20000 14246 20012
rect 14645 20009 14657 20012
rect 14691 20009 14703 20043
rect 14645 20003 14703 20009
rect 14918 20000 14924 20052
rect 14976 20040 14982 20052
rect 15013 20043 15071 20049
rect 15013 20040 15025 20043
rect 14976 20012 15025 20040
rect 14976 20000 14982 20012
rect 15013 20009 15025 20012
rect 15059 20009 15071 20043
rect 15013 20003 15071 20009
rect 17773 20043 17831 20049
rect 17773 20009 17785 20043
rect 17819 20040 17831 20043
rect 17862 20040 17868 20052
rect 17819 20012 17868 20040
rect 17819 20009 17831 20012
rect 17773 20003 17831 20009
rect 17862 20000 17868 20012
rect 17920 20000 17926 20052
rect 18506 20000 18512 20052
rect 18564 20040 18570 20052
rect 18966 20040 18972 20052
rect 18564 20012 18972 20040
rect 18564 20000 18570 20012
rect 18966 20000 18972 20012
rect 19024 20000 19030 20052
rect 20349 20043 20407 20049
rect 20349 20009 20361 20043
rect 20395 20040 20407 20043
rect 20901 20043 20959 20049
rect 20901 20040 20913 20043
rect 20395 20012 20913 20040
rect 20395 20009 20407 20012
rect 20349 20003 20407 20009
rect 20901 20009 20913 20012
rect 20947 20040 20959 20043
rect 21634 20040 21640 20052
rect 20947 20012 21640 20040
rect 20947 20009 20959 20012
rect 20901 20003 20959 20009
rect 21634 20000 21640 20012
rect 21692 20000 21698 20052
rect 22462 20040 22468 20052
rect 22423 20012 22468 20040
rect 22462 20000 22468 20012
rect 22520 20000 22526 20052
rect 23658 20000 23664 20052
rect 23716 20040 23722 20052
rect 24029 20043 24087 20049
rect 24029 20040 24041 20043
rect 23716 20012 24041 20040
rect 23716 20000 23722 20012
rect 24029 20009 24041 20012
rect 24075 20009 24087 20043
rect 24486 20040 24492 20052
rect 24447 20012 24492 20040
rect 24029 20003 24087 20009
rect 24486 20000 24492 20012
rect 24544 20040 24550 20052
rect 24854 20040 24860 20052
rect 24544 20012 24860 20040
rect 24544 20000 24550 20012
rect 24854 20000 24860 20012
rect 24912 20000 24918 20052
rect 25406 20040 25412 20052
rect 25367 20012 25412 20040
rect 25406 20000 25412 20012
rect 25464 20000 25470 20052
rect 10468 19944 11652 19972
rect 11885 19975 11943 19981
rect 10468 19932 10474 19944
rect 11885 19941 11897 19975
rect 11931 19972 11943 19975
rect 11974 19972 11980 19984
rect 11931 19944 11980 19972
rect 11931 19941 11943 19944
rect 11885 19935 11943 19941
rect 11974 19932 11980 19944
rect 12032 19932 12038 19984
rect 12986 19972 12992 19984
rect 12947 19944 12992 19972
rect 12986 19932 12992 19944
rect 13044 19932 13050 19984
rect 15648 19975 15706 19981
rect 15648 19941 15660 19975
rect 15694 19972 15706 19975
rect 16482 19972 16488 19984
rect 15694 19944 16488 19972
rect 15694 19941 15706 19944
rect 15648 19935 15706 19941
rect 16482 19932 16488 19944
rect 16540 19932 16546 19984
rect 18046 19932 18052 19984
rect 18104 19981 18110 19984
rect 18104 19975 18168 19981
rect 18104 19941 18122 19975
rect 18156 19972 18168 19975
rect 20530 19972 20536 19984
rect 18156 19944 20536 19972
rect 18156 19941 18168 19944
rect 18104 19935 18168 19941
rect 18104 19932 18110 19935
rect 20530 19932 20536 19944
rect 20588 19972 20594 19984
rect 20717 19975 20775 19981
rect 20717 19972 20729 19975
rect 20588 19944 20729 19972
rect 20588 19932 20594 19944
rect 20717 19941 20729 19944
rect 20763 19941 20775 19975
rect 21266 19972 21272 19984
rect 21227 19944 21272 19972
rect 20717 19935 20775 19941
rect 3329 19907 3387 19913
rect 3329 19873 3341 19907
rect 3375 19873 3387 19907
rect 3329 19867 3387 19873
rect 3513 19907 3571 19913
rect 3513 19873 3525 19907
rect 3559 19904 3571 19907
rect 4154 19904 4160 19916
rect 3559 19876 4160 19904
rect 3559 19873 3571 19876
rect 3513 19867 3571 19873
rect 4154 19864 4160 19876
rect 4212 19904 4218 19916
rect 4321 19907 4379 19913
rect 4321 19904 4333 19907
rect 4212 19876 4333 19904
rect 4212 19864 4218 19876
rect 4321 19873 4333 19876
rect 4367 19873 4379 19907
rect 4321 19867 4379 19873
rect 6914 19864 6920 19916
rect 6972 19904 6978 19916
rect 7081 19907 7139 19913
rect 7081 19904 7093 19907
rect 6972 19876 7093 19904
rect 6972 19864 6978 19876
rect 7081 19873 7093 19876
rect 7127 19873 7139 19907
rect 7081 19867 7139 19873
rect 11440 19876 12112 19904
rect 11440 19848 11468 19876
rect 2133 19839 2191 19845
rect 2133 19805 2145 19839
rect 2179 19836 2191 19839
rect 2682 19836 2688 19848
rect 2179 19808 2688 19836
rect 2179 19805 2191 19808
rect 2133 19799 2191 19805
rect 2682 19796 2688 19808
rect 2740 19836 2746 19848
rect 3050 19836 3056 19848
rect 2740 19808 3056 19836
rect 2740 19796 2746 19808
rect 3050 19796 3056 19808
rect 3108 19796 3114 19848
rect 3142 19796 3148 19848
rect 3200 19836 3206 19848
rect 3786 19836 3792 19848
rect 3200 19808 3792 19836
rect 3200 19796 3206 19808
rect 3786 19796 3792 19808
rect 3844 19796 3850 19848
rect 4062 19836 4068 19848
rect 4023 19808 4068 19836
rect 4062 19796 4068 19808
rect 4120 19796 4126 19848
rect 5074 19796 5080 19848
rect 5132 19836 5138 19848
rect 6638 19836 6644 19848
rect 5132 19808 6644 19836
rect 5132 19796 5138 19808
rect 6638 19796 6644 19808
rect 6696 19836 6702 19848
rect 6825 19839 6883 19845
rect 6825 19836 6837 19839
rect 6696 19808 6837 19836
rect 6696 19796 6702 19808
rect 6825 19805 6837 19808
rect 6871 19805 6883 19839
rect 6825 19799 6883 19805
rect 9766 19796 9772 19848
rect 9824 19836 9830 19848
rect 10413 19839 10471 19845
rect 10413 19836 10425 19839
rect 9824 19808 10425 19836
rect 9824 19796 9830 19808
rect 10413 19805 10425 19808
rect 10459 19805 10471 19839
rect 10413 19799 10471 19805
rect 10597 19839 10655 19845
rect 10597 19805 10609 19839
rect 10643 19836 10655 19839
rect 11422 19836 11428 19848
rect 10643 19808 11428 19836
rect 10643 19805 10655 19808
rect 10597 19799 10655 19805
rect 9493 19771 9551 19777
rect 9493 19737 9505 19771
rect 9539 19768 9551 19771
rect 10612 19768 10640 19799
rect 11422 19796 11428 19808
rect 11480 19796 11486 19848
rect 12084 19845 12112 19876
rect 12434 19864 12440 19916
rect 12492 19904 12498 19916
rect 12621 19907 12679 19913
rect 12621 19904 12633 19907
rect 12492 19876 12633 19904
rect 12492 19864 12498 19876
rect 12621 19873 12633 19876
rect 12667 19904 12679 19907
rect 13449 19907 13507 19913
rect 13449 19904 13461 19907
rect 12667 19876 13461 19904
rect 12667 19873 12679 19876
rect 12621 19867 12679 19873
rect 13449 19873 13461 19876
rect 13495 19873 13507 19907
rect 13449 19867 13507 19873
rect 13538 19864 13544 19916
rect 13596 19904 13602 19916
rect 14093 19907 14151 19913
rect 14093 19904 14105 19907
rect 13596 19876 14105 19904
rect 13596 19864 13602 19876
rect 14093 19873 14105 19876
rect 14139 19873 14151 19907
rect 14093 19867 14151 19873
rect 15194 19864 15200 19916
rect 15252 19904 15258 19916
rect 15381 19907 15439 19913
rect 15381 19904 15393 19907
rect 15252 19876 15393 19904
rect 15252 19864 15258 19876
rect 15381 19873 15393 19876
rect 15427 19904 15439 19907
rect 15470 19904 15476 19916
rect 15427 19876 15476 19904
rect 15427 19873 15439 19876
rect 15381 19867 15439 19873
rect 15470 19864 15476 19876
rect 15528 19904 15534 19916
rect 17865 19907 17923 19913
rect 17865 19904 17877 19907
rect 15528 19876 17877 19904
rect 15528 19864 15534 19876
rect 17865 19873 17877 19876
rect 17911 19873 17923 19907
rect 20732 19904 20760 19935
rect 21266 19932 21272 19944
rect 21324 19932 21330 19984
rect 21818 19932 21824 19984
rect 21876 19972 21882 19984
rect 22370 19972 22376 19984
rect 21876 19944 22376 19972
rect 21876 19932 21882 19944
rect 22370 19932 22376 19944
rect 22428 19932 22434 19984
rect 25222 19932 25228 19984
rect 25280 19972 25286 19984
rect 25777 19975 25835 19981
rect 25777 19972 25789 19975
rect 25280 19944 25789 19972
rect 25280 19932 25286 19944
rect 25777 19941 25789 19944
rect 25823 19941 25835 19975
rect 25777 19935 25835 19941
rect 22002 19904 22008 19916
rect 20732 19876 22008 19904
rect 17865 19867 17923 19873
rect 11977 19839 12035 19845
rect 11977 19805 11989 19839
rect 12023 19805 12035 19839
rect 11977 19799 12035 19805
rect 12069 19839 12127 19845
rect 12069 19805 12081 19839
rect 12115 19805 12127 19839
rect 12069 19799 12127 19805
rect 9539 19740 10640 19768
rect 9539 19737 9551 19740
rect 9493 19731 9551 19737
rect 11146 19728 11152 19780
rect 11204 19768 11210 19780
rect 11204 19740 11468 19768
rect 11204 19728 11210 19740
rect 1670 19700 1676 19712
rect 1631 19672 1676 19700
rect 1670 19660 1676 19672
rect 1728 19660 1734 19712
rect 2866 19660 2872 19712
rect 2924 19700 2930 19712
rect 3329 19703 3387 19709
rect 3329 19700 3341 19703
rect 2924 19672 3341 19700
rect 2924 19660 2930 19672
rect 3329 19669 3341 19672
rect 3375 19669 3387 19703
rect 3786 19700 3792 19712
rect 3747 19672 3792 19700
rect 3329 19663 3387 19669
rect 3786 19660 3792 19672
rect 3844 19660 3850 19712
rect 5442 19700 5448 19712
rect 5403 19672 5448 19700
rect 5442 19660 5448 19672
rect 5500 19660 5506 19712
rect 6362 19700 6368 19712
rect 6323 19672 6368 19700
rect 6362 19660 6368 19672
rect 6420 19660 6426 19712
rect 11054 19700 11060 19712
rect 11015 19672 11060 19700
rect 11054 19660 11060 19672
rect 11112 19700 11118 19712
rect 11333 19703 11391 19709
rect 11333 19700 11345 19703
rect 11112 19672 11345 19700
rect 11112 19660 11118 19672
rect 11333 19669 11345 19672
rect 11379 19669 11391 19703
rect 11440 19700 11468 19740
rect 11882 19728 11888 19780
rect 11940 19768 11946 19780
rect 11992 19768 12020 19799
rect 12802 19796 12808 19848
rect 12860 19836 12866 19848
rect 13633 19839 13691 19845
rect 13633 19836 13645 19839
rect 12860 19808 13645 19836
rect 12860 19796 12866 19808
rect 13633 19805 13645 19808
rect 13679 19805 13691 19839
rect 21358 19836 21364 19848
rect 21319 19808 21364 19836
rect 13633 19799 13691 19805
rect 21358 19796 21364 19808
rect 21416 19796 21422 19848
rect 21468 19845 21496 19876
rect 22002 19864 22008 19876
rect 22060 19864 22066 19916
rect 22278 19864 22284 19916
rect 22336 19864 22342 19916
rect 22830 19904 22836 19916
rect 22791 19876 22836 19904
rect 22830 19864 22836 19876
rect 22888 19864 22894 19916
rect 24026 19864 24032 19916
rect 24084 19904 24090 19916
rect 24397 19907 24455 19913
rect 24397 19904 24409 19907
rect 24084 19876 24409 19904
rect 24084 19864 24090 19876
rect 24397 19873 24409 19876
rect 24443 19873 24455 19907
rect 24397 19867 24455 19873
rect 21453 19839 21511 19845
rect 21453 19805 21465 19839
rect 21499 19805 21511 19839
rect 21453 19799 21511 19805
rect 21910 19796 21916 19848
rect 21968 19836 21974 19848
rect 22296 19836 22324 19864
rect 21968 19808 22324 19836
rect 21968 19796 21974 19808
rect 22738 19796 22744 19848
rect 22796 19836 22802 19848
rect 22922 19836 22928 19848
rect 22796 19808 22928 19836
rect 22796 19796 22802 19808
rect 22922 19796 22928 19808
rect 22980 19796 22986 19848
rect 23106 19836 23112 19848
rect 23067 19808 23112 19836
rect 23106 19796 23112 19808
rect 23164 19796 23170 19848
rect 23566 19796 23572 19848
rect 23624 19836 23630 19848
rect 24578 19836 24584 19848
rect 23624 19808 24584 19836
rect 23624 19796 23630 19808
rect 24578 19796 24584 19808
rect 24636 19796 24642 19848
rect 11940 19740 12020 19768
rect 11940 19728 11946 19740
rect 12158 19728 12164 19780
rect 12216 19768 12222 19780
rect 15286 19768 15292 19780
rect 12216 19740 15292 19768
rect 12216 19728 12222 19740
rect 15286 19728 15292 19740
rect 15344 19728 15350 19780
rect 21726 19728 21732 19780
rect 21784 19768 21790 19780
rect 21784 19740 24072 19768
rect 21784 19728 21790 19740
rect 12176 19700 12204 19728
rect 24044 19712 24072 19740
rect 11440 19672 12204 19700
rect 11333 19663 11391 19669
rect 16574 19660 16580 19712
rect 16632 19700 16638 19712
rect 16761 19703 16819 19709
rect 16761 19700 16773 19703
rect 16632 19672 16773 19700
rect 16632 19660 16638 19672
rect 16761 19669 16773 19672
rect 16807 19669 16819 19703
rect 17402 19700 17408 19712
rect 17363 19672 17408 19700
rect 16761 19663 16819 19669
rect 17402 19660 17408 19672
rect 17460 19660 17466 19712
rect 19242 19700 19248 19712
rect 19203 19672 19248 19700
rect 19242 19660 19248 19672
rect 19300 19700 19306 19712
rect 19797 19703 19855 19709
rect 19797 19700 19809 19703
rect 19300 19672 19809 19700
rect 19300 19660 19306 19672
rect 19797 19669 19809 19672
rect 19843 19700 19855 19703
rect 20162 19700 20168 19712
rect 19843 19672 20168 19700
rect 19843 19669 19855 19672
rect 19797 19663 19855 19669
rect 20162 19660 20168 19672
rect 20220 19660 20226 19712
rect 20530 19660 20536 19712
rect 20588 19700 20594 19712
rect 21450 19700 21456 19712
rect 20588 19672 21456 19700
rect 20588 19660 20594 19672
rect 21450 19660 21456 19672
rect 21508 19660 21514 19712
rect 21910 19700 21916 19712
rect 21871 19672 21916 19700
rect 21910 19660 21916 19672
rect 21968 19660 21974 19712
rect 22370 19700 22376 19712
rect 22331 19672 22376 19700
rect 22370 19660 22376 19672
rect 22428 19660 22434 19712
rect 22462 19660 22468 19712
rect 22520 19700 22526 19712
rect 23382 19700 23388 19712
rect 22520 19672 23388 19700
rect 22520 19660 22526 19672
rect 23382 19660 23388 19672
rect 23440 19700 23446 19712
rect 23661 19703 23719 19709
rect 23661 19700 23673 19703
rect 23440 19672 23673 19700
rect 23440 19660 23446 19672
rect 23661 19669 23673 19672
rect 23707 19669 23719 19703
rect 23661 19663 23719 19669
rect 24026 19660 24032 19712
rect 24084 19660 24090 19712
rect 24762 19660 24768 19712
rect 24820 19700 24826 19712
rect 25038 19700 25044 19712
rect 24820 19672 25044 19700
rect 24820 19660 24826 19672
rect 25038 19660 25044 19672
rect 25096 19660 25102 19712
rect 26237 19703 26295 19709
rect 26237 19669 26249 19703
rect 26283 19700 26295 19703
rect 26326 19700 26332 19712
rect 26283 19672 26332 19700
rect 26283 19669 26295 19672
rect 26237 19663 26295 19669
rect 26326 19660 26332 19672
rect 26384 19660 26390 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 3234 19456 3240 19508
rect 3292 19496 3298 19508
rect 3421 19499 3479 19505
rect 3421 19496 3433 19499
rect 3292 19468 3433 19496
rect 3292 19456 3298 19468
rect 3421 19465 3433 19468
rect 3467 19465 3479 19499
rect 3421 19459 3479 19465
rect 8938 19456 8944 19508
rect 8996 19496 9002 19508
rect 9309 19499 9367 19505
rect 9309 19496 9321 19499
rect 8996 19468 9321 19496
rect 8996 19456 9002 19468
rect 9309 19465 9321 19468
rect 9355 19465 9367 19499
rect 9766 19496 9772 19508
rect 9727 19468 9772 19496
rect 9309 19459 9367 19465
rect 9766 19456 9772 19468
rect 9824 19456 9830 19508
rect 12802 19496 12808 19508
rect 12763 19468 12808 19496
rect 12802 19456 12808 19468
rect 12860 19456 12866 19508
rect 14642 19456 14648 19508
rect 14700 19496 14706 19508
rect 15381 19499 15439 19505
rect 15381 19496 15393 19499
rect 14700 19468 15393 19496
rect 14700 19456 14706 19468
rect 15381 19465 15393 19468
rect 15427 19465 15439 19499
rect 16482 19496 16488 19508
rect 16443 19468 16488 19496
rect 15381 19459 15439 19465
rect 16482 19456 16488 19468
rect 16540 19456 16546 19508
rect 20993 19499 21051 19505
rect 20993 19465 21005 19499
rect 21039 19496 21051 19499
rect 21358 19496 21364 19508
rect 21039 19468 21364 19496
rect 21039 19465 21051 19468
rect 20993 19459 21051 19465
rect 21358 19456 21364 19468
rect 21416 19456 21422 19508
rect 22557 19499 22615 19505
rect 22557 19465 22569 19499
rect 22603 19496 22615 19499
rect 22830 19496 22836 19508
rect 22603 19468 22836 19496
rect 22603 19465 22615 19468
rect 22557 19459 22615 19465
rect 22830 19456 22836 19468
rect 22888 19456 22894 19508
rect 23477 19499 23535 19505
rect 23477 19465 23489 19499
rect 23523 19496 23535 19499
rect 23566 19496 23572 19508
rect 23523 19468 23572 19496
rect 23523 19465 23535 19468
rect 23477 19459 23535 19465
rect 23566 19456 23572 19468
rect 23624 19456 23630 19508
rect 23658 19456 23664 19508
rect 23716 19496 23722 19508
rect 26142 19496 26148 19508
rect 23716 19468 26148 19496
rect 23716 19456 23722 19468
rect 26142 19456 26148 19468
rect 26200 19456 26206 19508
rect 1670 19388 1676 19440
rect 1728 19428 1734 19440
rect 1728 19400 3280 19428
rect 1728 19388 1734 19400
rect 3252 19372 3280 19400
rect 2682 19360 2688 19372
rect 2643 19332 2688 19360
rect 2682 19320 2688 19332
rect 2740 19320 2746 19372
rect 3234 19320 3240 19372
rect 3292 19320 3298 19372
rect 4154 19360 4160 19372
rect 4115 19332 4160 19360
rect 4154 19320 4160 19332
rect 4212 19320 4218 19372
rect 5810 19360 5816 19372
rect 5771 19332 5816 19360
rect 5810 19320 5816 19332
rect 5868 19320 5874 19372
rect 7929 19363 7987 19369
rect 7929 19329 7941 19363
rect 7975 19360 7987 19363
rect 8110 19360 8116 19372
rect 7975 19332 8116 19360
rect 7975 19329 7987 19332
rect 7929 19323 7987 19329
rect 8110 19320 8116 19332
rect 8168 19360 8174 19372
rect 8846 19360 8852 19372
rect 8168 19332 8340 19360
rect 8807 19332 8852 19360
rect 8168 19320 8174 19332
rect 2409 19295 2467 19301
rect 2409 19292 2421 19295
rect 1872 19264 2421 19292
rect 934 19116 940 19168
rect 992 19156 998 19168
rect 1872 19165 1900 19264
rect 2409 19261 2421 19264
rect 2455 19261 2467 19295
rect 4062 19292 4068 19304
rect 4023 19264 4068 19292
rect 2409 19255 2467 19261
rect 4062 19252 4068 19264
rect 4120 19252 4126 19304
rect 4709 19295 4767 19301
rect 4709 19261 4721 19295
rect 4755 19292 4767 19295
rect 5537 19295 5595 19301
rect 5537 19292 5549 19295
rect 4755 19264 5549 19292
rect 4755 19261 4767 19264
rect 4709 19255 4767 19261
rect 5537 19261 5549 19264
rect 5583 19292 5595 19295
rect 6638 19292 6644 19304
rect 5583 19264 6644 19292
rect 5583 19261 5595 19264
rect 5537 19255 5595 19261
rect 6638 19252 6644 19264
rect 6696 19252 6702 19304
rect 7193 19295 7251 19301
rect 7193 19261 7205 19295
rect 7239 19292 7251 19295
rect 7466 19292 7472 19304
rect 7239 19264 7472 19292
rect 7239 19261 7251 19264
rect 7193 19255 7251 19261
rect 7466 19252 7472 19264
rect 7524 19292 7530 19304
rect 7745 19295 7803 19301
rect 7745 19292 7757 19295
rect 7524 19264 7757 19292
rect 7524 19252 7530 19264
rect 7745 19261 7757 19264
rect 7791 19261 7803 19295
rect 8312 19292 8340 19332
rect 8846 19320 8852 19332
rect 8904 19320 8910 19372
rect 9784 19360 9812 19456
rect 20806 19388 20812 19440
rect 20864 19428 20870 19440
rect 20864 19400 21772 19428
rect 20864 19388 20870 19400
rect 21744 19372 21772 19400
rect 22002 19388 22008 19440
rect 22060 19428 22066 19440
rect 23584 19428 23612 19456
rect 24673 19431 24731 19437
rect 24673 19428 24685 19431
rect 22060 19400 22600 19428
rect 23584 19400 24685 19428
rect 22060 19388 22066 19400
rect 22572 19372 22600 19400
rect 15933 19363 15991 19369
rect 15933 19360 15945 19363
rect 9784 19332 9996 19360
rect 8662 19292 8668 19304
rect 8312 19264 8432 19292
rect 8623 19264 8668 19292
rect 7745 19255 7803 19261
rect 2130 19184 2136 19236
rect 2188 19224 2194 19236
rect 2501 19227 2559 19233
rect 2501 19224 2513 19227
rect 2188 19196 2513 19224
rect 2188 19184 2194 19196
rect 2501 19193 2513 19196
rect 2547 19193 2559 19227
rect 2501 19187 2559 19193
rect 2774 19184 2780 19236
rect 2832 19224 2838 19236
rect 4080 19224 4108 19252
rect 5350 19224 5356 19236
rect 2832 19196 4108 19224
rect 5000 19196 5356 19224
rect 2832 19184 2838 19196
rect 1857 19159 1915 19165
rect 1857 19156 1869 19159
rect 992 19128 1869 19156
rect 992 19116 998 19128
rect 1857 19125 1869 19128
rect 1903 19125 1915 19159
rect 2038 19156 2044 19168
rect 1999 19128 2044 19156
rect 1857 19119 1915 19125
rect 2038 19116 2044 19128
rect 2096 19116 2102 19168
rect 2866 19116 2872 19168
rect 2924 19156 2930 19168
rect 3053 19159 3111 19165
rect 3053 19156 3065 19159
rect 2924 19128 3065 19156
rect 2924 19116 2930 19128
rect 3053 19125 3065 19128
rect 3099 19125 3111 19159
rect 3602 19156 3608 19168
rect 3563 19128 3608 19156
rect 3053 19119 3111 19125
rect 3602 19116 3608 19128
rect 3660 19116 3666 19168
rect 3970 19156 3976 19168
rect 3931 19128 3976 19156
rect 3970 19116 3976 19128
rect 4028 19116 4034 19168
rect 4890 19116 4896 19168
rect 4948 19156 4954 19168
rect 5000 19165 5028 19196
rect 5350 19184 5356 19196
rect 5408 19224 5414 19236
rect 5629 19227 5687 19233
rect 5629 19224 5641 19227
rect 5408 19196 5641 19224
rect 5408 19184 5414 19196
rect 5629 19193 5641 19196
rect 5675 19193 5687 19227
rect 5629 19187 5687 19193
rect 6362 19184 6368 19236
rect 6420 19224 6426 19236
rect 6420 19196 7328 19224
rect 6420 19184 6426 19196
rect 4985 19159 5043 19165
rect 4985 19156 4997 19159
rect 4948 19128 4997 19156
rect 4948 19116 4954 19128
rect 4985 19125 4997 19128
rect 5031 19125 5043 19159
rect 5166 19156 5172 19168
rect 5127 19128 5172 19156
rect 4985 19119 5043 19125
rect 5166 19116 5172 19128
rect 5224 19116 5230 19168
rect 5810 19116 5816 19168
rect 5868 19156 5874 19168
rect 6181 19159 6239 19165
rect 6181 19156 6193 19159
rect 5868 19128 6193 19156
rect 5868 19116 5874 19128
rect 6181 19125 6193 19128
rect 6227 19125 6239 19159
rect 6181 19119 6239 19125
rect 6546 19116 6552 19168
rect 6604 19156 6610 19168
rect 6641 19159 6699 19165
rect 6641 19156 6653 19159
rect 6604 19128 6653 19156
rect 6604 19116 6610 19128
rect 6641 19125 6653 19128
rect 6687 19156 6699 19159
rect 7190 19156 7196 19168
rect 6687 19128 7196 19156
rect 6687 19125 6699 19128
rect 6641 19119 6699 19125
rect 7190 19116 7196 19128
rect 7248 19116 7254 19168
rect 7300 19165 7328 19196
rect 7374 19184 7380 19236
rect 7432 19224 7438 19236
rect 7653 19227 7711 19233
rect 7653 19224 7665 19227
rect 7432 19196 7665 19224
rect 7432 19184 7438 19196
rect 7653 19193 7665 19196
rect 7699 19224 7711 19227
rect 8018 19224 8024 19236
rect 7699 19196 8024 19224
rect 7699 19193 7711 19196
rect 7653 19187 7711 19193
rect 8018 19184 8024 19196
rect 8076 19184 8082 19236
rect 8404 19165 8432 19264
rect 8662 19252 8668 19264
rect 8720 19252 8726 19304
rect 9861 19295 9919 19301
rect 9861 19261 9873 19295
rect 9907 19261 9919 19295
rect 9861 19255 9919 19261
rect 9582 19184 9588 19236
rect 9640 19224 9646 19236
rect 9876 19224 9904 19255
rect 9640 19196 9904 19224
rect 9640 19184 9646 19196
rect 9968 19168 9996 19332
rect 15120 19332 15945 19360
rect 10128 19295 10186 19301
rect 10128 19261 10140 19295
rect 10174 19261 10186 19295
rect 10128 19255 10186 19261
rect 12897 19295 12955 19301
rect 12897 19261 12909 19295
rect 12943 19261 12955 19295
rect 12897 19255 12955 19261
rect 7285 19159 7343 19165
rect 7285 19125 7297 19159
rect 7331 19125 7343 19159
rect 7285 19119 7343 19125
rect 8389 19159 8447 19165
rect 8389 19125 8401 19159
rect 8435 19156 8447 19159
rect 8846 19156 8852 19168
rect 8435 19128 8852 19156
rect 8435 19125 8447 19128
rect 8389 19119 8447 19125
rect 8846 19116 8852 19128
rect 8904 19116 8910 19168
rect 9950 19116 9956 19168
rect 10008 19116 10014 19168
rect 10042 19116 10048 19168
rect 10100 19156 10106 19168
rect 10152 19156 10180 19255
rect 10226 19184 10232 19236
rect 10284 19184 10290 19236
rect 12912 19224 12940 19255
rect 12986 19252 12992 19304
rect 13044 19292 13050 19304
rect 13153 19295 13211 19301
rect 13153 19292 13165 19295
rect 13044 19264 13165 19292
rect 13044 19252 13050 19264
rect 13153 19261 13165 19264
rect 13199 19261 13211 19295
rect 15120 19292 15148 19332
rect 15933 19329 15945 19332
rect 15979 19360 15991 19363
rect 16758 19360 16764 19372
rect 15979 19332 16764 19360
rect 15979 19329 15991 19332
rect 15933 19323 15991 19329
rect 16758 19320 16764 19332
rect 16816 19320 16822 19372
rect 20990 19360 20996 19372
rect 20640 19332 20996 19360
rect 16942 19292 16948 19304
rect 13153 19255 13211 19261
rect 14292 19264 15148 19292
rect 16903 19264 16948 19292
rect 13630 19224 13636 19236
rect 12912 19196 13636 19224
rect 13630 19184 13636 19196
rect 13688 19184 13694 19236
rect 10100 19128 10180 19156
rect 10244 19156 10272 19184
rect 11146 19156 11152 19168
rect 10244 19128 11152 19156
rect 10100 19116 10106 19128
rect 11146 19116 11152 19128
rect 11204 19116 11210 19168
rect 11241 19159 11299 19165
rect 11241 19125 11253 19159
rect 11287 19156 11299 19159
rect 11422 19156 11428 19168
rect 11287 19128 11428 19156
rect 11287 19125 11299 19128
rect 11241 19119 11299 19125
rect 11422 19116 11428 19128
rect 11480 19116 11486 19168
rect 11882 19156 11888 19168
rect 11843 19128 11888 19156
rect 11882 19116 11888 19128
rect 11940 19116 11946 19168
rect 11974 19116 11980 19168
rect 12032 19156 12038 19168
rect 12161 19159 12219 19165
rect 12161 19156 12173 19159
rect 12032 19128 12173 19156
rect 12032 19116 12038 19128
rect 12161 19125 12173 19128
rect 12207 19125 12219 19159
rect 12161 19119 12219 19125
rect 13814 19116 13820 19168
rect 13872 19156 13878 19168
rect 14292 19165 14320 19264
rect 16942 19252 16948 19264
rect 17000 19252 17006 19304
rect 17494 19292 17500 19304
rect 17455 19264 17500 19292
rect 17494 19252 17500 19264
rect 17552 19252 17558 19304
rect 18693 19295 18751 19301
rect 18693 19261 18705 19295
rect 18739 19292 18751 19295
rect 19426 19292 19432 19304
rect 18739 19264 19432 19292
rect 18739 19261 18751 19264
rect 18693 19255 18751 19261
rect 19426 19252 19432 19264
rect 19484 19252 19490 19304
rect 14921 19227 14979 19233
rect 14921 19193 14933 19227
rect 14967 19224 14979 19227
rect 15654 19224 15660 19236
rect 14967 19196 15660 19224
rect 14967 19193 14979 19196
rect 14921 19187 14979 19193
rect 15654 19184 15660 19196
rect 15712 19224 15718 19236
rect 15841 19227 15899 19233
rect 15841 19224 15853 19227
rect 15712 19196 15853 19224
rect 15712 19184 15718 19196
rect 15841 19193 15853 19196
rect 15887 19193 15899 19227
rect 15841 19187 15899 19193
rect 17865 19227 17923 19233
rect 17865 19193 17877 19227
rect 17911 19224 17923 19227
rect 18938 19227 18996 19233
rect 18938 19224 18950 19227
rect 17911 19196 18950 19224
rect 17911 19193 17923 19196
rect 17865 19187 17923 19193
rect 18938 19193 18950 19196
rect 18984 19224 18996 19227
rect 19242 19224 19248 19236
rect 18984 19196 19248 19224
rect 18984 19193 18996 19196
rect 18938 19187 18996 19193
rect 19242 19184 19248 19196
rect 19300 19184 19306 19236
rect 14277 19159 14335 19165
rect 14277 19156 14289 19159
rect 13872 19128 14289 19156
rect 13872 19116 13878 19128
rect 14277 19125 14289 19128
rect 14323 19125 14335 19159
rect 14277 19119 14335 19125
rect 15289 19159 15347 19165
rect 15289 19125 15301 19159
rect 15335 19156 15347 19159
rect 15746 19156 15752 19168
rect 15335 19128 15752 19156
rect 15335 19125 15347 19128
rect 15289 19119 15347 19125
rect 15746 19116 15752 19128
rect 15804 19116 15810 19168
rect 18046 19116 18052 19168
rect 18104 19156 18110 19168
rect 18322 19156 18328 19168
rect 18104 19128 18328 19156
rect 18104 19116 18110 19128
rect 18322 19116 18328 19128
rect 18380 19116 18386 19168
rect 19978 19116 19984 19168
rect 20036 19156 20042 19168
rect 20073 19159 20131 19165
rect 20073 19156 20085 19159
rect 20036 19128 20085 19156
rect 20036 19116 20042 19128
rect 20073 19125 20085 19128
rect 20119 19156 20131 19159
rect 20640 19156 20668 19332
rect 20990 19320 20996 19332
rect 21048 19320 21054 19372
rect 21726 19360 21732 19372
rect 21639 19332 21732 19360
rect 21726 19320 21732 19332
rect 21784 19320 21790 19372
rect 22554 19320 22560 19372
rect 22612 19320 22618 19372
rect 24320 19369 24348 19400
rect 24673 19397 24685 19400
rect 24719 19428 24731 19431
rect 25038 19428 25044 19440
rect 24719 19400 25044 19428
rect 24719 19397 24731 19400
rect 24673 19391 24731 19397
rect 25038 19388 25044 19400
rect 25096 19388 25102 19440
rect 24305 19363 24363 19369
rect 24305 19329 24317 19363
rect 24351 19360 24363 19363
rect 24351 19332 24385 19360
rect 24351 19329 24363 19332
rect 24305 19323 24363 19329
rect 24578 19320 24584 19372
rect 24636 19360 24642 19372
rect 25866 19360 25872 19372
rect 24636 19332 25872 19360
rect 24636 19320 24642 19332
rect 25866 19320 25872 19332
rect 25924 19320 25930 19372
rect 22738 19252 22744 19304
rect 22796 19292 22802 19304
rect 22833 19295 22891 19301
rect 22833 19292 22845 19295
rect 22796 19264 22845 19292
rect 22796 19252 22802 19264
rect 22833 19261 22845 19264
rect 22879 19261 22891 19295
rect 24026 19292 24032 19304
rect 23987 19264 24032 19292
rect 22833 19255 22891 19261
rect 24026 19252 24032 19264
rect 24084 19252 24090 19304
rect 24118 19252 24124 19304
rect 24176 19292 24182 19304
rect 25041 19295 25099 19301
rect 25041 19292 25053 19295
rect 24176 19264 25053 19292
rect 24176 19252 24182 19264
rect 25041 19261 25053 19264
rect 25087 19261 25099 19295
rect 25041 19255 25099 19261
rect 25225 19295 25283 19301
rect 25225 19261 25237 19295
rect 25271 19292 25283 19295
rect 25777 19295 25835 19301
rect 25777 19292 25789 19295
rect 25271 19264 25789 19292
rect 25271 19261 25283 19264
rect 25225 19255 25283 19261
rect 25777 19261 25789 19264
rect 25823 19292 25835 19295
rect 25958 19292 25964 19304
rect 25823 19264 25964 19292
rect 25823 19261 25835 19264
rect 25777 19255 25835 19261
rect 25958 19252 25964 19264
rect 26016 19252 26022 19304
rect 26234 19292 26240 19304
rect 26195 19264 26240 19292
rect 26234 19252 26240 19264
rect 26292 19252 26298 19304
rect 20990 19184 20996 19236
rect 21048 19224 21054 19236
rect 21637 19227 21695 19233
rect 21637 19224 21649 19227
rect 21048 19196 21649 19224
rect 21048 19184 21054 19196
rect 21637 19193 21649 19196
rect 21683 19224 21695 19227
rect 21910 19224 21916 19236
rect 21683 19196 21916 19224
rect 21683 19193 21695 19196
rect 21637 19187 21695 19193
rect 21910 19184 21916 19196
rect 21968 19184 21974 19236
rect 21174 19156 21180 19168
rect 20119 19128 20668 19156
rect 21135 19128 21180 19156
rect 20119 19125 20131 19128
rect 20073 19119 20131 19125
rect 21174 19116 21180 19128
rect 21232 19116 21238 19168
rect 21450 19116 21456 19168
rect 21508 19156 21514 19168
rect 21545 19159 21603 19165
rect 21545 19156 21557 19159
rect 21508 19128 21557 19156
rect 21508 19116 21514 19128
rect 21545 19125 21557 19128
rect 21591 19125 21603 19159
rect 21545 19119 21603 19125
rect 23474 19116 23480 19168
rect 23532 19156 23538 19168
rect 23661 19159 23719 19165
rect 23661 19156 23673 19159
rect 23532 19128 23673 19156
rect 23532 19116 23538 19128
rect 23661 19125 23673 19128
rect 23707 19125 23719 19159
rect 23661 19119 23719 19125
rect 25130 19116 25136 19168
rect 25188 19156 25194 19168
rect 25409 19159 25467 19165
rect 25409 19156 25421 19159
rect 25188 19128 25421 19156
rect 25188 19116 25194 19128
rect 25409 19125 25421 19128
rect 25455 19125 25467 19159
rect 25409 19119 25467 19125
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 2406 18952 2412 18964
rect 2367 18924 2412 18952
rect 2406 18912 2412 18924
rect 2464 18912 2470 18964
rect 2869 18955 2927 18961
rect 2869 18921 2881 18955
rect 2915 18952 2927 18955
rect 3602 18952 3608 18964
rect 2915 18924 3608 18952
rect 2915 18921 2927 18924
rect 2869 18915 2927 18921
rect 3602 18912 3608 18924
rect 3660 18912 3666 18964
rect 3878 18912 3884 18964
rect 3936 18952 3942 18964
rect 4249 18955 4307 18961
rect 4249 18952 4261 18955
rect 3936 18924 4261 18952
rect 3936 18912 3942 18924
rect 4249 18921 4261 18924
rect 4295 18921 4307 18955
rect 4249 18915 4307 18921
rect 6733 18955 6791 18961
rect 6733 18921 6745 18955
rect 6779 18952 6791 18955
rect 6822 18952 6828 18964
rect 6779 18924 6828 18952
rect 6779 18921 6791 18924
rect 6733 18915 6791 18921
rect 6822 18912 6828 18924
rect 6880 18912 6886 18964
rect 8386 18912 8392 18964
rect 8444 18952 8450 18964
rect 8573 18955 8631 18961
rect 8573 18952 8585 18955
rect 8444 18924 8585 18952
rect 8444 18912 8450 18924
rect 8573 18921 8585 18924
rect 8619 18921 8631 18955
rect 8573 18915 8631 18921
rect 9493 18955 9551 18961
rect 9493 18921 9505 18955
rect 9539 18952 9551 18955
rect 10042 18952 10048 18964
rect 9539 18924 10048 18952
rect 9539 18921 9551 18924
rect 9493 18915 9551 18921
rect 10042 18912 10048 18924
rect 10100 18952 10106 18964
rect 11057 18955 11115 18961
rect 11057 18952 11069 18955
rect 10100 18924 11069 18952
rect 10100 18912 10106 18924
rect 11057 18921 11069 18924
rect 11103 18952 11115 18955
rect 12802 18952 12808 18964
rect 11103 18924 12808 18952
rect 11103 18921 11115 18924
rect 11057 18915 11115 18921
rect 12802 18912 12808 18924
rect 12860 18912 12866 18964
rect 12986 18912 12992 18964
rect 13044 18952 13050 18964
rect 13541 18955 13599 18961
rect 13541 18952 13553 18955
rect 13044 18924 13553 18952
rect 13044 18912 13050 18924
rect 13541 18921 13553 18924
rect 13587 18921 13599 18955
rect 15102 18952 15108 18964
rect 15063 18924 15108 18952
rect 13541 18915 13599 18921
rect 15102 18912 15108 18924
rect 15160 18912 15166 18964
rect 16206 18912 16212 18964
rect 16264 18952 16270 18964
rect 16301 18955 16359 18961
rect 16301 18952 16313 18955
rect 16264 18924 16313 18952
rect 16264 18912 16270 18924
rect 16301 18921 16313 18924
rect 16347 18921 16359 18955
rect 16301 18915 16359 18921
rect 16853 18955 16911 18961
rect 16853 18921 16865 18955
rect 16899 18921 16911 18955
rect 16853 18915 16911 18921
rect 18141 18955 18199 18961
rect 18141 18921 18153 18955
rect 18187 18952 18199 18955
rect 18230 18952 18236 18964
rect 18187 18924 18236 18952
rect 18187 18921 18199 18924
rect 18141 18915 18199 18921
rect 2774 18844 2780 18896
rect 2832 18884 2838 18896
rect 4338 18884 4344 18896
rect 2832 18856 4344 18884
rect 2832 18844 2838 18856
rect 4338 18844 4344 18856
rect 4396 18844 4402 18896
rect 5534 18844 5540 18896
rect 5592 18884 5598 18896
rect 6914 18884 6920 18896
rect 5592 18856 6920 18884
rect 5592 18844 5598 18856
rect 6914 18844 6920 18856
rect 6972 18844 6978 18896
rect 7285 18887 7343 18893
rect 7285 18853 7297 18887
rect 7331 18884 7343 18887
rect 7650 18884 7656 18896
rect 7331 18856 7656 18884
rect 7331 18853 7343 18856
rect 7285 18847 7343 18853
rect 7650 18844 7656 18856
rect 7708 18844 7714 18896
rect 8938 18844 8944 18896
rect 8996 18884 9002 18896
rect 10226 18884 10232 18896
rect 8996 18856 10232 18884
rect 8996 18844 9002 18856
rect 10226 18844 10232 18856
rect 10284 18844 10290 18896
rect 11514 18844 11520 18896
rect 11572 18884 11578 18896
rect 11885 18887 11943 18893
rect 11885 18884 11897 18887
rect 11572 18856 11897 18884
rect 11572 18844 11578 18856
rect 11885 18853 11897 18856
rect 11931 18884 11943 18887
rect 11977 18887 12035 18893
rect 11977 18884 11989 18887
rect 11931 18856 11989 18884
rect 11931 18853 11943 18856
rect 11885 18847 11943 18853
rect 11977 18853 11989 18856
rect 12023 18853 12035 18887
rect 16868 18884 16896 18915
rect 18230 18912 18236 18924
rect 18288 18912 18294 18964
rect 18414 18952 18420 18964
rect 18375 18924 18420 18952
rect 18414 18912 18420 18924
rect 18472 18912 18478 18964
rect 18506 18912 18512 18964
rect 18564 18952 18570 18964
rect 18877 18955 18935 18961
rect 18877 18952 18889 18955
rect 18564 18924 18889 18952
rect 18564 18912 18570 18924
rect 18877 18921 18889 18924
rect 18923 18952 18935 18955
rect 19242 18952 19248 18964
rect 18923 18924 19248 18952
rect 18923 18921 18935 18924
rect 18877 18915 18935 18921
rect 19242 18912 19248 18924
rect 19300 18912 19306 18964
rect 19334 18912 19340 18964
rect 19392 18952 19398 18964
rect 19613 18955 19671 18961
rect 19613 18952 19625 18955
rect 19392 18924 19625 18952
rect 19392 18912 19398 18924
rect 19613 18921 19625 18924
rect 19659 18921 19671 18955
rect 19613 18915 19671 18921
rect 20717 18955 20775 18961
rect 20717 18921 20729 18955
rect 20763 18952 20775 18955
rect 21266 18952 21272 18964
rect 20763 18924 21272 18952
rect 20763 18921 20775 18924
rect 20717 18915 20775 18921
rect 21266 18912 21272 18924
rect 21324 18912 21330 18964
rect 21726 18912 21732 18964
rect 21784 18952 21790 18964
rect 21913 18955 21971 18961
rect 21913 18952 21925 18955
rect 21784 18924 21925 18952
rect 21784 18912 21790 18924
rect 21913 18921 21925 18924
rect 21959 18921 21971 18955
rect 21913 18915 21971 18921
rect 22370 18912 22376 18964
rect 22428 18952 22434 18964
rect 22465 18955 22523 18961
rect 22465 18952 22477 18955
rect 22428 18924 22477 18952
rect 22428 18912 22434 18924
rect 22465 18921 22477 18924
rect 22511 18921 22523 18955
rect 22465 18915 22523 18921
rect 24026 18912 24032 18964
rect 24084 18952 24090 18964
rect 25041 18955 25099 18961
rect 25041 18952 25053 18955
rect 24084 18924 25053 18952
rect 24084 18912 24090 18924
rect 25041 18921 25053 18924
rect 25087 18921 25099 18955
rect 25041 18915 25099 18921
rect 18046 18884 18052 18896
rect 16868 18856 18052 18884
rect 11977 18847 12035 18853
rect 18046 18844 18052 18856
rect 18104 18884 18110 18896
rect 18785 18887 18843 18893
rect 18785 18884 18797 18887
rect 18104 18856 18797 18884
rect 18104 18844 18110 18856
rect 18785 18853 18797 18856
rect 18831 18853 18843 18887
rect 18785 18847 18843 18853
rect 21174 18844 21180 18896
rect 21232 18884 21238 18896
rect 22554 18884 22560 18896
rect 21232 18856 22560 18884
rect 21232 18844 21238 18856
rect 22554 18844 22560 18856
rect 22612 18884 22618 18896
rect 22925 18887 22983 18893
rect 22925 18884 22937 18887
rect 22612 18856 22937 18884
rect 22612 18844 22618 18856
rect 22925 18853 22937 18856
rect 22971 18853 22983 18887
rect 22925 18847 22983 18853
rect 23753 18887 23811 18893
rect 23753 18853 23765 18887
rect 23799 18884 23811 18887
rect 24210 18884 24216 18896
rect 23799 18856 24216 18884
rect 23799 18853 23811 18856
rect 23753 18847 23811 18853
rect 24210 18844 24216 18856
rect 24268 18844 24274 18896
rect 24854 18844 24860 18896
rect 24912 18884 24918 18896
rect 25409 18887 25467 18893
rect 25409 18884 25421 18887
rect 24912 18856 25421 18884
rect 24912 18844 24918 18856
rect 25409 18853 25421 18856
rect 25455 18853 25467 18887
rect 25409 18847 25467 18853
rect 4065 18819 4123 18825
rect 4065 18785 4077 18819
rect 4111 18816 4123 18819
rect 4706 18816 4712 18828
rect 4111 18788 4712 18816
rect 4111 18785 4123 18788
rect 4065 18779 4123 18785
rect 4706 18776 4712 18788
rect 4764 18776 4770 18828
rect 4798 18776 4804 18828
rect 4856 18816 4862 18828
rect 5629 18819 5687 18825
rect 5629 18816 5641 18819
rect 4856 18788 5641 18816
rect 4856 18776 4862 18788
rect 5629 18785 5641 18788
rect 5675 18785 5687 18819
rect 5629 18779 5687 18785
rect 5721 18819 5779 18825
rect 5721 18785 5733 18819
rect 5767 18816 5779 18819
rect 6270 18816 6276 18828
rect 5767 18788 6276 18816
rect 5767 18785 5779 18788
rect 5721 18779 5779 18785
rect 6270 18776 6276 18788
rect 6328 18776 6334 18828
rect 7098 18776 7104 18828
rect 7156 18816 7162 18828
rect 7193 18819 7251 18825
rect 7193 18816 7205 18819
rect 7156 18788 7205 18816
rect 7156 18776 7162 18788
rect 7193 18785 7205 18788
rect 7239 18816 7251 18819
rect 7742 18816 7748 18828
rect 7239 18788 7748 18816
rect 7239 18785 7251 18788
rect 7193 18779 7251 18785
rect 7742 18776 7748 18788
rect 7800 18776 7806 18828
rect 8389 18819 8447 18825
rect 8389 18785 8401 18819
rect 8435 18816 8447 18819
rect 8478 18816 8484 18828
rect 8435 18788 8484 18816
rect 8435 18785 8447 18788
rect 8389 18779 8447 18785
rect 8478 18776 8484 18788
rect 8536 18776 8542 18828
rect 9122 18776 9128 18828
rect 9180 18816 9186 18828
rect 9933 18819 9991 18825
rect 9933 18816 9945 18819
rect 9180 18788 9945 18816
rect 9180 18776 9186 18788
rect 9933 18785 9945 18788
rect 9979 18816 9991 18819
rect 11054 18816 11060 18828
rect 9979 18788 11060 18816
rect 9979 18785 9991 18788
rect 9933 18779 9991 18785
rect 11054 18776 11060 18788
rect 11112 18776 11118 18828
rect 11790 18776 11796 18828
rect 11848 18816 11854 18828
rect 12250 18816 12256 18828
rect 11848 18788 12256 18816
rect 11848 18776 11854 18788
rect 12250 18776 12256 18788
rect 12308 18816 12314 18828
rect 12434 18825 12440 18828
rect 12428 18816 12440 18825
rect 12308 18788 12440 18816
rect 12308 18776 12314 18788
rect 12428 18779 12440 18788
rect 12492 18816 12498 18828
rect 15657 18819 15715 18825
rect 12492 18788 12576 18816
rect 12434 18776 12440 18779
rect 12492 18776 12498 18788
rect 15657 18785 15669 18819
rect 15703 18816 15715 18819
rect 15838 18816 15844 18828
rect 15703 18788 15844 18816
rect 15703 18785 15715 18788
rect 15657 18779 15715 18785
rect 15838 18776 15844 18788
rect 15896 18776 15902 18828
rect 16022 18776 16028 18828
rect 16080 18816 16086 18828
rect 16206 18816 16212 18828
rect 16080 18788 16212 18816
rect 16080 18776 16086 18788
rect 16206 18776 16212 18788
rect 16264 18816 16270 18828
rect 16942 18816 16948 18828
rect 16264 18788 16948 18816
rect 16264 18776 16270 18788
rect 16942 18776 16948 18788
rect 17000 18776 17006 18828
rect 17221 18819 17279 18825
rect 17221 18785 17233 18819
rect 17267 18816 17279 18819
rect 17494 18816 17500 18828
rect 17267 18788 17500 18816
rect 17267 18785 17279 18788
rect 17221 18779 17279 18785
rect 17494 18776 17500 18788
rect 17552 18776 17558 18828
rect 21082 18776 21088 18828
rect 21140 18816 21146 18828
rect 21269 18819 21327 18825
rect 21269 18816 21281 18819
rect 21140 18788 21281 18816
rect 21140 18776 21146 18788
rect 21269 18785 21281 18788
rect 21315 18816 21327 18819
rect 21634 18816 21640 18828
rect 21315 18788 21640 18816
rect 21315 18785 21327 18788
rect 21269 18779 21327 18785
rect 21634 18776 21640 18788
rect 21692 18776 21698 18828
rect 22186 18776 22192 18828
rect 22244 18816 22250 18828
rect 22833 18819 22891 18825
rect 22833 18816 22845 18819
rect 22244 18788 22845 18816
rect 22244 18776 22250 18788
rect 22833 18785 22845 18788
rect 22879 18785 22891 18819
rect 22833 18779 22891 18785
rect 24118 18776 24124 18828
rect 24176 18816 24182 18828
rect 24397 18819 24455 18825
rect 24397 18816 24409 18819
rect 24176 18788 24409 18816
rect 24176 18776 24182 18788
rect 24397 18785 24409 18788
rect 24443 18785 24455 18819
rect 24397 18779 24455 18785
rect 3053 18751 3111 18757
rect 3053 18717 3065 18751
rect 3099 18748 3111 18751
rect 3418 18748 3424 18760
rect 3099 18720 3424 18748
rect 3099 18717 3111 18720
rect 3053 18711 3111 18717
rect 3418 18708 3424 18720
rect 3476 18708 3482 18760
rect 5169 18751 5227 18757
rect 5169 18717 5181 18751
rect 5215 18748 5227 18751
rect 5350 18748 5356 18760
rect 5215 18720 5356 18748
rect 5215 18717 5227 18720
rect 5169 18711 5227 18717
rect 5350 18708 5356 18720
rect 5408 18748 5414 18760
rect 5810 18748 5816 18760
rect 5408 18720 5816 18748
rect 5408 18708 5414 18720
rect 5810 18708 5816 18720
rect 5868 18708 5874 18760
rect 7374 18748 7380 18760
rect 7335 18720 7380 18748
rect 7374 18708 7380 18720
rect 7432 18708 7438 18760
rect 9582 18708 9588 18760
rect 9640 18748 9646 18760
rect 9677 18751 9735 18757
rect 9677 18748 9689 18751
rect 9640 18720 9689 18748
rect 9640 18708 9646 18720
rect 9677 18717 9689 18720
rect 9723 18717 9735 18751
rect 9677 18711 9735 18717
rect 12161 18751 12219 18757
rect 12161 18717 12173 18751
rect 12207 18717 12219 18751
rect 12161 18711 12219 18717
rect 1765 18683 1823 18689
rect 1765 18649 1777 18683
rect 1811 18680 1823 18683
rect 2682 18680 2688 18692
rect 1811 18652 2688 18680
rect 1811 18649 1823 18652
rect 1765 18643 1823 18649
rect 2682 18640 2688 18652
rect 2740 18640 2746 18692
rect 3142 18640 3148 18692
rect 3200 18680 3206 18692
rect 3697 18683 3755 18689
rect 3697 18680 3709 18683
rect 3200 18652 3709 18680
rect 3200 18640 3206 18652
rect 3697 18649 3709 18652
rect 3743 18680 3755 18683
rect 4154 18680 4160 18692
rect 3743 18652 4160 18680
rect 3743 18649 3755 18652
rect 3697 18643 3755 18649
rect 4154 18640 4160 18652
rect 4212 18680 4218 18692
rect 4709 18683 4767 18689
rect 4709 18680 4721 18683
rect 4212 18652 4721 18680
rect 4212 18640 4218 18652
rect 4709 18649 4721 18652
rect 4755 18680 4767 18683
rect 5442 18680 5448 18692
rect 4755 18652 5448 18680
rect 4755 18649 4767 18652
rect 4709 18643 4767 18649
rect 5442 18640 5448 18652
rect 5500 18640 5506 18692
rect 2130 18612 2136 18624
rect 2091 18584 2136 18612
rect 2130 18572 2136 18584
rect 2188 18572 2194 18624
rect 5258 18612 5264 18624
rect 5219 18584 5264 18612
rect 5258 18572 5264 18584
rect 5316 18572 5322 18624
rect 5534 18572 5540 18624
rect 5592 18612 5598 18624
rect 6273 18615 6331 18621
rect 6273 18612 6285 18615
rect 5592 18584 6285 18612
rect 5592 18572 5598 18584
rect 6273 18581 6285 18584
rect 6319 18581 6331 18615
rect 6822 18612 6828 18624
rect 6783 18584 6828 18612
rect 6273 18575 6331 18581
rect 6822 18572 6828 18584
rect 6880 18572 6886 18624
rect 7929 18615 7987 18621
rect 7929 18581 7941 18615
rect 7975 18612 7987 18615
rect 8018 18612 8024 18624
rect 7975 18584 8024 18612
rect 7975 18581 7987 18584
rect 7929 18575 7987 18581
rect 8018 18572 8024 18584
rect 8076 18572 8082 18624
rect 8294 18612 8300 18624
rect 8255 18584 8300 18612
rect 8294 18572 8300 18584
rect 8352 18572 8358 18624
rect 9122 18612 9128 18624
rect 9083 18584 9128 18612
rect 9122 18572 9128 18584
rect 9180 18572 9186 18624
rect 9692 18612 9720 18711
rect 11790 18680 11796 18692
rect 10612 18652 11796 18680
rect 10612 18612 10640 18652
rect 11790 18640 11796 18652
rect 11848 18680 11854 18692
rect 12176 18680 12204 18711
rect 14182 18708 14188 18760
rect 14240 18748 14246 18760
rect 14642 18748 14648 18760
rect 14240 18720 14648 18748
rect 14240 18708 14246 18720
rect 14642 18708 14648 18720
rect 14700 18748 14706 18760
rect 15749 18751 15807 18757
rect 15749 18748 15761 18751
rect 14700 18720 15761 18748
rect 14700 18708 14706 18720
rect 15749 18717 15761 18720
rect 15795 18717 15807 18751
rect 15749 18711 15807 18717
rect 15933 18751 15991 18757
rect 15933 18717 15945 18751
rect 15979 18748 15991 18751
rect 16482 18748 16488 18760
rect 15979 18720 16488 18748
rect 15979 18717 15991 18720
rect 15933 18711 15991 18717
rect 11848 18652 12204 18680
rect 11848 18640 11854 18652
rect 13722 18640 13728 18692
rect 13780 18680 13786 18692
rect 14461 18683 14519 18689
rect 14461 18680 14473 18683
rect 13780 18652 14473 18680
rect 13780 18640 13786 18652
rect 14461 18649 14473 18652
rect 14507 18649 14519 18683
rect 14461 18643 14519 18649
rect 14734 18640 14740 18692
rect 14792 18680 14798 18692
rect 15948 18680 15976 18711
rect 16482 18708 16488 18720
rect 16540 18708 16546 18760
rect 17313 18751 17371 18757
rect 17313 18717 17325 18751
rect 17359 18717 17371 18751
rect 17313 18711 17371 18717
rect 17405 18751 17463 18757
rect 17405 18717 17417 18751
rect 17451 18717 17463 18751
rect 17405 18711 17463 18717
rect 14792 18652 15976 18680
rect 14792 18640 14798 18652
rect 16758 18640 16764 18692
rect 16816 18680 16822 18692
rect 17328 18680 17356 18711
rect 16816 18652 17356 18680
rect 16816 18640 16822 18652
rect 9692 18584 10640 18612
rect 11422 18572 11428 18624
rect 11480 18612 11486 18624
rect 11609 18615 11667 18621
rect 11609 18612 11621 18615
rect 11480 18584 11621 18612
rect 11480 18572 11486 18584
rect 11609 18581 11621 18584
rect 11655 18581 11667 18615
rect 11609 18575 11667 18581
rect 11885 18615 11943 18621
rect 11885 18581 11897 18615
rect 11931 18612 11943 18615
rect 12434 18612 12440 18624
rect 11931 18584 12440 18612
rect 11931 18581 11943 18584
rect 11885 18575 11943 18581
rect 12434 18572 12440 18584
rect 12492 18572 12498 18624
rect 14185 18615 14243 18621
rect 14185 18581 14197 18615
rect 14231 18612 14243 18615
rect 14752 18612 14780 18640
rect 15286 18612 15292 18624
rect 14231 18584 14780 18612
rect 15247 18584 15292 18612
rect 14231 18581 14243 18584
rect 14185 18575 14243 18581
rect 15286 18572 15292 18584
rect 15344 18572 15350 18624
rect 16666 18612 16672 18624
rect 16627 18584 16672 18612
rect 16666 18572 16672 18584
rect 16724 18612 16730 18624
rect 17420 18612 17448 18711
rect 18598 18708 18604 18760
rect 18656 18748 18662 18760
rect 19061 18751 19119 18757
rect 19061 18748 19073 18751
rect 18656 18720 19073 18748
rect 18656 18708 18662 18720
rect 19061 18717 19073 18720
rect 19107 18748 19119 18751
rect 19610 18748 19616 18760
rect 19107 18720 19616 18748
rect 19107 18717 19119 18720
rect 19061 18711 19119 18717
rect 19610 18708 19616 18720
rect 19668 18708 19674 18760
rect 21358 18748 21364 18760
rect 21319 18720 21364 18748
rect 21358 18708 21364 18720
rect 21416 18708 21422 18760
rect 21542 18748 21548 18760
rect 21503 18720 21548 18748
rect 21542 18708 21548 18720
rect 21600 18708 21606 18760
rect 23014 18748 23020 18760
rect 22975 18720 23020 18748
rect 23014 18708 23020 18720
rect 23072 18708 23078 18760
rect 23474 18708 23480 18760
rect 23532 18748 23538 18760
rect 24489 18751 24547 18757
rect 24489 18748 24501 18751
rect 23532 18720 24501 18748
rect 23532 18708 23538 18720
rect 24489 18717 24501 18720
rect 24535 18717 24547 18751
rect 24489 18711 24547 18717
rect 24581 18751 24639 18757
rect 24581 18717 24593 18751
rect 24627 18717 24639 18751
rect 24581 18711 24639 18717
rect 21450 18680 21456 18692
rect 20272 18652 21456 18680
rect 18598 18612 18604 18624
rect 16724 18584 18604 18612
rect 16724 18572 16730 18584
rect 18598 18572 18604 18584
rect 18656 18572 18662 18624
rect 19426 18572 19432 18624
rect 19484 18612 19490 18624
rect 20272 18621 20300 18652
rect 21450 18640 21456 18652
rect 21508 18640 21514 18692
rect 23934 18640 23940 18692
rect 23992 18680 23998 18692
rect 24596 18680 24624 18711
rect 24946 18680 24952 18692
rect 23992 18652 24952 18680
rect 23992 18640 23998 18652
rect 24946 18640 24952 18652
rect 25004 18640 25010 18692
rect 20257 18615 20315 18621
rect 20257 18612 20269 18615
rect 19484 18584 20269 18612
rect 19484 18572 19490 18584
rect 20257 18581 20269 18584
rect 20303 18581 20315 18615
rect 20898 18612 20904 18624
rect 20859 18584 20904 18612
rect 20257 18575 20315 18581
rect 20898 18572 20904 18584
rect 20956 18572 20962 18624
rect 22373 18615 22431 18621
rect 22373 18581 22385 18615
rect 22419 18612 22431 18615
rect 23106 18612 23112 18624
rect 22419 18584 23112 18612
rect 22419 18581 22431 18584
rect 22373 18575 22431 18581
rect 23106 18572 23112 18584
rect 23164 18572 23170 18624
rect 23382 18572 23388 18624
rect 23440 18612 23446 18624
rect 23658 18612 23664 18624
rect 23440 18584 23664 18612
rect 23440 18572 23446 18584
rect 23658 18572 23664 18584
rect 23716 18572 23722 18624
rect 24029 18615 24087 18621
rect 24029 18581 24041 18615
rect 24075 18612 24087 18615
rect 25130 18612 25136 18624
rect 24075 18584 25136 18612
rect 24075 18581 24087 18584
rect 24029 18575 24087 18581
rect 25130 18572 25136 18584
rect 25188 18572 25194 18624
rect 25869 18615 25927 18621
rect 25869 18581 25881 18615
rect 25915 18612 25927 18615
rect 26142 18612 26148 18624
rect 25915 18584 26148 18612
rect 25915 18581 25927 18584
rect 25869 18575 25927 18581
rect 26142 18572 26148 18584
rect 26200 18572 26206 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 2041 18411 2099 18417
rect 2041 18377 2053 18411
rect 2087 18408 2099 18411
rect 2774 18408 2780 18420
rect 2087 18380 2780 18408
rect 2087 18377 2099 18380
rect 2041 18371 2099 18377
rect 2774 18368 2780 18380
rect 2832 18368 2838 18420
rect 3142 18408 3148 18420
rect 3103 18380 3148 18408
rect 3142 18368 3148 18380
rect 3200 18368 3206 18420
rect 3510 18368 3516 18420
rect 3568 18408 3574 18420
rect 3605 18411 3663 18417
rect 3605 18408 3617 18411
rect 3568 18380 3617 18408
rect 3568 18368 3574 18380
rect 3605 18377 3617 18380
rect 3651 18377 3663 18411
rect 3605 18371 3663 18377
rect 6273 18411 6331 18417
rect 6273 18377 6285 18411
rect 6319 18408 6331 18411
rect 6730 18408 6736 18420
rect 6319 18380 6736 18408
rect 6319 18377 6331 18380
rect 6273 18371 6331 18377
rect 6730 18368 6736 18380
rect 6788 18408 6794 18420
rect 7374 18408 7380 18420
rect 6788 18380 7380 18408
rect 6788 18368 6794 18380
rect 7374 18368 7380 18380
rect 7432 18368 7438 18420
rect 10505 18411 10563 18417
rect 10505 18377 10517 18411
rect 10551 18408 10563 18411
rect 10686 18408 10692 18420
rect 10551 18380 10692 18408
rect 10551 18377 10563 18380
rect 10505 18371 10563 18377
rect 10686 18368 10692 18380
rect 10744 18368 10750 18420
rect 11514 18408 11520 18420
rect 11475 18380 11520 18408
rect 11514 18368 11520 18380
rect 11572 18368 11578 18420
rect 12621 18411 12679 18417
rect 12621 18377 12633 18411
rect 12667 18408 12679 18411
rect 12802 18408 12808 18420
rect 12667 18380 12808 18408
rect 12667 18377 12679 18380
rect 12621 18371 12679 18377
rect 12802 18368 12808 18380
rect 12860 18368 12866 18420
rect 13354 18408 13360 18420
rect 13315 18380 13360 18408
rect 13354 18368 13360 18380
rect 13412 18368 13418 18420
rect 18049 18411 18107 18417
rect 18049 18377 18061 18411
rect 18095 18408 18107 18411
rect 19058 18408 19064 18420
rect 18095 18380 19064 18408
rect 18095 18377 18107 18380
rect 18049 18371 18107 18377
rect 19058 18368 19064 18380
rect 19116 18368 19122 18420
rect 21542 18368 21548 18420
rect 21600 18408 21606 18420
rect 21637 18411 21695 18417
rect 21637 18408 21649 18411
rect 21600 18380 21649 18408
rect 21600 18368 21606 18380
rect 21637 18377 21649 18380
rect 21683 18377 21695 18411
rect 21637 18371 21695 18377
rect 22094 18368 22100 18420
rect 22152 18408 22158 18420
rect 22152 18380 24256 18408
rect 22152 18368 22158 18380
rect 2038 18232 2044 18284
rect 2096 18272 2102 18284
rect 2501 18275 2559 18281
rect 2501 18272 2513 18275
rect 2096 18244 2513 18272
rect 2096 18232 2102 18244
rect 2501 18241 2513 18244
rect 2547 18241 2559 18275
rect 2501 18235 2559 18241
rect 2685 18275 2743 18281
rect 2685 18241 2697 18275
rect 2731 18272 2743 18275
rect 3160 18272 3188 18368
rect 5169 18343 5227 18349
rect 5169 18340 5181 18343
rect 4080 18312 5181 18340
rect 2731 18244 3188 18272
rect 2731 18241 2743 18244
rect 2685 18235 2743 18241
rect 3694 18232 3700 18284
rect 3752 18272 3758 18284
rect 4080 18281 4108 18312
rect 5169 18309 5181 18312
rect 5215 18309 5227 18343
rect 12250 18340 12256 18352
rect 12163 18312 12256 18340
rect 5169 18303 5227 18309
rect 12250 18300 12256 18312
rect 12308 18340 12314 18352
rect 12894 18340 12900 18352
rect 12308 18312 12900 18340
rect 12308 18300 12314 18312
rect 12894 18300 12900 18312
rect 12952 18300 12958 18352
rect 4065 18275 4123 18281
rect 4065 18272 4077 18275
rect 3752 18244 4077 18272
rect 3752 18232 3758 18244
rect 4065 18241 4077 18244
rect 4111 18241 4123 18275
rect 4065 18235 4123 18241
rect 4157 18275 4215 18281
rect 4157 18241 4169 18275
rect 4203 18241 4215 18275
rect 4157 18235 4215 18241
rect 2409 18207 2467 18213
rect 2409 18173 2421 18207
rect 2455 18204 2467 18207
rect 2590 18204 2596 18216
rect 2455 18176 2596 18204
rect 2455 18173 2467 18176
rect 2409 18167 2467 18173
rect 2590 18164 2596 18176
rect 2648 18164 2654 18216
rect 3513 18207 3571 18213
rect 3513 18173 3525 18207
rect 3559 18204 3571 18207
rect 3970 18204 3976 18216
rect 3559 18176 3976 18204
rect 3559 18173 3571 18176
rect 3513 18167 3571 18173
rect 3970 18164 3976 18176
rect 4028 18204 4034 18216
rect 4172 18204 4200 18235
rect 4522 18232 4528 18284
rect 4580 18272 4586 18284
rect 4982 18272 4988 18284
rect 4580 18244 4988 18272
rect 4580 18232 4586 18244
rect 4982 18232 4988 18244
rect 5040 18232 5046 18284
rect 5350 18232 5356 18284
rect 5408 18272 5414 18284
rect 5810 18272 5816 18284
rect 5408 18244 5816 18272
rect 5408 18232 5414 18244
rect 5810 18232 5816 18244
rect 5868 18232 5874 18284
rect 10686 18232 10692 18284
rect 10744 18272 10750 18284
rect 11057 18275 11115 18281
rect 11057 18272 11069 18275
rect 10744 18244 11069 18272
rect 10744 18232 10750 18244
rect 11057 18241 11069 18244
rect 11103 18272 11115 18275
rect 11422 18272 11428 18284
rect 11103 18244 11428 18272
rect 11103 18241 11115 18244
rect 11057 18235 11115 18241
rect 11422 18232 11428 18244
rect 11480 18232 11486 18284
rect 13372 18272 13400 18368
rect 16850 18340 16856 18352
rect 16811 18312 16856 18340
rect 16850 18300 16856 18312
rect 16908 18300 16914 18352
rect 16942 18300 16948 18352
rect 17000 18340 17006 18352
rect 18877 18343 18935 18349
rect 18877 18340 18889 18343
rect 17000 18312 18889 18340
rect 17000 18300 17006 18312
rect 18877 18309 18889 18312
rect 18923 18309 18935 18343
rect 22922 18340 22928 18352
rect 22883 18312 22928 18340
rect 18877 18303 18935 18309
rect 22922 18300 22928 18312
rect 22980 18300 22986 18352
rect 14001 18275 14059 18281
rect 14001 18272 14013 18275
rect 13372 18244 14013 18272
rect 14001 18241 14013 18244
rect 14047 18241 14059 18275
rect 14001 18235 14059 18241
rect 14185 18275 14243 18281
rect 14185 18241 14197 18275
rect 14231 18272 14243 18275
rect 14734 18272 14740 18284
rect 14231 18244 14740 18272
rect 14231 18241 14243 18244
rect 14185 18235 14243 18241
rect 14734 18232 14740 18244
rect 14792 18232 14798 18284
rect 15470 18272 15476 18284
rect 15431 18244 15476 18272
rect 15470 18232 15476 18244
rect 15528 18232 15534 18284
rect 18598 18272 18604 18284
rect 18559 18244 18604 18272
rect 18598 18232 18604 18244
rect 18656 18272 18662 18284
rect 19061 18275 19119 18281
rect 19061 18272 19073 18275
rect 18656 18244 19073 18272
rect 18656 18232 18662 18244
rect 19061 18241 19073 18244
rect 19107 18241 19119 18275
rect 19061 18235 19119 18241
rect 19613 18275 19671 18281
rect 19613 18241 19625 18275
rect 19659 18272 19671 18275
rect 19659 18244 19840 18272
rect 19659 18241 19671 18244
rect 19613 18235 19671 18241
rect 4706 18204 4712 18216
rect 4028 18176 4200 18204
rect 4667 18176 4712 18204
rect 4028 18164 4034 18176
rect 4706 18164 4712 18176
rect 4764 18164 4770 18216
rect 5537 18207 5595 18213
rect 5537 18173 5549 18207
rect 5583 18204 5595 18207
rect 6362 18204 6368 18216
rect 5583 18176 6368 18204
rect 5583 18173 5595 18176
rect 5537 18167 5595 18173
rect 6362 18164 6368 18176
rect 6420 18164 6426 18216
rect 6641 18207 6699 18213
rect 6641 18173 6653 18207
rect 6687 18204 6699 18207
rect 7650 18204 7656 18216
rect 6687 18176 7656 18204
rect 6687 18173 6699 18176
rect 6641 18167 6699 18173
rect 7650 18164 7656 18176
rect 7708 18164 7714 18216
rect 7745 18207 7803 18213
rect 7745 18173 7757 18207
rect 7791 18204 7803 18207
rect 9582 18204 9588 18216
rect 7791 18176 9588 18204
rect 7791 18173 7803 18176
rect 7745 18167 7803 18173
rect 9582 18164 9588 18176
rect 9640 18164 9646 18216
rect 10413 18207 10471 18213
rect 10413 18173 10425 18207
rect 10459 18204 10471 18207
rect 10873 18207 10931 18213
rect 10873 18204 10885 18207
rect 10459 18176 10885 18204
rect 10459 18173 10471 18176
rect 10413 18167 10471 18173
rect 10873 18173 10885 18176
rect 10919 18204 10931 18207
rect 12425 18207 12483 18213
rect 10919 18176 11805 18204
rect 10919 18173 10931 18176
rect 10873 18167 10931 18173
rect 5629 18139 5687 18145
rect 5629 18105 5641 18139
rect 5675 18136 5687 18139
rect 6086 18136 6092 18148
rect 5675 18108 6092 18136
rect 5675 18105 5687 18108
rect 5629 18099 5687 18105
rect 6086 18096 6092 18108
rect 6144 18096 6150 18148
rect 8018 18145 8024 18148
rect 8012 18136 8024 18145
rect 7979 18108 8024 18136
rect 8012 18099 8024 18108
rect 8018 18096 8024 18099
rect 8076 18096 8082 18148
rect 11777 18136 11805 18176
rect 12425 18173 12437 18207
rect 12471 18173 12483 18207
rect 12425 18167 12483 18173
rect 12452 18136 12480 18167
rect 13538 18164 13544 18216
rect 13596 18204 13602 18216
rect 13909 18207 13967 18213
rect 13909 18204 13921 18207
rect 13596 18176 13921 18204
rect 13596 18164 13602 18176
rect 13909 18173 13921 18176
rect 13955 18204 13967 18207
rect 14553 18207 14611 18213
rect 14553 18204 14565 18207
rect 13955 18176 14565 18204
rect 13955 18173 13967 18176
rect 13909 18167 13967 18173
rect 14553 18173 14565 18176
rect 14599 18173 14611 18207
rect 15488 18204 15516 18232
rect 16482 18204 16488 18216
rect 15488 18176 16488 18204
rect 14553 18167 14611 18173
rect 16482 18164 16488 18176
rect 16540 18164 16546 18216
rect 18230 18164 18236 18216
rect 18288 18204 18294 18216
rect 18417 18207 18475 18213
rect 18417 18204 18429 18207
rect 18288 18176 18429 18204
rect 18288 18164 18294 18176
rect 18417 18173 18429 18176
rect 18463 18173 18475 18207
rect 18417 18167 18475 18173
rect 19705 18207 19763 18213
rect 19705 18173 19717 18207
rect 19751 18173 19763 18207
rect 19812 18204 19840 18244
rect 23658 18232 23664 18284
rect 23716 18272 23722 18284
rect 24228 18281 24256 18380
rect 24946 18368 24952 18420
rect 25004 18408 25010 18420
rect 25041 18411 25099 18417
rect 25041 18408 25053 18411
rect 25004 18380 25053 18408
rect 25004 18368 25010 18380
rect 25041 18377 25053 18380
rect 25087 18377 25099 18411
rect 25041 18371 25099 18377
rect 25409 18411 25467 18417
rect 25409 18377 25421 18411
rect 25455 18408 25467 18411
rect 25498 18408 25504 18420
rect 25455 18380 25504 18408
rect 25455 18377 25467 18380
rect 25409 18371 25467 18377
rect 25498 18368 25504 18380
rect 25556 18368 25562 18420
rect 24121 18275 24179 18281
rect 24121 18272 24133 18275
rect 23716 18244 24133 18272
rect 23716 18232 23722 18244
rect 24121 18241 24133 18244
rect 24167 18241 24179 18275
rect 24121 18235 24179 18241
rect 24213 18275 24271 18281
rect 24213 18241 24225 18275
rect 24259 18241 24271 18275
rect 24213 18235 24271 18241
rect 19978 18213 19984 18216
rect 19972 18204 19984 18213
rect 19812 18176 19984 18204
rect 19705 18167 19763 18173
rect 19972 18167 19984 18176
rect 15740 18139 15798 18145
rect 11777 18108 13032 18136
rect 13004 18080 13032 18108
rect 15740 18105 15752 18139
rect 15786 18136 15798 18139
rect 16298 18136 16304 18148
rect 15786 18108 16304 18136
rect 15786 18105 15798 18108
rect 15740 18099 15798 18105
rect 16298 18096 16304 18108
rect 16356 18096 16362 18148
rect 17494 18136 17500 18148
rect 17455 18108 17500 18136
rect 17494 18096 17500 18108
rect 17552 18096 17558 18148
rect 18598 18096 18604 18148
rect 18656 18136 18662 18148
rect 19334 18136 19340 18148
rect 18656 18108 19340 18136
rect 18656 18096 18662 18108
rect 19334 18096 19340 18108
rect 19392 18136 19398 18148
rect 19720 18136 19748 18167
rect 19978 18164 19984 18167
rect 20036 18164 20042 18216
rect 22189 18207 22247 18213
rect 22189 18173 22201 18207
rect 22235 18204 22247 18207
rect 22370 18204 22376 18216
rect 22235 18176 22376 18204
rect 22235 18173 22247 18176
rect 22189 18167 22247 18173
rect 22370 18164 22376 18176
rect 22428 18164 22434 18216
rect 23474 18164 23480 18216
rect 23532 18204 23538 18216
rect 25225 18207 25283 18213
rect 25225 18204 25237 18207
rect 23532 18176 25237 18204
rect 23532 18164 23538 18176
rect 25225 18173 25237 18176
rect 25271 18204 25283 18207
rect 25777 18207 25835 18213
rect 25777 18204 25789 18207
rect 25271 18176 25789 18204
rect 25271 18173 25283 18176
rect 25225 18167 25283 18173
rect 25777 18173 25789 18176
rect 25823 18173 25835 18207
rect 25777 18167 25835 18173
rect 20898 18136 20904 18148
rect 19392 18108 20904 18136
rect 19392 18096 19398 18108
rect 20898 18096 20904 18108
rect 20956 18096 20962 18148
rect 21818 18096 21824 18148
rect 21876 18136 21882 18148
rect 22465 18139 22523 18145
rect 22465 18136 22477 18139
rect 21876 18108 22477 18136
rect 21876 18096 21882 18108
rect 22465 18105 22477 18108
rect 22511 18105 22523 18139
rect 22465 18099 22523 18105
rect 24029 18139 24087 18145
rect 24029 18105 24041 18139
rect 24075 18136 24087 18139
rect 24210 18136 24216 18148
rect 24075 18108 24216 18136
rect 24075 18105 24087 18108
rect 24029 18099 24087 18105
rect 24210 18096 24216 18108
rect 24268 18136 24274 18148
rect 26418 18136 26424 18148
rect 24268 18108 26424 18136
rect 24268 18096 24274 18108
rect 26418 18096 26424 18108
rect 26476 18096 26482 18148
rect 1670 18068 1676 18080
rect 1631 18040 1676 18068
rect 1670 18028 1676 18040
rect 1728 18028 1734 18080
rect 3973 18071 4031 18077
rect 3973 18037 3985 18071
rect 4019 18068 4031 18071
rect 4154 18068 4160 18080
rect 4019 18040 4160 18068
rect 4019 18037 4031 18040
rect 3973 18031 4031 18037
rect 4154 18028 4160 18040
rect 4212 18028 4218 18080
rect 4798 18028 4804 18080
rect 4856 18068 4862 18080
rect 5077 18071 5135 18077
rect 5077 18068 5089 18071
rect 4856 18040 5089 18068
rect 4856 18028 4862 18040
rect 5077 18037 5089 18040
rect 5123 18068 5135 18071
rect 5166 18068 5172 18080
rect 5123 18040 5172 18068
rect 5123 18037 5135 18040
rect 5077 18031 5135 18037
rect 5166 18028 5172 18040
rect 5224 18028 5230 18080
rect 7098 18068 7104 18080
rect 7059 18040 7104 18068
rect 7098 18028 7104 18040
rect 7156 18028 7162 18080
rect 7653 18071 7711 18077
rect 7653 18037 7665 18071
rect 7699 18068 7711 18071
rect 8478 18068 8484 18080
rect 7699 18040 8484 18068
rect 7699 18037 7711 18040
rect 7653 18031 7711 18037
rect 8478 18028 8484 18040
rect 8536 18028 8542 18080
rect 9122 18068 9128 18080
rect 9083 18040 9128 18068
rect 9122 18028 9128 18040
rect 9180 18028 9186 18080
rect 10045 18071 10103 18077
rect 10045 18037 10057 18071
rect 10091 18068 10103 18071
rect 10962 18068 10968 18080
rect 10091 18040 10968 18068
rect 10091 18037 10103 18040
rect 10045 18031 10103 18037
rect 10962 18028 10968 18040
rect 11020 18028 11026 18080
rect 12986 18068 12992 18080
rect 12947 18040 12992 18068
rect 12986 18028 12992 18040
rect 13044 18028 13050 18080
rect 13538 18068 13544 18080
rect 13499 18040 13544 18068
rect 13538 18028 13544 18040
rect 13596 18028 13602 18080
rect 14642 18028 14648 18080
rect 14700 18068 14706 18080
rect 14921 18071 14979 18077
rect 14921 18068 14933 18071
rect 14700 18040 14933 18068
rect 14700 18028 14706 18040
rect 14921 18037 14933 18040
rect 14967 18037 14979 18071
rect 14921 18031 14979 18037
rect 15381 18071 15439 18077
rect 15381 18037 15393 18071
rect 15427 18068 15439 18071
rect 15838 18068 15844 18080
rect 15427 18040 15844 18068
rect 15427 18037 15439 18040
rect 15381 18031 15439 18037
rect 15838 18028 15844 18040
rect 15896 18068 15902 18080
rect 16390 18068 16396 18080
rect 15896 18040 16396 18068
rect 15896 18028 15902 18040
rect 16390 18028 16396 18040
rect 16448 18028 16454 18080
rect 17862 18068 17868 18080
rect 17823 18040 17868 18068
rect 17862 18028 17868 18040
rect 17920 18068 17926 18080
rect 18509 18071 18567 18077
rect 18509 18068 18521 18071
rect 17920 18040 18521 18068
rect 17920 18028 17926 18040
rect 18509 18037 18521 18040
rect 18555 18037 18567 18071
rect 18509 18031 18567 18037
rect 18877 18071 18935 18077
rect 18877 18037 18889 18071
rect 18923 18068 18935 18071
rect 20714 18068 20720 18080
rect 18923 18040 20720 18068
rect 18923 18037 18935 18040
rect 18877 18031 18935 18037
rect 20714 18028 20720 18040
rect 20772 18028 20778 18080
rect 21085 18071 21143 18077
rect 21085 18037 21097 18071
rect 21131 18068 21143 18071
rect 21266 18068 21272 18080
rect 21131 18040 21272 18068
rect 21131 18037 21143 18040
rect 21085 18031 21143 18037
rect 21266 18028 21272 18040
rect 21324 18028 21330 18080
rect 21450 18028 21456 18080
rect 21508 18068 21514 18080
rect 23474 18068 23480 18080
rect 21508 18040 23480 18068
rect 21508 18028 21514 18040
rect 23474 18028 23480 18040
rect 23532 18028 23538 18080
rect 23661 18071 23719 18077
rect 23661 18037 23673 18071
rect 23707 18068 23719 18071
rect 23750 18068 23756 18080
rect 23707 18040 23756 18068
rect 23707 18037 23719 18040
rect 23661 18031 23719 18037
rect 23750 18028 23756 18040
rect 23808 18028 23814 18080
rect 24118 18028 24124 18080
rect 24176 18068 24182 18080
rect 24673 18071 24731 18077
rect 24673 18068 24685 18071
rect 24176 18040 24685 18068
rect 24176 18028 24182 18040
rect 24673 18037 24685 18040
rect 24719 18037 24731 18071
rect 26234 18068 26240 18080
rect 26195 18040 26240 18068
rect 24673 18031 24731 18037
rect 26234 18028 26240 18040
rect 26292 18028 26298 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 2409 17867 2467 17873
rect 2409 17833 2421 17867
rect 2455 17864 2467 17867
rect 2590 17864 2596 17876
rect 2455 17836 2596 17864
rect 2455 17833 2467 17836
rect 2409 17827 2467 17833
rect 2590 17824 2596 17836
rect 2648 17824 2654 17876
rect 3418 17864 3424 17876
rect 3379 17836 3424 17864
rect 3418 17824 3424 17836
rect 3476 17824 3482 17876
rect 5442 17824 5448 17876
rect 5500 17864 5506 17876
rect 5537 17867 5595 17873
rect 5537 17864 5549 17867
rect 5500 17836 5549 17864
rect 5500 17824 5506 17836
rect 5537 17833 5549 17836
rect 5583 17833 5595 17867
rect 5537 17827 5595 17833
rect 6549 17867 6607 17873
rect 6549 17833 6561 17867
rect 6595 17864 6607 17867
rect 6822 17864 6828 17876
rect 6595 17836 6828 17864
rect 6595 17833 6607 17836
rect 6549 17827 6607 17833
rect 6822 17824 6828 17836
rect 6880 17864 6886 17876
rect 7101 17867 7159 17873
rect 7101 17864 7113 17867
rect 6880 17836 7113 17864
rect 6880 17824 6886 17836
rect 7101 17833 7113 17836
rect 7147 17833 7159 17867
rect 10686 17864 10692 17876
rect 10647 17836 10692 17864
rect 7101 17827 7159 17833
rect 10686 17824 10692 17836
rect 10744 17824 10750 17876
rect 11241 17867 11299 17873
rect 11241 17833 11253 17867
rect 11287 17864 11299 17867
rect 12342 17864 12348 17876
rect 11287 17836 12348 17864
rect 11287 17833 11299 17836
rect 11241 17827 11299 17833
rect 12342 17824 12348 17836
rect 12400 17824 12406 17876
rect 13538 17824 13544 17876
rect 13596 17864 13602 17876
rect 14093 17867 14151 17873
rect 14093 17864 14105 17867
rect 13596 17836 14105 17864
rect 13596 17824 13602 17836
rect 14093 17833 14105 17836
rect 14139 17833 14151 17867
rect 14093 17827 14151 17833
rect 14734 17824 14740 17876
rect 14792 17864 14798 17876
rect 15013 17867 15071 17873
rect 15013 17864 15025 17867
rect 14792 17836 15025 17864
rect 14792 17824 14798 17836
rect 15013 17833 15025 17836
rect 15059 17833 15071 17867
rect 15286 17864 15292 17876
rect 15247 17836 15292 17864
rect 15013 17827 15071 17833
rect 15286 17824 15292 17836
rect 15344 17824 15350 17876
rect 15930 17864 15936 17876
rect 15580 17836 15936 17864
rect 5810 17756 5816 17808
rect 5868 17796 5874 17808
rect 6181 17799 6239 17805
rect 6181 17796 6193 17799
rect 5868 17768 6193 17796
rect 5868 17756 5874 17768
rect 6181 17765 6193 17768
rect 6227 17796 6239 17799
rect 8018 17796 8024 17808
rect 6227 17768 8024 17796
rect 6227 17765 6239 17768
rect 6181 17759 6239 17765
rect 8018 17756 8024 17768
rect 8076 17756 8082 17808
rect 8481 17799 8539 17805
rect 8481 17765 8493 17799
rect 8527 17796 8539 17799
rect 10870 17796 10876 17808
rect 8527 17768 10876 17796
rect 8527 17765 8539 17768
rect 8481 17759 8539 17765
rect 10870 17756 10876 17768
rect 10928 17796 10934 17808
rect 11057 17799 11115 17805
rect 11057 17796 11069 17799
rect 10928 17768 11069 17796
rect 10928 17756 10934 17768
rect 11057 17765 11069 17768
rect 11103 17765 11115 17799
rect 11057 17759 11115 17765
rect 11514 17756 11520 17808
rect 11572 17796 11578 17808
rect 11609 17799 11667 17805
rect 11609 17796 11621 17799
rect 11572 17768 11621 17796
rect 11572 17756 11578 17768
rect 11609 17765 11621 17768
rect 11655 17765 11667 17799
rect 11609 17759 11667 17765
rect 11698 17756 11704 17808
rect 11756 17796 11762 17808
rect 11756 17768 11801 17796
rect 11756 17756 11762 17768
rect 12434 17756 12440 17808
rect 12492 17796 12498 17808
rect 12897 17799 12955 17805
rect 12897 17796 12909 17799
rect 12492 17768 12909 17796
rect 12492 17756 12498 17768
rect 12897 17765 12909 17768
rect 12943 17796 12955 17799
rect 13265 17799 13323 17805
rect 13265 17796 13277 17799
rect 12943 17768 13277 17796
rect 12943 17765 12955 17768
rect 12897 17759 12955 17765
rect 13265 17765 13277 17768
rect 13311 17796 13323 17799
rect 13722 17796 13728 17808
rect 13311 17768 13728 17796
rect 13311 17765 13323 17768
rect 13265 17759 13323 17765
rect 13722 17756 13728 17768
rect 13780 17756 13786 17808
rect 13998 17796 14004 17808
rect 13911 17768 14004 17796
rect 13998 17756 14004 17768
rect 14056 17796 14062 17808
rect 15102 17796 15108 17808
rect 14056 17768 15108 17796
rect 14056 17756 14062 17768
rect 15102 17756 15108 17768
rect 15160 17756 15166 17808
rect 15580 17796 15608 17836
rect 15930 17824 15936 17836
rect 15988 17864 15994 17876
rect 17402 17864 17408 17876
rect 15988 17836 17408 17864
rect 15988 17824 15994 17836
rect 17402 17824 17408 17836
rect 17460 17824 17466 17876
rect 18325 17867 18383 17873
rect 18325 17833 18337 17867
rect 18371 17864 18383 17867
rect 18414 17864 18420 17876
rect 18371 17836 18420 17864
rect 18371 17833 18383 17836
rect 18325 17827 18383 17833
rect 18414 17824 18420 17836
rect 18472 17824 18478 17876
rect 19334 17824 19340 17876
rect 19392 17864 19398 17876
rect 20257 17867 20315 17873
rect 20257 17864 20269 17867
rect 19392 17836 20269 17864
rect 19392 17824 19398 17836
rect 20257 17833 20269 17836
rect 20303 17833 20315 17867
rect 20257 17827 20315 17833
rect 22097 17867 22155 17873
rect 22097 17833 22109 17867
rect 22143 17864 22155 17867
rect 22186 17864 22192 17876
rect 22143 17836 22192 17864
rect 22143 17833 22155 17836
rect 22097 17827 22155 17833
rect 22186 17824 22192 17836
rect 22244 17824 22250 17876
rect 22465 17867 22523 17873
rect 22465 17833 22477 17867
rect 22511 17864 22523 17867
rect 22554 17864 22560 17876
rect 22511 17836 22560 17864
rect 22511 17833 22523 17836
rect 22465 17827 22523 17833
rect 22554 17824 22560 17836
rect 22612 17824 22618 17876
rect 24026 17864 24032 17876
rect 22664 17836 24032 17864
rect 15304 17768 15608 17796
rect 15304 17740 15332 17768
rect 16850 17756 16856 17808
rect 16908 17796 16914 17808
rect 17190 17799 17248 17805
rect 17190 17796 17202 17799
rect 16908 17768 17202 17796
rect 16908 17756 16914 17768
rect 17190 17765 17202 17768
rect 17236 17765 17248 17799
rect 17190 17759 17248 17765
rect 19242 17756 19248 17808
rect 19300 17796 19306 17808
rect 21450 17796 21456 17808
rect 19300 17768 21456 17796
rect 19300 17756 19306 17768
rect 21450 17756 21456 17768
rect 21508 17756 21514 17808
rect 22002 17756 22008 17808
rect 22060 17796 22066 17808
rect 22664 17796 22692 17836
rect 24026 17824 24032 17836
rect 24084 17864 24090 17876
rect 24581 17867 24639 17873
rect 24581 17864 24593 17867
rect 24084 17836 24593 17864
rect 24084 17824 24090 17836
rect 24581 17833 24593 17836
rect 24627 17833 24639 17867
rect 26326 17864 26332 17876
rect 26287 17836 26332 17864
rect 24581 17827 24639 17833
rect 26326 17824 26332 17836
rect 26384 17824 26390 17876
rect 23106 17796 23112 17808
rect 22060 17768 22692 17796
rect 22756 17768 23112 17796
rect 22060 17756 22066 17768
rect 2774 17688 2780 17740
rect 2832 17728 2838 17740
rect 4430 17737 4436 17740
rect 4424 17728 4436 17737
rect 2832 17700 2877 17728
rect 3068 17700 4436 17728
rect 2832 17688 2838 17700
rect 1397 17663 1455 17669
rect 1397 17629 1409 17663
rect 1443 17660 1455 17663
rect 2222 17660 2228 17672
rect 1443 17632 2228 17660
rect 1443 17629 1455 17632
rect 1397 17623 1455 17629
rect 2222 17620 2228 17632
rect 2280 17620 2286 17672
rect 2498 17620 2504 17672
rect 2556 17660 2562 17672
rect 3068 17669 3096 17700
rect 4424 17691 4436 17700
rect 4430 17688 4436 17691
rect 4488 17688 4494 17740
rect 6638 17688 6644 17740
rect 6696 17728 6702 17740
rect 6822 17728 6828 17740
rect 6696 17700 6828 17728
rect 6696 17688 6702 17700
rect 6822 17688 6828 17700
rect 6880 17688 6886 17740
rect 7006 17728 7012 17740
rect 6967 17700 7012 17728
rect 7006 17688 7012 17700
rect 7064 17688 7070 17740
rect 8110 17688 8116 17740
rect 8168 17728 8174 17740
rect 8205 17731 8263 17737
rect 8205 17728 8217 17731
rect 8168 17700 8217 17728
rect 8168 17688 8174 17700
rect 8205 17697 8217 17700
rect 8251 17697 8263 17731
rect 8205 17691 8263 17697
rect 9122 17688 9128 17740
rect 9180 17728 9186 17740
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 9180 17700 10057 17728
rect 9180 17688 9186 17700
rect 10045 17697 10057 17700
rect 10091 17697 10103 17731
rect 10045 17691 10103 17697
rect 10137 17731 10195 17737
rect 10137 17697 10149 17731
rect 10183 17728 10195 17731
rect 10410 17728 10416 17740
rect 10183 17700 10416 17728
rect 10183 17697 10195 17700
rect 10137 17691 10195 17697
rect 10410 17688 10416 17700
rect 10468 17688 10474 17740
rect 13630 17688 13636 17740
rect 13688 17688 13694 17740
rect 15286 17688 15292 17740
rect 15344 17688 15350 17740
rect 15470 17688 15476 17740
rect 15528 17728 15534 17740
rect 15657 17731 15715 17737
rect 15657 17728 15669 17731
rect 15528 17700 15669 17728
rect 15528 17688 15534 17700
rect 15657 17697 15669 17700
rect 15703 17697 15715 17731
rect 15657 17691 15715 17697
rect 16482 17688 16488 17740
rect 16540 17728 16546 17740
rect 16945 17731 17003 17737
rect 16945 17728 16957 17731
rect 16540 17700 16957 17728
rect 16540 17688 16546 17700
rect 16945 17697 16957 17700
rect 16991 17728 17003 17731
rect 17494 17728 17500 17740
rect 16991 17700 17500 17728
rect 16991 17697 17003 17700
rect 16945 17691 17003 17697
rect 17494 17688 17500 17700
rect 17552 17688 17558 17740
rect 19518 17728 19524 17740
rect 19479 17700 19524 17728
rect 19518 17688 19524 17700
rect 19576 17688 19582 17740
rect 20717 17731 20775 17737
rect 20717 17697 20729 17731
rect 20763 17728 20775 17731
rect 21361 17731 21419 17737
rect 21361 17728 21373 17731
rect 20763 17700 21373 17728
rect 20763 17697 20775 17700
rect 20717 17691 20775 17697
rect 21361 17697 21373 17700
rect 21407 17728 21419 17731
rect 21542 17728 21548 17740
rect 21407 17700 21548 17728
rect 21407 17697 21419 17700
rect 21361 17691 21419 17697
rect 21542 17688 21548 17700
rect 21600 17688 21606 17740
rect 22462 17688 22468 17740
rect 22520 17728 22526 17740
rect 22756 17728 22784 17768
rect 23106 17756 23112 17768
rect 23164 17756 23170 17808
rect 23658 17796 23664 17808
rect 23619 17768 23664 17796
rect 23658 17756 23664 17768
rect 23716 17756 23722 17808
rect 24670 17756 24676 17808
rect 24728 17796 24734 17808
rect 25222 17796 25228 17808
rect 24728 17768 25228 17796
rect 24728 17756 24734 17768
rect 25222 17756 25228 17768
rect 25280 17756 25286 17808
rect 22922 17728 22928 17740
rect 22520 17700 22784 17728
rect 22883 17700 22928 17728
rect 22520 17688 22526 17700
rect 22922 17688 22928 17700
rect 22980 17688 22986 17740
rect 24489 17731 24547 17737
rect 24489 17697 24501 17731
rect 24535 17728 24547 17731
rect 24762 17728 24768 17740
rect 24535 17700 24768 17728
rect 24535 17697 24547 17700
rect 24489 17691 24547 17697
rect 24762 17688 24768 17700
rect 24820 17688 24826 17740
rect 2869 17663 2927 17669
rect 2869 17660 2881 17663
rect 2556 17632 2881 17660
rect 2556 17620 2562 17632
rect 2869 17629 2881 17632
rect 2915 17629 2927 17663
rect 2869 17623 2927 17629
rect 3053 17663 3111 17669
rect 3053 17629 3065 17663
rect 3099 17629 3111 17663
rect 3053 17623 3111 17629
rect 4157 17663 4215 17669
rect 4157 17629 4169 17663
rect 4203 17629 4215 17663
rect 4157 17623 4215 17629
rect 2682 17552 2688 17604
rect 2740 17592 2746 17604
rect 3068 17592 3096 17623
rect 2740 17564 3096 17592
rect 2740 17552 2746 17564
rect 1946 17524 1952 17536
rect 1907 17496 1952 17524
rect 1946 17484 1952 17496
rect 2004 17484 2010 17536
rect 2317 17527 2375 17533
rect 2317 17493 2329 17527
rect 2363 17524 2375 17527
rect 2590 17524 2596 17536
rect 2363 17496 2596 17524
rect 2363 17493 2375 17496
rect 2317 17487 2375 17493
rect 2590 17484 2596 17496
rect 2648 17484 2654 17536
rect 3602 17484 3608 17536
rect 3660 17524 3666 17536
rect 3789 17527 3847 17533
rect 3789 17524 3801 17527
rect 3660 17496 3801 17524
rect 3660 17484 3666 17496
rect 3789 17493 3801 17496
rect 3835 17493 3847 17527
rect 4172 17524 4200 17623
rect 6086 17620 6092 17672
rect 6144 17660 6150 17672
rect 7193 17663 7251 17669
rect 7193 17660 7205 17663
rect 6144 17632 7205 17660
rect 6144 17620 6150 17632
rect 7193 17629 7205 17632
rect 7239 17660 7251 17663
rect 7466 17660 7472 17672
rect 7239 17632 7472 17660
rect 7239 17629 7251 17632
rect 7193 17623 7251 17629
rect 7466 17620 7472 17632
rect 7524 17620 7530 17672
rect 10226 17660 10232 17672
rect 10187 17632 10232 17660
rect 10226 17620 10232 17632
rect 10284 17620 10290 17672
rect 11054 17620 11060 17672
rect 11112 17660 11118 17672
rect 11793 17663 11851 17669
rect 11793 17660 11805 17663
rect 11112 17632 11805 17660
rect 11112 17620 11118 17632
rect 11793 17629 11805 17632
rect 11839 17629 11851 17663
rect 11793 17623 11851 17629
rect 12710 17620 12716 17672
rect 12768 17660 12774 17672
rect 12986 17660 12992 17672
rect 12768 17632 12992 17660
rect 12768 17620 12774 17632
rect 12986 17620 12992 17632
rect 13044 17620 13050 17672
rect 13648 17660 13676 17688
rect 14277 17663 14335 17669
rect 13648 17632 13860 17660
rect 7374 17552 7380 17604
rect 7432 17592 7438 17604
rect 7745 17595 7803 17601
rect 7745 17592 7757 17595
rect 7432 17564 7757 17592
rect 7432 17552 7438 17564
rect 7745 17561 7757 17564
rect 7791 17592 7803 17595
rect 8846 17592 8852 17604
rect 7791 17564 8852 17592
rect 7791 17561 7803 17564
rect 7745 17555 7803 17561
rect 8846 17552 8852 17564
rect 8904 17552 8910 17604
rect 9306 17592 9312 17604
rect 9267 17564 9312 17592
rect 9306 17552 9312 17564
rect 9364 17552 9370 17604
rect 13630 17592 13636 17604
rect 13591 17564 13636 17592
rect 13630 17552 13636 17564
rect 13688 17552 13694 17604
rect 13832 17536 13860 17632
rect 14277 17629 14289 17663
rect 14323 17660 14335 17663
rect 14458 17660 14464 17672
rect 14323 17632 14464 17660
rect 14323 17629 14335 17632
rect 14277 17623 14335 17629
rect 14458 17620 14464 17632
rect 14516 17620 14522 17672
rect 15746 17660 15752 17672
rect 15707 17632 15752 17660
rect 15746 17620 15752 17632
rect 15804 17620 15810 17672
rect 15933 17663 15991 17669
rect 15933 17629 15945 17663
rect 15979 17660 15991 17663
rect 16022 17660 16028 17672
rect 15979 17632 16028 17660
rect 15979 17629 15991 17632
rect 15933 17623 15991 17629
rect 16022 17620 16028 17632
rect 16080 17620 16086 17672
rect 19702 17660 19708 17672
rect 19663 17632 19708 17660
rect 19702 17620 19708 17632
rect 19760 17620 19766 17672
rect 21450 17660 21456 17672
rect 21411 17632 21456 17660
rect 21450 17620 21456 17632
rect 21508 17620 21514 17672
rect 21637 17663 21695 17669
rect 21637 17629 21649 17663
rect 21683 17660 21695 17663
rect 22002 17660 22008 17672
rect 21683 17632 22008 17660
rect 21683 17629 21695 17632
rect 21637 17623 21695 17629
rect 22002 17620 22008 17632
rect 22060 17620 22066 17672
rect 23014 17660 23020 17672
rect 22975 17632 23020 17660
rect 23014 17620 23020 17632
rect 23072 17620 23078 17672
rect 23106 17620 23112 17672
rect 23164 17660 23170 17672
rect 24670 17660 24676 17672
rect 23164 17632 23209 17660
rect 24631 17632 24676 17660
rect 23164 17620 23170 17632
rect 24670 17620 24676 17632
rect 24728 17620 24734 17672
rect 14737 17595 14795 17601
rect 14737 17561 14749 17595
rect 14783 17592 14795 17595
rect 16666 17592 16672 17604
rect 14783 17564 16672 17592
rect 14783 17561 14795 17564
rect 14737 17555 14795 17561
rect 16666 17552 16672 17564
rect 16724 17552 16730 17604
rect 19337 17595 19395 17601
rect 19337 17561 19349 17595
rect 19383 17592 19395 17595
rect 19610 17592 19616 17604
rect 19383 17564 19616 17592
rect 19383 17561 19395 17564
rect 19337 17555 19395 17561
rect 19610 17552 19616 17564
rect 19668 17592 19674 17604
rect 21174 17592 21180 17604
rect 19668 17564 21180 17592
rect 19668 17552 19674 17564
rect 21174 17552 21180 17564
rect 21232 17552 21238 17604
rect 21468 17592 21496 17620
rect 22557 17595 22615 17601
rect 22557 17592 22569 17595
rect 21468 17564 22569 17592
rect 22557 17561 22569 17564
rect 22603 17561 22615 17595
rect 22557 17555 22615 17561
rect 24121 17595 24179 17601
rect 24121 17561 24133 17595
rect 24167 17592 24179 17595
rect 24946 17592 24952 17604
rect 24167 17564 24952 17592
rect 24167 17561 24179 17564
rect 24121 17555 24179 17561
rect 24946 17552 24952 17564
rect 25004 17552 25010 17604
rect 5074 17524 5080 17536
rect 4172 17496 5080 17524
rect 3789 17487 3847 17493
rect 5074 17484 5080 17496
rect 5132 17484 5138 17536
rect 6638 17524 6644 17536
rect 6599 17496 6644 17524
rect 6638 17484 6644 17496
rect 6696 17484 6702 17536
rect 8113 17527 8171 17533
rect 8113 17493 8125 17527
rect 8159 17524 8171 17527
rect 8202 17524 8208 17536
rect 8159 17496 8208 17524
rect 8159 17493 8171 17496
rect 8113 17487 8171 17493
rect 8202 17484 8208 17496
rect 8260 17484 8266 17536
rect 8938 17524 8944 17536
rect 8899 17496 8944 17524
rect 8938 17484 8944 17496
rect 8996 17484 9002 17536
rect 9674 17524 9680 17536
rect 9635 17496 9680 17524
rect 9674 17484 9680 17496
rect 9732 17484 9738 17536
rect 12529 17527 12587 17533
rect 12529 17493 12541 17527
rect 12575 17524 12587 17527
rect 12710 17524 12716 17536
rect 12575 17496 12716 17524
rect 12575 17493 12587 17496
rect 12529 17487 12587 17493
rect 12710 17484 12716 17496
rect 12768 17484 12774 17536
rect 13078 17484 13084 17536
rect 13136 17524 13142 17536
rect 13354 17524 13360 17536
rect 13136 17496 13360 17524
rect 13136 17484 13142 17496
rect 13354 17484 13360 17496
rect 13412 17484 13418 17536
rect 13814 17484 13820 17536
rect 13872 17484 13878 17536
rect 16298 17524 16304 17536
rect 16259 17496 16304 17524
rect 16298 17484 16304 17496
rect 16356 17484 16362 17536
rect 16758 17524 16764 17536
rect 16719 17496 16764 17524
rect 16758 17484 16764 17496
rect 16816 17484 16822 17536
rect 18966 17524 18972 17536
rect 18927 17496 18972 17524
rect 18966 17484 18972 17496
rect 19024 17484 19030 17536
rect 20990 17524 20996 17536
rect 20951 17496 20996 17524
rect 20990 17484 20996 17496
rect 21048 17484 21054 17536
rect 24210 17484 24216 17536
rect 24268 17524 24274 17536
rect 25133 17527 25191 17533
rect 25133 17524 25145 17527
rect 24268 17496 25145 17524
rect 24268 17484 24274 17496
rect 25133 17493 25145 17496
rect 25179 17493 25191 17527
rect 25133 17487 25191 17493
rect 25593 17527 25651 17533
rect 25593 17493 25605 17527
rect 25639 17524 25651 17527
rect 25869 17527 25927 17533
rect 25869 17524 25881 17527
rect 25639 17496 25881 17524
rect 25639 17493 25651 17496
rect 25593 17487 25651 17493
rect 25869 17493 25881 17496
rect 25915 17524 25927 17527
rect 26142 17524 26148 17536
rect 25915 17496 26148 17524
rect 25915 17493 25927 17496
rect 25869 17487 25927 17493
rect 26142 17484 26148 17496
rect 26200 17484 26206 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 2774 17280 2780 17332
rect 2832 17320 2838 17332
rect 2832 17292 2877 17320
rect 2832 17280 2838 17292
rect 4430 17280 4436 17332
rect 4488 17320 4494 17332
rect 5721 17323 5779 17329
rect 5721 17320 5733 17323
rect 4488 17292 5733 17320
rect 4488 17280 4494 17292
rect 5721 17289 5733 17292
rect 5767 17289 5779 17323
rect 5721 17283 5779 17289
rect 6641 17323 6699 17329
rect 6641 17289 6653 17323
rect 6687 17320 6699 17323
rect 7006 17320 7012 17332
rect 6687 17292 7012 17320
rect 6687 17289 6699 17292
rect 6641 17283 6699 17289
rect 7006 17280 7012 17292
rect 7064 17280 7070 17332
rect 8018 17280 8024 17332
rect 8076 17320 8082 17332
rect 8205 17323 8263 17329
rect 8205 17320 8217 17323
rect 8076 17292 8217 17320
rect 8076 17280 8082 17292
rect 8205 17289 8217 17292
rect 8251 17289 8263 17323
rect 8205 17283 8263 17289
rect 9214 17280 9220 17332
rect 9272 17320 9278 17332
rect 9272 17292 11008 17320
rect 9272 17280 9278 17292
rect 4614 17252 4620 17264
rect 4575 17224 4620 17252
rect 4614 17212 4620 17224
rect 4672 17252 4678 17264
rect 4672 17224 5212 17252
rect 4672 17212 4678 17224
rect 1670 17144 1676 17196
rect 1728 17184 1734 17196
rect 2041 17187 2099 17193
rect 2041 17184 2053 17187
rect 1728 17156 2053 17184
rect 1728 17144 1734 17156
rect 2041 17153 2053 17156
rect 2087 17184 2099 17187
rect 2958 17184 2964 17196
rect 2087 17156 2964 17184
rect 2087 17153 2099 17156
rect 2041 17147 2099 17153
rect 2958 17144 2964 17156
rect 3016 17144 3022 17196
rect 3510 17144 3516 17196
rect 3568 17184 3574 17196
rect 3697 17187 3755 17193
rect 3697 17184 3709 17187
rect 3568 17156 3709 17184
rect 3568 17144 3574 17156
rect 3697 17153 3709 17156
rect 3743 17153 3755 17187
rect 3697 17147 3755 17153
rect 5074 17144 5080 17196
rect 5132 17144 5138 17196
rect 5184 17193 5212 17224
rect 9766 17212 9772 17264
rect 9824 17252 9830 17264
rect 9950 17252 9956 17264
rect 9824 17224 9956 17252
rect 9824 17212 9830 17224
rect 9950 17212 9956 17224
rect 10008 17212 10014 17264
rect 10410 17252 10416 17264
rect 10371 17224 10416 17252
rect 10410 17212 10416 17224
rect 10468 17212 10474 17264
rect 5169 17187 5227 17193
rect 5169 17153 5181 17187
rect 5215 17153 5227 17187
rect 5169 17147 5227 17153
rect 5258 17144 5264 17196
rect 5316 17184 5322 17196
rect 6086 17184 6092 17196
rect 5316 17156 6092 17184
rect 5316 17144 5322 17156
rect 6086 17144 6092 17156
rect 6144 17184 6150 17196
rect 6181 17187 6239 17193
rect 6181 17184 6193 17187
rect 6144 17156 6193 17184
rect 6144 17144 6150 17156
rect 6181 17153 6193 17156
rect 6227 17184 6239 17187
rect 6270 17184 6276 17196
rect 6227 17156 6276 17184
rect 6227 17153 6239 17156
rect 6181 17147 6239 17153
rect 6270 17144 6276 17156
rect 6328 17144 6334 17196
rect 8849 17187 8907 17193
rect 8849 17153 8861 17187
rect 8895 17184 8907 17187
rect 9582 17184 9588 17196
rect 8895 17156 9588 17184
rect 8895 17153 8907 17156
rect 8849 17147 8907 17153
rect 9582 17144 9588 17156
rect 9640 17184 9646 17196
rect 9861 17187 9919 17193
rect 9861 17184 9873 17187
rect 9640 17156 9873 17184
rect 9640 17144 9646 17156
rect 9861 17153 9873 17156
rect 9907 17184 9919 17187
rect 10226 17184 10232 17196
rect 9907 17156 10232 17184
rect 9907 17153 9919 17156
rect 9861 17147 9919 17153
rect 10226 17144 10232 17156
rect 10284 17184 10290 17196
rect 10689 17187 10747 17193
rect 10689 17184 10701 17187
rect 10284 17156 10701 17184
rect 10284 17144 10290 17156
rect 10689 17153 10701 17156
rect 10735 17153 10747 17187
rect 10980 17184 11008 17292
rect 11054 17280 11060 17332
rect 11112 17320 11118 17332
rect 11425 17323 11483 17329
rect 11425 17320 11437 17323
rect 11112 17292 11437 17320
rect 11112 17280 11118 17292
rect 11425 17289 11437 17292
rect 11471 17289 11483 17323
rect 11425 17283 11483 17289
rect 14182 17280 14188 17332
rect 14240 17320 14246 17332
rect 14553 17323 14611 17329
rect 14553 17320 14565 17323
rect 14240 17292 14565 17320
rect 14240 17280 14246 17292
rect 14553 17289 14565 17292
rect 14599 17320 14611 17323
rect 15470 17320 15476 17332
rect 14599 17292 15476 17320
rect 14599 17289 14611 17292
rect 14553 17283 14611 17289
rect 15470 17280 15476 17292
rect 15528 17280 15534 17332
rect 16117 17323 16175 17329
rect 16117 17289 16129 17323
rect 16163 17320 16175 17323
rect 16298 17320 16304 17332
rect 16163 17292 16304 17320
rect 16163 17289 16175 17292
rect 16117 17283 16175 17289
rect 16298 17280 16304 17292
rect 16356 17280 16362 17332
rect 16850 17280 16856 17332
rect 16908 17320 16914 17332
rect 16945 17323 17003 17329
rect 16945 17320 16957 17323
rect 16908 17292 16957 17320
rect 16908 17280 16914 17292
rect 16945 17289 16957 17292
rect 16991 17289 17003 17323
rect 16945 17283 17003 17289
rect 17954 17280 17960 17332
rect 18012 17320 18018 17332
rect 18049 17323 18107 17329
rect 18049 17320 18061 17323
rect 18012 17292 18061 17320
rect 18012 17280 18018 17292
rect 18049 17289 18061 17292
rect 18095 17289 18107 17323
rect 19702 17320 19708 17332
rect 19663 17292 19708 17320
rect 18049 17283 18107 17289
rect 19702 17280 19708 17292
rect 19760 17280 19766 17332
rect 19981 17323 20039 17329
rect 19981 17289 19993 17323
rect 20027 17320 20039 17323
rect 20070 17320 20076 17332
rect 20027 17292 20076 17320
rect 20027 17289 20039 17292
rect 19981 17283 20039 17289
rect 20070 17280 20076 17292
rect 20128 17280 20134 17332
rect 23566 17280 23572 17332
rect 23624 17320 23630 17332
rect 23661 17323 23719 17329
rect 23661 17320 23673 17323
rect 23624 17292 23673 17320
rect 23624 17280 23630 17292
rect 23661 17289 23673 17292
rect 23707 17289 23719 17323
rect 23661 17283 23719 17289
rect 23750 17280 23756 17332
rect 23808 17320 23814 17332
rect 24026 17320 24032 17332
rect 23808 17292 24032 17320
rect 23808 17280 23814 17292
rect 24026 17280 24032 17292
rect 24084 17320 24090 17332
rect 24673 17323 24731 17329
rect 24673 17320 24685 17323
rect 24084 17292 24685 17320
rect 24084 17280 24090 17292
rect 24673 17289 24685 17292
rect 24719 17289 24731 17323
rect 24673 17283 24731 17289
rect 24762 17280 24768 17332
rect 24820 17320 24826 17332
rect 25041 17323 25099 17329
rect 25041 17320 25053 17323
rect 24820 17292 25053 17320
rect 24820 17280 24826 17292
rect 25041 17289 25053 17292
rect 25087 17289 25099 17323
rect 25041 17283 25099 17289
rect 12526 17212 12532 17264
rect 12584 17252 12590 17264
rect 12802 17252 12808 17264
rect 12584 17224 12808 17252
rect 12584 17212 12590 17224
rect 12802 17212 12808 17224
rect 12860 17212 12866 17264
rect 13078 17212 13084 17264
rect 13136 17252 13142 17264
rect 13262 17252 13268 17264
rect 13136 17224 13268 17252
rect 13136 17212 13142 17224
rect 13262 17212 13268 17224
rect 13320 17212 13326 17264
rect 17221 17255 17279 17261
rect 17221 17221 17233 17255
rect 17267 17252 17279 17255
rect 17494 17252 17500 17264
rect 17267 17224 17500 17252
rect 17267 17221 17279 17224
rect 17221 17215 17279 17221
rect 11054 17184 11060 17196
rect 10980 17156 11060 17184
rect 10689 17147 10747 17153
rect 11054 17144 11060 17156
rect 11112 17144 11118 17196
rect 12250 17184 12256 17196
rect 12163 17156 12256 17184
rect 12250 17144 12256 17156
rect 12308 17184 12314 17196
rect 12989 17187 13047 17193
rect 12989 17184 13001 17187
rect 12308 17156 13001 17184
rect 12308 17144 12314 17156
rect 12989 17153 13001 17156
rect 13035 17153 13047 17187
rect 12989 17147 13047 17153
rect 13814 17144 13820 17196
rect 13872 17184 13878 17196
rect 14737 17187 14795 17193
rect 14737 17184 14749 17187
rect 13872 17156 14749 17184
rect 13872 17144 13878 17156
rect 14737 17153 14749 17156
rect 14783 17153 14795 17187
rect 14737 17147 14795 17153
rect 1765 17119 1823 17125
rect 1765 17085 1777 17119
rect 1811 17116 1823 17119
rect 2590 17116 2596 17128
rect 1811 17088 2596 17116
rect 1811 17085 1823 17088
rect 1765 17079 1823 17085
rect 2590 17076 2596 17088
rect 2648 17076 2654 17128
rect 3234 17076 3240 17128
rect 3292 17116 3298 17128
rect 3418 17116 3424 17128
rect 3292 17088 3424 17116
rect 3292 17076 3298 17088
rect 3418 17076 3424 17088
rect 3476 17076 3482 17128
rect 5092 17116 5120 17144
rect 6825 17119 6883 17125
rect 6825 17116 6837 17119
rect 5092 17088 6837 17116
rect 6825 17085 6837 17088
rect 6871 17085 6883 17119
rect 6825 17079 6883 17085
rect 7092 17119 7150 17125
rect 7092 17085 7104 17119
rect 7138 17116 7150 17119
rect 7374 17116 7380 17128
rect 7138 17088 7380 17116
rect 7138 17085 7150 17088
rect 7092 17079 7150 17085
rect 7374 17076 7380 17088
rect 7432 17076 7438 17128
rect 9306 17076 9312 17128
rect 9364 17116 9370 17128
rect 9677 17119 9735 17125
rect 9677 17116 9689 17119
rect 9364 17088 9689 17116
rect 9364 17076 9370 17088
rect 9677 17085 9689 17088
rect 9723 17085 9735 17119
rect 10870 17116 10876 17128
rect 10831 17088 10876 17116
rect 9677 17079 9735 17085
rect 10870 17076 10876 17088
rect 10928 17076 10934 17128
rect 12710 17076 12716 17128
rect 12768 17116 12774 17128
rect 12897 17119 12955 17125
rect 12897 17116 12909 17119
rect 12768 17088 12909 17116
rect 12768 17076 12774 17088
rect 12897 17085 12909 17088
rect 12943 17085 12955 17119
rect 14752 17116 14780 17147
rect 17236 17116 17264 17215
rect 17494 17212 17500 17224
rect 17552 17252 17558 17264
rect 17552 17224 19656 17252
rect 17552 17212 17558 17224
rect 18693 17187 18751 17193
rect 18693 17153 18705 17187
rect 18739 17184 18751 17187
rect 18966 17184 18972 17196
rect 18739 17156 18972 17184
rect 18739 17153 18751 17156
rect 18693 17147 18751 17153
rect 18966 17144 18972 17156
rect 19024 17144 19030 17196
rect 17402 17116 17408 17128
rect 14752 17088 17264 17116
rect 17363 17088 17408 17116
rect 12897 17079 12955 17085
rect 17402 17076 17408 17088
rect 17460 17076 17466 17128
rect 18417 17119 18475 17125
rect 18417 17085 18429 17119
rect 18463 17116 18475 17119
rect 19242 17116 19248 17128
rect 18463 17088 19248 17116
rect 18463 17085 18475 17088
rect 18417 17079 18475 17085
rect 1118 17008 1124 17060
rect 1176 17048 1182 17060
rect 2498 17048 2504 17060
rect 1176 17020 2504 17048
rect 1176 17008 1182 17020
rect 2498 17008 2504 17020
rect 2556 17008 2562 17060
rect 5077 17051 5135 17057
rect 5077 17048 5089 17051
rect 4356 17020 5089 17048
rect 4356 16992 4384 17020
rect 5077 17017 5089 17020
rect 5123 17017 5135 17051
rect 5077 17011 5135 17017
rect 8386 17008 8392 17060
rect 8444 17048 8450 17060
rect 9769 17051 9827 17057
rect 9769 17048 9781 17051
rect 8444 17020 9781 17048
rect 8444 17008 8450 17020
rect 9769 17017 9781 17020
rect 9815 17017 9827 17051
rect 9769 17011 9827 17017
rect 11885 17051 11943 17057
rect 11885 17017 11897 17051
rect 11931 17048 11943 17051
rect 12342 17048 12348 17060
rect 11931 17020 12348 17048
rect 11931 17017 11943 17020
rect 11885 17011 11943 17017
rect 12342 17008 12348 17020
rect 12400 17048 12406 17060
rect 12805 17051 12863 17057
rect 12805 17048 12817 17051
rect 12400 17020 12817 17048
rect 12400 17008 12406 17020
rect 12805 17017 12817 17020
rect 12851 17017 12863 17051
rect 12805 17011 12863 17017
rect 13725 17051 13783 17057
rect 13725 17017 13737 17051
rect 13771 17048 13783 17051
rect 14277 17051 14335 17057
rect 14277 17048 14289 17051
rect 13771 17020 14289 17048
rect 13771 17017 13783 17020
rect 13725 17011 13783 17017
rect 14277 17017 14289 17020
rect 14323 17048 14335 17051
rect 14458 17048 14464 17060
rect 14323 17020 14464 17048
rect 14323 17017 14335 17020
rect 14277 17011 14335 17017
rect 14458 17008 14464 17020
rect 14516 17048 14522 17060
rect 15004 17051 15062 17057
rect 15004 17048 15016 17051
rect 14516 17020 15016 17048
rect 14516 17008 14522 17020
rect 15004 17017 15016 17020
rect 15050 17048 15062 17051
rect 15102 17048 15108 17060
rect 15050 17020 15108 17048
rect 15050 17017 15062 17020
rect 15004 17011 15062 17017
rect 15102 17008 15108 17020
rect 15160 17008 15166 17060
rect 17865 17051 17923 17057
rect 17865 17017 17877 17051
rect 17911 17048 17923 17051
rect 17911 17020 18552 17048
rect 17911 17017 17923 17020
rect 17865 17011 17923 17017
rect 18524 16992 18552 17020
rect 18984 16992 19012 17088
rect 19242 17076 19248 17088
rect 19300 17076 19306 17128
rect 19628 17048 19656 17224
rect 19720 17116 19748 17280
rect 21910 17212 21916 17264
rect 21968 17252 21974 17264
rect 23477 17255 23535 17261
rect 23477 17252 23489 17255
rect 21968 17224 23489 17252
rect 21968 17212 21974 17224
rect 23477 17221 23489 17224
rect 23523 17221 23535 17255
rect 23477 17215 23535 17221
rect 19797 17119 19855 17125
rect 19797 17116 19809 17119
rect 19720 17088 19809 17116
rect 19797 17085 19809 17088
rect 19843 17085 19855 17119
rect 20898 17116 20904 17128
rect 20859 17088 20904 17116
rect 19797 17079 19855 17085
rect 20898 17076 20904 17088
rect 20956 17076 20962 17128
rect 22554 17076 22560 17128
rect 22612 17116 22618 17128
rect 23492 17116 23520 17215
rect 24210 17184 24216 17196
rect 24171 17156 24216 17184
rect 24210 17144 24216 17156
rect 24268 17144 24274 17196
rect 24118 17116 24124 17128
rect 22612 17088 23244 17116
rect 23492 17088 24124 17116
rect 22612 17076 22618 17088
rect 20809 17051 20867 17057
rect 19628 17020 20668 17048
rect 1397 16983 1455 16989
rect 1397 16949 1409 16983
rect 1443 16980 1455 16983
rect 1670 16980 1676 16992
rect 1443 16952 1676 16980
rect 1443 16949 1455 16952
rect 1397 16943 1455 16949
rect 1670 16940 1676 16952
rect 1728 16940 1734 16992
rect 1857 16983 1915 16989
rect 1857 16949 1869 16983
rect 1903 16980 1915 16983
rect 1946 16980 1952 16992
rect 1903 16952 1952 16980
rect 1903 16949 1915 16952
rect 1857 16943 1915 16949
rect 1946 16940 1952 16952
rect 2004 16940 2010 16992
rect 3050 16940 3056 16992
rect 3108 16980 3114 16992
rect 3145 16983 3203 16989
rect 3145 16980 3157 16983
rect 3108 16952 3157 16980
rect 3108 16940 3114 16952
rect 3145 16949 3157 16952
rect 3191 16949 3203 16983
rect 3145 16943 3203 16949
rect 3234 16940 3240 16992
rect 3292 16980 3298 16992
rect 3513 16983 3571 16989
rect 3513 16980 3525 16983
rect 3292 16952 3525 16980
rect 3292 16940 3298 16952
rect 3513 16949 3525 16952
rect 3559 16949 3571 16983
rect 3513 16943 3571 16949
rect 3602 16940 3608 16992
rect 3660 16980 3666 16992
rect 4249 16983 4307 16989
rect 3660 16952 3705 16980
rect 3660 16940 3666 16952
rect 4249 16949 4261 16983
rect 4295 16980 4307 16983
rect 4338 16980 4344 16992
rect 4295 16952 4344 16980
rect 4295 16949 4307 16952
rect 4249 16943 4307 16949
rect 4338 16940 4344 16952
rect 4396 16940 4402 16992
rect 4706 16980 4712 16992
rect 4667 16952 4712 16980
rect 4706 16940 4712 16952
rect 4764 16940 4770 16992
rect 8662 16940 8668 16992
rect 8720 16980 8726 16992
rect 9122 16980 9128 16992
rect 8720 16952 9128 16980
rect 8720 16940 8726 16952
rect 9122 16940 9128 16952
rect 9180 16940 9186 16992
rect 9214 16940 9220 16992
rect 9272 16980 9278 16992
rect 9309 16983 9367 16989
rect 9309 16980 9321 16983
rect 9272 16952 9321 16980
rect 9272 16940 9278 16952
rect 9309 16949 9321 16952
rect 9355 16949 9367 16983
rect 9309 16943 9367 16949
rect 10778 16940 10784 16992
rect 10836 16980 10842 16992
rect 11057 16983 11115 16989
rect 11057 16980 11069 16983
rect 10836 16952 11069 16980
rect 10836 16940 10842 16952
rect 11057 16949 11069 16952
rect 11103 16949 11115 16983
rect 11057 16943 11115 16949
rect 12434 16940 12440 16992
rect 12492 16980 12498 16992
rect 12492 16952 12537 16980
rect 12492 16940 12498 16952
rect 18506 16940 18512 16992
rect 18564 16980 18570 16992
rect 18564 16952 18609 16980
rect 18564 16940 18570 16952
rect 18966 16940 18972 16992
rect 19024 16980 19030 16992
rect 19061 16983 19119 16989
rect 19061 16980 19073 16983
rect 19024 16952 19073 16980
rect 19024 16940 19030 16952
rect 19061 16949 19073 16952
rect 19107 16949 19119 16983
rect 20438 16980 20444 16992
rect 20399 16952 20444 16980
rect 19061 16943 19119 16949
rect 20438 16940 20444 16952
rect 20496 16940 20502 16992
rect 20640 16980 20668 17020
rect 20809 17017 20821 17051
rect 20855 17048 20867 17051
rect 21146 17051 21204 17057
rect 21146 17048 21158 17051
rect 20855 17020 21158 17048
rect 20855 17017 20867 17020
rect 20809 17011 20867 17017
rect 21146 17017 21158 17020
rect 21192 17048 21204 17051
rect 22370 17048 22376 17060
rect 21192 17020 22376 17048
rect 21192 17017 21204 17020
rect 21146 17011 21204 17017
rect 22370 17008 22376 17020
rect 22428 17048 22434 17060
rect 23106 17048 23112 17060
rect 22428 17020 23112 17048
rect 22428 17008 22434 17020
rect 23106 17008 23112 17020
rect 23164 17008 23170 17060
rect 23216 17048 23244 17088
rect 24118 17076 24124 17088
rect 24176 17076 24182 17128
rect 25225 17119 25283 17125
rect 25225 17085 25237 17119
rect 25271 17116 25283 17119
rect 25271 17088 25544 17116
rect 25271 17085 25283 17088
rect 25225 17079 25283 17085
rect 24029 17051 24087 17057
rect 24029 17048 24041 17051
rect 23216 17020 24041 17048
rect 24029 17017 24041 17020
rect 24075 17048 24087 17051
rect 24394 17048 24400 17060
rect 24075 17020 24400 17048
rect 24075 17017 24087 17020
rect 24029 17011 24087 17017
rect 24394 17008 24400 17020
rect 24452 17008 24458 17060
rect 25516 16992 25544 17088
rect 21358 16980 21364 16992
rect 20640 16952 21364 16980
rect 21358 16940 21364 16952
rect 21416 16940 21422 16992
rect 22002 16940 22008 16992
rect 22060 16980 22066 16992
rect 22281 16983 22339 16989
rect 22281 16980 22293 16983
rect 22060 16952 22293 16980
rect 22060 16940 22066 16952
rect 22281 16949 22293 16952
rect 22327 16949 22339 16983
rect 22281 16943 22339 16949
rect 22554 16940 22560 16992
rect 22612 16980 22618 16992
rect 22830 16980 22836 16992
rect 22612 16952 22836 16980
rect 22612 16940 22618 16952
rect 22830 16940 22836 16952
rect 22888 16940 22894 16992
rect 22922 16940 22928 16992
rect 22980 16980 22986 16992
rect 22980 16952 23025 16980
rect 22980 16940 22986 16952
rect 24302 16940 24308 16992
rect 24360 16980 24366 16992
rect 25222 16980 25228 16992
rect 24360 16952 25228 16980
rect 24360 16940 24366 16952
rect 25222 16940 25228 16952
rect 25280 16940 25286 16992
rect 25406 16980 25412 16992
rect 25367 16952 25412 16980
rect 25406 16940 25412 16952
rect 25464 16940 25470 16992
rect 25498 16940 25504 16992
rect 25556 16980 25562 16992
rect 25777 16983 25835 16989
rect 25777 16980 25789 16983
rect 25556 16952 25789 16980
rect 25556 16940 25562 16952
rect 25777 16949 25789 16952
rect 25823 16949 25835 16983
rect 26142 16980 26148 16992
rect 26103 16952 26148 16980
rect 25777 16943 25835 16949
rect 26142 16940 26148 16952
rect 26200 16940 26206 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 2501 16779 2559 16785
rect 2501 16745 2513 16779
rect 2547 16776 2559 16779
rect 2682 16776 2688 16788
rect 2547 16748 2688 16776
rect 2547 16745 2559 16748
rect 2501 16739 2559 16745
rect 2682 16736 2688 16748
rect 2740 16736 2746 16788
rect 2774 16736 2780 16788
rect 2832 16776 2838 16788
rect 2961 16779 3019 16785
rect 2961 16776 2973 16779
rect 2832 16748 2973 16776
rect 2832 16736 2838 16748
rect 2961 16745 2973 16748
rect 3007 16745 3019 16779
rect 3510 16776 3516 16788
rect 3471 16748 3516 16776
rect 2961 16739 3019 16745
rect 3510 16736 3516 16748
rect 3568 16736 3574 16788
rect 4525 16779 4583 16785
rect 4525 16745 4537 16779
rect 4571 16776 4583 16779
rect 5629 16779 5687 16785
rect 5629 16776 5641 16779
rect 4571 16748 5641 16776
rect 4571 16745 4583 16748
rect 4525 16739 4583 16745
rect 5629 16745 5641 16748
rect 5675 16776 5687 16779
rect 6086 16776 6092 16788
rect 5675 16748 6092 16776
rect 5675 16745 5687 16748
rect 5629 16739 5687 16745
rect 6086 16736 6092 16748
rect 6144 16736 6150 16788
rect 7653 16779 7711 16785
rect 7653 16745 7665 16779
rect 7699 16776 7711 16779
rect 8018 16776 8024 16788
rect 7699 16748 8024 16776
rect 7699 16745 7711 16748
rect 7653 16739 7711 16745
rect 8018 16736 8024 16748
rect 8076 16776 8082 16788
rect 9677 16779 9735 16785
rect 9677 16776 9689 16779
rect 8076 16748 9689 16776
rect 8076 16736 8082 16748
rect 9677 16745 9689 16748
rect 9723 16745 9735 16779
rect 9677 16739 9735 16745
rect 9858 16736 9864 16788
rect 9916 16776 9922 16788
rect 10045 16779 10103 16785
rect 10045 16776 10057 16779
rect 9916 16748 10057 16776
rect 9916 16736 9922 16748
rect 10045 16745 10057 16748
rect 10091 16776 10103 16779
rect 10686 16776 10692 16788
rect 10091 16748 10692 16776
rect 10091 16745 10103 16748
rect 10045 16739 10103 16745
rect 10686 16736 10692 16748
rect 10744 16736 10750 16788
rect 11517 16779 11575 16785
rect 11517 16745 11529 16779
rect 11563 16776 11575 16779
rect 11698 16776 11704 16788
rect 11563 16748 11704 16776
rect 11563 16745 11575 16748
rect 11517 16739 11575 16745
rect 11698 16736 11704 16748
rect 11756 16736 11762 16788
rect 12894 16736 12900 16788
rect 12952 16776 12958 16788
rect 13081 16779 13139 16785
rect 13081 16776 13093 16779
rect 12952 16748 13093 16776
rect 12952 16736 12958 16748
rect 13081 16745 13093 16748
rect 13127 16745 13139 16779
rect 13081 16739 13139 16745
rect 13538 16736 13544 16788
rect 13596 16776 13602 16788
rect 13633 16779 13691 16785
rect 13633 16776 13645 16779
rect 13596 16748 13645 16776
rect 13596 16736 13602 16748
rect 13633 16745 13645 16748
rect 13679 16745 13691 16779
rect 13998 16776 14004 16788
rect 13959 16748 14004 16776
rect 13633 16739 13691 16745
rect 13998 16736 14004 16748
rect 14056 16736 14062 16788
rect 14182 16776 14188 16788
rect 14143 16748 14188 16776
rect 14182 16736 14188 16748
rect 14240 16736 14246 16788
rect 14737 16779 14795 16785
rect 14737 16745 14749 16779
rect 14783 16776 14795 16779
rect 15473 16779 15531 16785
rect 15473 16776 15485 16779
rect 14783 16748 15485 16776
rect 14783 16745 14795 16748
rect 14737 16739 14795 16745
rect 15473 16745 15485 16748
rect 15519 16776 15531 16779
rect 15746 16776 15752 16788
rect 15519 16748 15752 16776
rect 15519 16745 15531 16748
rect 15473 16739 15531 16745
rect 15746 16736 15752 16748
rect 15804 16736 15810 16788
rect 16577 16779 16635 16785
rect 16577 16745 16589 16779
rect 16623 16776 16635 16779
rect 16666 16776 16672 16788
rect 16623 16748 16672 16776
rect 16623 16745 16635 16748
rect 16577 16739 16635 16745
rect 16666 16736 16672 16748
rect 16724 16736 16730 16788
rect 17218 16776 17224 16788
rect 17179 16748 17224 16776
rect 17218 16736 17224 16748
rect 17276 16736 17282 16788
rect 18046 16776 18052 16788
rect 18007 16748 18052 16776
rect 18046 16736 18052 16748
rect 18104 16736 18110 16788
rect 19518 16736 19524 16788
rect 19576 16776 19582 16788
rect 20073 16779 20131 16785
rect 20073 16776 20085 16779
rect 19576 16748 20085 16776
rect 19576 16736 19582 16748
rect 20073 16745 20085 16748
rect 20119 16776 20131 16779
rect 20714 16776 20720 16788
rect 20119 16748 20720 16776
rect 20119 16745 20131 16748
rect 20073 16739 20131 16745
rect 20714 16736 20720 16748
rect 20772 16736 20778 16788
rect 21910 16736 21916 16788
rect 21968 16776 21974 16788
rect 22281 16779 22339 16785
rect 22281 16776 22293 16779
rect 21968 16748 22293 16776
rect 21968 16736 21974 16748
rect 22281 16745 22293 16748
rect 22327 16745 22339 16779
rect 22281 16739 22339 16745
rect 22925 16779 22983 16785
rect 22925 16745 22937 16779
rect 22971 16776 22983 16779
rect 23014 16776 23020 16788
rect 22971 16748 23020 16776
rect 22971 16745 22983 16748
rect 22925 16739 22983 16745
rect 23014 16736 23020 16748
rect 23072 16736 23078 16788
rect 23106 16736 23112 16788
rect 23164 16776 23170 16788
rect 23201 16779 23259 16785
rect 23201 16776 23213 16779
rect 23164 16748 23213 16776
rect 23164 16736 23170 16748
rect 23201 16745 23213 16748
rect 23247 16745 23259 16779
rect 23201 16739 23259 16745
rect 23385 16779 23443 16785
rect 23385 16745 23397 16779
rect 23431 16745 23443 16779
rect 23750 16776 23756 16788
rect 23385 16739 23443 16745
rect 23492 16748 23756 16776
rect 1762 16708 1768 16720
rect 1723 16680 1768 16708
rect 1762 16668 1768 16680
rect 1820 16668 1826 16720
rect 5442 16668 5448 16720
rect 5500 16708 5506 16720
rect 5537 16711 5595 16717
rect 5537 16708 5549 16711
rect 5500 16680 5549 16708
rect 5500 16668 5506 16680
rect 5537 16677 5549 16680
rect 5583 16708 5595 16711
rect 6638 16708 6644 16720
rect 5583 16680 6644 16708
rect 5583 16677 5595 16680
rect 5537 16671 5595 16677
rect 6638 16668 6644 16680
rect 6696 16668 6702 16720
rect 9306 16708 9312 16720
rect 9267 16680 9312 16708
rect 9306 16668 9312 16680
rect 9364 16668 9370 16720
rect 11606 16668 11612 16720
rect 11664 16708 11670 16720
rect 15102 16708 15108 16720
rect 11664 16680 14504 16708
rect 15015 16680 15108 16708
rect 11664 16668 11670 16680
rect 1857 16643 1915 16649
rect 1857 16609 1869 16643
rect 1903 16640 1915 16643
rect 2130 16640 2136 16652
rect 1903 16612 2136 16640
rect 1903 16609 1915 16612
rect 1857 16603 1915 16609
rect 2130 16600 2136 16612
rect 2188 16600 2194 16652
rect 2406 16600 2412 16652
rect 2464 16640 2470 16652
rect 2777 16643 2835 16649
rect 2777 16640 2789 16643
rect 2464 16612 2789 16640
rect 2464 16600 2470 16612
rect 2777 16609 2789 16612
rect 2823 16609 2835 16643
rect 2777 16603 2835 16609
rect 3234 16600 3240 16652
rect 3292 16640 3298 16652
rect 3789 16643 3847 16649
rect 3789 16640 3801 16643
rect 3292 16612 3801 16640
rect 3292 16600 3298 16612
rect 3789 16609 3801 16612
rect 3835 16609 3847 16643
rect 3789 16603 3847 16609
rect 4433 16643 4491 16649
rect 4433 16609 4445 16643
rect 4479 16640 4491 16643
rect 4706 16640 4712 16652
rect 4479 16612 4712 16640
rect 4479 16609 4491 16612
rect 4433 16603 4491 16609
rect 4706 16600 4712 16612
rect 4764 16640 4770 16652
rect 5350 16640 5356 16652
rect 4764 16612 5356 16640
rect 4764 16600 4770 16612
rect 5350 16600 5356 16612
rect 5408 16600 5414 16652
rect 5997 16643 6055 16649
rect 5997 16609 6009 16643
rect 6043 16609 6055 16643
rect 5997 16603 6055 16609
rect 6089 16643 6147 16649
rect 6089 16609 6101 16643
rect 6135 16640 6147 16643
rect 7098 16640 7104 16652
rect 6135 16612 7104 16640
rect 6135 16609 6147 16612
rect 6089 16603 6147 16609
rect 2038 16572 2044 16584
rect 1999 16544 2044 16572
rect 2038 16532 2044 16544
rect 2096 16532 2102 16584
rect 4614 16572 4620 16584
rect 4575 16544 4620 16572
rect 4614 16532 4620 16544
rect 4672 16532 4678 16584
rect 3418 16464 3424 16516
rect 3476 16504 3482 16516
rect 5077 16507 5135 16513
rect 5077 16504 5089 16507
rect 3476 16476 5089 16504
rect 3476 16464 3482 16476
rect 5077 16473 5089 16476
rect 5123 16504 5135 16507
rect 5258 16504 5264 16516
rect 5123 16476 5264 16504
rect 5123 16473 5135 16476
rect 5077 16467 5135 16473
rect 5258 16464 5264 16476
rect 5316 16464 5322 16516
rect 1397 16439 1455 16445
rect 1397 16405 1409 16439
rect 1443 16436 1455 16439
rect 2498 16436 2504 16448
rect 1443 16408 2504 16436
rect 1443 16405 1455 16408
rect 1397 16399 1455 16405
rect 2498 16396 2504 16408
rect 2556 16396 2562 16448
rect 4062 16436 4068 16448
rect 4023 16408 4068 16436
rect 4062 16396 4068 16408
rect 4120 16396 4126 16448
rect 6012 16436 6040 16603
rect 7098 16600 7104 16612
rect 7156 16600 7162 16652
rect 7561 16643 7619 16649
rect 7561 16609 7573 16643
rect 7607 16640 7619 16643
rect 8202 16640 8208 16652
rect 7607 16612 8208 16640
rect 7607 16609 7619 16612
rect 7561 16603 7619 16609
rect 8202 16600 8208 16612
rect 8260 16600 8266 16652
rect 8294 16600 8300 16652
rect 8352 16640 8358 16652
rect 10137 16643 10195 16649
rect 8352 16612 8397 16640
rect 8352 16600 8358 16612
rect 10137 16609 10149 16643
rect 10183 16640 10195 16643
rect 10226 16640 10232 16652
rect 10183 16612 10232 16640
rect 10183 16609 10195 16612
rect 10137 16603 10195 16609
rect 10226 16600 10232 16612
rect 10284 16640 10290 16652
rect 11422 16640 11428 16652
rect 10284 16612 11428 16640
rect 10284 16600 10290 16612
rect 11422 16600 11428 16612
rect 11480 16600 11486 16652
rect 11790 16640 11796 16652
rect 11716 16612 11796 16640
rect 6270 16572 6276 16584
rect 6231 16544 6276 16572
rect 6270 16532 6276 16544
rect 6328 16532 6334 16584
rect 6638 16532 6644 16584
rect 6696 16572 6702 16584
rect 6914 16572 6920 16584
rect 6696 16544 6920 16572
rect 6696 16532 6702 16544
rect 6914 16532 6920 16544
rect 6972 16532 6978 16584
rect 7745 16575 7803 16581
rect 7745 16572 7757 16575
rect 7024 16544 7757 16572
rect 6270 16436 6276 16448
rect 6012 16408 6276 16436
rect 6270 16396 6276 16408
rect 6328 16396 6334 16448
rect 6733 16439 6791 16445
rect 6733 16405 6745 16439
rect 6779 16436 6791 16439
rect 6914 16436 6920 16448
rect 6779 16408 6920 16436
rect 6779 16405 6791 16408
rect 6733 16399 6791 16405
rect 6914 16396 6920 16408
rect 6972 16436 6978 16448
rect 7024 16445 7052 16544
rect 7745 16541 7757 16544
rect 7791 16541 7803 16575
rect 10318 16572 10324 16584
rect 10279 16544 10324 16572
rect 7745 16535 7803 16541
rect 10318 16532 10324 16544
rect 10376 16532 10382 16584
rect 11716 16581 11744 16612
rect 11790 16600 11796 16612
rect 11848 16600 11854 16652
rect 11974 16649 11980 16652
rect 11968 16640 11980 16649
rect 11935 16612 11980 16640
rect 11968 16603 11980 16612
rect 12032 16640 12038 16652
rect 14476 16640 14504 16680
rect 15102 16668 15108 16680
rect 15160 16708 15166 16720
rect 16022 16708 16028 16720
rect 15160 16680 16028 16708
rect 15160 16668 15166 16680
rect 16022 16668 16028 16680
rect 16080 16668 16086 16720
rect 18138 16668 18144 16720
rect 18196 16708 18202 16720
rect 18598 16708 18604 16720
rect 18196 16680 18604 16708
rect 18196 16668 18202 16680
rect 18598 16668 18604 16680
rect 18656 16668 18662 16720
rect 20438 16668 20444 16720
rect 20496 16708 20502 16720
rect 21168 16711 21226 16717
rect 21168 16708 21180 16711
rect 20496 16680 21180 16708
rect 20496 16668 20502 16680
rect 21168 16677 21180 16680
rect 21214 16708 21226 16711
rect 22002 16708 22008 16720
rect 21214 16680 22008 16708
rect 21214 16677 21226 16680
rect 21168 16671 21226 16677
rect 22002 16668 22008 16680
rect 22060 16668 22066 16720
rect 15838 16640 15844 16652
rect 12032 16612 12756 16640
rect 14476 16612 15844 16640
rect 11974 16600 11980 16603
rect 12032 16600 12038 16612
rect 11701 16575 11759 16581
rect 11701 16541 11713 16575
rect 11747 16541 11759 16575
rect 12728 16572 12756 16612
rect 15838 16600 15844 16612
rect 15896 16600 15902 16652
rect 17034 16640 17040 16652
rect 16995 16612 17040 16640
rect 17034 16600 17040 16612
rect 17092 16600 17098 16652
rect 18408 16643 18466 16649
rect 18408 16640 18420 16643
rect 17880 16612 18420 16640
rect 13722 16572 13728 16584
rect 12728 16544 13728 16572
rect 11701 16535 11759 16541
rect 10594 16464 10600 16516
rect 10652 16504 10658 16516
rect 11057 16507 11115 16513
rect 11057 16504 11069 16507
rect 10652 16476 11069 16504
rect 10652 16464 10658 16476
rect 11057 16473 11069 16476
rect 11103 16473 11115 16507
rect 11057 16467 11115 16473
rect 7009 16439 7067 16445
rect 7009 16436 7021 16439
rect 6972 16408 7021 16436
rect 6972 16396 6978 16408
rect 7009 16405 7021 16408
rect 7055 16405 7067 16439
rect 7190 16436 7196 16448
rect 7151 16408 7196 16436
rect 7009 16399 7067 16405
rect 7190 16396 7196 16408
rect 7248 16396 7254 16448
rect 8757 16439 8815 16445
rect 8757 16405 8769 16439
rect 8803 16436 8815 16439
rect 9122 16436 9128 16448
rect 8803 16408 9128 16436
rect 8803 16405 8815 16408
rect 8757 16399 8815 16405
rect 9122 16396 9128 16408
rect 9180 16396 9186 16448
rect 10686 16436 10692 16448
rect 10647 16408 10692 16436
rect 10686 16396 10692 16408
rect 10744 16396 10750 16448
rect 11716 16436 11744 16535
rect 13722 16532 13728 16544
rect 13780 16532 13786 16584
rect 15930 16572 15936 16584
rect 15891 16544 15936 16572
rect 15930 16532 15936 16544
rect 15988 16532 15994 16584
rect 16025 16575 16083 16581
rect 16025 16541 16037 16575
rect 16071 16541 16083 16575
rect 16025 16535 16083 16541
rect 14734 16464 14740 16516
rect 14792 16504 14798 16516
rect 16040 16504 16068 16535
rect 17494 16532 17500 16584
rect 17552 16572 17558 16584
rect 17880 16572 17908 16612
rect 18408 16609 18420 16612
rect 18454 16640 18466 16643
rect 19242 16640 19248 16652
rect 18454 16612 19248 16640
rect 18454 16609 18466 16612
rect 18408 16603 18466 16609
rect 19242 16600 19248 16612
rect 19300 16600 19306 16652
rect 20717 16643 20775 16649
rect 20717 16609 20729 16643
rect 20763 16640 20775 16643
rect 21450 16640 21456 16652
rect 20763 16612 21456 16640
rect 20763 16609 20775 16612
rect 20717 16603 20775 16609
rect 21450 16600 21456 16612
rect 21508 16600 21514 16652
rect 21542 16600 21548 16652
rect 21600 16640 21606 16652
rect 23400 16640 23428 16739
rect 21600 16612 22968 16640
rect 21600 16600 21606 16612
rect 18138 16572 18144 16584
rect 17552 16544 17908 16572
rect 18099 16544 18144 16572
rect 17552 16532 17558 16544
rect 18138 16532 18144 16544
rect 18196 16532 18202 16584
rect 20898 16572 20904 16584
rect 20859 16544 20904 16572
rect 20898 16532 20904 16544
rect 20956 16532 20962 16584
rect 22940 16572 22968 16612
rect 23124 16612 23428 16640
rect 23124 16572 23152 16612
rect 22940 16544 23152 16572
rect 16390 16504 16396 16516
rect 14792 16476 16396 16504
rect 14792 16464 14798 16476
rect 16390 16464 16396 16476
rect 16448 16464 16454 16516
rect 16945 16507 17003 16513
rect 16945 16473 16957 16507
rect 16991 16504 17003 16507
rect 17402 16504 17408 16516
rect 16991 16476 17408 16504
rect 16991 16473 17003 16476
rect 16945 16467 17003 16473
rect 17402 16464 17408 16476
rect 17460 16464 17466 16516
rect 23106 16464 23112 16516
rect 23164 16504 23170 16516
rect 23492 16504 23520 16748
rect 23750 16736 23756 16748
rect 23808 16776 23814 16788
rect 23845 16779 23903 16785
rect 23845 16776 23857 16779
rect 23808 16748 23857 16776
rect 23808 16736 23814 16748
rect 23845 16745 23857 16748
rect 23891 16745 23903 16779
rect 24394 16776 24400 16788
rect 24355 16748 24400 16776
rect 23845 16739 23903 16745
rect 24394 16736 24400 16748
rect 24452 16736 24458 16788
rect 25222 16708 25228 16720
rect 25183 16680 25228 16708
rect 25222 16668 25228 16680
rect 25280 16668 25286 16720
rect 23750 16640 23756 16652
rect 23711 16612 23756 16640
rect 23750 16600 23756 16612
rect 23808 16600 23814 16652
rect 24949 16643 25007 16649
rect 24949 16609 24961 16643
rect 24995 16640 25007 16643
rect 25682 16640 25688 16652
rect 24995 16612 25688 16640
rect 24995 16609 25007 16612
rect 24949 16603 25007 16609
rect 25682 16600 25688 16612
rect 25740 16600 25746 16652
rect 24026 16572 24032 16584
rect 23987 16544 24032 16572
rect 24026 16532 24032 16544
rect 24084 16572 24090 16584
rect 24854 16572 24860 16584
rect 24084 16544 24860 16572
rect 24084 16532 24090 16544
rect 24854 16532 24860 16544
rect 24912 16532 24918 16584
rect 23164 16476 23520 16504
rect 23164 16464 23170 16476
rect 24118 16464 24124 16516
rect 24176 16504 24182 16516
rect 24302 16504 24308 16516
rect 24176 16476 24308 16504
rect 24176 16464 24182 16476
rect 24302 16464 24308 16476
rect 24360 16464 24366 16516
rect 16666 16436 16672 16448
rect 11716 16408 16672 16436
rect 16666 16396 16672 16408
rect 16724 16396 16730 16448
rect 17678 16436 17684 16448
rect 17639 16408 17684 16436
rect 17678 16396 17684 16408
rect 17736 16396 17742 16448
rect 19518 16436 19524 16448
rect 19479 16408 19524 16436
rect 19518 16396 19524 16408
rect 19576 16396 19582 16448
rect 23290 16396 23296 16448
rect 23348 16436 23354 16448
rect 23750 16436 23756 16448
rect 23348 16408 23756 16436
rect 23348 16396 23354 16408
rect 23750 16396 23756 16408
rect 23808 16396 23814 16448
rect 24670 16396 24676 16448
rect 24728 16436 24734 16448
rect 24765 16439 24823 16445
rect 24765 16436 24777 16439
rect 24728 16408 24777 16436
rect 24728 16396 24734 16408
rect 24765 16405 24777 16408
rect 24811 16405 24823 16439
rect 24765 16399 24823 16405
rect 25682 16396 25688 16448
rect 25740 16436 25746 16448
rect 26053 16439 26111 16445
rect 26053 16436 26065 16439
rect 25740 16408 26065 16436
rect 25740 16396 25746 16408
rect 26053 16405 26065 16408
rect 26099 16436 26111 16439
rect 26142 16436 26148 16448
rect 26099 16408 26148 16436
rect 26099 16405 26111 16408
rect 26053 16399 26111 16405
rect 26142 16396 26148 16408
rect 26200 16396 26206 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 5258 16192 5264 16244
rect 5316 16192 5322 16244
rect 8202 16192 8208 16244
rect 8260 16232 8266 16244
rect 8665 16235 8723 16241
rect 8665 16232 8677 16235
rect 8260 16204 8677 16232
rect 8260 16192 8266 16204
rect 8665 16201 8677 16204
rect 8711 16201 8723 16235
rect 8665 16195 8723 16201
rect 8846 16192 8852 16244
rect 8904 16192 8910 16244
rect 9769 16235 9827 16241
rect 9769 16201 9781 16235
rect 9815 16232 9827 16235
rect 9858 16232 9864 16244
rect 9815 16204 9864 16232
rect 9815 16201 9827 16204
rect 9769 16195 9827 16201
rect 9858 16192 9864 16204
rect 9916 16192 9922 16244
rect 9950 16192 9956 16244
rect 10008 16232 10014 16244
rect 10229 16235 10287 16241
rect 10229 16232 10241 16235
rect 10008 16204 10241 16232
rect 10008 16192 10014 16204
rect 10229 16201 10241 16204
rect 10275 16201 10287 16235
rect 10229 16195 10287 16201
rect 10318 16192 10324 16244
rect 10376 16232 10382 16244
rect 11241 16235 11299 16241
rect 11241 16232 11253 16235
rect 10376 16204 11253 16232
rect 10376 16192 10382 16204
rect 11241 16201 11253 16204
rect 11287 16201 11299 16235
rect 11241 16195 11299 16201
rect 12342 16192 12348 16244
rect 12400 16232 12406 16244
rect 12437 16235 12495 16241
rect 12437 16232 12449 16235
rect 12400 16204 12449 16232
rect 12400 16192 12406 16204
rect 12437 16201 12449 16204
rect 12483 16201 12495 16235
rect 12437 16195 12495 16201
rect 13541 16235 13599 16241
rect 13541 16201 13553 16235
rect 13587 16232 13599 16235
rect 13722 16232 13728 16244
rect 13587 16204 13728 16232
rect 13587 16201 13599 16204
rect 13541 16195 13599 16201
rect 13722 16192 13728 16204
rect 13780 16192 13786 16244
rect 14461 16235 14519 16241
rect 14461 16201 14473 16235
rect 14507 16232 14519 16235
rect 14734 16232 14740 16244
rect 14507 16204 14740 16232
rect 14507 16201 14519 16204
rect 14461 16195 14519 16201
rect 14734 16192 14740 16204
rect 14792 16192 14798 16244
rect 15933 16235 15991 16241
rect 15933 16201 15945 16235
rect 15979 16232 15991 16235
rect 16022 16232 16028 16244
rect 15979 16204 16028 16232
rect 15979 16201 15991 16204
rect 15933 16195 15991 16201
rect 16022 16192 16028 16204
rect 16080 16192 16086 16244
rect 16390 16192 16396 16244
rect 16448 16232 16454 16244
rect 16485 16235 16543 16241
rect 16485 16232 16497 16235
rect 16448 16204 16497 16232
rect 16448 16192 16454 16204
rect 16485 16201 16497 16204
rect 16531 16201 16543 16235
rect 17034 16232 17040 16244
rect 16995 16204 17040 16232
rect 16485 16195 16543 16201
rect 17034 16192 17040 16204
rect 17092 16192 17098 16244
rect 17494 16232 17500 16244
rect 17455 16204 17500 16232
rect 17494 16192 17500 16204
rect 17552 16192 17558 16244
rect 20714 16232 20720 16244
rect 20675 16204 20720 16232
rect 20714 16192 20720 16204
rect 20772 16192 20778 16244
rect 23106 16232 23112 16244
rect 23067 16204 23112 16232
rect 23106 16192 23112 16204
rect 23164 16192 23170 16244
rect 23750 16192 23756 16244
rect 23808 16232 23814 16244
rect 24673 16235 24731 16241
rect 24673 16232 24685 16235
rect 23808 16204 24685 16232
rect 23808 16192 23814 16204
rect 24673 16201 24685 16204
rect 24719 16201 24731 16235
rect 24673 16195 24731 16201
rect 24854 16192 24860 16244
rect 24912 16232 24918 16244
rect 25041 16235 25099 16241
rect 25041 16232 25053 16235
rect 24912 16204 25053 16232
rect 24912 16192 24918 16204
rect 25041 16201 25053 16204
rect 25087 16232 25099 16235
rect 25222 16232 25228 16244
rect 25087 16204 25228 16232
rect 25087 16201 25099 16204
rect 25041 16195 25099 16201
rect 25222 16192 25228 16204
rect 25280 16192 25286 16244
rect 2685 16167 2743 16173
rect 2685 16133 2697 16167
rect 2731 16164 2743 16167
rect 2866 16164 2872 16176
rect 2731 16136 2872 16164
rect 2731 16133 2743 16136
rect 2685 16127 2743 16133
rect 2866 16124 2872 16136
rect 2924 16164 2930 16176
rect 3878 16164 3884 16176
rect 2924 16136 3884 16164
rect 2924 16124 2930 16136
rect 3878 16124 3884 16136
rect 3936 16124 3942 16176
rect 4706 16164 4712 16176
rect 4667 16136 4712 16164
rect 4706 16124 4712 16136
rect 4764 16124 4770 16176
rect 5276 16164 5304 16192
rect 5718 16164 5724 16176
rect 5276 16136 5724 16164
rect 5718 16124 5724 16136
rect 5776 16124 5782 16176
rect 6181 16167 6239 16173
rect 6181 16133 6193 16167
rect 6227 16164 6239 16167
rect 6270 16164 6276 16176
rect 6227 16136 6276 16164
rect 6227 16133 6239 16136
rect 6181 16127 6239 16133
rect 6270 16124 6276 16136
rect 6328 16164 6334 16176
rect 8386 16164 8392 16176
rect 6328 16136 8392 16164
rect 6328 16124 6334 16136
rect 8386 16124 8392 16136
rect 8444 16164 8450 16176
rect 8754 16164 8760 16176
rect 8444 16136 8760 16164
rect 8444 16124 8450 16136
rect 8754 16124 8760 16136
rect 8812 16124 8818 16176
rect 2038 16096 2044 16108
rect 1999 16068 2044 16096
rect 2038 16056 2044 16068
rect 2096 16096 2102 16108
rect 2096 16068 3004 16096
rect 2096 16056 2102 16068
rect 2976 16028 3004 16068
rect 3418 16056 3424 16108
rect 3476 16096 3482 16108
rect 3697 16099 3755 16105
rect 3697 16096 3709 16099
rect 3476 16068 3709 16096
rect 3476 16056 3482 16068
rect 3697 16065 3709 16068
rect 3743 16065 3755 16099
rect 5261 16099 5319 16105
rect 5261 16096 5273 16099
rect 3697 16059 3755 16065
rect 4632 16068 5273 16096
rect 4632 16040 4660 16068
rect 5261 16065 5273 16068
rect 5307 16065 5319 16099
rect 5261 16059 5319 16065
rect 6914 16056 6920 16108
rect 6972 16096 6978 16108
rect 7653 16099 7711 16105
rect 7653 16096 7665 16099
rect 6972 16068 7665 16096
rect 6972 16056 6978 16068
rect 7653 16065 7665 16068
rect 7699 16065 7711 16099
rect 7653 16059 7711 16065
rect 4157 16031 4215 16037
rect 4157 16028 4169 16031
rect 2976 16000 4169 16028
rect 4157 15997 4169 16000
rect 4203 16028 4215 16031
rect 4525 16031 4583 16037
rect 4525 16028 4537 16031
rect 4203 16000 4537 16028
rect 4203 15997 4215 16000
rect 4157 15991 4215 15997
rect 4525 15997 4537 16000
rect 4571 16028 4583 16031
rect 4614 16028 4620 16040
rect 4571 16000 4620 16028
rect 4571 15997 4583 16000
rect 4525 15991 4583 15997
rect 4614 15988 4620 16000
rect 4672 15988 4678 16040
rect 5074 15988 5080 16040
rect 5132 15988 5138 16040
rect 5169 16031 5227 16037
rect 5169 15997 5181 16031
rect 5215 16028 5227 16031
rect 5442 16028 5448 16040
rect 5215 16000 5448 16028
rect 5215 15997 5227 16000
rect 5169 15991 5227 15997
rect 5442 15988 5448 16000
rect 5500 15988 5506 16040
rect 6457 16031 6515 16037
rect 6457 15997 6469 16031
rect 6503 16028 6515 16031
rect 6822 16028 6828 16040
rect 6503 16000 6828 16028
rect 6503 15997 6515 16000
rect 6457 15991 6515 15997
rect 6822 15988 6828 16000
rect 6880 15988 6886 16040
rect 7098 15988 7104 16040
rect 7156 15988 7162 16040
rect 8754 15988 8760 16040
rect 8812 16028 8818 16040
rect 8864 16028 8892 16192
rect 9122 16096 9128 16108
rect 9083 16068 9128 16096
rect 9122 16056 9128 16068
rect 9180 16056 9186 16108
rect 9214 16056 9220 16108
rect 9272 16096 9278 16108
rect 9309 16099 9367 16105
rect 9309 16096 9321 16099
rect 9272 16068 9321 16096
rect 9272 16056 9278 16068
rect 9309 16065 9321 16068
rect 9355 16096 9367 16099
rect 10336 16096 10364 16192
rect 11054 16124 11060 16176
rect 11112 16164 11118 16176
rect 11793 16167 11851 16173
rect 11793 16164 11805 16167
rect 11112 16136 11805 16164
rect 11112 16124 11118 16136
rect 11793 16133 11805 16136
rect 11839 16133 11851 16167
rect 11793 16127 11851 16133
rect 10778 16096 10784 16108
rect 9355 16068 10364 16096
rect 10739 16068 10784 16096
rect 9355 16065 9367 16068
rect 9309 16059 9367 16065
rect 10778 16056 10784 16068
rect 10836 16056 10842 16108
rect 8812 16000 8892 16028
rect 8812 15988 8818 16000
rect 9030 15988 9036 16040
rect 9088 15988 9094 16040
rect 10594 16028 10600 16040
rect 10428 16000 10600 16028
rect 1302 15920 1308 15972
rect 1360 15960 1366 15972
rect 1360 15932 1624 15960
rect 1360 15920 1366 15932
rect 1026 15852 1032 15904
rect 1084 15892 1090 15904
rect 1397 15895 1455 15901
rect 1397 15892 1409 15895
rect 1084 15864 1409 15892
rect 1084 15852 1090 15864
rect 1397 15861 1409 15864
rect 1443 15861 1455 15895
rect 1596 15892 1624 15932
rect 1670 15920 1676 15972
rect 1728 15960 1734 15972
rect 1765 15963 1823 15969
rect 1765 15960 1777 15963
rect 1728 15932 1777 15960
rect 1728 15920 1734 15932
rect 1765 15929 1777 15932
rect 1811 15960 1823 15963
rect 2314 15960 2320 15972
rect 1811 15932 2320 15960
rect 1811 15929 1823 15932
rect 1765 15923 1823 15929
rect 2314 15920 2320 15932
rect 2372 15920 2378 15972
rect 3053 15963 3111 15969
rect 3053 15929 3065 15963
rect 3099 15960 3111 15963
rect 5092 15960 5120 15988
rect 5813 15963 5871 15969
rect 3099 15932 3556 15960
rect 5092 15932 5212 15960
rect 3099 15929 3111 15932
rect 3053 15923 3111 15929
rect 3528 15904 3556 15932
rect 1857 15895 1915 15901
rect 1857 15892 1869 15895
rect 1596 15864 1869 15892
rect 1397 15855 1455 15861
rect 1857 15861 1869 15864
rect 1903 15892 1915 15895
rect 2590 15892 2596 15904
rect 1903 15864 2596 15892
rect 1903 15861 1915 15864
rect 1857 15855 1915 15861
rect 2590 15852 2596 15864
rect 2648 15852 2654 15904
rect 3142 15892 3148 15904
rect 3103 15864 3148 15892
rect 3142 15852 3148 15864
rect 3200 15852 3206 15904
rect 3510 15892 3516 15904
rect 3471 15864 3516 15892
rect 3510 15852 3516 15864
rect 3568 15852 3574 15904
rect 3605 15895 3663 15901
rect 3605 15861 3617 15895
rect 3651 15892 3663 15895
rect 3878 15892 3884 15904
rect 3651 15864 3884 15892
rect 3651 15861 3663 15864
rect 3605 15855 3663 15861
rect 3878 15852 3884 15864
rect 3936 15852 3942 15904
rect 5074 15892 5080 15904
rect 5035 15864 5080 15892
rect 5074 15852 5080 15864
rect 5132 15852 5138 15904
rect 5184 15892 5212 15932
rect 5813 15929 5825 15963
rect 5859 15960 5871 15963
rect 7116 15960 7144 15988
rect 5859 15932 7144 15960
rect 7469 15963 7527 15969
rect 5859 15929 5871 15932
rect 5813 15923 5871 15929
rect 6840 15904 6868 15932
rect 7469 15929 7481 15963
rect 7515 15960 7527 15963
rect 8205 15963 8263 15969
rect 8205 15960 8217 15963
rect 7515 15932 8217 15960
rect 7515 15929 7527 15932
rect 7469 15923 7527 15929
rect 8205 15929 8217 15932
rect 8251 15960 8263 15963
rect 8846 15960 8852 15972
rect 8251 15932 8852 15960
rect 8251 15929 8263 15932
rect 8205 15923 8263 15929
rect 8846 15920 8852 15932
rect 8904 15960 8910 15972
rect 9048 15960 9076 15988
rect 10042 15960 10048 15972
rect 8904 15932 9076 15960
rect 10003 15932 10048 15960
rect 8904 15920 8910 15932
rect 10042 15920 10048 15932
rect 10100 15960 10106 15972
rect 10226 15960 10232 15972
rect 10100 15932 10232 15960
rect 10100 15920 10106 15932
rect 10226 15920 10232 15932
rect 10284 15920 10290 15972
rect 5258 15892 5264 15904
rect 5171 15864 5264 15892
rect 5258 15852 5264 15864
rect 5316 15892 5322 15904
rect 6273 15895 6331 15901
rect 6273 15892 6285 15895
rect 5316 15864 6285 15892
rect 5316 15852 5322 15864
rect 6273 15861 6285 15864
rect 6319 15861 6331 15895
rect 6273 15855 6331 15861
rect 6822 15852 6828 15904
rect 6880 15852 6886 15904
rect 7098 15892 7104 15904
rect 7059 15864 7104 15892
rect 7098 15852 7104 15864
rect 7156 15852 7162 15904
rect 7558 15852 7564 15904
rect 7616 15892 7622 15904
rect 7616 15864 7661 15892
rect 7616 15852 7622 15864
rect 8478 15852 8484 15904
rect 8536 15892 8542 15904
rect 8573 15895 8631 15901
rect 8573 15892 8585 15895
rect 8536 15864 8585 15892
rect 8536 15852 8542 15864
rect 8573 15861 8585 15864
rect 8619 15892 8631 15895
rect 9030 15892 9036 15904
rect 8619 15864 9036 15892
rect 8619 15861 8631 15864
rect 8573 15855 8631 15861
rect 9030 15852 9036 15864
rect 9088 15852 9094 15904
rect 9490 15852 9496 15904
rect 9548 15892 9554 15904
rect 10428 15892 10456 16000
rect 10594 15988 10600 16000
rect 10652 15988 10658 16040
rect 11808 15960 11836 16127
rect 13814 16124 13820 16176
rect 13872 16164 13878 16176
rect 14090 16164 14096 16176
rect 13872 16136 14096 16164
rect 13872 16124 13878 16136
rect 14090 16124 14096 16136
rect 14148 16164 14154 16176
rect 23661 16167 23719 16173
rect 14148 16136 14596 16164
rect 14148 16124 14154 16136
rect 11977 16099 12035 16105
rect 11977 16065 11989 16099
rect 12023 16096 12035 16099
rect 12253 16099 12311 16105
rect 12253 16096 12265 16099
rect 12023 16068 12265 16096
rect 12023 16065 12035 16068
rect 11977 16059 12035 16065
rect 12253 16065 12265 16068
rect 12299 16096 12311 16099
rect 12299 16068 12848 16096
rect 12299 16065 12311 16068
rect 12253 16059 12311 16065
rect 12820 16028 12848 16068
rect 12894 16056 12900 16108
rect 12952 16096 12958 16108
rect 14568 16105 14596 16136
rect 23661 16133 23673 16167
rect 23707 16164 23719 16167
rect 26234 16164 26240 16176
rect 23707 16136 26240 16164
rect 23707 16133 23719 16136
rect 23661 16127 23719 16133
rect 26234 16124 26240 16136
rect 26292 16124 26298 16176
rect 12989 16099 13047 16105
rect 12989 16096 13001 16099
rect 12952 16068 13001 16096
rect 12952 16056 12958 16068
rect 12989 16065 13001 16068
rect 13035 16065 13047 16099
rect 12989 16059 13047 16065
rect 14553 16099 14611 16105
rect 14553 16065 14565 16099
rect 14599 16065 14611 16099
rect 14553 16059 14611 16065
rect 19242 16056 19248 16108
rect 19300 16096 19306 16108
rect 20625 16099 20683 16105
rect 20625 16096 20637 16099
rect 19300 16068 20637 16096
rect 19300 16056 19306 16068
rect 20625 16065 20637 16068
rect 20671 16096 20683 16099
rect 21361 16099 21419 16105
rect 21361 16096 21373 16099
rect 20671 16068 21373 16096
rect 20671 16065 20683 16068
rect 20625 16059 20683 16065
rect 21361 16065 21373 16068
rect 21407 16096 21419 16099
rect 21910 16096 21916 16108
rect 21407 16068 21916 16096
rect 21407 16065 21419 16068
rect 21361 16059 21419 16065
rect 21910 16056 21916 16068
rect 21968 16056 21974 16108
rect 22186 16056 22192 16108
rect 22244 16096 22250 16108
rect 22244 16068 23796 16096
rect 22244 16056 22250 16068
rect 13814 16028 13820 16040
rect 12820 16000 13032 16028
rect 13775 16000 13820 16028
rect 11808 15932 12296 15960
rect 9548 15864 10456 15892
rect 9548 15852 9554 15864
rect 10686 15852 10692 15904
rect 10744 15892 10750 15904
rect 10744 15864 10789 15892
rect 10744 15852 10750 15864
rect 11422 15852 11428 15904
rect 11480 15892 11486 15904
rect 11977 15895 12035 15901
rect 11977 15892 11989 15895
rect 11480 15864 11989 15892
rect 11480 15852 11486 15864
rect 11977 15861 11989 15864
rect 12023 15861 12035 15895
rect 12268 15892 12296 15932
rect 12805 15895 12863 15901
rect 12805 15892 12817 15895
rect 12268 15864 12817 15892
rect 11977 15855 12035 15861
rect 12805 15861 12817 15864
rect 12851 15861 12863 15895
rect 12805 15855 12863 15861
rect 12897 15895 12955 15901
rect 12897 15861 12909 15895
rect 12943 15892 12955 15895
rect 13004 15892 13032 16000
rect 13814 15988 13820 16000
rect 13872 15988 13878 16040
rect 16942 15988 16948 16040
rect 17000 16028 17006 16040
rect 17678 16028 17684 16040
rect 17000 16000 17684 16028
rect 17000 15988 17006 16000
rect 17678 15988 17684 16000
rect 17736 16028 17742 16040
rect 17773 16031 17831 16037
rect 17773 16028 17785 16031
rect 17736 16000 17785 16028
rect 17736 15988 17742 16000
rect 17773 15997 17785 16000
rect 17819 15997 17831 16031
rect 17773 15991 17831 15997
rect 18049 16031 18107 16037
rect 18049 15997 18061 16031
rect 18095 16028 18107 16031
rect 18138 16028 18144 16040
rect 18095 16000 18144 16028
rect 18095 15997 18107 16000
rect 18049 15991 18107 15997
rect 18138 15988 18144 16000
rect 18196 15988 18202 16040
rect 20990 15988 20996 16040
rect 21048 16028 21054 16040
rect 21085 16031 21143 16037
rect 21085 16028 21097 16031
rect 21048 16000 21097 16028
rect 21048 15988 21054 16000
rect 21085 15997 21097 16000
rect 21131 15997 21143 16031
rect 21085 15991 21143 15997
rect 21821 16031 21879 16037
rect 21821 15997 21833 16031
rect 21867 16028 21879 16031
rect 22002 16028 22008 16040
rect 21867 16000 22008 16028
rect 21867 15997 21879 16000
rect 21821 15991 21879 15997
rect 22002 15988 22008 16000
rect 22060 15988 22066 16040
rect 22465 16031 22523 16037
rect 22465 15997 22477 16031
rect 22511 16028 22523 16031
rect 22922 16028 22928 16040
rect 22511 16000 22928 16028
rect 22511 15997 22523 16000
rect 22465 15991 22523 15997
rect 14734 15920 14740 15972
rect 14792 15969 14798 15972
rect 14792 15963 14856 15969
rect 14792 15929 14810 15963
rect 14844 15929 14856 15963
rect 14792 15923 14856 15929
rect 18316 15963 18374 15969
rect 18316 15929 18328 15963
rect 18362 15960 18374 15963
rect 18598 15960 18604 15972
rect 18362 15932 18604 15960
rect 18362 15929 18374 15932
rect 18316 15923 18374 15929
rect 14792 15920 14798 15923
rect 18598 15920 18604 15932
rect 18656 15920 18662 15972
rect 20257 15963 20315 15969
rect 20257 15929 20269 15963
rect 20303 15960 20315 15963
rect 21177 15963 21235 15969
rect 21177 15960 21189 15963
rect 20303 15932 21189 15960
rect 20303 15929 20315 15932
rect 20257 15923 20315 15929
rect 21177 15929 21189 15932
rect 21223 15960 21235 15963
rect 22186 15960 22192 15972
rect 21223 15932 22192 15960
rect 21223 15929 21235 15932
rect 21177 15923 21235 15929
rect 22186 15920 22192 15932
rect 22244 15920 22250 15972
rect 17218 15892 17224 15904
rect 12943 15864 17224 15892
rect 12943 15861 12955 15864
rect 12897 15855 12955 15861
rect 17218 15852 17224 15864
rect 17276 15852 17282 15904
rect 17402 15852 17408 15904
rect 17460 15892 17466 15904
rect 17589 15895 17647 15901
rect 17589 15892 17601 15895
rect 17460 15864 17601 15892
rect 17460 15852 17466 15864
rect 17589 15861 17601 15864
rect 17635 15892 17647 15895
rect 17678 15892 17684 15904
rect 17635 15864 17684 15892
rect 17635 15861 17647 15864
rect 17589 15855 17647 15861
rect 17678 15852 17684 15864
rect 17736 15852 17742 15904
rect 19334 15852 19340 15904
rect 19392 15892 19398 15904
rect 19429 15895 19487 15901
rect 19429 15892 19441 15895
rect 19392 15864 19441 15892
rect 19392 15852 19398 15864
rect 19429 15861 19441 15864
rect 19475 15861 19487 15895
rect 19429 15855 19487 15861
rect 20622 15852 20628 15904
rect 20680 15892 20686 15904
rect 22281 15895 22339 15901
rect 22281 15892 22293 15895
rect 20680 15864 22293 15892
rect 20680 15852 20686 15864
rect 22281 15861 22293 15864
rect 22327 15892 22339 15895
rect 22480 15892 22508 15991
rect 22922 15988 22928 16000
rect 22980 15988 22986 16040
rect 23768 16028 23796 16068
rect 23842 16056 23848 16108
rect 23900 16096 23906 16108
rect 24213 16099 24271 16105
rect 24213 16096 24225 16099
rect 23900 16068 24225 16096
rect 23900 16056 23906 16068
rect 24213 16065 24225 16068
rect 24259 16096 24271 16099
rect 25038 16096 25044 16108
rect 24259 16068 25044 16096
rect 24259 16065 24271 16068
rect 24213 16059 24271 16065
rect 25038 16056 25044 16068
rect 25096 16056 25102 16108
rect 24670 16028 24676 16040
rect 23768 16000 24676 16028
rect 24670 15988 24676 16000
rect 24728 15988 24734 16040
rect 25225 16031 25283 16037
rect 25225 15997 25237 16031
rect 25271 16028 25283 16031
rect 25590 16028 25596 16040
rect 25271 16000 25596 16028
rect 25271 15997 25283 16000
rect 25225 15991 25283 15997
rect 25590 15988 25596 16000
rect 25648 16028 25654 16040
rect 25961 16031 26019 16037
rect 25961 16028 25973 16031
rect 25648 16000 25973 16028
rect 25648 15988 25654 16000
rect 25961 15997 25973 16000
rect 26007 15997 26019 16031
rect 25961 15991 26019 15997
rect 24029 15963 24087 15969
rect 24029 15960 24041 15963
rect 23584 15932 24041 15960
rect 23584 15904 23612 15932
rect 24029 15929 24041 15932
rect 24075 15929 24087 15963
rect 24029 15923 24087 15929
rect 24854 15920 24860 15972
rect 24912 15960 24918 15972
rect 25501 15963 25559 15969
rect 25501 15960 25513 15963
rect 24912 15932 25513 15960
rect 24912 15920 24918 15932
rect 25501 15929 25513 15932
rect 25547 15929 25559 15963
rect 25501 15923 25559 15929
rect 22327 15864 22508 15892
rect 22327 15861 22339 15864
rect 22281 15855 22339 15861
rect 22554 15852 22560 15904
rect 22612 15892 22618 15904
rect 22649 15895 22707 15901
rect 22649 15892 22661 15895
rect 22612 15864 22661 15892
rect 22612 15852 22618 15864
rect 22649 15861 22661 15864
rect 22695 15861 22707 15895
rect 22649 15855 22707 15861
rect 23477 15895 23535 15901
rect 23477 15861 23489 15895
rect 23523 15892 23535 15895
rect 23566 15892 23572 15904
rect 23523 15864 23572 15892
rect 23523 15861 23535 15864
rect 23477 15855 23535 15861
rect 23566 15852 23572 15864
rect 23624 15852 23630 15904
rect 23842 15852 23848 15904
rect 23900 15892 23906 15904
rect 24121 15895 24179 15901
rect 24121 15892 24133 15895
rect 23900 15864 24133 15892
rect 23900 15852 23906 15864
rect 24121 15861 24133 15864
rect 24167 15861 24179 15895
rect 24121 15855 24179 15861
rect 26234 15852 26240 15904
rect 26292 15892 26298 15904
rect 26329 15895 26387 15901
rect 26329 15892 26341 15895
rect 26292 15864 26341 15892
rect 26292 15852 26298 15864
rect 26329 15861 26341 15864
rect 26375 15861 26387 15895
rect 26329 15855 26387 15861
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 2682 15688 2688 15700
rect 2643 15660 2688 15688
rect 2682 15648 2688 15660
rect 2740 15648 2746 15700
rect 3142 15648 3148 15700
rect 3200 15688 3206 15700
rect 4525 15691 4583 15697
rect 4525 15688 4537 15691
rect 3200 15660 4537 15688
rect 3200 15648 3206 15660
rect 4525 15657 4537 15660
rect 4571 15688 4583 15691
rect 5074 15688 5080 15700
rect 4571 15660 5080 15688
rect 4571 15657 4583 15660
rect 4525 15651 4583 15657
rect 5074 15648 5080 15660
rect 5132 15648 5138 15700
rect 5169 15691 5227 15697
rect 5169 15657 5181 15691
rect 5215 15688 5227 15691
rect 5442 15688 5448 15700
rect 5215 15660 5448 15688
rect 5215 15657 5227 15660
rect 5169 15651 5227 15657
rect 5442 15648 5448 15660
rect 5500 15648 5506 15700
rect 5718 15688 5724 15700
rect 5679 15660 5724 15688
rect 5718 15648 5724 15660
rect 5776 15648 5782 15700
rect 6086 15688 6092 15700
rect 6047 15660 6092 15688
rect 6086 15648 6092 15660
rect 6144 15648 6150 15700
rect 8573 15691 8631 15697
rect 8573 15688 8585 15691
rect 6196 15660 8585 15688
rect 2593 15623 2651 15629
rect 2593 15589 2605 15623
rect 2639 15620 2651 15623
rect 3697 15623 3755 15629
rect 3697 15620 3709 15623
rect 2639 15592 3709 15620
rect 2639 15589 2651 15592
rect 2593 15583 2651 15589
rect 3697 15589 3709 15592
rect 3743 15620 3755 15623
rect 4062 15620 4068 15632
rect 3743 15592 4068 15620
rect 3743 15589 3755 15592
rect 3697 15583 3755 15589
rect 4062 15580 4068 15592
rect 4120 15580 4126 15632
rect 4890 15580 4896 15632
rect 4948 15620 4954 15632
rect 5258 15620 5264 15632
rect 4948 15592 5264 15620
rect 4948 15580 4954 15592
rect 5258 15580 5264 15592
rect 5316 15580 5322 15632
rect 6196 15620 6224 15660
rect 8573 15657 8585 15660
rect 8619 15657 8631 15691
rect 8573 15651 8631 15657
rect 8938 15648 8944 15700
rect 8996 15688 9002 15700
rect 9214 15688 9220 15700
rect 8996 15660 9220 15688
rect 8996 15648 9002 15660
rect 9214 15648 9220 15660
rect 9272 15648 9278 15700
rect 9674 15688 9680 15700
rect 9635 15660 9680 15688
rect 9674 15648 9680 15660
rect 9732 15648 9738 15700
rect 9858 15648 9864 15700
rect 9916 15688 9922 15700
rect 10321 15691 10379 15697
rect 10321 15688 10333 15691
rect 9916 15660 10333 15688
rect 9916 15648 9922 15660
rect 10321 15657 10333 15660
rect 10367 15688 10379 15691
rect 10778 15688 10784 15700
rect 10367 15660 10784 15688
rect 10367 15657 10379 15660
rect 10321 15651 10379 15657
rect 10778 15648 10784 15660
rect 10836 15648 10842 15700
rect 11974 15648 11980 15700
rect 12032 15688 12038 15700
rect 12069 15691 12127 15697
rect 12069 15688 12081 15691
rect 12032 15660 12081 15688
rect 12032 15648 12038 15660
rect 12069 15657 12081 15660
rect 12115 15657 12127 15691
rect 12069 15651 12127 15657
rect 12710 15648 12716 15700
rect 12768 15688 12774 15700
rect 13173 15691 13231 15697
rect 13173 15688 13185 15691
rect 12768 15660 13185 15688
rect 12768 15648 12774 15660
rect 13173 15657 13185 15660
rect 13219 15657 13231 15691
rect 13173 15651 13231 15657
rect 14277 15691 14335 15697
rect 14277 15657 14289 15691
rect 14323 15688 14335 15691
rect 14366 15688 14372 15700
rect 14323 15660 14372 15688
rect 14323 15657 14335 15660
rect 14277 15651 14335 15657
rect 14366 15648 14372 15660
rect 14424 15648 14430 15700
rect 16482 15648 16488 15700
rect 16540 15688 16546 15700
rect 16577 15691 16635 15697
rect 16577 15688 16589 15691
rect 16540 15660 16589 15688
rect 16540 15648 16546 15660
rect 16577 15657 16589 15660
rect 16623 15657 16635 15691
rect 16577 15651 16635 15657
rect 19426 15648 19432 15700
rect 19484 15688 19490 15700
rect 19613 15691 19671 15697
rect 19613 15688 19625 15691
rect 19484 15660 19625 15688
rect 19484 15648 19490 15660
rect 19613 15657 19625 15660
rect 19659 15657 19671 15691
rect 19613 15651 19671 15657
rect 20349 15691 20407 15697
rect 20349 15657 20361 15691
rect 20395 15688 20407 15691
rect 20990 15688 20996 15700
rect 20395 15660 20996 15688
rect 20395 15657 20407 15660
rect 20349 15651 20407 15657
rect 20990 15648 20996 15660
rect 21048 15648 21054 15700
rect 21634 15648 21640 15700
rect 21692 15688 21698 15700
rect 21913 15691 21971 15697
rect 21913 15688 21925 15691
rect 21692 15660 21925 15688
rect 21692 15648 21698 15660
rect 21913 15657 21925 15660
rect 21959 15657 21971 15691
rect 21913 15651 21971 15657
rect 22186 15648 22192 15700
rect 22244 15688 22250 15700
rect 22465 15691 22523 15697
rect 22465 15688 22477 15691
rect 22244 15660 22477 15688
rect 22244 15648 22250 15660
rect 22465 15657 22477 15660
rect 22511 15657 22523 15691
rect 22465 15651 22523 15657
rect 22833 15691 22891 15697
rect 22833 15657 22845 15691
rect 22879 15688 22891 15691
rect 24029 15691 24087 15697
rect 24029 15688 24041 15691
rect 22879 15660 24041 15688
rect 22879 15657 22891 15660
rect 22833 15651 22891 15657
rect 24029 15657 24041 15660
rect 24075 15657 24087 15691
rect 25038 15688 25044 15700
rect 24999 15660 25044 15688
rect 24029 15651 24087 15657
rect 5460 15592 6224 15620
rect 5077 15555 5135 15561
rect 5077 15521 5089 15555
rect 5123 15552 5135 15555
rect 5166 15552 5172 15564
rect 5123 15524 5172 15552
rect 5123 15521 5135 15524
rect 5077 15515 5135 15521
rect 5166 15512 5172 15524
rect 5224 15512 5230 15564
rect 2314 15444 2320 15496
rect 2372 15484 2378 15496
rect 2777 15487 2835 15493
rect 2777 15484 2789 15487
rect 2372 15456 2789 15484
rect 2372 15444 2378 15456
rect 2777 15453 2789 15456
rect 2823 15453 2835 15487
rect 2777 15447 2835 15453
rect 2958 15444 2964 15496
rect 3016 15484 3022 15496
rect 3237 15487 3295 15493
rect 3237 15484 3249 15487
rect 3016 15456 3249 15484
rect 3016 15444 3022 15456
rect 3237 15453 3249 15456
rect 3283 15484 3295 15487
rect 3418 15484 3424 15496
rect 3283 15456 3424 15484
rect 3283 15453 3295 15456
rect 3237 15447 3295 15453
rect 3418 15444 3424 15456
rect 3476 15444 3482 15496
rect 5258 15444 5264 15496
rect 5316 15484 5322 15496
rect 5316 15456 5361 15484
rect 5316 15444 5322 15456
rect 1854 15376 1860 15428
rect 1912 15416 1918 15428
rect 2225 15419 2283 15425
rect 2225 15416 2237 15419
rect 1912 15388 2237 15416
rect 1912 15376 1918 15388
rect 2225 15385 2237 15388
rect 2271 15385 2283 15419
rect 2225 15379 2283 15385
rect 2498 15376 2504 15428
rect 2556 15416 2562 15428
rect 3142 15416 3148 15428
rect 2556 15388 3148 15416
rect 2556 15376 2562 15388
rect 3142 15376 3148 15388
rect 3200 15376 3206 15428
rect 4706 15416 4712 15428
rect 4667 15388 4712 15416
rect 4706 15376 4712 15388
rect 4764 15376 4770 15428
rect 1673 15351 1731 15357
rect 1673 15317 1685 15351
rect 1719 15348 1731 15351
rect 2038 15348 2044 15360
rect 1719 15320 2044 15348
rect 1719 15317 1731 15320
rect 1673 15311 1731 15317
rect 2038 15308 2044 15320
rect 2096 15308 2102 15360
rect 2590 15308 2596 15360
rect 2648 15348 2654 15360
rect 5460 15348 5488 15592
rect 6270 15580 6276 15632
rect 6328 15620 6334 15632
rect 6518 15623 6576 15629
rect 6518 15620 6530 15623
rect 6328 15592 6530 15620
rect 6328 15580 6334 15592
rect 6518 15589 6530 15592
rect 6564 15589 6576 15623
rect 8294 15620 8300 15632
rect 8255 15592 8300 15620
rect 6518 15583 6576 15589
rect 8294 15580 8300 15592
rect 8352 15580 8358 15632
rect 10956 15623 11014 15629
rect 10956 15589 10968 15623
rect 11002 15620 11014 15623
rect 11146 15620 11152 15632
rect 11002 15592 11152 15620
rect 11002 15589 11014 15592
rect 10956 15583 11014 15589
rect 11146 15580 11152 15592
rect 11204 15580 11210 15632
rect 13541 15623 13599 15629
rect 13541 15589 13553 15623
rect 13587 15620 13599 15623
rect 13722 15620 13728 15632
rect 13587 15592 13728 15620
rect 13587 15589 13599 15592
rect 13541 15583 13599 15589
rect 13722 15580 13728 15592
rect 13780 15580 13786 15632
rect 15838 15620 15844 15632
rect 15799 15592 15844 15620
rect 15838 15580 15844 15592
rect 15896 15580 15902 15632
rect 20714 15580 20720 15632
rect 20772 15620 20778 15632
rect 21361 15623 21419 15629
rect 21361 15620 21373 15623
rect 20772 15592 21373 15620
rect 20772 15580 20778 15592
rect 21361 15589 21373 15592
rect 21407 15589 21419 15623
rect 21361 15583 21419 15589
rect 22373 15623 22431 15629
rect 22373 15589 22385 15623
rect 22419 15620 22431 15623
rect 22848 15620 22876 15651
rect 25038 15648 25044 15660
rect 25096 15648 25102 15700
rect 26237 15691 26295 15697
rect 26237 15657 26249 15691
rect 26283 15688 26295 15691
rect 26326 15688 26332 15700
rect 26283 15660 26332 15688
rect 26283 15657 26295 15660
rect 26237 15651 26295 15657
rect 26326 15648 26332 15660
rect 26384 15648 26390 15700
rect 22419 15592 22876 15620
rect 22419 15589 22431 15592
rect 22373 15583 22431 15589
rect 23750 15580 23756 15632
rect 23808 15620 23814 15632
rect 24397 15623 24455 15629
rect 24397 15620 24409 15623
rect 23808 15592 24409 15620
rect 23808 15580 23814 15592
rect 24397 15589 24409 15592
rect 24443 15620 24455 15623
rect 24670 15620 24676 15632
rect 24443 15592 24676 15620
rect 24443 15589 24455 15592
rect 24397 15583 24455 15589
rect 24670 15580 24676 15592
rect 24728 15580 24734 15632
rect 6086 15512 6092 15564
rect 6144 15552 6150 15564
rect 6362 15552 6368 15564
rect 6144 15524 6368 15552
rect 6144 15512 6150 15524
rect 6362 15512 6368 15524
rect 6420 15512 6426 15564
rect 8941 15555 8999 15561
rect 8941 15521 8953 15555
rect 8987 15552 8999 15555
rect 9122 15552 9128 15564
rect 8987 15524 9128 15552
rect 8987 15521 8999 15524
rect 8941 15515 8999 15521
rect 9122 15512 9128 15524
rect 9180 15512 9186 15564
rect 10689 15555 10747 15561
rect 10689 15521 10701 15555
rect 10735 15552 10747 15555
rect 11790 15552 11796 15564
rect 10735 15524 11796 15552
rect 10735 15521 10747 15524
rect 10689 15515 10747 15521
rect 6273 15487 6331 15493
rect 6273 15453 6285 15487
rect 6319 15453 6331 15487
rect 6273 15447 6331 15453
rect 2648 15320 5488 15348
rect 6288 15348 6316 15447
rect 8757 15419 8815 15425
rect 8757 15385 8769 15419
rect 8803 15416 8815 15419
rect 9766 15416 9772 15428
rect 8803 15388 9772 15416
rect 8803 15385 8815 15388
rect 8757 15379 8815 15385
rect 9766 15376 9772 15388
rect 9824 15416 9830 15428
rect 10704 15416 10732 15515
rect 11790 15512 11796 15524
rect 11848 15512 11854 15564
rect 16482 15552 16488 15564
rect 16443 15524 16488 15552
rect 16482 15512 16488 15524
rect 16540 15512 16546 15564
rect 18049 15555 18107 15561
rect 18049 15552 18061 15555
rect 17144 15524 18061 15552
rect 13630 15484 13636 15496
rect 13591 15456 13636 15484
rect 13630 15444 13636 15456
rect 13688 15444 13694 15496
rect 13725 15487 13783 15493
rect 13725 15453 13737 15487
rect 13771 15453 13783 15487
rect 16666 15484 16672 15496
rect 16627 15456 16672 15484
rect 13725 15447 13783 15453
rect 9824 15388 10732 15416
rect 9824 15376 9830 15388
rect 7282 15348 7288 15360
rect 6288 15320 7288 15348
rect 2648 15308 2654 15320
rect 7282 15308 7288 15320
rect 7340 15308 7346 15360
rect 7650 15348 7656 15360
rect 7611 15320 7656 15348
rect 7650 15308 7656 15320
rect 7708 15308 7714 15360
rect 8294 15308 8300 15360
rect 8352 15348 8358 15360
rect 9490 15348 9496 15360
rect 8352 15320 9496 15348
rect 8352 15308 8358 15320
rect 9490 15308 9496 15320
rect 9548 15308 9554 15360
rect 12713 15351 12771 15357
rect 12713 15317 12725 15351
rect 12759 15348 12771 15351
rect 12802 15348 12808 15360
rect 12759 15320 12808 15348
rect 12759 15317 12771 15320
rect 12713 15311 12771 15317
rect 12802 15308 12808 15320
rect 12860 15348 12866 15360
rect 12989 15351 13047 15357
rect 12989 15348 13001 15351
rect 12860 15320 13001 15348
rect 12860 15308 12866 15320
rect 12989 15317 13001 15320
rect 13035 15348 13047 15351
rect 13740 15348 13768 15447
rect 16666 15444 16672 15456
rect 16724 15444 16730 15496
rect 17144 15425 17172 15524
rect 18049 15521 18061 15524
rect 18095 15521 18107 15555
rect 18049 15515 18107 15521
rect 21269 15555 21327 15561
rect 21269 15521 21281 15555
rect 21315 15552 21327 15555
rect 21542 15552 21548 15564
rect 21315 15524 21548 15552
rect 21315 15521 21327 15524
rect 21269 15515 21327 15521
rect 21542 15512 21548 15524
rect 21600 15512 21606 15564
rect 22922 15552 22928 15564
rect 22883 15524 22928 15552
rect 22922 15512 22928 15524
rect 22980 15512 22986 15564
rect 17589 15487 17647 15493
rect 17589 15453 17601 15487
rect 17635 15484 17647 15487
rect 17954 15484 17960 15496
rect 17635 15456 17960 15484
rect 17635 15453 17647 15456
rect 17589 15447 17647 15453
rect 17954 15444 17960 15456
rect 18012 15484 18018 15496
rect 18141 15487 18199 15493
rect 18141 15484 18153 15487
rect 18012 15456 18153 15484
rect 18012 15444 18018 15456
rect 18141 15453 18153 15456
rect 18187 15453 18199 15487
rect 18141 15447 18199 15453
rect 18325 15487 18383 15493
rect 18325 15453 18337 15487
rect 18371 15484 18383 15487
rect 18414 15484 18420 15496
rect 18371 15456 18420 15484
rect 18371 15453 18383 15456
rect 18325 15447 18383 15453
rect 18414 15444 18420 15456
rect 18472 15444 18478 15496
rect 19702 15484 19708 15496
rect 19663 15456 19708 15484
rect 19702 15444 19708 15456
rect 19760 15444 19766 15496
rect 19797 15487 19855 15493
rect 19797 15453 19809 15487
rect 19843 15453 19855 15487
rect 19797 15447 19855 15453
rect 21453 15487 21511 15493
rect 21453 15453 21465 15487
rect 21499 15453 21511 15487
rect 21453 15447 21511 15453
rect 16117 15419 16175 15425
rect 16117 15385 16129 15419
rect 16163 15416 16175 15419
rect 17129 15419 17187 15425
rect 17129 15416 17141 15419
rect 16163 15388 17141 15416
rect 16163 15385 16175 15388
rect 16117 15379 16175 15385
rect 17129 15385 17141 15388
rect 17175 15385 17187 15419
rect 17129 15379 17187 15385
rect 17494 15376 17500 15428
rect 17552 15416 17558 15428
rect 19245 15419 19303 15425
rect 19245 15416 19257 15419
rect 17552 15388 19257 15416
rect 17552 15376 17558 15388
rect 19245 15385 19257 15388
rect 19291 15385 19303 15419
rect 19812 15416 19840 15447
rect 19245 15379 19303 15385
rect 19536 15388 19840 15416
rect 20717 15419 20775 15425
rect 19536 15360 19564 15388
rect 20717 15385 20729 15419
rect 20763 15416 20775 15419
rect 21174 15416 21180 15428
rect 20763 15388 21180 15416
rect 20763 15385 20775 15388
rect 20717 15379 20775 15385
rect 21174 15376 21180 15388
rect 21232 15416 21238 15428
rect 21468 15416 21496 15447
rect 22002 15444 22008 15496
rect 22060 15484 22066 15496
rect 23014 15484 23020 15496
rect 22060 15456 23020 15484
rect 22060 15444 22066 15456
rect 23014 15444 23020 15456
rect 23072 15444 23078 15496
rect 23753 15487 23811 15493
rect 23753 15453 23765 15487
rect 23799 15484 23811 15487
rect 23842 15484 23848 15496
rect 23799 15456 23848 15484
rect 23799 15453 23811 15456
rect 23753 15447 23811 15453
rect 23842 15444 23848 15456
rect 23900 15444 23906 15496
rect 24026 15444 24032 15496
rect 24084 15484 24090 15496
rect 24489 15487 24547 15493
rect 24489 15484 24501 15487
rect 24084 15456 24501 15484
rect 24084 15444 24090 15456
rect 24489 15453 24501 15456
rect 24535 15453 24547 15487
rect 24489 15447 24547 15453
rect 24673 15487 24731 15493
rect 24673 15453 24685 15487
rect 24719 15484 24731 15487
rect 25222 15484 25228 15496
rect 24719 15456 25228 15484
rect 24719 15453 24731 15456
rect 24673 15447 24731 15453
rect 21232 15388 21496 15416
rect 24504 15416 24532 15447
rect 25222 15444 25228 15456
rect 25280 15444 25286 15496
rect 25409 15419 25467 15425
rect 25409 15416 25421 15419
rect 24504 15388 25421 15416
rect 21232 15376 21238 15388
rect 25409 15385 25421 15388
rect 25455 15385 25467 15419
rect 25409 15379 25467 15385
rect 14642 15348 14648 15360
rect 13035 15320 13768 15348
rect 14603 15320 14648 15348
rect 13035 15317 13047 15320
rect 12989 15311 13047 15317
rect 14642 15308 14648 15320
rect 14700 15348 14706 15360
rect 14921 15351 14979 15357
rect 14921 15348 14933 15351
rect 14700 15320 14933 15348
rect 14700 15308 14706 15320
rect 14921 15317 14933 15320
rect 14967 15317 14979 15351
rect 14921 15311 14979 15317
rect 15286 15308 15292 15360
rect 15344 15348 15350 15360
rect 15473 15351 15531 15357
rect 15473 15348 15485 15351
rect 15344 15320 15485 15348
rect 15344 15308 15350 15320
rect 15473 15317 15485 15320
rect 15519 15348 15531 15351
rect 15930 15348 15936 15360
rect 15519 15320 15936 15348
rect 15519 15317 15531 15320
rect 15473 15311 15531 15317
rect 15930 15308 15936 15320
rect 15988 15308 15994 15360
rect 17681 15351 17739 15357
rect 17681 15317 17693 15351
rect 17727 15348 17739 15351
rect 17862 15348 17868 15360
rect 17727 15320 17868 15348
rect 17727 15317 17739 15320
rect 17681 15311 17739 15317
rect 17862 15308 17868 15320
rect 17920 15308 17926 15360
rect 18598 15308 18604 15360
rect 18656 15348 18662 15360
rect 18785 15351 18843 15357
rect 18785 15348 18797 15351
rect 18656 15320 18797 15348
rect 18656 15308 18662 15320
rect 18785 15317 18797 15320
rect 18831 15348 18843 15351
rect 19153 15351 19211 15357
rect 19153 15348 19165 15351
rect 18831 15320 19165 15348
rect 18831 15317 18843 15320
rect 18785 15311 18843 15317
rect 19153 15317 19165 15320
rect 19199 15348 19211 15351
rect 19518 15348 19524 15360
rect 19199 15320 19524 15348
rect 19199 15317 19211 15320
rect 19153 15311 19211 15317
rect 19518 15308 19524 15320
rect 19576 15308 19582 15360
rect 20898 15348 20904 15360
rect 20859 15320 20904 15348
rect 20898 15308 20904 15320
rect 20956 15308 20962 15360
rect 23106 15308 23112 15360
rect 23164 15348 23170 15360
rect 23382 15348 23388 15360
rect 23164 15320 23388 15348
rect 23164 15308 23170 15320
rect 23382 15308 23388 15320
rect 23440 15308 23446 15360
rect 25682 15308 25688 15360
rect 25740 15348 25746 15360
rect 25777 15351 25835 15357
rect 25777 15348 25789 15351
rect 25740 15320 25789 15348
rect 25740 15308 25746 15320
rect 25777 15317 25789 15320
rect 25823 15317 25835 15351
rect 25777 15311 25835 15317
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 3050 15144 3056 15156
rect 1504 15116 3056 15144
rect 1504 14949 1532 15116
rect 3050 15104 3056 15116
rect 3108 15104 3114 15156
rect 4801 15147 4859 15153
rect 4801 15113 4813 15147
rect 4847 15144 4859 15147
rect 5258 15144 5264 15156
rect 4847 15116 5264 15144
rect 4847 15113 4859 15116
rect 4801 15107 4859 15113
rect 5258 15104 5264 15116
rect 5316 15104 5322 15156
rect 8754 15104 8760 15156
rect 8812 15144 8818 15156
rect 11054 15144 11060 15156
rect 8812 15116 11060 15144
rect 8812 15104 8818 15116
rect 11054 15104 11060 15116
rect 11112 15104 11118 15156
rect 11146 15104 11152 15156
rect 11204 15144 11210 15156
rect 11241 15147 11299 15153
rect 11241 15144 11253 15147
rect 11204 15116 11253 15144
rect 11204 15104 11210 15116
rect 11241 15113 11253 15116
rect 11287 15113 11299 15147
rect 11241 15107 11299 15113
rect 12342 15104 12348 15156
rect 12400 15144 12406 15156
rect 12437 15147 12495 15153
rect 12437 15144 12449 15147
rect 12400 15116 12449 15144
rect 12400 15104 12406 15116
rect 12437 15113 12449 15116
rect 12483 15113 12495 15147
rect 12437 15107 12495 15113
rect 16209 15147 16267 15153
rect 16209 15113 16221 15147
rect 16255 15144 16267 15147
rect 16390 15144 16396 15156
rect 16255 15116 16396 15144
rect 16255 15113 16267 15116
rect 16209 15107 16267 15113
rect 16390 15104 16396 15116
rect 16448 15104 16454 15156
rect 18230 15144 18236 15156
rect 18064 15116 18236 15144
rect 2314 15076 2320 15088
rect 2275 15048 2320 15076
rect 2314 15036 2320 15048
rect 2372 15036 2378 15088
rect 9122 15076 9128 15088
rect 9083 15048 9128 15076
rect 9122 15036 9128 15048
rect 9180 15036 9186 15088
rect 12526 15036 12532 15088
rect 12584 15076 12590 15088
rect 13814 15076 13820 15088
rect 12584 15048 13820 15076
rect 12584 15036 12590 15048
rect 13814 15036 13820 15048
rect 13872 15036 13878 15088
rect 9140 15008 9168 15036
rect 12989 15011 13047 15017
rect 9140 14980 9444 15008
rect 1489 14943 1547 14949
rect 1489 14909 1501 14943
rect 1535 14909 1547 14943
rect 1489 14903 1547 14909
rect 1578 14900 1584 14952
rect 1636 14940 1642 14952
rect 2777 14943 2835 14949
rect 2777 14940 2789 14943
rect 1636 14912 2789 14940
rect 1636 14900 1642 14912
rect 2777 14909 2789 14912
rect 2823 14940 2835 14943
rect 3786 14940 3792 14952
rect 2823 14912 3792 14940
rect 2823 14909 2835 14912
rect 2777 14903 2835 14909
rect 3786 14900 3792 14912
rect 3844 14900 3850 14952
rect 5261 14943 5319 14949
rect 5261 14940 5273 14943
rect 5092 14912 5273 14940
rect 1762 14872 1768 14884
rect 1723 14844 1768 14872
rect 1762 14832 1768 14844
rect 1820 14832 1826 14884
rect 2498 14832 2504 14884
rect 2556 14872 2562 14884
rect 2685 14875 2743 14881
rect 2685 14872 2697 14875
rect 2556 14844 2697 14872
rect 2556 14832 2562 14844
rect 2685 14841 2697 14844
rect 2731 14872 2743 14875
rect 3022 14875 3080 14881
rect 3022 14872 3034 14875
rect 2731 14844 3034 14872
rect 2731 14841 2743 14844
rect 2685 14835 2743 14841
rect 3022 14841 3034 14844
rect 3068 14841 3080 14875
rect 3022 14835 3080 14841
rect 5092 14816 5120 14912
rect 5261 14909 5273 14912
rect 5307 14909 5319 14943
rect 6822 14940 6828 14952
rect 6783 14912 6828 14940
rect 5261 14903 5319 14909
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 6914 14900 6920 14952
rect 6972 14940 6978 14952
rect 7081 14943 7139 14949
rect 7081 14940 7093 14943
rect 6972 14912 7093 14940
rect 6972 14900 6978 14912
rect 7081 14909 7093 14912
rect 7127 14909 7139 14943
rect 7081 14903 7139 14909
rect 9309 14943 9367 14949
rect 9309 14909 9321 14943
rect 9355 14909 9367 14943
rect 9416 14940 9444 14980
rect 12989 14977 13001 15011
rect 13035 14977 13047 15011
rect 12989 14971 13047 14977
rect 9565 14943 9623 14949
rect 9565 14940 9577 14943
rect 9416 14912 9577 14940
rect 9309 14903 9367 14909
rect 9565 14909 9577 14912
rect 9611 14909 9623 14943
rect 9565 14903 9623 14909
rect 5537 14875 5595 14881
rect 5537 14841 5549 14875
rect 5583 14872 5595 14875
rect 5583 14844 7052 14872
rect 5583 14841 5595 14844
rect 5537 14835 5595 14841
rect 4157 14807 4215 14813
rect 4157 14773 4169 14807
rect 4203 14804 4215 14807
rect 4706 14804 4712 14816
rect 4203 14776 4712 14804
rect 4203 14773 4215 14776
rect 4157 14767 4215 14773
rect 4706 14764 4712 14776
rect 4764 14764 4770 14816
rect 5074 14804 5080 14816
rect 5035 14776 5080 14804
rect 5074 14764 5080 14776
rect 5132 14764 5138 14816
rect 6270 14804 6276 14816
rect 6231 14776 6276 14804
rect 6270 14764 6276 14776
rect 6328 14764 6334 14816
rect 6362 14764 6368 14816
rect 6420 14804 6426 14816
rect 6549 14807 6607 14813
rect 6549 14804 6561 14807
rect 6420 14776 6561 14804
rect 6420 14764 6426 14776
rect 6549 14773 6561 14776
rect 6595 14804 6607 14807
rect 6914 14804 6920 14816
rect 6595 14776 6920 14804
rect 6595 14773 6607 14776
rect 6549 14767 6607 14773
rect 6914 14764 6920 14776
rect 6972 14764 6978 14816
rect 7024 14804 7052 14844
rect 7558 14832 7564 14884
rect 7616 14872 7622 14884
rect 8757 14875 8815 14881
rect 8757 14872 8769 14875
rect 7616 14844 8769 14872
rect 7616 14832 7622 14844
rect 8757 14841 8769 14844
rect 8803 14841 8815 14875
rect 9324 14872 9352 14903
rect 10042 14900 10048 14952
rect 10100 14940 10106 14952
rect 10778 14940 10784 14952
rect 10100 14912 10784 14940
rect 10100 14900 10106 14912
rect 10778 14900 10784 14912
rect 10836 14900 10842 14952
rect 11054 14900 11060 14952
rect 11112 14940 11118 14952
rect 12161 14943 12219 14949
rect 12161 14940 12173 14943
rect 11112 14912 12173 14940
rect 11112 14900 11118 14912
rect 12161 14909 12173 14912
rect 12207 14940 12219 14943
rect 13004 14940 13032 14971
rect 17034 14968 17040 15020
rect 17092 15008 17098 15020
rect 17402 15008 17408 15020
rect 17092 14980 17408 15008
rect 17092 14968 17098 14980
rect 17402 14968 17408 14980
rect 17460 14968 17466 15020
rect 18064 15017 18092 15116
rect 18230 15104 18236 15116
rect 18288 15104 18294 15156
rect 18414 15104 18420 15156
rect 18472 15144 18478 15156
rect 19429 15147 19487 15153
rect 19429 15144 19441 15147
rect 18472 15116 19441 15144
rect 18472 15104 18478 15116
rect 19429 15113 19441 15116
rect 19475 15113 19487 15147
rect 20438 15144 20444 15156
rect 20351 15116 20444 15144
rect 19429 15107 19487 15113
rect 20438 15104 20444 15116
rect 20496 15144 20502 15156
rect 20714 15144 20720 15156
rect 20496 15116 20720 15144
rect 20496 15104 20502 15116
rect 20714 15104 20720 15116
rect 20772 15104 20778 15156
rect 22370 15144 22376 15156
rect 22331 15116 22376 15144
rect 22370 15104 22376 15116
rect 22428 15104 22434 15156
rect 23014 15144 23020 15156
rect 22975 15116 23020 15144
rect 23014 15104 23020 15116
rect 23072 15104 23078 15156
rect 24670 15144 24676 15156
rect 24631 15116 24676 15144
rect 24670 15104 24676 15116
rect 24728 15104 24734 15156
rect 26326 15144 26332 15156
rect 26287 15116 26332 15144
rect 26326 15104 26332 15116
rect 26384 15104 26390 15156
rect 22388 15076 22416 15104
rect 23385 15079 23443 15085
rect 23385 15076 23397 15079
rect 22388 15048 23397 15076
rect 23385 15045 23397 15048
rect 23431 15076 23443 15079
rect 23566 15076 23572 15088
rect 23431 15048 23572 15076
rect 23431 15045 23443 15048
rect 23385 15039 23443 15045
rect 23566 15036 23572 15048
rect 23624 15076 23630 15088
rect 23624 15048 24256 15076
rect 23624 15036 23630 15048
rect 18049 15011 18107 15017
rect 18049 14977 18061 15011
rect 18095 14977 18107 15011
rect 18049 14971 18107 14977
rect 19242 14968 19248 15020
rect 19300 14968 19306 15020
rect 19426 14968 19432 15020
rect 19484 15008 19490 15020
rect 19981 15011 20039 15017
rect 19981 15008 19993 15011
rect 19484 14980 19993 15008
rect 19484 14968 19490 14980
rect 19981 14977 19993 14980
rect 20027 14977 20039 15011
rect 24118 15008 24124 15020
rect 24079 14980 24124 15008
rect 19981 14971 20039 14977
rect 24118 14968 24124 14980
rect 24176 14968 24182 15020
rect 24228 15017 24256 15048
rect 24213 15011 24271 15017
rect 24213 14977 24225 15011
rect 24259 14977 24271 15011
rect 24213 14971 24271 14977
rect 12207 14912 13032 14940
rect 12207 14909 12219 14912
rect 12161 14903 12219 14909
rect 13906 14900 13912 14952
rect 13964 14940 13970 14952
rect 14001 14943 14059 14949
rect 14001 14940 14013 14943
rect 13964 14912 14013 14940
rect 13964 14900 13970 14912
rect 14001 14909 14013 14912
rect 14047 14940 14059 14943
rect 14090 14940 14096 14952
rect 14047 14912 14096 14940
rect 14047 14909 14059 14912
rect 14001 14903 14059 14909
rect 14090 14900 14096 14912
rect 14148 14900 14154 14952
rect 15562 14900 15568 14952
rect 15620 14940 15626 14952
rect 15930 14940 15936 14952
rect 15620 14912 15936 14940
rect 15620 14900 15626 14912
rect 15930 14900 15936 14912
rect 15988 14900 15994 14952
rect 16390 14900 16396 14952
rect 16448 14940 16454 14952
rect 16853 14943 16911 14949
rect 16853 14940 16865 14943
rect 16448 14912 16865 14940
rect 16448 14900 16454 14912
rect 16853 14909 16865 14912
rect 16899 14940 16911 14943
rect 17497 14943 17555 14949
rect 17497 14940 17509 14943
rect 16899 14912 17509 14940
rect 16899 14909 16911 14912
rect 16853 14903 16911 14909
rect 17497 14909 17509 14912
rect 17543 14940 17555 14943
rect 17678 14940 17684 14952
rect 17543 14912 17684 14940
rect 17543 14909 17555 14912
rect 17497 14903 17555 14909
rect 17678 14900 17684 14912
rect 17736 14900 17742 14952
rect 17865 14943 17923 14949
rect 17865 14909 17877 14943
rect 17911 14940 17923 14943
rect 18316 14943 18374 14949
rect 18316 14940 18328 14943
rect 17911 14912 18328 14940
rect 17911 14909 17923 14912
rect 17865 14903 17923 14909
rect 18316 14909 18328 14912
rect 18362 14940 18374 14943
rect 18598 14940 18604 14952
rect 18362 14912 18604 14940
rect 18362 14909 18374 14912
rect 18316 14903 18374 14909
rect 18598 14900 18604 14912
rect 18656 14940 18662 14952
rect 19260 14940 19288 14968
rect 18656 14912 19288 14940
rect 18656 14900 18662 14912
rect 20622 14900 20628 14952
rect 20680 14940 20686 14952
rect 20717 14943 20775 14949
rect 20717 14940 20729 14943
rect 20680 14912 20729 14940
rect 20680 14900 20686 14912
rect 20717 14909 20729 14912
rect 20763 14909 20775 14943
rect 20717 14903 20775 14909
rect 20993 14943 21051 14949
rect 20993 14909 21005 14943
rect 21039 14940 21051 14943
rect 22002 14940 22008 14952
rect 21039 14912 22008 14940
rect 21039 14909 21051 14912
rect 20993 14903 21051 14909
rect 9766 14872 9772 14884
rect 9324 14844 9772 14872
rect 8757 14835 8815 14841
rect 9766 14832 9772 14844
rect 9824 14832 9830 14884
rect 12897 14875 12955 14881
rect 12897 14872 12909 14875
rect 11808 14844 12909 14872
rect 11808 14816 11836 14844
rect 12897 14841 12909 14844
rect 12943 14841 12955 14875
rect 12897 14835 12955 14841
rect 14268 14875 14326 14881
rect 14268 14841 14280 14875
rect 14314 14872 14326 14875
rect 14366 14872 14372 14884
rect 14314 14844 14372 14872
rect 14314 14841 14326 14844
rect 14268 14835 14326 14841
rect 14366 14832 14372 14844
rect 14424 14832 14430 14884
rect 19334 14832 19340 14884
rect 19392 14872 19398 14884
rect 19702 14872 19708 14884
rect 19392 14844 19708 14872
rect 19392 14832 19398 14844
rect 19702 14832 19708 14844
rect 19760 14832 19766 14884
rect 8110 14804 8116 14816
rect 7024 14776 8116 14804
rect 8110 14764 8116 14776
rect 8168 14764 8174 14816
rect 8202 14764 8208 14816
rect 8260 14804 8266 14816
rect 10686 14804 10692 14816
rect 8260 14776 8305 14804
rect 10647 14776 10692 14804
rect 8260 14764 8266 14776
rect 10686 14764 10692 14776
rect 10744 14764 10750 14816
rect 11790 14804 11796 14816
rect 11751 14776 11796 14804
rect 11790 14764 11796 14776
rect 11848 14764 11854 14816
rect 12434 14764 12440 14816
rect 12492 14804 12498 14816
rect 12805 14807 12863 14813
rect 12805 14804 12817 14807
rect 12492 14776 12817 14804
rect 12492 14764 12498 14776
rect 12805 14773 12817 14776
rect 12851 14773 12863 14807
rect 12805 14767 12863 14773
rect 13541 14807 13599 14813
rect 13541 14773 13553 14807
rect 13587 14804 13599 14807
rect 13630 14804 13636 14816
rect 13587 14776 13636 14804
rect 13587 14773 13599 14776
rect 13541 14767 13599 14773
rect 13630 14764 13636 14776
rect 13688 14764 13694 14816
rect 13722 14764 13728 14816
rect 13780 14804 13786 14816
rect 13909 14807 13967 14813
rect 13909 14804 13921 14807
rect 13780 14776 13921 14804
rect 13780 14764 13786 14776
rect 13909 14773 13921 14776
rect 13955 14804 13967 14807
rect 14090 14804 14096 14816
rect 13955 14776 14096 14804
rect 13955 14773 13967 14776
rect 13909 14767 13967 14773
rect 14090 14764 14096 14776
rect 14148 14764 14154 14816
rect 15381 14807 15439 14813
rect 15381 14773 15393 14807
rect 15427 14804 15439 14807
rect 15562 14804 15568 14816
rect 15427 14776 15568 14804
rect 15427 14773 15439 14776
rect 15381 14767 15439 14773
rect 15562 14764 15568 14776
rect 15620 14764 15626 14816
rect 16482 14804 16488 14816
rect 16443 14776 16488 14804
rect 16482 14764 16488 14776
rect 16540 14764 16546 14816
rect 17034 14804 17040 14816
rect 16995 14776 17040 14804
rect 17034 14764 17040 14776
rect 17092 14764 17098 14816
rect 18230 14764 18236 14816
rect 18288 14804 18294 14816
rect 20533 14807 20591 14813
rect 20533 14804 20545 14807
rect 18288 14776 20545 14804
rect 18288 14764 18294 14776
rect 20533 14773 20545 14776
rect 20579 14804 20591 14807
rect 21008 14804 21036 14903
rect 22002 14900 22008 14912
rect 22060 14900 22066 14952
rect 24136 14940 24164 14968
rect 25041 14943 25099 14949
rect 25041 14940 25053 14943
rect 24136 14912 25053 14940
rect 25041 14909 25053 14912
rect 25087 14909 25099 14943
rect 25041 14903 25099 14909
rect 25225 14943 25283 14949
rect 25225 14909 25237 14943
rect 25271 14940 25283 14943
rect 25406 14940 25412 14952
rect 25271 14912 25412 14940
rect 25271 14909 25283 14912
rect 25225 14903 25283 14909
rect 25406 14900 25412 14912
rect 25464 14940 25470 14952
rect 25961 14943 26019 14949
rect 25961 14940 25973 14943
rect 25464 14912 25973 14940
rect 25464 14900 25470 14912
rect 25961 14909 25973 14912
rect 26007 14909 26019 14943
rect 25961 14903 26019 14909
rect 21174 14832 21180 14884
rect 21232 14881 21238 14884
rect 21232 14875 21296 14881
rect 21232 14841 21250 14875
rect 21284 14841 21296 14875
rect 21232 14835 21296 14841
rect 21232 14832 21238 14835
rect 23014 14832 23020 14884
rect 23072 14872 23078 14884
rect 23072 14844 24900 14872
rect 23072 14832 23078 14844
rect 20579 14776 21036 14804
rect 20579 14773 20591 14776
rect 20533 14767 20591 14773
rect 22922 14764 22928 14816
rect 22980 14804 22986 14816
rect 23661 14807 23719 14813
rect 23661 14804 23673 14807
rect 22980 14776 23673 14804
rect 22980 14764 22986 14776
rect 23661 14773 23673 14776
rect 23707 14773 23719 14807
rect 24026 14804 24032 14816
rect 23987 14776 24032 14804
rect 23661 14767 23719 14773
rect 24026 14764 24032 14776
rect 24084 14764 24090 14816
rect 24872 14804 24900 14844
rect 24946 14832 24952 14884
rect 25004 14872 25010 14884
rect 25501 14875 25559 14881
rect 25501 14872 25513 14875
rect 25004 14844 25513 14872
rect 25004 14832 25010 14844
rect 25501 14841 25513 14844
rect 25547 14841 25559 14875
rect 25501 14835 25559 14841
rect 25682 14804 25688 14816
rect 24872 14776 25688 14804
rect 25682 14764 25688 14776
rect 25740 14764 25746 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1394 14600 1400 14612
rect 1355 14572 1400 14600
rect 1394 14560 1400 14572
rect 1452 14560 1458 14612
rect 2498 14600 2504 14612
rect 2459 14572 2504 14600
rect 2498 14560 2504 14572
rect 2556 14560 2562 14612
rect 3050 14560 3056 14612
rect 3108 14600 3114 14612
rect 3421 14603 3479 14609
rect 3421 14600 3433 14603
rect 3108 14572 3433 14600
rect 3108 14560 3114 14572
rect 3421 14569 3433 14572
rect 3467 14569 3479 14603
rect 3421 14563 3479 14569
rect 5350 14560 5356 14612
rect 5408 14600 5414 14612
rect 5997 14603 6055 14609
rect 5997 14600 6009 14603
rect 5408 14572 6009 14600
rect 5408 14560 5414 14572
rect 5997 14569 6009 14572
rect 6043 14569 6055 14603
rect 5997 14563 6055 14569
rect 6917 14603 6975 14609
rect 6917 14569 6929 14603
rect 6963 14600 6975 14603
rect 7098 14600 7104 14612
rect 6963 14572 7104 14600
rect 6963 14569 6975 14572
rect 6917 14563 6975 14569
rect 7098 14560 7104 14572
rect 7156 14600 7162 14612
rect 9033 14603 9091 14609
rect 9033 14600 9045 14603
rect 7156 14572 9045 14600
rect 7156 14560 7162 14572
rect 9033 14569 9045 14572
rect 9079 14569 9091 14603
rect 9214 14600 9220 14612
rect 9175 14572 9220 14600
rect 9033 14563 9091 14569
rect 9214 14560 9220 14572
rect 9272 14560 9278 14612
rect 9582 14560 9588 14612
rect 9640 14600 9646 14612
rect 10045 14603 10103 14609
rect 10045 14600 10057 14603
rect 9640 14572 10057 14600
rect 9640 14560 9646 14572
rect 10045 14569 10057 14572
rect 10091 14600 10103 14603
rect 11793 14603 11851 14609
rect 11793 14600 11805 14603
rect 10091 14572 11805 14600
rect 10091 14569 10103 14572
rect 10045 14563 10103 14569
rect 11793 14569 11805 14572
rect 11839 14569 11851 14603
rect 11793 14563 11851 14569
rect 13262 14560 13268 14612
rect 13320 14600 13326 14612
rect 13357 14603 13415 14609
rect 13357 14600 13369 14603
rect 13320 14572 13369 14600
rect 13320 14560 13326 14572
rect 13357 14569 13369 14572
rect 13403 14600 13415 14603
rect 13538 14600 13544 14612
rect 13403 14572 13544 14600
rect 13403 14569 13415 14572
rect 13357 14563 13415 14569
rect 13538 14560 13544 14572
rect 13596 14560 13602 14612
rect 15381 14603 15439 14609
rect 15381 14569 15393 14603
rect 15427 14600 15439 14603
rect 16482 14600 16488 14612
rect 15427 14572 16488 14600
rect 15427 14569 15439 14572
rect 15381 14563 15439 14569
rect 16482 14560 16488 14572
rect 16540 14560 16546 14612
rect 16853 14603 16911 14609
rect 16853 14569 16865 14603
rect 16899 14600 16911 14603
rect 17494 14600 17500 14612
rect 16899 14572 17500 14600
rect 16899 14569 16911 14572
rect 16853 14563 16911 14569
rect 17494 14560 17500 14572
rect 17552 14560 17558 14612
rect 17954 14600 17960 14612
rect 17915 14572 17960 14600
rect 17954 14560 17960 14572
rect 18012 14560 18018 14612
rect 19334 14600 19340 14612
rect 19295 14572 19340 14600
rect 19334 14560 19340 14572
rect 19392 14560 19398 14612
rect 19889 14603 19947 14609
rect 19889 14569 19901 14603
rect 19935 14600 19947 14603
rect 19978 14600 19984 14612
rect 19935 14572 19984 14600
rect 19935 14569 19947 14572
rect 19889 14563 19947 14569
rect 19978 14560 19984 14572
rect 20036 14560 20042 14612
rect 20349 14603 20407 14609
rect 20349 14569 20361 14603
rect 20395 14600 20407 14603
rect 20622 14600 20628 14612
rect 20395 14572 20628 14600
rect 20395 14569 20407 14572
rect 20349 14563 20407 14569
rect 20622 14560 20628 14572
rect 20680 14560 20686 14612
rect 20717 14603 20775 14609
rect 20717 14569 20729 14603
rect 20763 14600 20775 14603
rect 21174 14600 21180 14612
rect 20763 14572 21180 14600
rect 20763 14569 20775 14572
rect 20717 14563 20775 14569
rect 21174 14560 21180 14572
rect 21232 14560 21238 14612
rect 21729 14603 21787 14609
rect 21729 14569 21741 14603
rect 21775 14600 21787 14603
rect 21910 14600 21916 14612
rect 21775 14572 21916 14600
rect 21775 14569 21787 14572
rect 21729 14563 21787 14569
rect 21910 14560 21916 14572
rect 21968 14560 21974 14612
rect 22557 14603 22615 14609
rect 22557 14569 22569 14603
rect 22603 14600 22615 14603
rect 22922 14600 22928 14612
rect 22603 14572 22928 14600
rect 22603 14569 22615 14572
rect 22557 14563 22615 14569
rect 22922 14560 22928 14572
rect 22980 14560 22986 14612
rect 23385 14603 23443 14609
rect 23385 14569 23397 14603
rect 23431 14600 23443 14603
rect 24026 14600 24032 14612
rect 23431 14572 24032 14600
rect 23431 14569 23443 14572
rect 23385 14563 23443 14569
rect 1670 14492 1676 14544
rect 1728 14532 1734 14544
rect 1765 14535 1823 14541
rect 1765 14532 1777 14535
rect 1728 14504 1777 14532
rect 1728 14492 1734 14504
rect 1765 14501 1777 14504
rect 1811 14532 1823 14535
rect 2406 14532 2412 14544
rect 1811 14504 2412 14532
rect 1811 14501 1823 14504
rect 1765 14495 1823 14501
rect 2406 14492 2412 14504
rect 2464 14492 2470 14544
rect 3786 14492 3792 14544
rect 3844 14532 3850 14544
rect 4890 14532 4896 14544
rect 3844 14504 4896 14532
rect 3844 14492 3850 14504
rect 4080 14473 4108 14504
rect 4890 14492 4896 14504
rect 4948 14532 4954 14544
rect 5442 14532 5448 14544
rect 4948 14504 5448 14532
rect 4948 14492 4954 14504
rect 5442 14492 5448 14504
rect 5500 14492 5506 14544
rect 7009 14535 7067 14541
rect 7009 14501 7021 14535
rect 7055 14532 7067 14535
rect 7190 14532 7196 14544
rect 7055 14504 7196 14532
rect 7055 14501 7067 14504
rect 7009 14495 7067 14501
rect 7190 14492 7196 14504
rect 7248 14492 7254 14544
rect 7374 14492 7380 14544
rect 7432 14532 7438 14544
rect 7561 14535 7619 14541
rect 7561 14532 7573 14535
rect 7432 14504 7573 14532
rect 7432 14492 7438 14504
rect 7561 14501 7573 14504
rect 7607 14501 7619 14535
rect 8018 14532 8024 14544
rect 7979 14504 8024 14532
rect 7561 14495 7619 14501
rect 8018 14492 8024 14504
rect 8076 14492 8082 14544
rect 10686 14541 10692 14544
rect 10680 14532 10692 14541
rect 10647 14504 10692 14532
rect 10680 14495 10692 14504
rect 10686 14492 10692 14495
rect 10744 14492 10750 14544
rect 15470 14492 15476 14544
rect 15528 14532 15534 14544
rect 15746 14532 15752 14544
rect 15528 14504 15752 14532
rect 15528 14492 15534 14504
rect 15746 14492 15752 14504
rect 15804 14532 15810 14544
rect 17218 14532 17224 14544
rect 15804 14504 17224 14532
rect 15804 14492 15810 14504
rect 17218 14492 17224 14504
rect 17276 14492 17282 14544
rect 17773 14535 17831 14541
rect 17773 14501 17785 14535
rect 17819 14532 17831 14535
rect 18138 14532 18144 14544
rect 17819 14504 18144 14532
rect 17819 14501 17831 14504
rect 17773 14495 17831 14501
rect 18138 14492 18144 14504
rect 18196 14532 18202 14544
rect 18414 14532 18420 14544
rect 18196 14504 18420 14532
rect 18196 14492 18202 14504
rect 18414 14492 18420 14504
rect 18472 14492 18478 14544
rect 21192 14532 21220 14560
rect 21358 14532 21364 14544
rect 21192 14504 21364 14532
rect 21358 14492 21364 14504
rect 21416 14532 21422 14544
rect 22833 14535 22891 14541
rect 21416 14504 21772 14532
rect 21416 14492 21422 14504
rect 4065 14467 4123 14473
rect 4065 14433 4077 14467
rect 4111 14433 4123 14467
rect 4065 14427 4123 14433
rect 4332 14467 4390 14473
rect 4332 14433 4344 14467
rect 4378 14464 4390 14467
rect 4706 14464 4712 14476
rect 4378 14436 4712 14464
rect 4378 14433 4390 14436
rect 4332 14427 4390 14433
rect 4706 14424 4712 14436
rect 4764 14424 4770 14476
rect 8110 14464 8116 14476
rect 8071 14436 8116 14464
rect 8110 14424 8116 14436
rect 8168 14424 8174 14476
rect 9306 14424 9312 14476
rect 9364 14464 9370 14476
rect 9401 14467 9459 14473
rect 9401 14464 9413 14467
rect 9364 14436 9413 14464
rect 9364 14424 9370 14436
rect 9401 14433 9413 14436
rect 9447 14464 9459 14467
rect 11698 14464 11704 14476
rect 9447 14436 11704 14464
rect 9447 14433 9459 14436
rect 9401 14427 9459 14433
rect 11698 14424 11704 14436
rect 11756 14424 11762 14476
rect 12526 14424 12532 14476
rect 12584 14464 12590 14476
rect 13265 14467 13323 14473
rect 13265 14464 13277 14467
rect 12584 14436 13277 14464
rect 12584 14424 12590 14436
rect 13265 14433 13277 14436
rect 13311 14464 13323 14467
rect 16390 14464 16396 14476
rect 13311 14436 16396 14464
rect 13311 14433 13323 14436
rect 13265 14427 13323 14433
rect 16390 14424 16396 14436
rect 16448 14424 16454 14476
rect 16761 14467 16819 14473
rect 16761 14433 16773 14467
rect 16807 14464 16819 14467
rect 16850 14464 16856 14476
rect 16807 14436 16856 14464
rect 16807 14433 16819 14436
rect 16761 14427 16819 14433
rect 16850 14424 16856 14436
rect 16908 14424 16914 14476
rect 17954 14424 17960 14476
rect 18012 14464 18018 14476
rect 18325 14467 18383 14473
rect 18325 14464 18337 14467
rect 18012 14436 18337 14464
rect 18012 14424 18018 14436
rect 18325 14433 18337 14436
rect 18371 14464 18383 14467
rect 18966 14464 18972 14476
rect 18371 14436 18972 14464
rect 18371 14433 18383 14436
rect 18325 14427 18383 14433
rect 18966 14424 18972 14436
rect 19024 14424 19030 14476
rect 19705 14467 19763 14473
rect 19705 14433 19717 14467
rect 19751 14464 19763 14467
rect 20070 14464 20076 14476
rect 19751 14436 20076 14464
rect 19751 14433 19763 14436
rect 19705 14427 19763 14433
rect 20070 14424 20076 14436
rect 20128 14424 20134 14476
rect 21634 14464 21640 14476
rect 21595 14436 21640 14464
rect 21634 14424 21640 14436
rect 21692 14424 21698 14476
rect 21744 14464 21772 14504
rect 22833 14501 22845 14535
rect 22879 14532 22891 14535
rect 23290 14532 23296 14544
rect 22879 14504 23296 14532
rect 22879 14501 22891 14504
rect 22833 14495 22891 14501
rect 23290 14492 23296 14504
rect 23348 14492 23354 14544
rect 21744 14436 21864 14464
rect 1854 14396 1860 14408
rect 1815 14368 1860 14396
rect 1854 14356 1860 14368
rect 1912 14356 1918 14408
rect 2041 14399 2099 14405
rect 2041 14365 2053 14399
rect 2087 14396 2099 14399
rect 2498 14396 2504 14408
rect 2087 14368 2504 14396
rect 2087 14365 2099 14368
rect 2041 14359 2099 14365
rect 2498 14356 2504 14368
rect 2556 14356 2562 14408
rect 2961 14399 3019 14405
rect 2961 14365 2973 14399
rect 3007 14396 3019 14399
rect 3970 14396 3976 14408
rect 3007 14368 3976 14396
rect 3007 14365 3019 14368
rect 2961 14359 3019 14365
rect 3970 14356 3976 14368
rect 4028 14356 4034 14408
rect 6270 14356 6276 14408
rect 6328 14396 6334 14408
rect 6457 14399 6515 14405
rect 6457 14396 6469 14399
rect 6328 14368 6469 14396
rect 6328 14356 6334 14368
rect 6457 14365 6469 14368
rect 6503 14396 6515 14399
rect 7193 14399 7251 14405
rect 7193 14396 7205 14399
rect 6503 14368 7205 14396
rect 6503 14365 6515 14368
rect 6457 14359 6515 14365
rect 7193 14365 7205 14368
rect 7239 14396 7251 14399
rect 8202 14396 8208 14408
rect 7239 14368 8208 14396
rect 7239 14365 7251 14368
rect 7193 14359 7251 14365
rect 8202 14356 8208 14368
rect 8260 14356 8266 14408
rect 8754 14356 8760 14408
rect 8812 14356 8818 14408
rect 9766 14356 9772 14408
rect 9824 14396 9830 14408
rect 10413 14399 10471 14405
rect 10413 14396 10425 14399
rect 9824 14368 10425 14396
rect 9824 14356 9830 14368
rect 10413 14365 10425 14368
rect 10459 14365 10471 14399
rect 10413 14359 10471 14365
rect 12434 14356 12440 14408
rect 12492 14396 12498 14408
rect 13449 14399 13507 14405
rect 12492 14368 12537 14396
rect 12492 14356 12498 14368
rect 13449 14365 13461 14399
rect 13495 14365 13507 14399
rect 15838 14396 15844 14408
rect 13449 14359 13507 14365
rect 13556 14368 15844 14396
rect 1026 14288 1032 14340
rect 1084 14328 1090 14340
rect 3789 14331 3847 14337
rect 3789 14328 3801 14331
rect 1084 14300 3801 14328
rect 1084 14288 1090 14300
rect 3789 14297 3801 14300
rect 3835 14297 3847 14331
rect 3789 14291 3847 14297
rect 5534 14288 5540 14340
rect 5592 14328 5598 14340
rect 6549 14331 6607 14337
rect 6549 14328 6561 14331
rect 5592 14300 6561 14328
rect 5592 14288 5598 14300
rect 6549 14297 6561 14300
rect 6595 14297 6607 14331
rect 6549 14291 6607 14297
rect 7006 14288 7012 14340
rect 7064 14328 7070 14340
rect 7926 14328 7932 14340
rect 7064 14300 7932 14328
rect 7064 14288 7070 14300
rect 7926 14288 7932 14300
rect 7984 14288 7990 14340
rect 8018 14288 8024 14340
rect 8076 14328 8082 14340
rect 8772 14328 8800 14356
rect 12802 14328 12808 14340
rect 8076 14300 8800 14328
rect 12715 14300 12808 14328
rect 8076 14288 8082 14300
rect 12802 14288 12808 14300
rect 12860 14328 12866 14340
rect 13464 14328 13492 14359
rect 13556 14340 13584 14368
rect 15838 14356 15844 14368
rect 15896 14356 15902 14408
rect 16209 14399 16267 14405
rect 16209 14365 16221 14399
rect 16255 14396 16267 14399
rect 17037 14399 17095 14405
rect 16255 14368 16712 14396
rect 16255 14365 16267 14368
rect 16209 14359 16267 14365
rect 16684 14340 16712 14368
rect 17037 14365 17049 14399
rect 17083 14365 17095 14399
rect 17037 14359 17095 14365
rect 12860 14300 13492 14328
rect 12860 14288 12866 14300
rect 13538 14288 13544 14340
rect 13596 14288 13602 14340
rect 15470 14288 15476 14340
rect 15528 14328 15534 14340
rect 16393 14331 16451 14337
rect 16393 14328 16405 14331
rect 15528 14300 16405 14328
rect 15528 14288 15534 14300
rect 16393 14297 16405 14300
rect 16439 14297 16451 14331
rect 16393 14291 16451 14297
rect 16666 14288 16672 14340
rect 16724 14328 16730 14340
rect 17052 14328 17080 14359
rect 17218 14356 17224 14408
rect 17276 14396 17282 14408
rect 18417 14399 18475 14405
rect 18417 14396 18429 14399
rect 17276 14368 18429 14396
rect 17276 14356 17282 14368
rect 18417 14365 18429 14368
rect 18463 14365 18475 14399
rect 18598 14396 18604 14408
rect 18559 14368 18604 14396
rect 18417 14359 18475 14365
rect 18598 14356 18604 14368
rect 18656 14356 18662 14408
rect 21836 14405 21864 14436
rect 21821 14399 21879 14405
rect 21821 14365 21833 14399
rect 21867 14396 21879 14399
rect 22278 14396 22284 14408
rect 21867 14368 22284 14396
rect 21867 14365 21879 14368
rect 21821 14359 21879 14365
rect 22278 14356 22284 14368
rect 22336 14356 22342 14408
rect 18616 14328 18644 14356
rect 16724 14300 18644 14328
rect 21269 14331 21327 14337
rect 16724 14288 16730 14300
rect 21269 14297 21281 14331
rect 21315 14328 21327 14331
rect 23400 14328 23428 14563
rect 24026 14560 24032 14572
rect 24084 14560 24090 14612
rect 24578 14560 24584 14612
rect 24636 14600 24642 14612
rect 25869 14603 25927 14609
rect 25869 14600 25881 14603
rect 24636 14572 25881 14600
rect 24636 14560 24642 14572
rect 25869 14569 25881 14572
rect 25915 14600 25927 14603
rect 26142 14600 26148 14612
rect 25915 14572 26148 14600
rect 25915 14569 25927 14572
rect 25869 14563 25927 14569
rect 26142 14560 26148 14572
rect 26200 14560 26206 14612
rect 26237 14603 26295 14609
rect 26237 14569 26249 14603
rect 26283 14600 26295 14603
rect 26326 14600 26332 14612
rect 26283 14572 26332 14600
rect 26283 14569 26295 14572
rect 26237 14563 26295 14569
rect 23566 14492 23572 14544
rect 23624 14532 23630 14544
rect 24118 14541 24124 14544
rect 23661 14535 23719 14541
rect 23661 14532 23673 14535
rect 23624 14504 23673 14532
rect 23624 14492 23630 14504
rect 23661 14501 23673 14504
rect 23707 14501 23719 14535
rect 24112 14532 24124 14541
rect 24079 14504 24124 14532
rect 23661 14495 23719 14501
rect 24112 14495 24124 14504
rect 24176 14532 24182 14544
rect 24854 14532 24860 14544
rect 24176 14504 24860 14532
rect 24118 14492 24124 14495
rect 24176 14492 24182 14504
rect 24854 14492 24860 14504
rect 24912 14492 24918 14544
rect 26252 14464 26280 14563
rect 26326 14560 26332 14572
rect 26384 14560 26390 14612
rect 23860 14436 26280 14464
rect 23860 14408 23888 14436
rect 23842 14396 23848 14408
rect 23755 14368 23848 14396
rect 23842 14356 23848 14368
rect 23900 14356 23906 14408
rect 21315 14300 23428 14328
rect 21315 14297 21327 14300
rect 21269 14291 21327 14297
rect 2869 14263 2927 14269
rect 2869 14229 2881 14263
rect 2915 14260 2927 14263
rect 2958 14260 2964 14272
rect 2915 14232 2964 14260
rect 2915 14229 2927 14232
rect 2869 14223 2927 14229
rect 2958 14220 2964 14232
rect 3016 14220 3022 14272
rect 5350 14220 5356 14272
rect 5408 14260 5414 14272
rect 5445 14263 5503 14269
rect 5445 14260 5457 14263
rect 5408 14232 5457 14260
rect 5408 14220 5414 14232
rect 5445 14229 5457 14232
rect 5491 14260 5503 14263
rect 6362 14260 6368 14272
rect 5491 14232 6368 14260
rect 5491 14229 5503 14232
rect 5445 14223 5503 14229
rect 6362 14220 6368 14232
rect 6420 14220 6426 14272
rect 7834 14220 7840 14272
rect 7892 14260 7898 14272
rect 8297 14263 8355 14269
rect 8297 14260 8309 14263
rect 7892 14232 8309 14260
rect 7892 14220 7898 14232
rect 8297 14229 8309 14232
rect 8343 14229 8355 14263
rect 8754 14260 8760 14272
rect 8715 14232 8760 14260
rect 8297 14223 8355 14229
rect 8754 14220 8760 14232
rect 8812 14220 8818 14272
rect 9766 14220 9772 14272
rect 9824 14260 9830 14272
rect 9950 14260 9956 14272
rect 9824 14232 9956 14260
rect 9824 14220 9830 14232
rect 9950 14220 9956 14232
rect 10008 14220 10014 14272
rect 12894 14260 12900 14272
rect 12855 14232 12900 14260
rect 12894 14220 12900 14232
rect 12952 14220 12958 14272
rect 13998 14260 14004 14272
rect 13959 14232 14004 14260
rect 13998 14220 14004 14232
rect 14056 14220 14062 14272
rect 14090 14220 14096 14272
rect 14148 14260 14154 14272
rect 14277 14263 14335 14269
rect 14277 14260 14289 14263
rect 14148 14232 14289 14260
rect 14148 14220 14154 14232
rect 14277 14229 14289 14232
rect 14323 14260 14335 14263
rect 14642 14260 14648 14272
rect 14323 14232 14648 14260
rect 14323 14229 14335 14232
rect 14277 14223 14335 14229
rect 14642 14220 14648 14232
rect 14700 14220 14706 14272
rect 15105 14263 15163 14269
rect 15105 14229 15117 14263
rect 15151 14260 15163 14263
rect 15286 14260 15292 14272
rect 15151 14232 15292 14260
rect 15151 14229 15163 14232
rect 15105 14223 15163 14229
rect 15286 14220 15292 14232
rect 15344 14220 15350 14272
rect 21177 14263 21235 14269
rect 21177 14229 21189 14263
rect 21223 14260 21235 14263
rect 21542 14260 21548 14272
rect 21223 14232 21548 14260
rect 21223 14229 21235 14232
rect 21177 14223 21235 14229
rect 21542 14220 21548 14232
rect 21600 14220 21606 14272
rect 25222 14260 25228 14272
rect 25183 14232 25228 14260
rect 25222 14220 25228 14232
rect 25280 14220 25286 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 2498 14016 2504 14068
rect 2556 14056 2562 14068
rect 2961 14059 3019 14065
rect 2961 14056 2973 14059
rect 2556 14028 2973 14056
rect 2556 14016 2562 14028
rect 2961 14025 2973 14028
rect 3007 14025 3019 14059
rect 2961 14019 3019 14025
rect 3142 14016 3148 14068
rect 3200 14056 3206 14068
rect 3513 14059 3571 14065
rect 3513 14056 3525 14059
rect 3200 14028 3525 14056
rect 3200 14016 3206 14028
rect 3513 14025 3525 14028
rect 3559 14025 3571 14059
rect 4246 14056 4252 14068
rect 4207 14028 4252 14056
rect 3513 14019 3571 14025
rect 4246 14016 4252 14028
rect 4304 14016 4310 14068
rect 5166 14056 5172 14068
rect 5127 14028 5172 14056
rect 5166 14016 5172 14028
rect 5224 14016 5230 14068
rect 8478 14056 8484 14068
rect 8439 14028 8484 14056
rect 8478 14016 8484 14028
rect 8536 14016 8542 14068
rect 10042 14056 10048 14068
rect 10003 14028 10048 14056
rect 10042 14016 10048 14028
rect 10100 14016 10106 14068
rect 10686 14016 10692 14068
rect 10744 14056 10750 14068
rect 11057 14059 11115 14065
rect 11057 14056 11069 14059
rect 10744 14028 11069 14056
rect 10744 14016 10750 14028
rect 11057 14025 11069 14028
rect 11103 14056 11115 14059
rect 11790 14056 11796 14068
rect 11103 14028 11796 14056
rect 11103 14025 11115 14028
rect 11057 14019 11115 14025
rect 11790 14016 11796 14028
rect 11848 14016 11854 14068
rect 12989 14059 13047 14065
rect 12989 14025 13001 14059
rect 13035 14056 13047 14059
rect 13262 14056 13268 14068
rect 13035 14028 13268 14056
rect 13035 14025 13047 14028
rect 12989 14019 13047 14025
rect 13262 14016 13268 14028
rect 13320 14016 13326 14068
rect 13722 14016 13728 14068
rect 13780 14056 13786 14068
rect 14366 14056 14372 14068
rect 13780 14028 14372 14056
rect 13780 14016 13786 14028
rect 14366 14016 14372 14028
rect 14424 14056 14430 14068
rect 14461 14059 14519 14065
rect 14461 14056 14473 14059
rect 14424 14028 14473 14056
rect 14424 14016 14430 14028
rect 14461 14025 14473 14028
rect 14507 14025 14519 14059
rect 14461 14019 14519 14025
rect 15197 14059 15255 14065
rect 15197 14025 15209 14059
rect 15243 14056 15255 14059
rect 16850 14056 16856 14068
rect 15243 14028 16856 14056
rect 15243 14025 15255 14028
rect 15197 14019 15255 14025
rect 16850 14016 16856 14028
rect 16908 14016 16914 14068
rect 17218 14016 17224 14068
rect 17276 14056 17282 14068
rect 17405 14059 17463 14065
rect 17405 14056 17417 14059
rect 17276 14028 17417 14056
rect 17276 14016 17282 14028
rect 17405 14025 17417 14028
rect 17451 14025 17463 14059
rect 17405 14019 17463 14025
rect 18046 14016 18052 14068
rect 18104 14056 18110 14068
rect 18230 14056 18236 14068
rect 18104 14028 18236 14056
rect 18104 14016 18110 14028
rect 18230 14016 18236 14028
rect 18288 14016 18294 14068
rect 20806 14056 20812 14068
rect 20767 14028 20812 14056
rect 20806 14016 20812 14028
rect 20864 14016 20870 14068
rect 22649 14059 22707 14065
rect 22649 14025 22661 14059
rect 22695 14056 22707 14059
rect 23106 14056 23112 14068
rect 22695 14028 23112 14056
rect 22695 14025 22707 14028
rect 22649 14019 22707 14025
rect 23106 14016 23112 14028
rect 23164 14016 23170 14068
rect 23477 14059 23535 14065
rect 23477 14025 23489 14059
rect 23523 14056 23535 14059
rect 24854 14056 24860 14068
rect 23523 14028 24860 14056
rect 23523 14025 23535 14028
rect 23477 14019 23535 14025
rect 24854 14016 24860 14028
rect 24912 14056 24918 14068
rect 25041 14059 25099 14065
rect 25041 14056 25053 14059
rect 24912 14028 25053 14056
rect 24912 14016 24918 14028
rect 25041 14025 25053 14028
rect 25087 14025 25099 14059
rect 25682 14056 25688 14068
rect 25643 14028 25688 14056
rect 25041 14019 25099 14025
rect 25682 14016 25688 14028
rect 25740 14016 25746 14068
rect 26053 14059 26111 14065
rect 26053 14025 26065 14059
rect 26099 14056 26111 14059
rect 26326 14056 26332 14068
rect 26099 14028 26332 14056
rect 26099 14025 26111 14028
rect 26053 14019 26111 14025
rect 26326 14016 26332 14028
rect 26384 14016 26390 14068
rect 2682 13948 2688 14000
rect 2740 13988 2746 14000
rect 3160 13988 3188 14016
rect 4706 13988 4712 14000
rect 2740 13960 3188 13988
rect 4667 13960 4712 13988
rect 2740 13948 2746 13960
rect 4706 13948 4712 13960
rect 4764 13948 4770 14000
rect 6822 13988 6828 14000
rect 5644 13960 6828 13988
rect 1578 13920 1584 13932
rect 1539 13892 1584 13920
rect 1578 13880 1584 13892
rect 1636 13880 1642 13932
rect 2774 13880 2780 13932
rect 2832 13920 2838 13932
rect 5644 13929 5672 13960
rect 6822 13948 6828 13960
rect 6880 13948 6886 14000
rect 6914 13948 6920 14000
rect 6972 13988 6978 14000
rect 8294 13988 8300 14000
rect 6972 13960 8300 13988
rect 6972 13948 6978 13960
rect 8294 13948 8300 13960
rect 8352 13948 8358 14000
rect 8389 13991 8447 13997
rect 8389 13957 8401 13991
rect 8435 13988 8447 13991
rect 9582 13988 9588 14000
rect 8435 13960 9588 13988
rect 8435 13957 8447 13960
rect 8389 13951 8447 13957
rect 5629 13923 5687 13929
rect 2832 13892 4752 13920
rect 2832 13880 2838 13892
rect 4724 13864 4752 13892
rect 5629 13889 5641 13923
rect 5675 13889 5687 13923
rect 5629 13883 5687 13889
rect 5813 13923 5871 13929
rect 5813 13889 5825 13923
rect 5859 13920 5871 13923
rect 6270 13920 6276 13932
rect 5859 13892 6276 13920
rect 5859 13889 5871 13892
rect 5813 13883 5871 13889
rect 1848 13855 1906 13861
rect 1848 13821 1860 13855
rect 1894 13852 1906 13855
rect 2314 13852 2320 13864
rect 1894 13824 2320 13852
rect 1894 13821 1906 13824
rect 1848 13815 1906 13821
rect 2314 13812 2320 13824
rect 2372 13852 2378 13864
rect 2958 13852 2964 13864
rect 2372 13824 2964 13852
rect 2372 13812 2378 13824
rect 2958 13812 2964 13824
rect 3016 13812 3022 13864
rect 4065 13855 4123 13861
rect 4065 13852 4077 13855
rect 3896 13824 4077 13852
rect 2498 13744 2504 13796
rect 2556 13784 2562 13796
rect 3896 13793 3924 13824
rect 4065 13821 4077 13824
rect 4111 13821 4123 13855
rect 4065 13815 4123 13821
rect 4706 13812 4712 13864
rect 4764 13812 4770 13864
rect 5077 13855 5135 13861
rect 5077 13821 5089 13855
rect 5123 13852 5135 13855
rect 5828 13852 5856 13883
rect 6270 13880 6276 13892
rect 6328 13880 6334 13932
rect 6641 13923 6699 13929
rect 6641 13889 6653 13923
rect 6687 13920 6699 13923
rect 7282 13920 7288 13932
rect 6687 13892 7288 13920
rect 6687 13889 6699 13892
rect 6641 13883 6699 13889
rect 7282 13880 7288 13892
rect 7340 13880 7346 13932
rect 7377 13923 7435 13929
rect 7377 13889 7389 13923
rect 7423 13920 7435 13923
rect 7837 13923 7895 13929
rect 7837 13920 7849 13923
rect 7423 13892 7849 13920
rect 7423 13889 7435 13892
rect 7377 13883 7435 13889
rect 7837 13889 7849 13892
rect 7883 13889 7895 13923
rect 8938 13920 8944 13932
rect 8899 13892 8944 13920
rect 7837 13883 7895 13889
rect 5123 13824 5856 13852
rect 5123 13821 5135 13824
rect 5077 13815 5135 13821
rect 5902 13812 5908 13864
rect 5960 13852 5966 13864
rect 6181 13855 6239 13861
rect 6181 13852 6193 13855
rect 5960 13824 6193 13852
rect 5960 13812 5966 13824
rect 3881 13787 3939 13793
rect 3881 13784 3893 13787
rect 2556 13756 3893 13784
rect 2556 13744 2562 13756
rect 3881 13753 3893 13756
rect 3927 13753 3939 13787
rect 3881 13747 3939 13753
rect 2774 13676 2780 13728
rect 2832 13716 2838 13728
rect 3234 13716 3240 13728
rect 2832 13688 3240 13716
rect 2832 13676 2838 13688
rect 3234 13676 3240 13688
rect 3292 13676 3298 13728
rect 5534 13716 5540 13728
rect 5495 13688 5540 13716
rect 5534 13676 5540 13688
rect 5592 13676 5598 13728
rect 6012 13716 6040 13824
rect 6181 13821 6193 13824
rect 6227 13821 6239 13855
rect 6181 13815 6239 13821
rect 6362 13812 6368 13864
rect 6420 13852 6426 13864
rect 7392 13852 7420 13883
rect 8938 13880 8944 13892
rect 8996 13880 9002 13932
rect 9140 13929 9168 13960
rect 9582 13948 9588 13960
rect 9640 13988 9646 14000
rect 9950 13988 9956 14000
rect 9640 13960 9956 13988
rect 9640 13948 9646 13960
rect 9950 13948 9956 13960
rect 10008 13988 10014 14000
rect 10008 13960 10640 13988
rect 10008 13948 10014 13960
rect 10612 13929 10640 13960
rect 15378 13948 15384 14000
rect 15436 13948 15442 14000
rect 15838 13948 15844 14000
rect 15896 13988 15902 14000
rect 16117 13991 16175 13997
rect 16117 13988 16129 13991
rect 15896 13960 16129 13988
rect 15896 13948 15902 13960
rect 16117 13957 16129 13960
rect 16163 13988 16175 13991
rect 16209 13991 16267 13997
rect 16209 13988 16221 13991
rect 16163 13960 16221 13988
rect 16163 13957 16175 13960
rect 16117 13951 16175 13957
rect 16209 13957 16221 13960
rect 16255 13957 16267 13991
rect 17954 13988 17960 14000
rect 16209 13951 16267 13957
rect 17604 13960 17960 13988
rect 9125 13923 9183 13929
rect 9125 13889 9137 13923
rect 9171 13889 9183 13923
rect 9125 13883 9183 13889
rect 10597 13923 10655 13929
rect 10597 13889 10609 13923
rect 10643 13889 10655 13923
rect 10597 13883 10655 13889
rect 11698 13880 11704 13932
rect 11756 13920 11762 13932
rect 11793 13923 11851 13929
rect 11793 13920 11805 13923
rect 11756 13892 11805 13920
rect 11756 13880 11762 13892
rect 11793 13889 11805 13892
rect 11839 13920 11851 13923
rect 12250 13920 12256 13932
rect 11839 13892 12256 13920
rect 11839 13889 11851 13892
rect 11793 13883 11851 13889
rect 12250 13880 12256 13892
rect 12308 13880 12314 13932
rect 15396 13920 15424 13948
rect 15304 13892 15424 13920
rect 15565 13923 15623 13929
rect 6420 13824 7420 13852
rect 9585 13855 9643 13861
rect 6420 13812 6426 13824
rect 9585 13821 9597 13855
rect 9631 13852 9643 13855
rect 10505 13855 10563 13861
rect 10505 13852 10517 13855
rect 9631 13824 10517 13852
rect 9631 13821 9643 13824
rect 9585 13815 9643 13821
rect 10505 13821 10517 13824
rect 10551 13852 10563 13855
rect 10962 13852 10968 13864
rect 10551 13824 10968 13852
rect 10551 13821 10563 13824
rect 10505 13815 10563 13821
rect 10962 13812 10968 13824
rect 11020 13812 11026 13864
rect 11422 13852 11428 13864
rect 11383 13824 11428 13852
rect 11422 13812 11428 13824
rect 11480 13812 11486 13864
rect 13081 13855 13139 13861
rect 13081 13821 13093 13855
rect 13127 13852 13139 13855
rect 13348 13855 13406 13861
rect 13127 13824 13308 13852
rect 13127 13821 13139 13824
rect 13081 13815 13139 13821
rect 6086 13744 6092 13796
rect 6144 13784 6150 13796
rect 6270 13784 6276 13796
rect 6144 13756 6276 13784
rect 6144 13744 6150 13756
rect 6270 13744 6276 13756
rect 6328 13744 6334 13796
rect 9398 13744 9404 13796
rect 9456 13784 9462 13796
rect 12161 13787 12219 13793
rect 12161 13784 12173 13787
rect 9456 13756 12173 13784
rect 9456 13744 9462 13756
rect 12161 13753 12173 13756
rect 12207 13784 12219 13787
rect 12526 13784 12532 13796
rect 12207 13756 12532 13784
rect 12207 13753 12219 13756
rect 12161 13747 12219 13753
rect 12526 13744 12532 13756
rect 12584 13744 12590 13796
rect 13280 13784 13308 13824
rect 13348 13821 13360 13855
rect 13394 13852 13406 13855
rect 13394 13824 14044 13852
rect 13394 13821 13406 13824
rect 13348 13815 13406 13821
rect 14016 13796 14044 13824
rect 13906 13784 13912 13796
rect 13280 13756 13912 13784
rect 13906 13744 13912 13756
rect 13964 13744 13970 13796
rect 13998 13744 14004 13796
rect 14056 13744 14062 13796
rect 7193 13719 7251 13725
rect 7193 13716 7205 13719
rect 6012 13688 7205 13716
rect 7193 13685 7205 13688
rect 7239 13685 7251 13719
rect 7193 13679 7251 13685
rect 8754 13676 8760 13728
rect 8812 13716 8818 13728
rect 8849 13719 8907 13725
rect 8849 13716 8861 13719
rect 8812 13688 8861 13716
rect 8812 13676 8818 13688
rect 8849 13685 8861 13688
rect 8895 13716 8907 13719
rect 9674 13716 9680 13728
rect 8895 13688 9680 13716
rect 8895 13685 8907 13688
rect 8849 13679 8907 13685
rect 9674 13676 9680 13688
rect 9732 13676 9738 13728
rect 9953 13719 10011 13725
rect 9953 13685 9965 13719
rect 9999 13716 10011 13719
rect 10413 13719 10471 13725
rect 10413 13716 10425 13719
rect 9999 13688 10425 13716
rect 9999 13685 10011 13688
rect 9953 13679 10011 13685
rect 10413 13685 10425 13688
rect 10459 13716 10471 13719
rect 10686 13716 10692 13728
rect 10459 13688 10692 13716
rect 10459 13685 10471 13688
rect 10413 13679 10471 13685
rect 10686 13676 10692 13688
rect 10744 13716 10750 13728
rect 14182 13716 14188 13728
rect 10744 13688 14188 13716
rect 10744 13676 10750 13688
rect 14182 13676 14188 13688
rect 14240 13676 14246 13728
rect 15304 13716 15332 13892
rect 15565 13889 15577 13923
rect 15611 13920 15623 13923
rect 15933 13923 15991 13929
rect 15933 13920 15945 13923
rect 15611 13892 15945 13920
rect 15611 13889 15623 13892
rect 15565 13883 15623 13889
rect 15933 13889 15945 13892
rect 15979 13920 15991 13923
rect 16666 13920 16672 13932
rect 15979 13892 16672 13920
rect 15979 13889 15991 13892
rect 15933 13883 15991 13889
rect 16666 13880 16672 13892
rect 16724 13920 16730 13932
rect 16945 13923 17003 13929
rect 16945 13920 16957 13923
rect 16724 13892 16957 13920
rect 16724 13880 16730 13892
rect 16945 13889 16957 13892
rect 16991 13889 17003 13923
rect 16945 13883 17003 13889
rect 16850 13852 16856 13864
rect 16811 13824 16856 13852
rect 16850 13812 16856 13824
rect 16908 13812 16914 13864
rect 17218 13812 17224 13864
rect 17276 13852 17282 13864
rect 17604 13852 17632 13960
rect 17954 13948 17960 13960
rect 18012 13948 18018 14000
rect 20349 13991 20407 13997
rect 20349 13957 20361 13991
rect 20395 13988 20407 13991
rect 22278 13988 22284 14000
rect 20395 13960 21496 13988
rect 22239 13960 22284 13988
rect 20395 13957 20407 13960
rect 20349 13951 20407 13957
rect 17678 13880 17684 13932
rect 17736 13920 17742 13932
rect 20714 13920 20720 13932
rect 17736 13892 18184 13920
rect 20675 13892 20720 13920
rect 17736 13880 17742 13892
rect 18156 13864 18184 13892
rect 20714 13880 20720 13892
rect 20772 13920 20778 13932
rect 21358 13920 21364 13932
rect 20772 13892 21220 13920
rect 21319 13892 21364 13920
rect 20772 13880 20778 13892
rect 17773 13855 17831 13861
rect 17773 13852 17785 13855
rect 17276 13824 17785 13852
rect 17276 13812 17282 13824
rect 17773 13821 17785 13824
rect 17819 13821 17831 13855
rect 18046 13852 18052 13864
rect 18007 13824 18052 13852
rect 17773 13815 17831 13821
rect 18046 13812 18052 13824
rect 18104 13812 18110 13864
rect 18138 13812 18144 13864
rect 18196 13852 18202 13864
rect 21192 13861 21220 13892
rect 21358 13880 21364 13892
rect 21416 13880 21422 13932
rect 18305 13855 18363 13861
rect 18305 13852 18317 13855
rect 18196 13824 18317 13852
rect 18196 13812 18202 13824
rect 18305 13821 18317 13824
rect 18351 13821 18363 13855
rect 18305 13815 18363 13821
rect 21177 13855 21235 13861
rect 21177 13821 21189 13855
rect 21223 13821 21235 13855
rect 21177 13815 21235 13821
rect 21269 13855 21327 13861
rect 21269 13821 21281 13855
rect 21315 13852 21327 13855
rect 21468 13852 21496 13960
rect 22278 13948 22284 13960
rect 22336 13948 22342 14000
rect 25700 13920 25728 14016
rect 26234 13920 26240 13932
rect 25700 13892 26240 13920
rect 26234 13880 26240 13892
rect 26292 13880 26298 13932
rect 21726 13852 21732 13864
rect 21315 13824 21732 13852
rect 21315 13821 21327 13824
rect 21269 13815 21327 13821
rect 21726 13812 21732 13824
rect 21784 13812 21790 13864
rect 21910 13852 21916 13864
rect 21871 13824 21916 13852
rect 21910 13812 21916 13824
rect 21968 13812 21974 13864
rect 22094 13812 22100 13864
rect 22152 13852 22158 13864
rect 23934 13861 23940 13864
rect 22465 13855 22523 13861
rect 22465 13852 22477 13855
rect 22152 13824 22477 13852
rect 22152 13812 22158 13824
rect 22465 13821 22477 13824
rect 22511 13852 22523 13855
rect 23661 13855 23719 13861
rect 22511 13824 23152 13852
rect 22511 13821 22523 13824
rect 22465 13815 22523 13821
rect 16117 13787 16175 13793
rect 16117 13753 16129 13787
rect 16163 13784 16175 13787
rect 16163 13756 16528 13784
rect 16163 13753 16175 13756
rect 16117 13747 16175 13753
rect 15838 13716 15844 13728
rect 15304 13688 15844 13716
rect 15838 13676 15844 13688
rect 15896 13676 15902 13728
rect 16390 13716 16396 13728
rect 16351 13688 16396 13716
rect 16390 13676 16396 13688
rect 16448 13676 16454 13728
rect 16500 13716 16528 13756
rect 16761 13719 16819 13725
rect 16761 13716 16773 13719
rect 16500 13688 16773 13716
rect 16761 13685 16773 13688
rect 16807 13685 16819 13719
rect 16761 13679 16819 13685
rect 18414 13676 18420 13728
rect 18472 13716 18478 13728
rect 23124 13725 23152 13824
rect 23661 13821 23673 13855
rect 23707 13821 23719 13855
rect 23928 13852 23940 13861
rect 23895 13824 23940 13852
rect 23661 13815 23719 13821
rect 23928 13815 23940 13824
rect 23566 13744 23572 13796
rect 23624 13784 23630 13796
rect 23676 13784 23704 13815
rect 23934 13812 23940 13815
rect 23992 13812 23998 13864
rect 23842 13784 23848 13796
rect 23624 13756 23848 13784
rect 23624 13744 23630 13756
rect 23842 13744 23848 13756
rect 23900 13744 23906 13796
rect 19429 13719 19487 13725
rect 19429 13716 19441 13719
rect 18472 13688 19441 13716
rect 18472 13676 18478 13688
rect 19429 13685 19441 13688
rect 19475 13685 19487 13719
rect 19429 13679 19487 13685
rect 23109 13719 23167 13725
rect 23109 13685 23121 13719
rect 23155 13716 23167 13719
rect 23750 13716 23756 13728
rect 23155 13688 23756 13716
rect 23155 13685 23167 13688
rect 23109 13679 23167 13685
rect 23750 13676 23756 13688
rect 23808 13676 23814 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 4709 13515 4767 13521
rect 4709 13481 4721 13515
rect 4755 13512 4767 13515
rect 5534 13512 5540 13524
rect 4755 13484 5540 13512
rect 4755 13481 4767 13484
rect 4709 13475 4767 13481
rect 5534 13472 5540 13484
rect 5592 13472 5598 13524
rect 5718 13512 5724 13524
rect 5679 13484 5724 13512
rect 5718 13472 5724 13484
rect 5776 13472 5782 13524
rect 6181 13515 6239 13521
rect 6181 13481 6193 13515
rect 6227 13512 6239 13515
rect 7190 13512 7196 13524
rect 6227 13484 7196 13512
rect 6227 13481 6239 13484
rect 6181 13475 6239 13481
rect 7190 13472 7196 13484
rect 7248 13472 7254 13524
rect 7466 13472 7472 13524
rect 7524 13512 7530 13524
rect 7653 13515 7711 13521
rect 7653 13512 7665 13515
rect 7524 13484 7665 13512
rect 7524 13472 7530 13484
rect 7653 13481 7665 13484
rect 7699 13481 7711 13515
rect 7653 13475 7711 13481
rect 8573 13515 8631 13521
rect 8573 13481 8585 13515
rect 8619 13512 8631 13515
rect 8938 13512 8944 13524
rect 8619 13484 8944 13512
rect 8619 13481 8631 13484
rect 8573 13475 8631 13481
rect 8938 13472 8944 13484
rect 8996 13472 9002 13524
rect 9214 13512 9220 13524
rect 9175 13484 9220 13512
rect 9214 13472 9220 13484
rect 9272 13472 9278 13524
rect 10962 13472 10968 13524
rect 11020 13512 11026 13524
rect 12161 13515 12219 13521
rect 12161 13512 12173 13515
rect 11020 13484 12173 13512
rect 11020 13472 11026 13484
rect 12161 13481 12173 13484
rect 12207 13481 12219 13515
rect 12161 13475 12219 13481
rect 12526 13472 12532 13524
rect 12584 13512 12590 13524
rect 12621 13515 12679 13521
rect 12621 13512 12633 13515
rect 12584 13484 12633 13512
rect 12584 13472 12590 13484
rect 12621 13481 12633 13484
rect 12667 13481 12679 13515
rect 12621 13475 12679 13481
rect 13262 13472 13268 13524
rect 13320 13512 13326 13524
rect 13357 13515 13415 13521
rect 13357 13512 13369 13515
rect 13320 13484 13369 13512
rect 13320 13472 13326 13484
rect 13357 13481 13369 13484
rect 13403 13512 13415 13515
rect 16022 13512 16028 13524
rect 13403 13484 16028 13512
rect 13403 13481 13415 13484
rect 13357 13475 13415 13481
rect 16022 13472 16028 13484
rect 16080 13472 16086 13524
rect 17313 13515 17371 13521
rect 17313 13481 17325 13515
rect 17359 13512 17371 13515
rect 17494 13512 17500 13524
rect 17359 13484 17500 13512
rect 17359 13481 17371 13484
rect 17313 13475 17371 13481
rect 17494 13472 17500 13484
rect 17552 13472 17558 13524
rect 17586 13472 17592 13524
rect 17644 13512 17650 13524
rect 17773 13515 17831 13521
rect 17773 13512 17785 13515
rect 17644 13484 17785 13512
rect 17644 13472 17650 13484
rect 17773 13481 17785 13484
rect 17819 13481 17831 13515
rect 17773 13475 17831 13481
rect 17954 13472 17960 13524
rect 18012 13512 18018 13524
rect 18141 13515 18199 13521
rect 18141 13512 18153 13515
rect 18012 13484 18153 13512
rect 18012 13472 18018 13484
rect 18141 13481 18153 13484
rect 18187 13512 18199 13515
rect 19521 13515 19579 13521
rect 19521 13512 19533 13515
rect 18187 13484 19533 13512
rect 18187 13481 18199 13484
rect 18141 13475 18199 13481
rect 19521 13481 19533 13484
rect 19567 13481 19579 13515
rect 19521 13475 19579 13481
rect 19889 13515 19947 13521
rect 19889 13481 19901 13515
rect 19935 13512 19947 13515
rect 20346 13512 20352 13524
rect 19935 13484 20352 13512
rect 19935 13481 19947 13484
rect 19889 13475 19947 13481
rect 20346 13472 20352 13484
rect 20404 13472 20410 13524
rect 21082 13472 21088 13524
rect 21140 13512 21146 13524
rect 21177 13515 21235 13521
rect 21177 13512 21189 13515
rect 21140 13484 21189 13512
rect 21140 13472 21146 13484
rect 21177 13481 21189 13484
rect 21223 13481 21235 13515
rect 21634 13512 21640 13524
rect 21595 13484 21640 13512
rect 21177 13475 21235 13481
rect 21634 13472 21640 13484
rect 21692 13472 21698 13524
rect 23477 13515 23535 13521
rect 23477 13481 23489 13515
rect 23523 13512 23535 13515
rect 23934 13512 23940 13524
rect 23523 13484 23940 13512
rect 23523 13481 23535 13484
rect 23477 13475 23535 13481
rect 23934 13472 23940 13484
rect 23992 13512 23998 13524
rect 24029 13515 24087 13521
rect 24029 13512 24041 13515
rect 23992 13484 24041 13512
rect 23992 13472 23998 13484
rect 24029 13481 24041 13484
rect 24075 13481 24087 13515
rect 24029 13475 24087 13481
rect 24949 13515 25007 13521
rect 24949 13481 24961 13515
rect 24995 13512 25007 13515
rect 25038 13512 25044 13524
rect 24995 13484 25044 13512
rect 24995 13481 25007 13484
rect 24949 13475 25007 13481
rect 25038 13472 25044 13484
rect 25096 13472 25102 13524
rect 26053 13515 26111 13521
rect 26053 13481 26065 13515
rect 26099 13512 26111 13515
rect 26326 13512 26332 13524
rect 26099 13484 26332 13512
rect 26099 13481 26111 13484
rect 26053 13475 26111 13481
rect 26326 13472 26332 13484
rect 26384 13472 26390 13524
rect 2038 13444 2044 13456
rect 1688 13416 2044 13444
rect 1688 13388 1716 13416
rect 2038 13404 2044 13416
rect 2096 13404 2102 13456
rect 3970 13404 3976 13456
rect 4028 13444 4034 13456
rect 5077 13447 5135 13453
rect 5077 13444 5089 13447
rect 4028 13416 5089 13444
rect 4028 13404 4034 13416
rect 5077 13413 5089 13416
rect 5123 13413 5135 13447
rect 5077 13407 5135 13413
rect 6540 13447 6598 13453
rect 6540 13413 6552 13447
rect 6586 13444 6598 13447
rect 6730 13444 6736 13456
rect 6586 13416 6736 13444
rect 6586 13413 6598 13416
rect 6540 13407 6598 13413
rect 6730 13404 6736 13416
rect 6788 13404 6794 13456
rect 8294 13404 8300 13456
rect 8352 13444 8358 13456
rect 9950 13453 9956 13456
rect 8849 13447 8907 13453
rect 8849 13444 8861 13447
rect 8352 13416 8861 13444
rect 8352 13404 8358 13416
rect 8849 13413 8861 13416
rect 8895 13413 8907 13447
rect 9944 13444 9956 13453
rect 9911 13416 9956 13444
rect 8849 13407 8907 13413
rect 9944 13407 9956 13416
rect 9950 13404 9956 13407
rect 10008 13404 10014 13456
rect 10594 13404 10600 13456
rect 10652 13444 10658 13456
rect 10778 13444 10784 13456
rect 10652 13416 10784 13444
rect 10652 13404 10658 13416
rect 10778 13404 10784 13416
rect 10836 13404 10842 13456
rect 11790 13404 11796 13456
rect 11848 13444 11854 13456
rect 11977 13447 12035 13453
rect 11977 13444 11989 13447
rect 11848 13416 11989 13444
rect 11848 13404 11854 13416
rect 11977 13413 11989 13416
rect 12023 13413 12035 13447
rect 11977 13407 12035 13413
rect 13538 13404 13544 13456
rect 13596 13444 13602 13456
rect 13633 13447 13691 13453
rect 13633 13444 13645 13447
rect 13596 13416 13645 13444
rect 13596 13404 13602 13416
rect 13633 13413 13645 13416
rect 13679 13413 13691 13447
rect 13633 13407 13691 13413
rect 13814 13404 13820 13456
rect 13872 13444 13878 13456
rect 14458 13444 14464 13456
rect 13872 13416 14464 13444
rect 13872 13404 13878 13416
rect 14458 13404 14464 13416
rect 14516 13404 14522 13456
rect 14921 13447 14979 13453
rect 14921 13413 14933 13447
rect 14967 13444 14979 13447
rect 15378 13444 15384 13456
rect 14967 13416 15384 13444
rect 14967 13413 14979 13416
rect 14921 13407 14979 13413
rect 15378 13404 15384 13416
rect 15436 13444 15442 13456
rect 17678 13444 17684 13456
rect 15436 13416 17684 13444
rect 15436 13404 15442 13416
rect 17678 13404 17684 13416
rect 17736 13404 17742 13456
rect 18598 13404 18604 13456
rect 18656 13444 18662 13456
rect 18785 13447 18843 13453
rect 18785 13444 18797 13447
rect 18656 13416 18797 13444
rect 18656 13404 18662 13416
rect 18785 13413 18797 13416
rect 18831 13413 18843 13447
rect 18785 13407 18843 13413
rect 20070 13404 20076 13456
rect 20128 13444 20134 13456
rect 20257 13447 20315 13453
rect 20257 13444 20269 13447
rect 20128 13416 20269 13444
rect 20128 13404 20134 13416
rect 20257 13413 20269 13416
rect 20303 13413 20315 13447
rect 20257 13407 20315 13413
rect 21358 13404 21364 13456
rect 21416 13444 21422 13456
rect 21913 13447 21971 13453
rect 21913 13444 21925 13447
rect 21416 13416 21925 13444
rect 21416 13404 21422 13416
rect 21913 13413 21925 13416
rect 21959 13413 21971 13447
rect 21913 13407 21971 13413
rect 22278 13404 22284 13456
rect 22336 13453 22342 13456
rect 22336 13447 22400 13453
rect 22336 13413 22354 13447
rect 22388 13444 22400 13447
rect 22554 13444 22560 13456
rect 22388 13416 22560 13444
rect 22388 13413 22400 13416
rect 22336 13407 22400 13413
rect 22336 13404 22342 13407
rect 22554 13404 22560 13416
rect 22612 13404 22618 13456
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 1486 13376 1492 13388
rect 1443 13348 1492 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 1486 13336 1492 13348
rect 1544 13336 1550 13388
rect 1670 13385 1676 13388
rect 1664 13376 1676 13385
rect 1631 13348 1676 13376
rect 1664 13339 1676 13348
rect 1670 13336 1676 13339
rect 1728 13336 1734 13388
rect 4617 13379 4675 13385
rect 4617 13345 4629 13379
rect 4663 13376 4675 13379
rect 5350 13376 5356 13388
rect 4663 13348 5356 13376
rect 4663 13345 4675 13348
rect 4617 13339 4675 13345
rect 4706 13268 4712 13320
rect 4764 13308 4770 13320
rect 5276 13317 5304 13348
rect 5350 13336 5356 13348
rect 5408 13336 5414 13388
rect 5442 13336 5448 13388
rect 5500 13376 5506 13388
rect 6273 13379 6331 13385
rect 6273 13376 6285 13379
rect 5500 13348 6285 13376
rect 5500 13336 5506 13348
rect 6273 13345 6285 13348
rect 6319 13345 6331 13379
rect 6273 13339 6331 13345
rect 8386 13336 8392 13388
rect 8444 13376 8450 13388
rect 8754 13376 8760 13388
rect 8444 13348 8760 13376
rect 8444 13336 8450 13348
rect 8754 13336 8760 13348
rect 8812 13336 8818 13388
rect 9214 13336 9220 13388
rect 9272 13376 9278 13388
rect 9582 13376 9588 13388
rect 9272 13348 9588 13376
rect 9272 13336 9278 13348
rect 9582 13336 9588 13348
rect 9640 13376 9646 13388
rect 9677 13379 9735 13385
rect 9677 13376 9689 13379
rect 9640 13348 9689 13376
rect 9640 13336 9646 13348
rect 9677 13345 9689 13348
rect 9723 13345 9735 13379
rect 9677 13339 9735 13345
rect 12158 13336 12164 13388
rect 12216 13376 12222 13388
rect 12529 13379 12587 13385
rect 12529 13376 12541 13379
rect 12216 13348 12541 13376
rect 12216 13336 12222 13348
rect 12529 13345 12541 13348
rect 12575 13345 12587 13379
rect 13906 13376 13912 13388
rect 12529 13339 12587 13345
rect 12636 13348 13912 13376
rect 5169 13311 5227 13317
rect 5169 13308 5181 13311
rect 4764 13280 5181 13308
rect 4764 13268 4770 13280
rect 5169 13277 5181 13280
rect 5215 13277 5227 13311
rect 5169 13271 5227 13277
rect 5261 13311 5319 13317
rect 5261 13277 5273 13311
rect 5307 13277 5319 13311
rect 5261 13271 5319 13277
rect 7926 13268 7932 13320
rect 7984 13308 7990 13320
rect 12636 13308 12664 13348
rect 13906 13336 13912 13348
rect 13964 13376 13970 13388
rect 14001 13379 14059 13385
rect 14001 13376 14013 13379
rect 13964 13348 14013 13376
rect 13964 13336 13970 13348
rect 14001 13345 14013 13348
rect 14047 13345 14059 13379
rect 14001 13339 14059 13345
rect 15194 13336 15200 13388
rect 15252 13376 15258 13388
rect 15562 13385 15568 13388
rect 15289 13379 15347 13385
rect 15289 13376 15301 13379
rect 15252 13348 15301 13376
rect 15252 13336 15258 13348
rect 15289 13345 15301 13348
rect 15335 13345 15347 13379
rect 15556 13376 15568 13385
rect 15523 13348 15568 13376
rect 15289 13339 15347 13345
rect 15556 13339 15568 13348
rect 15562 13336 15568 13339
rect 15620 13336 15626 13388
rect 18230 13376 18236 13388
rect 18191 13348 18236 13376
rect 18230 13336 18236 13348
rect 18288 13376 18294 13388
rect 19153 13379 19211 13385
rect 19153 13376 19165 13379
rect 18288 13348 19165 13376
rect 18288 13336 18294 13348
rect 19153 13345 19165 13348
rect 19199 13345 19211 13379
rect 19153 13339 19211 13345
rect 19705 13379 19763 13385
rect 19705 13345 19717 13379
rect 19751 13345 19763 13379
rect 19705 13339 19763 13345
rect 12802 13308 12808 13320
rect 7984 13280 9168 13308
rect 7984 13268 7990 13280
rect 3142 13200 3148 13252
rect 3200 13240 3206 13252
rect 8386 13240 8392 13252
rect 3200 13212 5304 13240
rect 3200 13200 3206 13212
rect 2777 13175 2835 13181
rect 2777 13141 2789 13175
rect 2823 13172 2835 13175
rect 2958 13172 2964 13184
rect 2823 13144 2964 13172
rect 2823 13141 2835 13144
rect 2777 13135 2835 13141
rect 2958 13132 2964 13144
rect 3016 13132 3022 13184
rect 3326 13172 3332 13184
rect 3287 13144 3332 13172
rect 3326 13132 3332 13144
rect 3384 13132 3390 13184
rect 3694 13172 3700 13184
rect 3655 13144 3700 13172
rect 3694 13132 3700 13144
rect 3752 13132 3758 13184
rect 5276 13172 5304 13212
rect 7208 13212 8392 13240
rect 7208 13172 7236 13212
rect 8386 13200 8392 13212
rect 8444 13200 8450 13252
rect 9140 13240 9168 13280
rect 11624 13280 12664 13308
rect 12763 13280 12808 13308
rect 9582 13240 9588 13252
rect 9140 13212 9588 13240
rect 9582 13200 9588 13212
rect 9640 13200 9646 13252
rect 10778 13200 10784 13252
rect 10836 13240 10842 13252
rect 11624 13249 11652 13280
rect 12802 13268 12808 13280
rect 12860 13268 12866 13320
rect 14182 13308 14188 13320
rect 14143 13280 14188 13308
rect 14182 13268 14188 13280
rect 14240 13268 14246 13320
rect 18414 13308 18420 13320
rect 18375 13280 18420 13308
rect 18414 13268 18420 13280
rect 18472 13268 18478 13320
rect 19720 13308 19748 13339
rect 20806 13336 20812 13388
rect 20864 13376 20870 13388
rect 20993 13379 21051 13385
rect 20993 13376 21005 13379
rect 20864 13348 21005 13376
rect 20864 13336 20870 13348
rect 20993 13345 21005 13348
rect 21039 13345 21051 13379
rect 20993 13339 21051 13345
rect 22002 13336 22008 13388
rect 22060 13376 22066 13388
rect 22097 13379 22155 13385
rect 22097 13376 22109 13379
rect 22060 13348 22109 13376
rect 22060 13336 22066 13348
rect 22097 13345 22109 13348
rect 22143 13376 22155 13379
rect 23566 13376 23572 13388
rect 22143 13348 23572 13376
rect 22143 13345 22155 13348
rect 22097 13339 22155 13345
rect 23566 13336 23572 13348
rect 23624 13336 23630 13388
rect 20717 13311 20775 13317
rect 20717 13308 20729 13311
rect 19720 13280 20729 13308
rect 20717 13277 20729 13280
rect 20763 13308 20775 13311
rect 21818 13308 21824 13320
rect 20763 13280 21824 13308
rect 20763 13277 20775 13280
rect 20717 13271 20775 13277
rect 21818 13268 21824 13280
rect 21876 13268 21882 13320
rect 25038 13308 25044 13320
rect 24999 13280 25044 13308
rect 25038 13268 25044 13280
rect 25096 13268 25102 13320
rect 25133 13311 25191 13317
rect 25133 13277 25145 13311
rect 25179 13277 25191 13311
rect 25133 13271 25191 13277
rect 11609 13243 11667 13249
rect 11609 13240 11621 13243
rect 10836 13212 11621 13240
rect 10836 13200 10842 13212
rect 11609 13209 11621 13212
rect 11655 13209 11667 13243
rect 11609 13203 11667 13209
rect 11790 13200 11796 13252
rect 11848 13240 11854 13252
rect 12820 13240 12848 13268
rect 11848 13212 12848 13240
rect 11848 13200 11854 13212
rect 24762 13200 24768 13252
rect 24820 13240 24826 13252
rect 25148 13240 25176 13271
rect 24820 13212 25176 13240
rect 24820 13200 24826 13212
rect 5276 13144 7236 13172
rect 8294 13132 8300 13184
rect 8352 13172 8358 13184
rect 11054 13172 11060 13184
rect 8352 13144 11060 13172
rect 8352 13132 8358 13144
rect 11054 13132 11060 13144
rect 11112 13132 11118 13184
rect 11146 13132 11152 13184
rect 11204 13172 11210 13184
rect 11808 13172 11836 13200
rect 16666 13172 16672 13184
rect 11204 13144 11836 13172
rect 16627 13144 16672 13172
rect 11204 13132 11210 13144
rect 16666 13132 16672 13144
rect 16724 13132 16730 13184
rect 24118 13132 24124 13184
rect 24176 13172 24182 13184
rect 24489 13175 24547 13181
rect 24489 13172 24501 13175
rect 24176 13144 24501 13172
rect 24176 13132 24182 13144
rect 24489 13141 24501 13144
rect 24535 13172 24547 13175
rect 24581 13175 24639 13181
rect 24581 13172 24593 13175
rect 24535 13144 24593 13172
rect 24535 13141 24547 13144
rect 24489 13135 24547 13141
rect 24581 13141 24593 13144
rect 24627 13141 24639 13175
rect 25590 13172 25596 13184
rect 25551 13144 25596 13172
rect 24581 13135 24639 13141
rect 25590 13132 25596 13144
rect 25648 13132 25654 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1854 12928 1860 12980
rect 1912 12968 1918 12980
rect 3970 12968 3976 12980
rect 1912 12940 3096 12968
rect 3931 12940 3976 12968
rect 1912 12928 1918 12940
rect 1578 12832 1584 12844
rect 1539 12804 1584 12832
rect 1578 12792 1584 12804
rect 1636 12792 1642 12844
rect 3068 12832 3096 12940
rect 3970 12928 3976 12940
rect 4028 12928 4034 12980
rect 4890 12968 4896 12980
rect 4851 12940 4896 12968
rect 4890 12928 4896 12940
rect 4948 12928 4954 12980
rect 6638 12968 6644 12980
rect 6599 12940 6644 12968
rect 6638 12928 6644 12940
rect 6696 12968 6702 12980
rect 6825 12971 6883 12977
rect 6825 12968 6837 12971
rect 6696 12940 6837 12968
rect 6696 12928 6702 12940
rect 6825 12937 6837 12940
rect 6871 12937 6883 12971
rect 6825 12931 6883 12937
rect 6917 12971 6975 12977
rect 6917 12937 6929 12971
rect 6963 12968 6975 12971
rect 7558 12968 7564 12980
rect 6963 12940 7564 12968
rect 6963 12937 6975 12940
rect 6917 12931 6975 12937
rect 7558 12928 7564 12940
rect 7616 12928 7622 12980
rect 9582 12928 9588 12980
rect 9640 12968 9646 12980
rect 9858 12968 9864 12980
rect 9640 12940 9864 12968
rect 9640 12928 9646 12940
rect 9858 12928 9864 12940
rect 9916 12928 9922 12980
rect 9950 12928 9956 12980
rect 10008 12968 10014 12980
rect 10413 12971 10471 12977
rect 10413 12968 10425 12971
rect 10008 12940 10425 12968
rect 10008 12928 10014 12940
rect 10413 12937 10425 12940
rect 10459 12937 10471 12971
rect 10413 12931 10471 12937
rect 11698 12928 11704 12980
rect 11756 12968 11762 12980
rect 11793 12971 11851 12977
rect 11793 12968 11805 12971
rect 11756 12940 11805 12968
rect 11756 12928 11762 12940
rect 11793 12937 11805 12940
rect 11839 12968 11851 12971
rect 12158 12968 12164 12980
rect 11839 12940 12164 12968
rect 11839 12937 11851 12940
rect 11793 12931 11851 12937
rect 12158 12928 12164 12940
rect 12216 12928 12222 12980
rect 12253 12971 12311 12977
rect 12253 12937 12265 12971
rect 12299 12968 12311 12971
rect 12526 12968 12532 12980
rect 12299 12940 12532 12968
rect 12299 12937 12311 12940
rect 12253 12931 12311 12937
rect 12526 12928 12532 12940
rect 12584 12928 12590 12980
rect 13004 12940 13860 12968
rect 4341 12903 4399 12909
rect 4341 12900 4353 12903
rect 4172 12872 4353 12900
rect 4172 12832 4200 12872
rect 4341 12869 4353 12872
rect 4387 12900 4399 12903
rect 4617 12903 4675 12909
rect 4617 12900 4629 12903
rect 4387 12872 4629 12900
rect 4387 12869 4399 12872
rect 4341 12863 4399 12869
rect 4617 12869 4629 12872
rect 4663 12869 4675 12903
rect 4617 12863 4675 12869
rect 4816 12872 6224 12900
rect 4816 12832 4844 12872
rect 3068 12804 4200 12832
rect 4264 12804 4844 12832
rect 3602 12724 3608 12776
rect 3660 12764 3666 12776
rect 3878 12764 3884 12776
rect 3660 12736 3884 12764
rect 3660 12724 3666 12736
rect 3878 12724 3884 12736
rect 3936 12724 3942 12776
rect 1848 12699 1906 12705
rect 1848 12665 1860 12699
rect 1894 12696 1906 12699
rect 1946 12696 1952 12708
rect 1894 12668 1952 12696
rect 1894 12665 1906 12668
rect 1848 12659 1906 12665
rect 1946 12656 1952 12668
rect 2004 12696 2010 12708
rect 3050 12696 3056 12708
rect 2004 12668 3056 12696
rect 2004 12656 2010 12668
rect 3050 12656 3056 12668
rect 3108 12656 3114 12708
rect 4264 12696 4292 12804
rect 5350 12792 5356 12844
rect 5408 12832 5414 12844
rect 5445 12835 5503 12841
rect 5445 12832 5457 12835
rect 5408 12804 5457 12832
rect 5408 12792 5414 12804
rect 5445 12801 5457 12804
rect 5491 12801 5503 12835
rect 5445 12795 5503 12801
rect 3620 12668 4292 12696
rect 4617 12699 4675 12705
rect 3620 12640 3648 12668
rect 4617 12665 4629 12699
rect 4663 12696 4675 12699
rect 4663 12668 4936 12696
rect 4663 12665 4675 12668
rect 4617 12659 4675 12665
rect 1210 12588 1216 12640
rect 1268 12628 1274 12640
rect 1394 12628 1400 12640
rect 1268 12600 1400 12628
rect 1268 12588 1274 12600
rect 1394 12588 1400 12600
rect 1452 12588 1458 12640
rect 1670 12588 1676 12640
rect 1728 12628 1734 12640
rect 2682 12628 2688 12640
rect 1728 12600 2688 12628
rect 1728 12588 1734 12600
rect 2682 12588 2688 12600
rect 2740 12628 2746 12640
rect 2961 12631 3019 12637
rect 2961 12628 2973 12631
rect 2740 12600 2973 12628
rect 2740 12588 2746 12600
rect 2961 12597 2973 12600
rect 3007 12597 3019 12631
rect 3510 12628 3516 12640
rect 3471 12600 3516 12628
rect 2961 12591 3019 12597
rect 3510 12588 3516 12600
rect 3568 12588 3574 12640
rect 3602 12588 3608 12640
rect 3660 12588 3666 12640
rect 4430 12588 4436 12640
rect 4488 12628 4494 12640
rect 4706 12628 4712 12640
rect 4488 12600 4712 12628
rect 4488 12588 4494 12600
rect 4706 12588 4712 12600
rect 4764 12588 4770 12640
rect 4908 12628 4936 12668
rect 4982 12656 4988 12708
rect 5040 12696 5046 12708
rect 5353 12699 5411 12705
rect 5353 12696 5365 12699
rect 5040 12668 5365 12696
rect 5040 12656 5046 12668
rect 5353 12665 5365 12668
rect 5399 12665 5411 12699
rect 6196 12696 6224 12872
rect 6730 12860 6736 12912
rect 6788 12900 6794 12912
rect 7929 12903 7987 12909
rect 7929 12900 7941 12903
rect 6788 12872 7941 12900
rect 6788 12860 6794 12872
rect 7929 12869 7941 12872
rect 7975 12869 7987 12903
rect 13004 12900 13032 12940
rect 7929 12863 7987 12869
rect 11164 12872 13032 12900
rect 7561 12835 7619 12841
rect 7561 12801 7573 12835
rect 7607 12832 7619 12835
rect 7650 12832 7656 12844
rect 7607 12804 7656 12832
rect 7607 12801 7619 12804
rect 7561 12795 7619 12801
rect 7650 12792 7656 12804
rect 7708 12792 7714 12844
rect 9950 12792 9956 12844
rect 10008 12832 10014 12844
rect 10686 12832 10692 12844
rect 10008 12804 10692 12832
rect 10008 12792 10014 12804
rect 10686 12792 10692 12804
rect 10744 12792 10750 12844
rect 6273 12767 6331 12773
rect 6273 12733 6285 12767
rect 6319 12764 6331 12767
rect 7285 12767 7343 12773
rect 7285 12764 7297 12767
rect 6319 12736 7297 12764
rect 6319 12733 6331 12736
rect 6273 12727 6331 12733
rect 7285 12733 7297 12736
rect 7331 12764 7343 12767
rect 7374 12764 7380 12776
rect 7331 12736 7380 12764
rect 7331 12733 7343 12736
rect 7285 12727 7343 12733
rect 7374 12724 7380 12736
rect 7432 12724 7438 12776
rect 8294 12764 8300 12776
rect 8255 12736 8300 12764
rect 8294 12724 8300 12736
rect 8352 12724 8358 12776
rect 8481 12767 8539 12773
rect 8481 12733 8493 12767
rect 8527 12764 8539 12767
rect 9214 12764 9220 12776
rect 8527 12736 9220 12764
rect 8527 12733 8539 12736
rect 8481 12727 8539 12733
rect 9214 12724 9220 12736
rect 9272 12724 9278 12776
rect 10042 12724 10048 12776
rect 10100 12764 10106 12776
rect 10594 12764 10600 12776
rect 10100 12736 10600 12764
rect 10100 12724 10106 12736
rect 10594 12724 10600 12736
rect 10652 12724 10658 12776
rect 6638 12696 6644 12708
rect 6196 12668 6644 12696
rect 5353 12659 5411 12665
rect 6638 12656 6644 12668
rect 6696 12656 6702 12708
rect 8312 12696 8340 12724
rect 8726 12699 8784 12705
rect 8726 12696 8738 12699
rect 8312 12668 8738 12696
rect 8726 12665 8738 12668
rect 8772 12665 8784 12699
rect 8726 12659 8784 12665
rect 10686 12656 10692 12708
rect 10744 12696 10750 12708
rect 11164 12705 11192 12872
rect 11330 12832 11336 12844
rect 11291 12804 11336 12832
rect 11330 12792 11336 12804
rect 11388 12792 11394 12844
rect 12710 12792 12716 12844
rect 12768 12832 12774 12844
rect 13004 12841 13032 12872
rect 12897 12835 12955 12841
rect 12897 12832 12909 12835
rect 12768 12804 12909 12832
rect 12768 12792 12774 12804
rect 12897 12801 12909 12804
rect 12943 12801 12955 12835
rect 12897 12795 12955 12801
rect 12989 12835 13047 12841
rect 12989 12801 13001 12835
rect 13035 12801 13047 12835
rect 12989 12795 13047 12801
rect 13262 12792 13268 12844
rect 13320 12832 13326 12844
rect 13832 12841 13860 12940
rect 14734 12928 14740 12980
rect 14792 12968 14798 12980
rect 14829 12971 14887 12977
rect 14829 12968 14841 12971
rect 14792 12940 14841 12968
rect 14792 12928 14798 12940
rect 14829 12937 14841 12940
rect 14875 12937 14887 12971
rect 14829 12931 14887 12937
rect 15286 12928 15292 12980
rect 15344 12968 15350 12980
rect 16298 12968 16304 12980
rect 15344 12940 16304 12968
rect 15344 12928 15350 12940
rect 16298 12928 16304 12940
rect 16356 12968 16362 12980
rect 16393 12971 16451 12977
rect 16393 12968 16405 12971
rect 16356 12940 16405 12968
rect 16356 12928 16362 12940
rect 16393 12937 16405 12940
rect 16439 12937 16451 12971
rect 17494 12968 17500 12980
rect 17455 12940 17500 12968
rect 16393 12931 16451 12937
rect 17494 12928 17500 12940
rect 17552 12928 17558 12980
rect 17865 12971 17923 12977
rect 17865 12937 17877 12971
rect 17911 12968 17923 12971
rect 18414 12968 18420 12980
rect 17911 12940 18420 12968
rect 17911 12937 17923 12940
rect 17865 12931 17923 12937
rect 18414 12928 18420 12940
rect 18472 12928 18478 12980
rect 20990 12968 20996 12980
rect 20951 12940 20996 12968
rect 20990 12928 20996 12940
rect 21048 12928 21054 12980
rect 23750 12928 23756 12980
rect 23808 12968 23814 12980
rect 24762 12968 24768 12980
rect 23808 12940 24768 12968
rect 23808 12928 23814 12940
rect 24762 12928 24768 12940
rect 24820 12928 24826 12980
rect 25130 12928 25136 12980
rect 25188 12968 25194 12980
rect 25961 12971 26019 12977
rect 25961 12968 25973 12971
rect 25188 12940 25973 12968
rect 25188 12928 25194 12940
rect 25961 12937 25973 12940
rect 26007 12937 26019 12971
rect 25961 12931 26019 12937
rect 26234 12928 26240 12980
rect 26292 12968 26298 12980
rect 26329 12971 26387 12977
rect 26329 12968 26341 12971
rect 26292 12940 26341 12968
rect 26292 12928 26298 12940
rect 26329 12937 26341 12940
rect 26375 12937 26387 12971
rect 26329 12931 26387 12937
rect 14645 12903 14703 12909
rect 14645 12869 14657 12903
rect 14691 12900 14703 12903
rect 15562 12900 15568 12912
rect 14691 12872 15568 12900
rect 14691 12869 14703 12872
rect 14645 12863 14703 12869
rect 15562 12860 15568 12872
rect 15620 12860 15626 12912
rect 15654 12860 15660 12912
rect 15712 12900 15718 12912
rect 15838 12900 15844 12912
rect 15712 12872 15844 12900
rect 15712 12860 15718 12872
rect 15838 12860 15844 12872
rect 15896 12860 15902 12912
rect 13725 12835 13783 12841
rect 13725 12832 13737 12835
rect 13320 12804 13737 12832
rect 13320 12792 13326 12804
rect 13725 12801 13737 12804
rect 13771 12801 13783 12835
rect 13725 12795 13783 12801
rect 13817 12835 13875 12841
rect 13817 12801 13829 12835
rect 13863 12832 13875 12835
rect 14277 12835 14335 12841
rect 14277 12832 14289 12835
rect 13863 12804 14289 12832
rect 13863 12801 13875 12804
rect 13817 12795 13875 12801
rect 14277 12801 14289 12804
rect 14323 12801 14335 12835
rect 15378 12832 15384 12844
rect 15339 12804 15384 12832
rect 14277 12795 14335 12801
rect 15378 12792 15384 12804
rect 15436 12792 15442 12844
rect 16206 12832 16212 12844
rect 16167 12804 16212 12832
rect 16206 12792 16212 12804
rect 16264 12832 16270 12844
rect 17037 12835 17095 12841
rect 16264 12804 16804 12832
rect 16264 12792 16270 12804
rect 12434 12724 12440 12776
rect 12492 12764 12498 12776
rect 12805 12767 12863 12773
rect 12805 12764 12817 12767
rect 12492 12736 12817 12764
rect 12492 12724 12498 12736
rect 12805 12733 12817 12736
rect 12851 12733 12863 12767
rect 12805 12727 12863 12733
rect 11149 12699 11207 12705
rect 11149 12696 11161 12699
rect 10744 12668 11161 12696
rect 10744 12656 10750 12668
rect 11149 12665 11161 12668
rect 11195 12665 11207 12699
rect 12618 12696 12624 12708
rect 11149 12659 11207 12665
rect 12452 12668 12624 12696
rect 5261 12631 5319 12637
rect 5261 12628 5273 12631
rect 4908 12600 5273 12628
rect 5261 12597 5273 12600
rect 5307 12597 5319 12631
rect 5261 12591 5319 12597
rect 6825 12631 6883 12637
rect 6825 12597 6837 12631
rect 6871 12628 6883 12631
rect 7377 12631 7435 12637
rect 7377 12628 7389 12631
rect 6871 12600 7389 12628
rect 6871 12597 6883 12600
rect 6825 12591 6883 12597
rect 7377 12597 7389 12600
rect 7423 12597 7435 12631
rect 10778 12628 10784 12640
rect 10739 12600 10784 12628
rect 7377 12591 7435 12597
rect 10778 12588 10784 12600
rect 10836 12588 10842 12640
rect 12452 12637 12480 12668
rect 12618 12656 12624 12668
rect 12676 12656 12682 12708
rect 12820 12696 12848 12727
rect 13538 12724 13544 12776
rect 13596 12764 13602 12776
rect 13633 12767 13691 12773
rect 13633 12764 13645 12767
rect 13596 12736 13645 12764
rect 13596 12724 13602 12736
rect 13633 12733 13645 12736
rect 13679 12733 13691 12767
rect 13633 12727 13691 12733
rect 15102 12724 15108 12776
rect 15160 12764 15166 12776
rect 15289 12767 15347 12773
rect 15289 12764 15301 12767
rect 15160 12736 15301 12764
rect 15160 12724 15166 12736
rect 15289 12733 15301 12736
rect 15335 12764 15347 12767
rect 15470 12764 15476 12776
rect 15335 12736 15476 12764
rect 15335 12733 15347 12736
rect 15289 12727 15347 12733
rect 15470 12724 15476 12736
rect 15528 12724 15534 12776
rect 16776 12773 16804 12804
rect 17037 12801 17049 12835
rect 17083 12832 17095 12835
rect 17512 12832 17540 12928
rect 17083 12804 17540 12832
rect 18432 12832 18460 12928
rect 20070 12860 20076 12912
rect 20128 12900 20134 12912
rect 20441 12903 20499 12909
rect 20441 12900 20453 12903
rect 20128 12872 20453 12900
rect 20128 12860 20134 12872
rect 20441 12869 20453 12872
rect 20487 12869 20499 12903
rect 20441 12863 20499 12869
rect 23661 12903 23719 12909
rect 23661 12869 23673 12903
rect 23707 12900 23719 12903
rect 24670 12900 24676 12912
rect 23707 12872 24676 12900
rect 23707 12869 23719 12872
rect 23661 12863 23719 12869
rect 20456 12832 20484 12863
rect 24670 12860 24676 12872
rect 24728 12860 24734 12912
rect 21453 12835 21511 12841
rect 21453 12832 21465 12835
rect 18432 12804 18644 12832
rect 20456 12804 21465 12832
rect 17083 12801 17095 12804
rect 17037 12795 17095 12801
rect 16761 12767 16819 12773
rect 16761 12733 16773 12767
rect 16807 12733 16819 12767
rect 16761 12727 16819 12733
rect 18230 12724 18236 12776
rect 18288 12764 18294 12776
rect 18509 12767 18567 12773
rect 18509 12764 18521 12767
rect 18288 12736 18521 12764
rect 18288 12724 18294 12736
rect 18509 12733 18521 12736
rect 18555 12733 18567 12767
rect 18616 12764 18644 12804
rect 21453 12801 21465 12804
rect 21499 12801 21511 12835
rect 21634 12832 21640 12844
rect 21547 12804 21640 12832
rect 21453 12795 21511 12801
rect 21634 12792 21640 12804
rect 21692 12832 21698 12844
rect 22373 12835 22431 12841
rect 22373 12832 22385 12835
rect 21692 12804 22385 12832
rect 21692 12792 21698 12804
rect 22373 12801 22385 12804
rect 22419 12801 22431 12835
rect 22373 12795 22431 12801
rect 22557 12835 22615 12841
rect 22557 12801 22569 12835
rect 22603 12832 22615 12835
rect 23198 12832 23204 12844
rect 22603 12804 23204 12832
rect 22603 12801 22615 12804
rect 22557 12795 22615 12801
rect 23198 12792 23204 12804
rect 23256 12792 23262 12844
rect 24213 12835 24271 12841
rect 24213 12801 24225 12835
rect 24259 12801 24271 12835
rect 25038 12832 25044 12844
rect 24999 12804 25044 12832
rect 24213 12795 24271 12801
rect 18765 12767 18823 12773
rect 18765 12764 18777 12767
rect 18616 12736 18777 12764
rect 18509 12727 18567 12733
rect 18765 12733 18777 12736
rect 18811 12733 18823 12767
rect 18765 12727 18823 12733
rect 20254 12724 20260 12776
rect 20312 12764 20318 12776
rect 20990 12764 20996 12776
rect 20312 12736 20996 12764
rect 20312 12724 20318 12736
rect 20990 12724 20996 12736
rect 21048 12724 21054 12776
rect 22278 12724 22284 12776
rect 22336 12764 22342 12776
rect 23106 12764 23112 12776
rect 22336 12736 23112 12764
rect 22336 12724 22342 12736
rect 23106 12724 23112 12736
rect 23164 12724 23170 12776
rect 24029 12767 24087 12773
rect 24029 12733 24041 12767
rect 24075 12764 24087 12767
rect 24118 12764 24124 12776
rect 24075 12736 24124 12764
rect 24075 12733 24087 12736
rect 24029 12727 24087 12733
rect 24118 12724 24124 12736
rect 24176 12724 24182 12776
rect 15933 12699 15991 12705
rect 12820 12668 15884 12696
rect 12437 12631 12495 12637
rect 12437 12597 12449 12631
rect 12483 12597 12495 12631
rect 13262 12628 13268 12640
rect 13223 12600 13268 12628
rect 12437 12591 12495 12597
rect 13262 12588 13268 12600
rect 13320 12588 13326 12640
rect 15194 12628 15200 12640
rect 15155 12600 15200 12628
rect 15194 12588 15200 12600
rect 15252 12588 15258 12640
rect 15856 12628 15884 12668
rect 15933 12665 15945 12699
rect 15979 12696 15991 12699
rect 16298 12696 16304 12708
rect 15979 12668 16304 12696
rect 15979 12665 15991 12668
rect 15933 12659 15991 12665
rect 16298 12656 16304 12668
rect 16356 12696 16362 12708
rect 16853 12699 16911 12705
rect 16853 12696 16865 12699
rect 16356 12668 16865 12696
rect 16356 12656 16362 12668
rect 16853 12665 16865 12668
rect 16899 12665 16911 12699
rect 16853 12659 16911 12665
rect 23477 12699 23535 12705
rect 23477 12665 23489 12699
rect 23523 12696 23535 12699
rect 23566 12696 23572 12708
rect 23523 12668 23572 12696
rect 23523 12665 23535 12668
rect 23477 12659 23535 12665
rect 23566 12656 23572 12668
rect 23624 12696 23630 12708
rect 24228 12696 24256 12795
rect 25038 12792 25044 12804
rect 25096 12792 25102 12844
rect 25498 12832 25504 12844
rect 25459 12804 25504 12832
rect 25498 12792 25504 12804
rect 25556 12792 25562 12844
rect 25130 12724 25136 12776
rect 25188 12764 25194 12776
rect 25225 12767 25283 12773
rect 25225 12764 25237 12767
rect 25188 12736 25237 12764
rect 25188 12724 25194 12736
rect 25225 12733 25237 12736
rect 25271 12764 25283 12767
rect 25590 12764 25596 12776
rect 25271 12736 25596 12764
rect 25271 12733 25283 12736
rect 25225 12727 25283 12733
rect 25590 12724 25596 12736
rect 25648 12724 25654 12776
rect 23624 12668 24256 12696
rect 23624 12656 23630 12668
rect 18046 12628 18052 12640
rect 15856 12600 18052 12628
rect 18046 12588 18052 12600
rect 18104 12588 18110 12640
rect 19889 12631 19947 12637
rect 19889 12597 19901 12631
rect 19935 12628 19947 12631
rect 20530 12628 20536 12640
rect 19935 12600 20536 12628
rect 19935 12597 19947 12600
rect 19889 12591 19947 12597
rect 20530 12588 20536 12600
rect 20588 12588 20594 12640
rect 20806 12628 20812 12640
rect 20767 12600 20812 12628
rect 20806 12588 20812 12600
rect 20864 12588 20870 12640
rect 21174 12588 21180 12640
rect 21232 12628 21238 12640
rect 21361 12631 21419 12637
rect 21361 12628 21373 12631
rect 21232 12600 21373 12628
rect 21232 12588 21238 12600
rect 21361 12597 21373 12600
rect 21407 12628 21419 12631
rect 22005 12631 22063 12637
rect 22005 12628 22017 12631
rect 21407 12600 22017 12628
rect 21407 12597 21419 12600
rect 21361 12591 21419 12597
rect 22005 12597 22017 12600
rect 22051 12597 22063 12631
rect 22005 12591 22063 12597
rect 23109 12631 23167 12637
rect 23109 12597 23121 12631
rect 23155 12628 23167 12631
rect 23382 12628 23388 12640
rect 23155 12600 23388 12628
rect 23155 12597 23167 12600
rect 23109 12591 23167 12597
rect 23382 12588 23388 12600
rect 23440 12628 23446 12640
rect 24121 12631 24179 12637
rect 24121 12628 24133 12631
rect 23440 12600 24133 12628
rect 23440 12588 23446 12600
rect 24121 12597 24133 12600
rect 24167 12597 24179 12631
rect 24121 12591 24179 12597
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1394 12424 1400 12436
rect 1355 12396 1400 12424
rect 1394 12384 1400 12396
rect 1452 12384 1458 12436
rect 2130 12384 2136 12436
rect 2188 12384 2194 12436
rect 2869 12427 2927 12433
rect 2869 12393 2881 12427
rect 2915 12424 2927 12427
rect 3418 12424 3424 12436
rect 2915 12396 3424 12424
rect 2915 12393 2927 12396
rect 2869 12387 2927 12393
rect 3418 12384 3424 12396
rect 3476 12384 3482 12436
rect 4154 12384 4160 12436
rect 4212 12424 4218 12436
rect 4249 12427 4307 12433
rect 4249 12424 4261 12427
rect 4212 12396 4261 12424
rect 4212 12384 4218 12396
rect 4249 12393 4261 12396
rect 4295 12393 4307 12427
rect 4249 12387 4307 12393
rect 6730 12384 6736 12436
rect 6788 12424 6794 12436
rect 6825 12427 6883 12433
rect 6825 12424 6837 12427
rect 6788 12396 6837 12424
rect 6788 12384 6794 12396
rect 6825 12393 6837 12396
rect 6871 12393 6883 12427
rect 6825 12387 6883 12393
rect 7457 12384 7463 12436
rect 7515 12424 7521 12436
rect 7745 12427 7803 12433
rect 7745 12424 7757 12427
rect 7515 12396 7757 12424
rect 7515 12384 7521 12396
rect 7745 12393 7757 12396
rect 7791 12393 7803 12427
rect 7745 12387 7803 12393
rect 8018 12384 8024 12436
rect 8076 12424 8082 12436
rect 9122 12424 9128 12436
rect 8076 12396 8616 12424
rect 9083 12396 9128 12424
rect 8076 12384 8082 12396
rect 1670 12112 1676 12164
rect 1728 12152 1734 12164
rect 1857 12155 1915 12161
rect 1857 12152 1869 12155
rect 1728 12124 1869 12152
rect 1728 12112 1734 12124
rect 1857 12121 1869 12124
rect 1903 12152 1915 12155
rect 2038 12152 2044 12164
rect 1903 12124 2044 12152
rect 1903 12121 1915 12124
rect 1857 12115 1915 12121
rect 2038 12112 2044 12124
rect 2096 12112 2102 12164
rect 1394 12044 1400 12096
rect 1452 12084 1458 12096
rect 2148 12084 2176 12384
rect 2317 12359 2375 12365
rect 2317 12325 2329 12359
rect 2363 12356 2375 12359
rect 2682 12356 2688 12368
rect 2363 12328 2688 12356
rect 2363 12325 2375 12328
rect 2317 12319 2375 12325
rect 2682 12316 2688 12328
rect 2740 12316 2746 12368
rect 5534 12316 5540 12368
rect 5592 12356 5598 12368
rect 5712 12359 5770 12365
rect 5712 12356 5724 12359
rect 5592 12328 5724 12356
rect 5592 12316 5598 12328
rect 5712 12325 5724 12328
rect 5758 12356 5770 12359
rect 6270 12356 6276 12368
rect 5758 12328 6276 12356
rect 5758 12325 5770 12328
rect 5712 12319 5770 12325
rect 6270 12316 6276 12328
rect 6328 12316 6334 12368
rect 8588 12356 8616 12396
rect 9122 12384 9128 12396
rect 9180 12384 9186 12436
rect 9674 12384 9680 12436
rect 9732 12424 9738 12436
rect 10873 12427 10931 12433
rect 10873 12424 10885 12427
rect 9732 12396 10885 12424
rect 9732 12384 9738 12396
rect 10873 12393 10885 12396
rect 10919 12393 10931 12427
rect 10873 12387 10931 12393
rect 11238 12384 11244 12436
rect 11296 12424 11302 12436
rect 12069 12427 12127 12433
rect 12069 12424 12081 12427
rect 11296 12396 12081 12424
rect 11296 12384 11302 12396
rect 12069 12393 12081 12396
rect 12115 12424 12127 12427
rect 12434 12424 12440 12436
rect 12115 12396 12440 12424
rect 12115 12393 12127 12396
rect 12069 12387 12127 12393
rect 12434 12384 12440 12396
rect 12492 12384 12498 12436
rect 12529 12427 12587 12433
rect 12529 12393 12541 12427
rect 12575 12424 12587 12427
rect 12710 12424 12716 12436
rect 12575 12396 12716 12424
rect 12575 12393 12587 12396
rect 12529 12387 12587 12393
rect 12710 12384 12716 12396
rect 12768 12384 12774 12436
rect 15102 12424 15108 12436
rect 15063 12396 15108 12424
rect 15102 12384 15108 12396
rect 15160 12384 15166 12436
rect 15194 12384 15200 12436
rect 15252 12424 15258 12436
rect 15565 12427 15623 12433
rect 15565 12424 15577 12427
rect 15252 12396 15577 12424
rect 15252 12384 15258 12396
rect 15565 12393 15577 12396
rect 15611 12424 15623 12427
rect 16390 12424 16396 12436
rect 15611 12396 16396 12424
rect 15611 12393 15623 12396
rect 15565 12387 15623 12393
rect 16390 12384 16396 12396
rect 16448 12384 16454 12436
rect 16666 12384 16672 12436
rect 16724 12424 16730 12436
rect 17494 12424 17500 12436
rect 16724 12396 17500 12424
rect 16724 12384 16730 12396
rect 17494 12384 17500 12396
rect 17552 12384 17558 12436
rect 21358 12384 21364 12436
rect 21416 12424 21422 12436
rect 22189 12427 22247 12433
rect 21416 12396 21588 12424
rect 21416 12384 21422 12396
rect 9030 12356 9036 12368
rect 8588 12328 9036 12356
rect 9030 12316 9036 12328
rect 9088 12316 9094 12368
rect 9858 12356 9864 12368
rect 9819 12328 9864 12356
rect 9858 12316 9864 12328
rect 9916 12316 9922 12368
rect 9950 12316 9956 12368
rect 10008 12356 10014 12368
rect 10226 12356 10232 12368
rect 10008 12328 10232 12356
rect 10008 12316 10014 12328
rect 10226 12316 10232 12328
rect 10284 12316 10290 12368
rect 10413 12359 10471 12365
rect 10413 12325 10425 12359
rect 10459 12356 10471 12359
rect 10778 12356 10784 12368
rect 10459 12328 10784 12356
rect 10459 12325 10471 12328
rect 10413 12319 10471 12325
rect 2777 12291 2835 12297
rect 2777 12257 2789 12291
rect 2823 12288 2835 12291
rect 3789 12291 3847 12297
rect 3789 12288 3801 12291
rect 2823 12260 3801 12288
rect 2823 12257 2835 12260
rect 2777 12251 2835 12257
rect 3789 12257 3801 12260
rect 3835 12288 3847 12291
rect 3878 12288 3884 12300
rect 3835 12260 3884 12288
rect 3835 12257 3847 12260
rect 3789 12251 3847 12257
rect 3878 12248 3884 12260
rect 3936 12248 3942 12300
rect 4065 12291 4123 12297
rect 4065 12257 4077 12291
rect 4111 12288 4123 12291
rect 4246 12288 4252 12300
rect 4111 12260 4252 12288
rect 4111 12257 4123 12260
rect 4065 12251 4123 12257
rect 4246 12248 4252 12260
rect 4304 12248 4310 12300
rect 5442 12288 5448 12300
rect 5403 12260 5448 12288
rect 5442 12248 5448 12260
rect 5500 12248 5506 12300
rect 6914 12288 6920 12300
rect 5552 12260 6920 12288
rect 3050 12220 3056 12232
rect 2963 12192 3056 12220
rect 3050 12180 3056 12192
rect 3108 12220 3114 12232
rect 3602 12220 3608 12232
rect 3108 12192 3608 12220
rect 3108 12180 3114 12192
rect 3602 12180 3608 12192
rect 3660 12180 3666 12232
rect 5552 12220 5580 12260
rect 6914 12248 6920 12260
rect 6972 12248 6978 12300
rect 7834 12248 7840 12300
rect 7892 12288 7898 12300
rect 8389 12291 8447 12297
rect 8389 12288 8401 12291
rect 7892 12260 8401 12288
rect 7892 12248 7898 12260
rect 8389 12257 8401 12260
rect 8435 12257 8447 12291
rect 8389 12251 8447 12257
rect 9122 12248 9128 12300
rect 9180 12288 9186 12300
rect 9493 12291 9551 12297
rect 9493 12288 9505 12291
rect 9180 12260 9505 12288
rect 9180 12248 9186 12260
rect 9493 12257 9505 12260
rect 9539 12288 9551 12291
rect 10428 12288 10456 12319
rect 10778 12316 10784 12328
rect 10836 12316 10842 12368
rect 11422 12316 11428 12368
rect 11480 12356 11486 12368
rect 16292 12359 16350 12365
rect 11480 12328 14228 12356
rect 11480 12316 11486 12328
rect 11238 12288 11244 12300
rect 9539 12260 10456 12288
rect 11199 12260 11244 12288
rect 9539 12257 9551 12260
rect 9493 12251 9551 12257
rect 11238 12248 11244 12260
rect 11296 12248 11302 12300
rect 11333 12291 11391 12297
rect 11333 12257 11345 12291
rect 11379 12288 11391 12291
rect 11379 12260 11928 12288
rect 11379 12257 11391 12260
rect 11333 12251 11391 12257
rect 11900 12232 11928 12260
rect 12158 12248 12164 12300
rect 12216 12288 12222 12300
rect 12621 12291 12679 12297
rect 12621 12288 12633 12291
rect 12216 12260 12633 12288
rect 12216 12248 12222 12260
rect 12621 12257 12633 12260
rect 12667 12257 12679 12291
rect 12621 12251 12679 12257
rect 13998 12248 14004 12300
rect 14056 12288 14062 12300
rect 14056 12260 14136 12288
rect 14056 12248 14062 12260
rect 5460 12192 5580 12220
rect 2409 12155 2467 12161
rect 2409 12121 2421 12155
rect 2455 12152 2467 12155
rect 5460 12152 5488 12192
rect 7098 12180 7104 12232
rect 7156 12220 7162 12232
rect 7558 12220 7564 12232
rect 7156 12192 7564 12220
rect 7156 12180 7162 12192
rect 7558 12180 7564 12192
rect 7616 12180 7622 12232
rect 7742 12180 7748 12232
rect 7800 12220 7806 12232
rect 8478 12220 8484 12232
rect 7800 12192 8484 12220
rect 7800 12180 7806 12192
rect 8478 12180 8484 12192
rect 8536 12180 8542 12232
rect 8662 12220 8668 12232
rect 8623 12192 8668 12220
rect 8662 12180 8668 12192
rect 8720 12180 8726 12232
rect 9858 12180 9864 12232
rect 9916 12220 9922 12232
rect 10134 12220 10140 12232
rect 9916 12192 10140 12220
rect 9916 12180 9922 12192
rect 10134 12180 10140 12192
rect 10192 12180 10198 12232
rect 11425 12223 11483 12229
rect 11425 12189 11437 12223
rect 11471 12189 11483 12223
rect 11425 12183 11483 12189
rect 8680 12152 8708 12180
rect 2455 12124 5488 12152
rect 6932 12124 8708 12152
rect 10781 12155 10839 12161
rect 2455 12121 2467 12124
rect 2409 12115 2467 12121
rect 4982 12084 4988 12096
rect 1452 12056 2176 12084
rect 4943 12056 4988 12084
rect 1452 12044 1458 12056
rect 4982 12044 4988 12056
rect 5040 12044 5046 12096
rect 5350 12084 5356 12096
rect 5263 12056 5356 12084
rect 5350 12044 5356 12056
rect 5408 12084 5414 12096
rect 6932 12084 6960 12124
rect 10781 12121 10793 12155
rect 10827 12152 10839 12155
rect 11146 12152 11152 12164
rect 10827 12124 11152 12152
rect 10827 12121 10839 12124
rect 10781 12115 10839 12121
rect 11146 12112 11152 12124
rect 11204 12152 11210 12164
rect 11440 12152 11468 12183
rect 11882 12180 11888 12232
rect 11940 12180 11946 12232
rect 11204 12124 11468 12152
rect 11204 12112 11210 12124
rect 12250 12112 12256 12164
rect 12308 12152 12314 12164
rect 13722 12152 13728 12164
rect 12308 12124 13728 12152
rect 12308 12112 12314 12124
rect 13722 12112 13728 12124
rect 13780 12152 13786 12164
rect 13909 12155 13967 12161
rect 13909 12152 13921 12155
rect 13780 12124 13921 12152
rect 13780 12112 13786 12124
rect 13909 12121 13921 12124
rect 13955 12121 13967 12155
rect 13909 12115 13967 12121
rect 14108 12096 14136 12260
rect 14200 12220 14228 12328
rect 16292 12325 16304 12359
rect 16338 12356 16350 12359
rect 16684 12356 16712 12384
rect 16338 12328 16712 12356
rect 16338 12325 16350 12328
rect 16292 12319 16350 12325
rect 17862 12316 17868 12368
rect 17920 12356 17926 12368
rect 18414 12356 18420 12368
rect 17920 12328 18420 12356
rect 17920 12316 17926 12328
rect 18414 12316 18420 12328
rect 18472 12316 18478 12368
rect 14461 12291 14519 12297
rect 14461 12257 14473 12291
rect 14507 12288 14519 12291
rect 14734 12288 14740 12300
rect 14507 12260 14740 12288
rect 14507 12257 14519 12260
rect 14461 12251 14519 12257
rect 14734 12248 14740 12260
rect 14792 12248 14798 12300
rect 15378 12248 15384 12300
rect 15436 12288 15442 12300
rect 16025 12291 16083 12297
rect 16025 12288 16037 12291
rect 15436 12260 16037 12288
rect 15436 12248 15442 12260
rect 16025 12257 16037 12260
rect 16071 12257 16083 12291
rect 16025 12251 16083 12257
rect 16850 12248 16856 12300
rect 16908 12288 16914 12300
rect 18049 12291 18107 12297
rect 18049 12288 18061 12291
rect 16908 12260 18061 12288
rect 16908 12248 16914 12260
rect 18049 12257 18061 12260
rect 18095 12257 18107 12291
rect 18049 12251 18107 12257
rect 18693 12291 18751 12297
rect 18693 12257 18705 12291
rect 18739 12288 18751 12291
rect 19518 12288 19524 12300
rect 18739 12260 19524 12288
rect 18739 12257 18751 12260
rect 18693 12251 18751 12257
rect 19518 12248 19524 12260
rect 19576 12248 19582 12300
rect 21269 12291 21327 12297
rect 21269 12257 21281 12291
rect 21315 12288 21327 12291
rect 21315 12260 21496 12288
rect 21315 12257 21327 12260
rect 21269 12251 21327 12257
rect 15930 12220 15936 12232
rect 14200 12192 15936 12220
rect 15930 12180 15936 12192
rect 15988 12180 15994 12232
rect 19613 12223 19671 12229
rect 19613 12220 19625 12223
rect 18984 12192 19625 12220
rect 18984 12096 19012 12192
rect 19613 12189 19625 12192
rect 19659 12189 19671 12223
rect 19613 12183 19671 12189
rect 19797 12223 19855 12229
rect 19797 12189 19809 12223
rect 19843 12220 19855 12223
rect 20070 12220 20076 12232
rect 19843 12192 20076 12220
rect 19843 12189 19855 12192
rect 19797 12183 19855 12189
rect 20070 12180 20076 12192
rect 20128 12180 20134 12232
rect 20717 12223 20775 12229
rect 20717 12189 20729 12223
rect 20763 12220 20775 12223
rect 20898 12220 20904 12232
rect 20763 12192 20904 12220
rect 20763 12189 20775 12192
rect 20717 12183 20775 12189
rect 20898 12180 20904 12192
rect 20956 12180 20962 12232
rect 21174 12180 21180 12232
rect 21232 12220 21238 12232
rect 21361 12223 21419 12229
rect 21361 12220 21373 12223
rect 21232 12192 21373 12220
rect 21232 12180 21238 12192
rect 21361 12189 21373 12192
rect 21407 12189 21419 12223
rect 21361 12183 21419 12189
rect 21468 12164 21496 12260
rect 21560 12229 21588 12396
rect 22189 12393 22201 12427
rect 22235 12424 22247 12427
rect 22278 12424 22284 12436
rect 22235 12396 22284 12424
rect 22235 12393 22247 12396
rect 22189 12387 22247 12393
rect 22278 12384 22284 12396
rect 22336 12384 22342 12436
rect 22830 12424 22836 12436
rect 22791 12396 22836 12424
rect 22830 12384 22836 12396
rect 22888 12384 22894 12436
rect 23290 12384 23296 12436
rect 23348 12424 23354 12436
rect 24302 12424 24308 12436
rect 23348 12396 24308 12424
rect 23348 12384 23354 12396
rect 24302 12384 24308 12396
rect 24360 12384 24366 12436
rect 25038 12384 25044 12436
rect 25096 12424 25102 12436
rect 25133 12427 25191 12433
rect 25133 12424 25145 12427
rect 25096 12396 25145 12424
rect 25096 12384 25102 12396
rect 25133 12393 25145 12396
rect 25179 12393 25191 12427
rect 25133 12387 25191 12393
rect 26145 12427 26203 12433
rect 26145 12393 26157 12427
rect 26191 12424 26203 12427
rect 26326 12424 26332 12436
rect 26191 12396 26332 12424
rect 26191 12393 26203 12396
rect 26145 12387 26203 12393
rect 26326 12384 26332 12396
rect 26384 12384 26390 12436
rect 23198 12356 23204 12368
rect 22664 12328 23204 12356
rect 22664 12297 22692 12328
rect 23198 12316 23204 12328
rect 23256 12356 23262 12368
rect 24946 12356 24952 12368
rect 23256 12328 24952 12356
rect 23256 12316 23262 12328
rect 24946 12316 24952 12328
rect 25004 12316 25010 12368
rect 22649 12291 22707 12297
rect 22649 12257 22661 12291
rect 22695 12257 22707 12291
rect 22649 12251 22707 12257
rect 23753 12291 23811 12297
rect 23753 12257 23765 12291
rect 23799 12288 23811 12291
rect 23842 12288 23848 12300
rect 23799 12260 23848 12288
rect 23799 12257 23811 12260
rect 23753 12251 23811 12257
rect 23842 12248 23848 12260
rect 23900 12248 23906 12300
rect 24020 12291 24078 12297
rect 24020 12257 24032 12291
rect 24066 12288 24078 12291
rect 24854 12288 24860 12300
rect 24066 12260 24860 12288
rect 24066 12257 24078 12260
rect 24020 12251 24078 12257
rect 24854 12248 24860 12260
rect 24912 12248 24918 12300
rect 21545 12223 21603 12229
rect 21545 12189 21557 12223
rect 21591 12189 21603 12223
rect 21545 12183 21603 12189
rect 22370 12180 22376 12232
rect 22428 12220 22434 12232
rect 22557 12223 22615 12229
rect 22557 12220 22569 12223
rect 22428 12192 22569 12220
rect 22428 12180 22434 12192
rect 22557 12189 22569 12192
rect 22603 12220 22615 12223
rect 23201 12223 23259 12229
rect 23201 12220 23213 12223
rect 22603 12192 23213 12220
rect 22603 12189 22615 12192
rect 22557 12183 22615 12189
rect 23201 12189 23213 12192
rect 23247 12189 23259 12223
rect 23201 12183 23259 12189
rect 21450 12152 21456 12164
rect 21363 12124 21456 12152
rect 21450 12112 21456 12124
rect 21508 12152 21514 12164
rect 22738 12152 22744 12164
rect 21508 12124 22744 12152
rect 21508 12112 21514 12124
rect 22738 12112 22744 12124
rect 22796 12112 22802 12164
rect 5408 12056 6960 12084
rect 5408 12044 5414 12056
rect 7098 12044 7104 12096
rect 7156 12084 7162 12096
rect 7377 12087 7435 12093
rect 7377 12084 7389 12087
rect 7156 12056 7389 12084
rect 7156 12044 7162 12056
rect 7377 12053 7389 12056
rect 7423 12053 7435 12087
rect 8018 12084 8024 12096
rect 7979 12056 8024 12084
rect 7377 12047 7435 12053
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 9766 12044 9772 12096
rect 9824 12084 9830 12096
rect 12986 12084 12992 12096
rect 9824 12056 12992 12084
rect 9824 12044 9830 12056
rect 12986 12044 12992 12056
rect 13044 12044 13050 12096
rect 14090 12044 14096 12096
rect 14148 12044 14154 12096
rect 14458 12044 14464 12096
rect 14516 12084 14522 12096
rect 14645 12087 14703 12093
rect 14645 12084 14657 12087
rect 14516 12056 14657 12084
rect 14516 12044 14522 12056
rect 14645 12053 14657 12056
rect 14691 12053 14703 12087
rect 15930 12084 15936 12096
rect 15891 12056 15936 12084
rect 14645 12047 14703 12053
rect 15930 12044 15936 12056
rect 15988 12044 15994 12096
rect 16666 12044 16672 12096
rect 16724 12084 16730 12096
rect 17402 12084 17408 12096
rect 16724 12056 17408 12084
rect 16724 12044 16730 12056
rect 17402 12044 17408 12056
rect 17460 12044 17466 12096
rect 18966 12084 18972 12096
rect 18927 12056 18972 12084
rect 18966 12044 18972 12056
rect 19024 12044 19030 12096
rect 19153 12087 19211 12093
rect 19153 12053 19165 12087
rect 19199 12084 19211 12087
rect 20165 12087 20223 12093
rect 20165 12084 20177 12087
rect 19199 12056 20177 12084
rect 19199 12053 19211 12056
rect 19153 12047 19211 12053
rect 20165 12053 20177 12056
rect 20211 12084 20223 12087
rect 20438 12084 20444 12096
rect 20211 12056 20444 12084
rect 20211 12053 20223 12056
rect 20165 12047 20223 12053
rect 20438 12044 20444 12056
rect 20496 12044 20502 12096
rect 20901 12087 20959 12093
rect 20901 12053 20913 12087
rect 20947 12084 20959 12087
rect 22002 12084 22008 12096
rect 20947 12056 22008 12084
rect 20947 12053 20959 12056
rect 20901 12047 20959 12053
rect 22002 12044 22008 12056
rect 22060 12044 22066 12096
rect 23661 12087 23719 12093
rect 23661 12053 23673 12087
rect 23707 12084 23719 12087
rect 24762 12084 24768 12096
rect 23707 12056 24768 12084
rect 23707 12053 23719 12056
rect 23661 12047 23719 12053
rect 24762 12044 24768 12056
rect 24820 12044 24826 12096
rect 25498 12044 25504 12096
rect 25556 12084 25562 12096
rect 25685 12087 25743 12093
rect 25685 12084 25697 12087
rect 25556 12056 25697 12084
rect 25556 12044 25562 12056
rect 25685 12053 25697 12056
rect 25731 12053 25743 12087
rect 25685 12047 25743 12053
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1581 11883 1639 11889
rect 1581 11849 1593 11883
rect 1627 11880 1639 11883
rect 3234 11880 3240 11892
rect 1627 11852 3240 11880
rect 1627 11849 1639 11852
rect 1581 11843 1639 11849
rect 3234 11840 3240 11852
rect 3292 11840 3298 11892
rect 5534 11880 5540 11892
rect 5495 11852 5540 11880
rect 5534 11840 5540 11852
rect 5592 11840 5598 11892
rect 9122 11880 9128 11892
rect 8404 11852 9128 11880
rect 2501 11815 2559 11821
rect 2501 11781 2513 11815
rect 2547 11812 2559 11815
rect 3418 11812 3424 11824
rect 2547 11784 3424 11812
rect 2547 11781 2559 11784
rect 2501 11775 2559 11781
rect 3068 11753 3096 11784
rect 3418 11772 3424 11784
rect 3476 11772 3482 11824
rect 8404 11812 8432 11852
rect 9122 11840 9128 11852
rect 9180 11840 9186 11892
rect 9217 11883 9275 11889
rect 9217 11849 9229 11883
rect 9263 11880 9275 11883
rect 9766 11880 9772 11892
rect 9263 11852 9772 11880
rect 9263 11849 9275 11852
rect 9217 11843 9275 11849
rect 9766 11840 9772 11852
rect 9824 11840 9830 11892
rect 10318 11880 10324 11892
rect 10279 11852 10324 11880
rect 10318 11840 10324 11852
rect 10376 11840 10382 11892
rect 10413 11883 10471 11889
rect 10413 11849 10425 11883
rect 10459 11880 10471 11883
rect 10870 11880 10876 11892
rect 10459 11852 10876 11880
rect 10459 11849 10471 11852
rect 10413 11843 10471 11849
rect 10870 11840 10876 11852
rect 10928 11840 10934 11892
rect 11882 11880 11888 11892
rect 11843 11852 11888 11880
rect 11882 11840 11888 11852
rect 11940 11840 11946 11892
rect 13630 11840 13636 11892
rect 13688 11880 13694 11892
rect 16206 11880 16212 11892
rect 13688 11852 16212 11880
rect 13688 11840 13694 11852
rect 16206 11840 16212 11852
rect 16264 11840 16270 11892
rect 16390 11880 16396 11892
rect 16351 11852 16396 11880
rect 16390 11840 16396 11852
rect 16448 11840 16454 11892
rect 17494 11880 17500 11892
rect 17455 11852 17500 11880
rect 17494 11840 17500 11852
rect 17552 11840 17558 11892
rect 22557 11883 22615 11889
rect 22557 11880 22569 11883
rect 21468 11852 22569 11880
rect 5460 11784 8432 11812
rect 13909 11815 13967 11821
rect 3053 11747 3111 11753
rect 3053 11713 3065 11747
rect 3099 11713 3111 11747
rect 3053 11707 3111 11713
rect 3145 11747 3203 11753
rect 3145 11713 3157 11747
rect 3191 11744 3203 11747
rect 3602 11744 3608 11756
rect 3191 11716 3608 11744
rect 3191 11713 3203 11716
rect 3145 11707 3203 11713
rect 3602 11704 3608 11716
rect 3660 11704 3666 11756
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11676 1455 11679
rect 1949 11679 2007 11685
rect 1949 11676 1961 11679
rect 1443 11648 1961 11676
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 1949 11645 1961 11648
rect 1995 11676 2007 11679
rect 2222 11676 2228 11688
rect 1995 11648 2228 11676
rect 1995 11645 2007 11648
rect 1949 11639 2007 11645
rect 2222 11636 2228 11648
rect 2280 11636 2286 11688
rect 4154 11676 4160 11688
rect 4067 11648 4160 11676
rect 4154 11636 4160 11648
rect 4212 11676 4218 11688
rect 5460 11676 5488 11784
rect 13909 11781 13921 11815
rect 13955 11812 13967 11815
rect 14090 11812 14096 11824
rect 13955 11784 14096 11812
rect 13955 11781 13967 11784
rect 13909 11775 13967 11781
rect 14090 11772 14096 11784
rect 14148 11812 14154 11824
rect 16574 11812 16580 11824
rect 14148 11784 16580 11812
rect 14148 11772 14154 11784
rect 16574 11772 16580 11784
rect 16632 11772 16638 11824
rect 21266 11772 21272 11824
rect 21324 11812 21330 11824
rect 21468 11812 21496 11852
rect 22557 11849 22569 11852
rect 22603 11849 22615 11883
rect 22557 11843 22615 11849
rect 23566 11840 23572 11892
rect 23624 11880 23630 11892
rect 23661 11883 23719 11889
rect 23661 11880 23673 11883
rect 23624 11852 23673 11880
rect 23624 11840 23630 11852
rect 23661 11849 23673 11852
rect 23707 11849 23719 11883
rect 23661 11843 23719 11849
rect 25314 11840 25320 11892
rect 25372 11880 25378 11892
rect 25409 11883 25467 11889
rect 25409 11880 25421 11883
rect 25372 11852 25421 11880
rect 25372 11840 25378 11852
rect 25409 11849 25421 11852
rect 25455 11849 25467 11883
rect 25409 11843 25467 11849
rect 21324 11784 21496 11812
rect 21324 11772 21330 11784
rect 21910 11772 21916 11824
rect 21968 11812 21974 11824
rect 23477 11815 23535 11821
rect 21968 11784 22140 11812
rect 21968 11772 21974 11784
rect 6641 11747 6699 11753
rect 6641 11713 6653 11747
rect 6687 11744 6699 11747
rect 7282 11744 7288 11756
rect 6687 11716 7288 11744
rect 6687 11713 6699 11716
rect 6641 11707 6699 11713
rect 7282 11704 7288 11716
rect 7340 11704 7346 11756
rect 7377 11747 7435 11753
rect 7377 11713 7389 11747
rect 7423 11713 7435 11747
rect 7377 11707 7435 11713
rect 8941 11747 8999 11753
rect 8941 11713 8953 11747
rect 8987 11713 8999 11747
rect 8941 11707 8999 11713
rect 4212 11648 5488 11676
rect 4212 11636 4218 11648
rect 7098 11636 7104 11688
rect 7156 11676 7162 11688
rect 7392 11676 7420 11707
rect 8956 11676 8984 11707
rect 9674 11704 9680 11756
rect 9732 11744 9738 11756
rect 10689 11747 10747 11753
rect 10689 11744 10701 11747
rect 9732 11716 10701 11744
rect 9732 11704 9738 11716
rect 10689 11713 10701 11716
rect 10735 11713 10747 11747
rect 10689 11707 10747 11713
rect 9401 11679 9459 11685
rect 9401 11676 9413 11679
rect 7156 11648 9413 11676
rect 7156 11636 7162 11648
rect 9401 11645 9413 11648
rect 9447 11676 9459 11679
rect 9490 11676 9496 11688
rect 9447 11648 9496 11676
rect 9447 11645 9459 11648
rect 9401 11639 9459 11645
rect 9490 11636 9496 11648
rect 9548 11636 9554 11688
rect 9766 11636 9772 11688
rect 9824 11676 9830 11688
rect 10413 11679 10471 11685
rect 10413 11676 10425 11679
rect 9824 11648 10425 11676
rect 9824 11636 9830 11648
rect 10413 11645 10425 11648
rect 10459 11645 10471 11679
rect 10704 11676 10732 11707
rect 10870 11704 10876 11756
rect 10928 11744 10934 11756
rect 11333 11747 11391 11753
rect 11333 11744 11345 11747
rect 10928 11716 11345 11744
rect 10928 11704 10934 11716
rect 11333 11713 11345 11716
rect 11379 11713 11391 11747
rect 11333 11707 11391 11713
rect 15930 11704 15936 11756
rect 15988 11744 15994 11756
rect 16850 11744 16856 11756
rect 15988 11716 16856 11744
rect 15988 11704 15994 11716
rect 16850 11704 16856 11716
rect 16908 11744 16914 11756
rect 16945 11747 17003 11753
rect 16945 11744 16957 11747
rect 16908 11716 16957 11744
rect 16908 11704 16914 11716
rect 16945 11713 16957 11716
rect 16991 11744 17003 11747
rect 18598 11744 18604 11756
rect 16991 11716 18604 11744
rect 16991 11713 17003 11716
rect 16945 11707 17003 11713
rect 18598 11704 18604 11716
rect 18656 11704 18662 11756
rect 20254 11744 20260 11756
rect 18708 11716 20260 11744
rect 11149 11679 11207 11685
rect 11149 11676 11161 11679
rect 10704 11648 11161 11676
rect 10413 11639 10471 11645
rect 11149 11645 11161 11648
rect 11195 11676 11207 11679
rect 11606 11676 11612 11688
rect 11195 11648 11612 11676
rect 11195 11645 11207 11648
rect 11149 11639 11207 11645
rect 11606 11636 11612 11648
rect 11664 11636 11670 11688
rect 11882 11636 11888 11688
rect 11940 11676 11946 11688
rect 12066 11676 12072 11688
rect 11940 11648 12072 11676
rect 11940 11636 11946 11648
rect 12066 11636 12072 11648
rect 12124 11636 12130 11688
rect 12250 11636 12256 11688
rect 12308 11676 12314 11688
rect 12529 11679 12587 11685
rect 12529 11676 12541 11679
rect 12308 11648 12541 11676
rect 12308 11636 12314 11648
rect 12529 11645 12541 11648
rect 12575 11676 12587 11679
rect 13906 11676 13912 11688
rect 12575 11648 13912 11676
rect 12575 11645 12587 11648
rect 12529 11639 12587 11645
rect 13906 11636 13912 11648
rect 13964 11676 13970 11688
rect 14550 11676 14556 11688
rect 13964 11648 14556 11676
rect 13964 11636 13970 11648
rect 14550 11636 14556 11648
rect 14608 11636 14614 11688
rect 15289 11679 15347 11685
rect 15289 11645 15301 11679
rect 15335 11676 15347 11679
rect 15335 11648 15369 11676
rect 15335 11645 15347 11648
rect 15289 11639 15347 11645
rect 3878 11568 3884 11620
rect 3936 11608 3942 11620
rect 4424 11611 4482 11617
rect 4424 11608 4436 11611
rect 3936 11580 4436 11608
rect 3936 11568 3942 11580
rect 4424 11577 4436 11580
rect 4470 11608 4482 11611
rect 5442 11608 5448 11620
rect 4470 11580 5448 11608
rect 4470 11577 4482 11580
rect 4424 11571 4482 11577
rect 5442 11568 5448 11580
rect 5500 11568 5506 11620
rect 7193 11611 7251 11617
rect 7193 11608 7205 11611
rect 6196 11580 7205 11608
rect 6196 11552 6224 11580
rect 7193 11577 7205 11580
rect 7239 11608 7251 11611
rect 8110 11608 8116 11620
rect 7239 11580 8116 11608
rect 7239 11577 7251 11580
rect 7193 11571 7251 11577
rect 8110 11568 8116 11580
rect 8168 11568 8174 11620
rect 8757 11611 8815 11617
rect 8757 11608 8769 11611
rect 8220 11580 8769 11608
rect 8220 11552 8248 11580
rect 8757 11577 8769 11580
rect 8803 11577 8815 11611
rect 8757 11571 8815 11577
rect 8849 11611 8907 11617
rect 8849 11577 8861 11611
rect 8895 11608 8907 11611
rect 9217 11611 9275 11617
rect 9217 11608 9229 11611
rect 8895 11580 9229 11608
rect 8895 11577 8907 11580
rect 8849 11571 8907 11577
rect 9217 11577 9229 11580
rect 9263 11577 9275 11611
rect 9217 11571 9275 11577
rect 9953 11611 10011 11617
rect 9953 11577 9965 11611
rect 9999 11608 10011 11611
rect 10870 11608 10876 11620
rect 9999 11580 10876 11608
rect 9999 11577 10011 11580
rect 9953 11571 10011 11577
rect 2590 11540 2596 11552
rect 2551 11512 2596 11540
rect 2590 11500 2596 11512
rect 2648 11500 2654 11552
rect 2961 11543 3019 11549
rect 2961 11509 2973 11543
rect 3007 11540 3019 11543
rect 3418 11540 3424 11552
rect 3007 11512 3424 11540
rect 3007 11509 3019 11512
rect 2961 11503 3019 11509
rect 3418 11500 3424 11512
rect 3476 11540 3482 11552
rect 3605 11543 3663 11549
rect 3605 11540 3617 11543
rect 3476 11512 3617 11540
rect 3476 11500 3482 11512
rect 3605 11509 3617 11512
rect 3651 11509 3663 11543
rect 3605 11503 3663 11509
rect 4065 11543 4123 11549
rect 4065 11509 4077 11543
rect 4111 11540 4123 11543
rect 4246 11540 4252 11552
rect 4111 11512 4252 11540
rect 4111 11509 4123 11512
rect 4065 11503 4123 11509
rect 4246 11500 4252 11512
rect 4304 11500 4310 11552
rect 6178 11540 6184 11552
rect 6139 11512 6184 11540
rect 6178 11500 6184 11512
rect 6236 11500 6242 11552
rect 6822 11540 6828 11552
rect 6783 11512 6828 11540
rect 6822 11500 6828 11512
rect 6880 11500 6886 11552
rect 7006 11500 7012 11552
rect 7064 11540 7070 11552
rect 7650 11540 7656 11552
rect 7064 11512 7656 11540
rect 7064 11500 7070 11512
rect 7650 11500 7656 11512
rect 7708 11500 7714 11552
rect 7834 11540 7840 11552
rect 7795 11512 7840 11540
rect 7834 11500 7840 11512
rect 7892 11500 7898 11552
rect 8202 11540 8208 11552
rect 8163 11512 8208 11540
rect 8202 11500 8208 11512
rect 8260 11500 8266 11552
rect 8294 11500 8300 11552
rect 8352 11540 8358 11552
rect 8389 11543 8447 11549
rect 8389 11540 8401 11543
rect 8352 11512 8401 11540
rect 8352 11500 8358 11512
rect 8389 11509 8401 11512
rect 8435 11509 8447 11543
rect 8389 11503 8447 11509
rect 8478 11500 8484 11552
rect 8536 11540 8542 11552
rect 8864 11540 8892 11571
rect 10870 11568 10876 11580
rect 10928 11568 10934 11620
rect 11054 11568 11060 11620
rect 11112 11608 11118 11620
rect 11241 11611 11299 11617
rect 11241 11608 11253 11611
rect 11112 11580 11253 11608
rect 11112 11568 11118 11580
rect 11241 11577 11253 11580
rect 11287 11577 11299 11611
rect 12158 11608 12164 11620
rect 11241 11571 11299 11577
rect 11348 11580 12164 11608
rect 10778 11540 10784 11552
rect 8536 11512 8892 11540
rect 10739 11512 10784 11540
rect 8536 11500 8542 11512
rect 10778 11500 10784 11512
rect 10836 11500 10842 11552
rect 11146 11500 11152 11552
rect 11204 11540 11210 11552
rect 11348 11540 11376 11580
rect 12158 11568 12164 11580
rect 12216 11568 12222 11620
rect 12796 11611 12854 11617
rect 12796 11577 12808 11611
rect 12842 11608 12854 11611
rect 13170 11608 13176 11620
rect 12842 11580 13176 11608
rect 12842 11577 12854 11580
rect 12796 11571 12854 11577
rect 13170 11568 13176 11580
rect 13228 11568 13234 11620
rect 15197 11611 15255 11617
rect 15197 11577 15209 11611
rect 15243 11608 15255 11611
rect 15304 11608 15332 11639
rect 16758 11636 16764 11688
rect 16816 11676 16822 11688
rect 17773 11679 17831 11685
rect 17773 11676 17785 11679
rect 16816 11648 17785 11676
rect 16816 11636 16822 11648
rect 17773 11645 17785 11648
rect 17819 11676 17831 11679
rect 18509 11679 18567 11685
rect 18509 11676 18521 11679
rect 17819 11648 18521 11676
rect 17819 11645 17831 11648
rect 17773 11639 17831 11645
rect 18509 11645 18521 11648
rect 18555 11676 18567 11679
rect 18708 11676 18736 11716
rect 20254 11704 20260 11716
rect 20312 11704 20318 11756
rect 20438 11744 20444 11756
rect 20399 11716 20444 11744
rect 20438 11704 20444 11716
rect 20496 11704 20502 11756
rect 20533 11747 20591 11753
rect 20533 11713 20545 11747
rect 20579 11713 20591 11747
rect 21450 11744 21456 11756
rect 21411 11716 21456 11744
rect 20533 11707 20591 11713
rect 18555 11648 18736 11676
rect 19889 11679 19947 11685
rect 18555 11645 18567 11648
rect 18509 11639 18567 11645
rect 19889 11645 19901 11679
rect 19935 11676 19947 11679
rect 19978 11676 19984 11688
rect 19935 11648 19984 11676
rect 19935 11645 19947 11648
rect 19889 11639 19947 11645
rect 19978 11636 19984 11648
rect 20036 11676 20042 11688
rect 20548 11676 20576 11707
rect 21450 11704 21456 11716
rect 21508 11704 21514 11756
rect 22002 11744 22008 11756
rect 21963 11716 22008 11744
rect 22002 11704 22008 11716
rect 22060 11704 22066 11756
rect 22112 11753 22140 11784
rect 23477 11781 23489 11815
rect 23523 11812 23535 11815
rect 23750 11812 23756 11824
rect 23523 11784 23756 11812
rect 23523 11781 23535 11784
rect 23477 11775 23535 11781
rect 23750 11772 23756 11784
rect 23808 11812 23814 11824
rect 23808 11784 24256 11812
rect 23808 11772 23814 11784
rect 24228 11753 24256 11784
rect 22097 11747 22155 11753
rect 22097 11713 22109 11747
rect 22143 11713 22155 11747
rect 22097 11707 22155 11713
rect 24213 11747 24271 11753
rect 24213 11713 24225 11747
rect 24259 11713 24271 11747
rect 24213 11707 24271 11713
rect 20036 11648 20576 11676
rect 20036 11636 20042 11648
rect 20898 11636 20904 11688
rect 20956 11676 20962 11688
rect 21913 11679 21971 11685
rect 21913 11676 21925 11679
rect 20956 11648 21925 11676
rect 20956 11636 20962 11648
rect 21913 11645 21925 11648
rect 21959 11645 21971 11679
rect 21913 11639 21971 11645
rect 22462 11636 22468 11688
rect 22520 11676 22526 11688
rect 23109 11679 23167 11685
rect 23109 11676 23121 11679
rect 22520 11648 23121 11676
rect 22520 11636 22526 11648
rect 23109 11645 23121 11648
rect 23155 11676 23167 11679
rect 24854 11676 24860 11688
rect 23155 11648 24860 11676
rect 23155 11645 23167 11648
rect 23109 11639 23167 11645
rect 24854 11636 24860 11648
rect 24912 11636 24918 11688
rect 25222 11676 25228 11688
rect 25183 11648 25228 11676
rect 25222 11636 25228 11648
rect 25280 11676 25286 11688
rect 25777 11679 25835 11685
rect 25777 11676 25789 11679
rect 25280 11648 25789 11676
rect 25280 11636 25286 11648
rect 25777 11645 25789 11648
rect 25823 11645 25835 11679
rect 25777 11639 25835 11645
rect 15654 11608 15660 11620
rect 15243 11580 15660 11608
rect 15243 11577 15255 11580
rect 15197 11571 15255 11577
rect 15654 11568 15660 11580
rect 15712 11568 15718 11620
rect 15933 11611 15991 11617
rect 15933 11608 15945 11611
rect 15764 11580 15945 11608
rect 11204 11512 11376 11540
rect 14553 11543 14611 11549
rect 11204 11500 11210 11512
rect 14553 11509 14565 11543
rect 14599 11540 14611 11543
rect 14734 11540 14740 11552
rect 14599 11512 14740 11540
rect 14599 11509 14611 11512
rect 14553 11503 14611 11509
rect 14734 11500 14740 11512
rect 14792 11500 14798 11552
rect 15470 11540 15476 11552
rect 15431 11512 15476 11540
rect 15470 11500 15476 11512
rect 15528 11500 15534 11552
rect 15562 11500 15568 11552
rect 15620 11540 15626 11552
rect 15764 11540 15792 11580
rect 15933 11577 15945 11580
rect 15979 11608 15991 11611
rect 16666 11608 16672 11620
rect 15979 11580 16672 11608
rect 15979 11577 15991 11580
rect 15933 11571 15991 11577
rect 16666 11568 16672 11580
rect 16724 11608 16730 11620
rect 16853 11611 16911 11617
rect 16853 11608 16865 11611
rect 16724 11580 16865 11608
rect 16724 11568 16730 11580
rect 16853 11577 16865 11580
rect 16899 11577 16911 11611
rect 17218 11608 17224 11620
rect 16853 11571 16911 11577
rect 16960 11580 17224 11608
rect 15620 11512 15792 11540
rect 15620 11500 15626 11512
rect 15838 11500 15844 11552
rect 15896 11540 15902 11552
rect 16301 11543 16359 11549
rect 16301 11540 16313 11543
rect 15896 11512 16313 11540
rect 15896 11500 15902 11512
rect 16301 11509 16313 11512
rect 16347 11540 16359 11543
rect 16761 11543 16819 11549
rect 16761 11540 16773 11543
rect 16347 11512 16773 11540
rect 16347 11509 16359 11512
rect 16301 11503 16359 11509
rect 16761 11509 16773 11512
rect 16807 11540 16819 11543
rect 16960 11540 16988 11580
rect 17218 11568 17224 11580
rect 17276 11568 17282 11620
rect 17310 11568 17316 11620
rect 17368 11608 17374 11620
rect 17494 11608 17500 11620
rect 17368 11580 17500 11608
rect 17368 11568 17374 11580
rect 17494 11568 17500 11580
rect 17552 11568 17558 11620
rect 17954 11568 17960 11620
rect 18012 11608 18018 11620
rect 18417 11611 18475 11617
rect 18417 11608 18429 11611
rect 18012 11580 18429 11608
rect 18012 11568 18018 11580
rect 18417 11577 18429 11580
rect 18463 11577 18475 11611
rect 18417 11571 18475 11577
rect 19245 11611 19303 11617
rect 19245 11577 19257 11611
rect 19291 11608 19303 11611
rect 20070 11608 20076 11620
rect 19291 11580 20076 11608
rect 19291 11577 19303 11580
rect 19245 11571 19303 11577
rect 20070 11568 20076 11580
rect 20128 11568 20134 11620
rect 20349 11611 20407 11617
rect 20349 11577 20361 11611
rect 20395 11608 20407 11611
rect 20622 11608 20628 11620
rect 20395 11580 20628 11608
rect 20395 11577 20407 11580
rect 20349 11571 20407 11577
rect 20622 11568 20628 11580
rect 20680 11608 20686 11620
rect 20680 11580 21588 11608
rect 20680 11568 20686 11580
rect 18046 11540 18052 11552
rect 16807 11512 16988 11540
rect 18007 11512 18052 11540
rect 16807 11509 16819 11512
rect 16761 11503 16819 11509
rect 18046 11500 18052 11512
rect 18104 11500 18110 11552
rect 19981 11543 20039 11549
rect 19981 11509 19993 11543
rect 20027 11540 20039 11543
rect 20806 11540 20812 11552
rect 20027 11512 20812 11540
rect 20027 11509 20039 11512
rect 19981 11503 20039 11509
rect 20806 11500 20812 11512
rect 20864 11500 20870 11552
rect 21085 11543 21143 11549
rect 21085 11509 21097 11543
rect 21131 11540 21143 11543
rect 21174 11540 21180 11552
rect 21131 11512 21180 11540
rect 21131 11509 21143 11512
rect 21085 11503 21143 11509
rect 21174 11500 21180 11512
rect 21232 11500 21238 11552
rect 21560 11549 21588 11580
rect 23750 11568 23756 11620
rect 23808 11608 23814 11620
rect 24121 11611 24179 11617
rect 24121 11608 24133 11611
rect 23808 11580 24133 11608
rect 23808 11568 23814 11580
rect 24121 11577 24133 11580
rect 24167 11608 24179 11611
rect 24673 11611 24731 11617
rect 24673 11608 24685 11611
rect 24167 11580 24685 11608
rect 24167 11577 24179 11580
rect 24121 11571 24179 11577
rect 24673 11577 24685 11580
rect 24719 11577 24731 11611
rect 24673 11571 24731 11577
rect 21545 11543 21603 11549
rect 21545 11509 21557 11543
rect 21591 11509 21603 11543
rect 21545 11503 21603 11509
rect 23566 11500 23572 11552
rect 23624 11540 23630 11552
rect 24029 11543 24087 11549
rect 24029 11540 24041 11543
rect 23624 11512 24041 11540
rect 23624 11500 23630 11512
rect 24029 11509 24041 11512
rect 24075 11540 24087 11543
rect 25041 11543 25099 11549
rect 25041 11540 25053 11543
rect 24075 11512 25053 11540
rect 24075 11509 24087 11512
rect 24029 11503 24087 11509
rect 25041 11509 25053 11512
rect 25087 11509 25099 11543
rect 25041 11503 25099 11509
rect 25498 11500 25504 11552
rect 25556 11540 25562 11552
rect 26145 11543 26203 11549
rect 26145 11540 26157 11543
rect 25556 11512 26157 11540
rect 25556 11500 25562 11512
rect 26145 11509 26157 11512
rect 26191 11509 26203 11543
rect 26145 11503 26203 11509
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 2409 11339 2467 11345
rect 2409 11305 2421 11339
rect 2455 11336 2467 11339
rect 2682 11336 2688 11348
rect 2455 11308 2688 11336
rect 2455 11305 2467 11308
rect 2409 11299 2467 11305
rect 2682 11296 2688 11308
rect 2740 11296 2746 11348
rect 2774 11296 2780 11348
rect 2832 11336 2838 11348
rect 2869 11339 2927 11345
rect 2869 11336 2881 11339
rect 2832 11308 2881 11336
rect 2832 11296 2838 11308
rect 2869 11305 2881 11308
rect 2915 11336 2927 11339
rect 3326 11336 3332 11348
rect 2915 11308 3332 11336
rect 2915 11305 2927 11308
rect 2869 11299 2927 11305
rect 3326 11296 3332 11308
rect 3384 11296 3390 11348
rect 3878 11336 3884 11348
rect 3839 11308 3884 11336
rect 3878 11296 3884 11308
rect 3936 11296 3942 11348
rect 5534 11296 5540 11348
rect 5592 11336 5598 11348
rect 5997 11339 6055 11345
rect 5997 11336 6009 11339
rect 5592 11308 6009 11336
rect 5592 11296 5598 11308
rect 5997 11305 6009 11308
rect 6043 11305 6055 11339
rect 5997 11299 6055 11305
rect 6362 11296 6368 11348
rect 6420 11336 6426 11348
rect 6549 11339 6607 11345
rect 6549 11336 6561 11339
rect 6420 11308 6561 11336
rect 6420 11296 6426 11308
rect 6549 11305 6561 11308
rect 6595 11305 6607 11339
rect 7742 11336 7748 11348
rect 7703 11308 7748 11336
rect 6549 11299 6607 11305
rect 7742 11296 7748 11308
rect 7800 11296 7806 11348
rect 8570 11336 8576 11348
rect 8531 11308 8576 11336
rect 8570 11296 8576 11308
rect 8628 11296 8634 11348
rect 9306 11296 9312 11348
rect 9364 11336 9370 11348
rect 9401 11339 9459 11345
rect 9401 11336 9413 11339
rect 9364 11308 9413 11336
rect 9364 11296 9370 11308
rect 9401 11305 9413 11308
rect 9447 11305 9459 11339
rect 9401 11299 9459 11305
rect 10689 11339 10747 11345
rect 10689 11305 10701 11339
rect 10735 11336 10747 11339
rect 11054 11336 11060 11348
rect 10735 11308 11060 11336
rect 10735 11305 10747 11308
rect 10689 11299 10747 11305
rect 11054 11296 11060 11308
rect 11112 11336 11118 11348
rect 11514 11336 11520 11348
rect 11112 11308 11520 11336
rect 11112 11296 11118 11308
rect 11514 11296 11520 11308
rect 11572 11296 11578 11348
rect 12434 11296 12440 11348
rect 12492 11336 12498 11348
rect 12802 11336 12808 11348
rect 12492 11308 12808 11336
rect 12492 11296 12498 11308
rect 12802 11296 12808 11308
rect 12860 11296 12866 11348
rect 13170 11336 13176 11348
rect 13131 11308 13176 11336
rect 13170 11296 13176 11308
rect 13228 11296 13234 11348
rect 16482 11296 16488 11348
rect 16540 11336 16546 11348
rect 17037 11339 17095 11345
rect 17037 11336 17049 11339
rect 16540 11308 17049 11336
rect 16540 11296 16546 11308
rect 17037 11305 17049 11308
rect 17083 11305 17095 11339
rect 17037 11299 17095 11305
rect 18230 11296 18236 11348
rect 18288 11336 18294 11348
rect 20162 11336 20168 11348
rect 18288 11308 20168 11336
rect 18288 11296 18294 11308
rect 20162 11296 20168 11308
rect 20220 11296 20226 11348
rect 20349 11339 20407 11345
rect 20349 11305 20361 11339
rect 20395 11336 20407 11339
rect 20622 11336 20628 11348
rect 20395 11308 20628 11336
rect 20395 11305 20407 11308
rect 20349 11299 20407 11305
rect 20622 11296 20628 11308
rect 20680 11296 20686 11348
rect 21910 11336 21916 11348
rect 21871 11308 21916 11336
rect 21910 11296 21916 11308
rect 21968 11296 21974 11348
rect 22002 11296 22008 11348
rect 22060 11336 22066 11348
rect 22281 11339 22339 11345
rect 22281 11336 22293 11339
rect 22060 11308 22293 11336
rect 22060 11296 22066 11308
rect 22281 11305 22293 11308
rect 22327 11305 22339 11339
rect 22646 11336 22652 11348
rect 22607 11308 22652 11336
rect 22281 11299 22339 11305
rect 22646 11296 22652 11308
rect 22704 11296 22710 11348
rect 23109 11339 23167 11345
rect 23109 11305 23121 11339
rect 23155 11336 23167 11339
rect 23198 11336 23204 11348
rect 23155 11308 23204 11336
rect 23155 11305 23167 11308
rect 23109 11299 23167 11305
rect 23198 11296 23204 11308
rect 23256 11296 23262 11348
rect 23842 11336 23848 11348
rect 23676 11308 23848 11336
rect 2317 11271 2375 11277
rect 2317 11237 2329 11271
rect 2363 11268 2375 11271
rect 3050 11268 3056 11280
rect 2363 11240 3056 11268
rect 2363 11237 2375 11240
rect 2317 11231 2375 11237
rect 3050 11228 3056 11240
rect 3108 11228 3114 11280
rect 3513 11271 3571 11277
rect 3513 11237 3525 11271
rect 3559 11268 3571 11271
rect 3602 11268 3608 11280
rect 3559 11240 3608 11268
rect 3559 11237 3571 11240
rect 3513 11231 3571 11237
rect 3602 11228 3608 11240
rect 3660 11268 3666 11280
rect 5350 11268 5356 11280
rect 3660 11240 5356 11268
rect 3660 11228 3666 11240
rect 5350 11228 5356 11240
rect 5408 11228 5414 11280
rect 6917 11271 6975 11277
rect 6917 11237 6929 11271
rect 6963 11268 6975 11271
rect 7006 11268 7012 11280
rect 6963 11240 7012 11268
rect 6963 11237 6975 11240
rect 6917 11231 6975 11237
rect 7006 11228 7012 11240
rect 7064 11228 7070 11280
rect 8478 11268 8484 11280
rect 8439 11240 8484 11268
rect 8478 11228 8484 11240
rect 8536 11228 8542 11280
rect 12250 11268 12256 11280
rect 11808 11240 12256 11268
rect 2777 11203 2835 11209
rect 2777 11169 2789 11203
rect 2823 11200 2835 11203
rect 3142 11200 3148 11212
rect 2823 11172 3148 11200
rect 2823 11169 2835 11172
rect 2777 11163 2835 11169
rect 3142 11160 3148 11172
rect 3200 11200 3206 11212
rect 3694 11200 3700 11212
rect 3200 11172 3700 11200
rect 3200 11160 3206 11172
rect 3694 11160 3700 11172
rect 3752 11160 3758 11212
rect 4065 11203 4123 11209
rect 4065 11169 4077 11203
rect 4111 11200 4123 11203
rect 4154 11200 4160 11212
rect 4111 11172 4160 11200
rect 4111 11169 4123 11172
rect 4065 11163 4123 11169
rect 1394 11132 1400 11144
rect 1355 11104 1400 11132
rect 1394 11092 1400 11104
rect 1452 11092 1458 11144
rect 2498 11092 2504 11144
rect 2556 11132 2562 11144
rect 3053 11135 3111 11141
rect 3053 11132 3065 11135
rect 2556 11104 3065 11132
rect 2556 11092 2562 11104
rect 3053 11101 3065 11104
rect 3099 11132 3111 11135
rect 3878 11132 3884 11144
rect 3099 11104 3884 11132
rect 3099 11101 3111 11104
rect 3053 11095 3111 11101
rect 3878 11092 3884 11104
rect 3936 11092 3942 11144
rect 1949 11067 2007 11073
rect 1949 11033 1961 11067
rect 1995 11064 2007 11067
rect 2682 11064 2688 11076
rect 1995 11036 2688 11064
rect 1995 11033 2007 11036
rect 1949 11027 2007 11033
rect 2682 11024 2688 11036
rect 2740 11024 2746 11076
rect 2866 11024 2872 11076
rect 2924 11064 2930 11076
rect 3326 11064 3332 11076
rect 2924 11036 3332 11064
rect 2924 11024 2930 11036
rect 3326 11024 3332 11036
rect 3384 11024 3390 11076
rect 3694 11024 3700 11076
rect 3752 11064 3758 11076
rect 4080 11064 4108 11163
rect 4154 11160 4160 11172
rect 4212 11160 4218 11212
rect 4332 11203 4390 11209
rect 4332 11169 4344 11203
rect 4378 11200 4390 11203
rect 4706 11200 4712 11212
rect 4378 11172 4712 11200
rect 4378 11169 4390 11172
rect 4332 11163 4390 11169
rect 4706 11160 4712 11172
rect 4764 11160 4770 11212
rect 9033 11203 9091 11209
rect 9033 11200 9045 11203
rect 7024 11172 9045 11200
rect 6638 11092 6644 11144
rect 6696 11132 6702 11144
rect 7024 11141 7052 11172
rect 9033 11169 9045 11172
rect 9079 11169 9091 11203
rect 10594 11200 10600 11212
rect 10555 11172 10600 11200
rect 9033 11163 9091 11169
rect 10594 11160 10600 11172
rect 10652 11160 10658 11212
rect 11514 11160 11520 11212
rect 11572 11200 11578 11212
rect 11808 11209 11836 11240
rect 12250 11228 12256 11240
rect 12308 11228 12314 11280
rect 13998 11268 14004 11280
rect 13959 11240 14004 11268
rect 13998 11228 14004 11240
rect 14056 11228 14062 11280
rect 14550 11228 14556 11280
rect 14608 11268 14614 11280
rect 18598 11277 18604 11280
rect 18592 11268 18604 11277
rect 14608 11240 17724 11268
rect 18559 11240 18604 11268
rect 14608 11228 14614 11240
rect 12066 11209 12072 11212
rect 11793 11203 11851 11209
rect 11793 11200 11805 11203
rect 11572 11172 11805 11200
rect 11572 11160 11578 11172
rect 11793 11169 11805 11172
rect 11839 11169 11851 11203
rect 12060 11200 12072 11209
rect 12027 11172 12072 11200
rect 11793 11163 11851 11169
rect 12060 11163 12072 11172
rect 12066 11160 12072 11163
rect 12124 11160 12130 11212
rect 15562 11160 15568 11212
rect 15620 11200 15626 11212
rect 15924 11203 15982 11209
rect 15924 11200 15936 11203
rect 15620 11172 15936 11200
rect 15620 11160 15626 11172
rect 15924 11169 15936 11172
rect 15970 11200 15982 11203
rect 17402 11200 17408 11212
rect 15970 11172 17408 11200
rect 15970 11169 15982 11172
rect 15924 11163 15982 11169
rect 17402 11160 17408 11172
rect 17460 11160 17466 11212
rect 17696 11209 17724 11240
rect 18592 11231 18604 11240
rect 18598 11228 18604 11231
rect 18656 11228 18662 11280
rect 20438 11228 20444 11280
rect 20496 11268 20502 11280
rect 20714 11268 20720 11280
rect 20496 11240 20720 11268
rect 20496 11228 20502 11240
rect 20714 11228 20720 11240
rect 20772 11228 20778 11280
rect 17681 11203 17739 11209
rect 17681 11169 17693 11203
rect 17727 11200 17739 11203
rect 18874 11200 18880 11212
rect 17727 11172 18880 11200
rect 17727 11169 17739 11172
rect 17681 11163 17739 11169
rect 18874 11160 18880 11172
rect 18932 11160 18938 11212
rect 19886 11160 19892 11212
rect 19944 11200 19950 11212
rect 21269 11203 21327 11209
rect 21269 11200 21281 11203
rect 19944 11172 21281 11200
rect 19944 11160 19950 11172
rect 21269 11169 21281 11172
rect 21315 11169 21327 11203
rect 21269 11163 21327 11169
rect 21358 11160 21364 11212
rect 21416 11200 21422 11212
rect 21416 11172 22324 11200
rect 21416 11160 21422 11172
rect 7009 11135 7067 11141
rect 7009 11132 7021 11135
rect 6696 11104 7021 11132
rect 6696 11092 6702 11104
rect 7009 11101 7021 11104
rect 7055 11101 7067 11135
rect 7009 11095 7067 11101
rect 7101 11135 7159 11141
rect 7101 11101 7113 11135
rect 7147 11101 7159 11135
rect 7101 11095 7159 11101
rect 5442 11064 5448 11076
rect 3752 11036 4108 11064
rect 5355 11036 5448 11064
rect 3752 11024 3758 11036
rect 5442 11024 5448 11036
rect 5500 11064 5506 11076
rect 6270 11064 6276 11076
rect 5500 11036 6276 11064
rect 5500 11024 5506 11036
rect 6270 11024 6276 11036
rect 6328 11064 6334 11076
rect 7116 11064 7144 11095
rect 7834 11092 7840 11144
rect 7892 11132 7898 11144
rect 8478 11132 8484 11144
rect 7892 11104 8484 11132
rect 7892 11092 7898 11104
rect 8478 11092 8484 11104
rect 8536 11092 8542 11144
rect 8662 11092 8668 11144
rect 8720 11092 8726 11144
rect 10870 11132 10876 11144
rect 10831 11104 10876 11132
rect 10870 11092 10876 11104
rect 10928 11132 10934 11144
rect 11330 11132 11336 11144
rect 10928 11104 11336 11132
rect 10928 11092 10934 11104
rect 11330 11092 11336 11104
rect 11388 11092 11394 11144
rect 12986 11092 12992 11144
rect 13044 11132 13050 11144
rect 15286 11132 15292 11144
rect 13044 11104 15292 11132
rect 13044 11092 13050 11104
rect 15286 11092 15292 11104
rect 15344 11092 15350 11144
rect 15378 11092 15384 11144
rect 15436 11132 15442 11144
rect 15657 11135 15715 11141
rect 15657 11132 15669 11135
rect 15436 11104 15669 11132
rect 15436 11092 15442 11104
rect 15657 11101 15669 11104
rect 15703 11101 15715 11135
rect 15657 11095 15715 11101
rect 18230 11092 18236 11144
rect 18288 11132 18294 11144
rect 18325 11135 18383 11141
rect 18325 11132 18337 11135
rect 18288 11104 18337 11132
rect 18288 11092 18294 11104
rect 18325 11101 18337 11104
rect 18371 11101 18383 11135
rect 20070 11132 20076 11144
rect 18325 11095 18383 11101
rect 19720 11104 20076 11132
rect 6328 11036 7144 11064
rect 8113 11067 8171 11073
rect 6328 11024 6334 11036
rect 8113 11033 8125 11067
rect 8159 11064 8171 11067
rect 8680 11064 8708 11092
rect 9398 11064 9404 11076
rect 8159 11036 9404 11064
rect 8159 11033 8171 11036
rect 8113 11027 8171 11033
rect 9398 11024 9404 11036
rect 9456 11024 9462 11076
rect 9861 11067 9919 11073
rect 9861 11064 9873 11067
rect 9600 11036 9873 11064
rect 6362 10996 6368 11008
rect 6323 10968 6368 10996
rect 6362 10956 6368 10968
rect 6420 10956 6426 11008
rect 8662 10956 8668 11008
rect 8720 10996 8726 11008
rect 9600 10996 9628 11036
rect 9861 11033 9873 11036
rect 9907 11033 9919 11067
rect 10226 11064 10232 11076
rect 10187 11036 10232 11064
rect 9861 11027 9919 11033
rect 10226 11024 10232 11036
rect 10284 11024 10290 11076
rect 11238 11064 11244 11076
rect 11199 11036 11244 11064
rect 11238 11024 11244 11036
rect 11296 11024 11302 11076
rect 15473 11067 15531 11073
rect 15473 11064 15485 11067
rect 14752 11036 15485 11064
rect 8720 10968 9628 10996
rect 11701 10999 11759 11005
rect 8720 10956 8726 10968
rect 11701 10965 11713 10999
rect 11747 10996 11759 10999
rect 12158 10996 12164 11008
rect 11747 10968 12164 10996
rect 11747 10965 11759 10968
rect 11701 10959 11759 10965
rect 12158 10956 12164 10968
rect 12216 10996 12222 11008
rect 13170 10996 13176 11008
rect 12216 10968 13176 10996
rect 12216 10956 12222 10968
rect 13170 10956 13176 10968
rect 13228 10956 13234 11008
rect 14182 10956 14188 11008
rect 14240 10996 14246 11008
rect 14752 11005 14780 11036
rect 15473 11033 15485 11036
rect 15519 11033 15531 11067
rect 15473 11027 15531 11033
rect 17954 11024 17960 11076
rect 18012 11064 18018 11076
rect 19720 11073 19748 11104
rect 20070 11092 20076 11104
rect 20128 11132 20134 11144
rect 21545 11135 21603 11141
rect 21545 11132 21557 11135
rect 20128 11104 21557 11132
rect 20128 11092 20134 11104
rect 21545 11101 21557 11104
rect 21591 11132 21603 11135
rect 21910 11132 21916 11144
rect 21591 11104 21916 11132
rect 21591 11101 21603 11104
rect 21545 11095 21603 11101
rect 21910 11092 21916 11104
rect 21968 11092 21974 11144
rect 22296 11132 22324 11172
rect 22370 11160 22376 11212
rect 22428 11200 22434 11212
rect 23676 11209 23704 11308
rect 23842 11296 23848 11308
rect 23900 11336 23906 11348
rect 24026 11336 24032 11348
rect 23900 11308 24032 11336
rect 23900 11296 23906 11308
rect 24026 11296 24032 11308
rect 24084 11296 24090 11348
rect 24854 11296 24860 11348
rect 24912 11336 24918 11348
rect 25041 11339 25099 11345
rect 25041 11336 25053 11339
rect 24912 11308 25053 11336
rect 24912 11296 24918 11308
rect 25041 11305 25053 11308
rect 25087 11305 25099 11339
rect 25041 11299 25099 11305
rect 25685 11339 25743 11345
rect 25685 11305 25697 11339
rect 25731 11336 25743 11339
rect 26053 11339 26111 11345
rect 26053 11336 26065 11339
rect 25731 11308 26065 11336
rect 25731 11305 25743 11308
rect 25685 11299 25743 11305
rect 26053 11305 26065 11308
rect 26099 11336 26111 11339
rect 26326 11336 26332 11348
rect 26099 11308 26332 11336
rect 26099 11305 26111 11308
rect 26053 11299 26111 11305
rect 26326 11296 26332 11308
rect 26384 11296 26390 11348
rect 23934 11277 23940 11280
rect 23928 11268 23940 11277
rect 23895 11240 23940 11268
rect 23928 11231 23940 11240
rect 23934 11228 23940 11231
rect 23992 11228 23998 11280
rect 22465 11203 22523 11209
rect 22465 11200 22477 11203
rect 22428 11172 22477 11200
rect 22428 11160 22434 11172
rect 22465 11169 22477 11172
rect 22511 11169 22523 11203
rect 22465 11163 22523 11169
rect 23661 11203 23719 11209
rect 23661 11169 23673 11203
rect 23707 11169 23719 11203
rect 25958 11200 25964 11212
rect 23661 11163 23719 11169
rect 23768 11172 25964 11200
rect 23768 11132 23796 11172
rect 25958 11160 25964 11172
rect 26016 11160 26022 11212
rect 22296 11104 23796 11132
rect 18049 11067 18107 11073
rect 18049 11064 18061 11067
rect 18012 11036 18061 11064
rect 18012 11024 18018 11036
rect 18049 11033 18061 11036
rect 18095 11033 18107 11067
rect 18049 11027 18107 11033
rect 19705 11067 19763 11073
rect 19705 11033 19717 11067
rect 19751 11033 19763 11067
rect 19705 11027 19763 11033
rect 20346 11024 20352 11076
rect 20404 11064 20410 11076
rect 20901 11067 20959 11073
rect 20901 11064 20913 11067
rect 20404 11036 20913 11064
rect 20404 11024 20410 11036
rect 20901 11033 20913 11036
rect 20947 11033 20959 11067
rect 20901 11027 20959 11033
rect 21174 11024 21180 11076
rect 21232 11064 21238 11076
rect 22462 11064 22468 11076
rect 21232 11036 22468 11064
rect 21232 11024 21238 11036
rect 22462 11024 22468 11036
rect 22520 11024 22526 11076
rect 14369 10999 14427 11005
rect 14369 10996 14381 10999
rect 14240 10968 14381 10996
rect 14240 10956 14246 10968
rect 14369 10965 14381 10968
rect 14415 10996 14427 10999
rect 14737 10999 14795 11005
rect 14737 10996 14749 10999
rect 14415 10968 14749 10996
rect 14415 10965 14427 10968
rect 14369 10959 14427 10965
rect 14737 10965 14749 10968
rect 14783 10965 14795 10999
rect 20714 10996 20720 11008
rect 20675 10968 20720 10996
rect 14737 10959 14795 10965
rect 20714 10956 20720 10968
rect 20772 10956 20778 11008
rect 23106 10956 23112 11008
rect 23164 10996 23170 11008
rect 23382 10996 23388 11008
rect 23164 10968 23388 10996
rect 23164 10956 23170 10968
rect 23382 10956 23388 10968
rect 23440 10956 23446 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1397 10795 1455 10801
rect 1397 10761 1409 10795
rect 1443 10792 1455 10795
rect 1762 10792 1768 10804
rect 1443 10764 1768 10792
rect 1443 10761 1455 10764
rect 1397 10755 1455 10761
rect 1762 10752 1768 10764
rect 1820 10752 1826 10804
rect 2498 10792 2504 10804
rect 2459 10764 2504 10792
rect 2498 10752 2504 10764
rect 2556 10752 2562 10804
rect 5258 10752 5264 10804
rect 5316 10792 5322 10804
rect 5353 10795 5411 10801
rect 5353 10792 5365 10795
rect 5316 10764 5365 10792
rect 5316 10752 5322 10764
rect 5353 10761 5365 10764
rect 5399 10761 5411 10795
rect 6270 10792 6276 10804
rect 6231 10764 6276 10792
rect 5353 10755 5411 10761
rect 1946 10616 1952 10668
rect 2004 10656 2010 10668
rect 2041 10659 2099 10665
rect 2041 10656 2053 10659
rect 2004 10628 2053 10656
rect 2004 10616 2010 10628
rect 2041 10625 2053 10628
rect 2087 10656 2099 10659
rect 2958 10656 2964 10668
rect 2087 10628 2964 10656
rect 2087 10625 2099 10628
rect 2041 10619 2099 10625
rect 2958 10616 2964 10628
rect 3016 10616 3022 10668
rect 1026 10548 1032 10600
rect 1084 10588 1090 10600
rect 1765 10591 1823 10597
rect 1765 10588 1777 10591
rect 1084 10560 1777 10588
rect 1084 10548 1090 10560
rect 1765 10557 1777 10560
rect 1811 10557 1823 10591
rect 1765 10551 1823 10557
rect 1857 10591 1915 10597
rect 1857 10557 1869 10591
rect 1903 10588 1915 10591
rect 2406 10588 2412 10600
rect 1903 10560 2412 10588
rect 1903 10557 1915 10560
rect 1857 10551 1915 10557
rect 2406 10548 2412 10560
rect 2464 10548 2470 10600
rect 3053 10591 3111 10597
rect 3053 10557 3065 10591
rect 3099 10588 3111 10591
rect 3694 10588 3700 10600
rect 3099 10560 3700 10588
rect 3099 10557 3111 10560
rect 3053 10551 3111 10557
rect 3694 10548 3700 10560
rect 3752 10548 3758 10600
rect 4430 10588 4436 10600
rect 3896 10560 4436 10588
rect 2961 10523 3019 10529
rect 2961 10489 2973 10523
rect 3007 10520 3019 10523
rect 3320 10523 3378 10529
rect 3320 10520 3332 10523
rect 3007 10492 3332 10520
rect 3007 10489 3019 10492
rect 2961 10483 3019 10489
rect 3320 10489 3332 10492
rect 3366 10520 3378 10523
rect 3602 10520 3608 10532
rect 3366 10492 3608 10520
rect 3366 10489 3378 10492
rect 3320 10483 3378 10489
rect 3602 10480 3608 10492
rect 3660 10480 3666 10532
rect 2498 10412 2504 10464
rect 2556 10452 2562 10464
rect 3896 10452 3924 10560
rect 4430 10548 4436 10560
rect 4488 10548 4494 10600
rect 5368 10588 5396 10755
rect 6270 10752 6276 10764
rect 6328 10752 6334 10804
rect 7929 10795 7987 10801
rect 7929 10761 7941 10795
rect 7975 10792 7987 10795
rect 8110 10792 8116 10804
rect 7975 10764 8116 10792
rect 7975 10761 7987 10764
rect 7929 10755 7987 10761
rect 8110 10752 8116 10764
rect 8168 10752 8174 10804
rect 9674 10752 9680 10804
rect 9732 10792 9738 10804
rect 10413 10795 10471 10801
rect 10413 10792 10425 10795
rect 9732 10764 10425 10792
rect 9732 10752 9738 10764
rect 10413 10761 10425 10764
rect 10459 10792 10471 10795
rect 10502 10792 10508 10804
rect 10459 10764 10508 10792
rect 10459 10761 10471 10764
rect 10413 10755 10471 10761
rect 10502 10752 10508 10764
rect 10560 10752 10566 10804
rect 11054 10792 11060 10804
rect 11015 10764 11060 10792
rect 11054 10752 11060 10764
rect 11112 10752 11118 10804
rect 11330 10792 11336 10804
rect 11291 10764 11336 10792
rect 11330 10752 11336 10764
rect 11388 10752 11394 10804
rect 12158 10792 12164 10804
rect 12119 10764 12164 10792
rect 12158 10752 12164 10764
rect 12216 10752 12222 10804
rect 13446 10792 13452 10804
rect 13407 10764 13452 10792
rect 13446 10752 13452 10764
rect 13504 10752 13510 10804
rect 14550 10792 14556 10804
rect 13832 10764 14556 10792
rect 5718 10724 5724 10736
rect 5679 10696 5724 10724
rect 5718 10684 5724 10696
rect 5776 10684 5782 10736
rect 8205 10727 8263 10733
rect 8205 10724 8217 10727
rect 7300 10696 8217 10724
rect 6914 10616 6920 10668
rect 6972 10656 6978 10668
rect 7300 10665 7328 10696
rect 8205 10693 8217 10696
rect 8251 10693 8263 10727
rect 8205 10687 8263 10693
rect 11885 10727 11943 10733
rect 11885 10693 11897 10727
rect 11931 10724 11943 10727
rect 12066 10724 12072 10736
rect 11931 10696 12072 10724
rect 11931 10693 11943 10696
rect 11885 10687 11943 10693
rect 12066 10684 12072 10696
rect 12124 10724 12130 10736
rect 12802 10724 12808 10736
rect 12124 10696 12808 10724
rect 12124 10684 12130 10696
rect 12802 10684 12808 10696
rect 12860 10724 12866 10736
rect 13832 10733 13860 10764
rect 14550 10752 14556 10764
rect 14608 10752 14614 10804
rect 15562 10792 15568 10804
rect 15523 10764 15568 10792
rect 15562 10752 15568 10764
rect 15620 10752 15626 10804
rect 16390 10792 16396 10804
rect 16351 10764 16396 10792
rect 16390 10752 16396 10764
rect 16448 10752 16454 10804
rect 18690 10752 18696 10804
rect 18748 10792 18754 10804
rect 19058 10792 19064 10804
rect 18748 10764 19064 10792
rect 18748 10752 18754 10764
rect 19058 10752 19064 10764
rect 19116 10752 19122 10804
rect 19518 10792 19524 10804
rect 19479 10764 19524 10792
rect 19518 10752 19524 10764
rect 19576 10752 19582 10804
rect 20993 10795 21051 10801
rect 20993 10761 21005 10795
rect 21039 10792 21051 10795
rect 21358 10792 21364 10804
rect 21039 10764 21364 10792
rect 21039 10761 21051 10764
rect 20993 10755 21051 10761
rect 21358 10752 21364 10764
rect 21416 10752 21422 10804
rect 22370 10752 22376 10804
rect 22428 10792 22434 10804
rect 22465 10795 22523 10801
rect 22465 10792 22477 10795
rect 22428 10764 22477 10792
rect 22428 10752 22434 10764
rect 22465 10761 22477 10764
rect 22511 10761 22523 10795
rect 22465 10755 22523 10761
rect 22830 10752 22836 10804
rect 22888 10792 22894 10804
rect 23017 10795 23075 10801
rect 23017 10792 23029 10795
rect 22888 10764 23029 10792
rect 22888 10752 22894 10764
rect 23017 10761 23029 10764
rect 23063 10761 23075 10795
rect 23017 10755 23075 10761
rect 23477 10795 23535 10801
rect 23477 10761 23489 10795
rect 23523 10792 23535 10795
rect 23934 10792 23940 10804
rect 23523 10764 23940 10792
rect 23523 10761 23535 10764
rect 23477 10755 23535 10761
rect 13817 10727 13875 10733
rect 13817 10724 13829 10727
rect 12860 10696 13829 10724
rect 12860 10684 12866 10696
rect 13817 10693 13829 10696
rect 13863 10693 13875 10727
rect 13817 10687 13875 10693
rect 14001 10727 14059 10733
rect 14001 10693 14013 10727
rect 14047 10724 14059 10727
rect 15013 10727 15071 10733
rect 15013 10724 15025 10727
rect 14047 10696 15025 10724
rect 14047 10693 14059 10696
rect 14001 10687 14059 10693
rect 15013 10693 15025 10696
rect 15059 10693 15071 10727
rect 15013 10687 15071 10693
rect 7285 10659 7343 10665
rect 7285 10656 7297 10659
rect 6972 10628 7297 10656
rect 6972 10616 6978 10628
rect 7285 10625 7297 10628
rect 7331 10625 7343 10659
rect 7285 10619 7343 10625
rect 7377 10659 7435 10665
rect 7377 10625 7389 10659
rect 7423 10625 7435 10659
rect 7377 10619 7435 10625
rect 8941 10659 8999 10665
rect 8941 10625 8953 10659
rect 8987 10656 8999 10659
rect 13081 10659 13139 10665
rect 8987 10628 9168 10656
rect 8987 10625 8999 10628
rect 8941 10619 8999 10625
rect 5537 10591 5595 10597
rect 5537 10588 5549 10591
rect 5368 10560 5549 10588
rect 5537 10557 5549 10560
rect 5583 10557 5595 10591
rect 5537 10551 5595 10557
rect 6270 10548 6276 10600
rect 6328 10588 6334 10600
rect 6641 10591 6699 10597
rect 6641 10588 6653 10591
rect 6328 10560 6653 10588
rect 6328 10548 6334 10560
rect 6641 10557 6653 10560
rect 6687 10588 6699 10591
rect 7392 10588 7420 10619
rect 6687 10560 7420 10588
rect 9033 10591 9091 10597
rect 6687 10557 6699 10560
rect 6641 10551 6699 10557
rect 9033 10557 9045 10591
rect 9079 10557 9091 10591
rect 9140 10588 9168 10628
rect 13081 10625 13093 10659
rect 13127 10656 13139 10659
rect 13170 10656 13176 10668
rect 13127 10628 13176 10656
rect 13127 10625 13139 10628
rect 13081 10619 13139 10625
rect 13170 10616 13176 10628
rect 13228 10616 13234 10668
rect 9300 10591 9358 10597
rect 9300 10588 9312 10591
rect 9140 10560 9312 10588
rect 9033 10551 9091 10557
rect 9300 10557 9312 10560
rect 9346 10588 9358 10591
rect 9582 10588 9588 10600
rect 9346 10560 9588 10588
rect 9346 10557 9358 10560
rect 9300 10551 9358 10557
rect 4706 10520 4712 10532
rect 4448 10492 4712 10520
rect 2556 10424 3924 10452
rect 2556 10412 2562 10424
rect 3970 10412 3976 10464
rect 4028 10452 4034 10464
rect 4448 10461 4476 10492
rect 4706 10480 4712 10492
rect 4764 10520 4770 10532
rect 5077 10523 5135 10529
rect 5077 10520 5089 10523
rect 4764 10492 5089 10520
rect 4764 10480 4770 10492
rect 5077 10489 5089 10492
rect 5123 10520 5135 10523
rect 6288 10520 6316 10548
rect 5123 10492 6316 10520
rect 7193 10523 7251 10529
rect 5123 10489 5135 10492
rect 5077 10483 5135 10489
rect 7193 10489 7205 10523
rect 7239 10520 7251 10523
rect 8570 10520 8576 10532
rect 7239 10492 8576 10520
rect 7239 10489 7251 10492
rect 7193 10483 7251 10489
rect 8570 10480 8576 10492
rect 8628 10480 8634 10532
rect 9048 10520 9076 10551
rect 9582 10548 9588 10560
rect 9640 10548 9646 10600
rect 12805 10591 12863 10597
rect 12805 10557 12817 10591
rect 12851 10588 12863 10591
rect 14016 10588 14044 10687
rect 15286 10684 15292 10736
rect 15344 10724 15350 10736
rect 19337 10727 19395 10733
rect 19337 10724 19349 10727
rect 15344 10696 19349 10724
rect 15344 10684 15350 10696
rect 19337 10693 19349 10696
rect 19383 10724 19395 10727
rect 19794 10724 19800 10736
rect 19383 10696 19800 10724
rect 19383 10693 19395 10696
rect 19337 10687 19395 10693
rect 19794 10684 19800 10696
rect 19852 10684 19858 10736
rect 19886 10684 19892 10736
rect 19944 10724 19950 10736
rect 20533 10727 20591 10733
rect 20533 10724 20545 10727
rect 19944 10696 20545 10724
rect 19944 10684 19950 10696
rect 20533 10693 20545 10696
rect 20579 10693 20591 10727
rect 21082 10724 21088 10736
rect 21043 10696 21088 10724
rect 20533 10687 20591 10693
rect 21082 10684 21088 10696
rect 21140 10684 21146 10736
rect 14090 10616 14096 10668
rect 14148 10656 14154 10668
rect 14461 10659 14519 10665
rect 14461 10656 14473 10659
rect 14148 10628 14473 10656
rect 14148 10616 14154 10628
rect 14461 10625 14473 10628
rect 14507 10625 14519 10659
rect 14461 10619 14519 10625
rect 14550 10616 14556 10668
rect 14608 10656 14614 10668
rect 14608 10628 14653 10656
rect 14608 10616 14614 10628
rect 16298 10616 16304 10668
rect 16356 10616 16362 10668
rect 16850 10616 16856 10668
rect 16908 10656 16914 10668
rect 16945 10659 17003 10665
rect 16945 10656 16957 10659
rect 16908 10628 16957 10656
rect 16908 10616 16914 10628
rect 16945 10625 16957 10628
rect 16991 10656 17003 10659
rect 17405 10659 17463 10665
rect 17405 10656 17417 10659
rect 16991 10628 17417 10656
rect 16991 10625 17003 10628
rect 16945 10619 17003 10625
rect 17405 10625 17417 10628
rect 17451 10656 17463 10659
rect 18233 10659 18291 10665
rect 18233 10656 18245 10659
rect 17451 10628 18245 10656
rect 17451 10625 17463 10628
rect 17405 10619 17463 10625
rect 18233 10625 18245 10628
rect 18279 10656 18291 10659
rect 20073 10659 20131 10665
rect 20073 10656 20085 10659
rect 18279 10628 20085 10656
rect 18279 10625 18291 10628
rect 18233 10619 18291 10625
rect 20073 10625 20085 10628
rect 20119 10656 20131 10659
rect 20254 10656 20260 10668
rect 20119 10628 20260 10656
rect 20119 10625 20131 10628
rect 20073 10619 20131 10625
rect 20254 10616 20260 10628
rect 20312 10616 20318 10668
rect 20806 10616 20812 10668
rect 20864 10656 20870 10668
rect 21545 10659 21603 10665
rect 21545 10656 21557 10659
rect 20864 10628 21557 10656
rect 20864 10616 20870 10628
rect 21545 10625 21557 10628
rect 21591 10656 21603 10659
rect 21634 10656 21640 10668
rect 21591 10628 21640 10656
rect 21591 10625 21603 10628
rect 21545 10619 21603 10625
rect 21634 10616 21640 10628
rect 21692 10616 21698 10668
rect 21729 10659 21787 10665
rect 21729 10625 21741 10659
rect 21775 10656 21787 10659
rect 22094 10656 22100 10668
rect 21775 10628 22100 10656
rect 21775 10625 21787 10628
rect 21729 10619 21787 10625
rect 22094 10616 22100 10628
rect 22152 10656 22158 10668
rect 23032 10656 23060 10755
rect 23934 10752 23940 10764
rect 23992 10792 23998 10804
rect 25041 10795 25099 10801
rect 25041 10792 25053 10795
rect 23992 10764 25053 10792
rect 23992 10752 23998 10764
rect 25041 10761 25053 10764
rect 25087 10761 25099 10795
rect 25041 10755 25099 10761
rect 22152 10628 22245 10656
rect 23032 10628 23796 10656
rect 22152 10616 22158 10628
rect 12851 10560 14044 10588
rect 15933 10591 15991 10597
rect 12851 10557 12863 10560
rect 12805 10551 12863 10557
rect 15933 10557 15945 10591
rect 15979 10588 15991 10591
rect 16316 10588 16344 10616
rect 17865 10591 17923 10597
rect 15979 10560 16896 10588
rect 15979 10557 15991 10560
rect 15933 10551 15991 10557
rect 9122 10520 9128 10532
rect 9048 10492 9128 10520
rect 9122 10480 9128 10492
rect 9180 10480 9186 10532
rect 11238 10480 11244 10532
rect 11296 10520 11302 10532
rect 11296 10492 13124 10520
rect 11296 10480 11302 10492
rect 4433 10455 4491 10461
rect 4433 10452 4445 10455
rect 4028 10424 4445 10452
rect 4028 10412 4034 10424
rect 4433 10421 4445 10424
rect 4479 10421 4491 10455
rect 6822 10452 6828 10464
rect 6783 10424 6828 10452
rect 4433 10415 4491 10421
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 12437 10455 12495 10461
rect 12437 10421 12449 10455
rect 12483 10452 12495 10455
rect 12710 10452 12716 10464
rect 12483 10424 12716 10452
rect 12483 10421 12495 10424
rect 12437 10415 12495 10421
rect 12710 10412 12716 10424
rect 12768 10412 12774 10464
rect 12894 10452 12900 10464
rect 12855 10424 12900 10452
rect 12894 10412 12900 10424
rect 12952 10412 12958 10464
rect 13096 10452 13124 10492
rect 13446 10480 13452 10532
rect 13504 10520 13510 10532
rect 14369 10523 14427 10529
rect 14369 10520 14381 10523
rect 13504 10492 14381 10520
rect 13504 10480 13510 10492
rect 14369 10489 14381 10492
rect 14415 10489 14427 10523
rect 16761 10523 16819 10529
rect 16761 10520 16773 10523
rect 14369 10483 14427 10489
rect 16224 10492 16773 10520
rect 16224 10464 16252 10492
rect 16761 10489 16773 10492
rect 16807 10489 16819 10523
rect 16761 10483 16819 10489
rect 16868 10464 16896 10560
rect 17865 10557 17877 10591
rect 17911 10588 17923 10591
rect 18417 10591 18475 10597
rect 18417 10588 18429 10591
rect 17911 10560 18429 10588
rect 17911 10557 17923 10560
rect 17865 10551 17923 10557
rect 18417 10557 18429 10560
rect 18463 10588 18475 10591
rect 18506 10588 18512 10600
rect 18463 10560 18512 10588
rect 18463 10557 18475 10560
rect 18417 10551 18475 10557
rect 18506 10548 18512 10560
rect 18564 10548 18570 10600
rect 19794 10548 19800 10600
rect 19852 10588 19858 10600
rect 19981 10591 20039 10597
rect 19981 10588 19993 10591
rect 19852 10560 19993 10588
rect 19852 10548 19858 10560
rect 19981 10557 19993 10560
rect 20027 10557 20039 10591
rect 19981 10551 20039 10557
rect 20714 10548 20720 10600
rect 20772 10588 20778 10600
rect 21453 10591 21511 10597
rect 21453 10588 21465 10591
rect 20772 10560 21465 10588
rect 20772 10548 20778 10560
rect 21453 10557 21465 10560
rect 21499 10557 21511 10591
rect 21453 10551 21511 10557
rect 23661 10591 23719 10597
rect 23661 10557 23673 10591
rect 23707 10557 23719 10591
rect 23768 10588 23796 10628
rect 23917 10591 23975 10597
rect 23917 10588 23929 10591
rect 23768 10560 23929 10588
rect 23661 10551 23719 10557
rect 23917 10557 23929 10560
rect 23963 10588 23975 10591
rect 24854 10588 24860 10600
rect 23963 10560 24860 10588
rect 23963 10557 23975 10560
rect 23917 10551 23975 10557
rect 19061 10523 19119 10529
rect 19061 10489 19073 10523
rect 19107 10520 19119 10523
rect 19889 10523 19947 10529
rect 19889 10520 19901 10523
rect 19107 10492 19901 10520
rect 19107 10489 19119 10492
rect 19061 10483 19119 10489
rect 19889 10489 19901 10492
rect 19935 10520 19947 10523
rect 22554 10520 22560 10532
rect 19935 10492 22560 10520
rect 19935 10489 19947 10492
rect 19889 10483 19947 10489
rect 22554 10480 22560 10492
rect 22612 10480 22618 10532
rect 15930 10452 15936 10464
rect 13096 10424 15936 10452
rect 15930 10412 15936 10424
rect 15988 10412 15994 10464
rect 16206 10452 16212 10464
rect 16167 10424 16212 10452
rect 16206 10412 16212 10424
rect 16264 10412 16270 10464
rect 16850 10452 16856 10464
rect 16811 10424 16856 10452
rect 16850 10412 16856 10424
rect 16908 10412 16914 10464
rect 18601 10455 18659 10461
rect 18601 10421 18613 10455
rect 18647 10452 18659 10455
rect 18966 10452 18972 10464
rect 18647 10424 18972 10452
rect 18647 10421 18659 10424
rect 18601 10415 18659 10421
rect 18966 10412 18972 10424
rect 19024 10412 19030 10464
rect 23676 10452 23704 10551
rect 24854 10548 24860 10560
rect 24912 10548 24918 10600
rect 24026 10452 24032 10464
rect 23676 10424 24032 10452
rect 24026 10412 24032 10424
rect 24084 10452 24090 10464
rect 25498 10452 25504 10464
rect 24084 10424 25504 10452
rect 24084 10412 24090 10424
rect 25498 10412 25504 10424
rect 25556 10452 25562 10464
rect 25593 10455 25651 10461
rect 25593 10452 25605 10455
rect 25556 10424 25605 10452
rect 25556 10412 25562 10424
rect 25593 10421 25605 10424
rect 25639 10452 25651 10455
rect 25961 10455 26019 10461
rect 25961 10452 25973 10455
rect 25639 10424 25973 10452
rect 25639 10421 25651 10424
rect 25593 10415 25651 10421
rect 25961 10421 25973 10424
rect 26007 10452 26019 10455
rect 26329 10455 26387 10461
rect 26329 10452 26341 10455
rect 26007 10424 26341 10452
rect 26007 10421 26019 10424
rect 25961 10415 26019 10421
rect 26329 10421 26341 10424
rect 26375 10421 26387 10455
rect 26329 10415 26387 10421
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1946 10248 1952 10260
rect 1907 10220 1952 10248
rect 1946 10208 1952 10220
rect 2004 10208 2010 10260
rect 2409 10251 2467 10257
rect 2409 10217 2421 10251
rect 2455 10248 2467 10251
rect 2774 10248 2780 10260
rect 2455 10220 2780 10248
rect 2455 10217 2467 10220
rect 2409 10211 2467 10217
rect 2774 10208 2780 10220
rect 2832 10208 2838 10260
rect 3142 10208 3148 10260
rect 3200 10248 3206 10260
rect 4065 10251 4123 10257
rect 4065 10248 4077 10251
rect 3200 10220 4077 10248
rect 3200 10208 3206 10220
rect 4065 10217 4077 10220
rect 4111 10217 4123 10251
rect 4065 10211 4123 10217
rect 6089 10251 6147 10257
rect 6089 10217 6101 10251
rect 6135 10248 6147 10251
rect 6362 10248 6368 10260
rect 6135 10220 6368 10248
rect 6135 10217 6147 10220
rect 6089 10211 6147 10217
rect 6362 10208 6368 10220
rect 6420 10208 6426 10260
rect 7561 10251 7619 10257
rect 7561 10217 7573 10251
rect 7607 10248 7619 10251
rect 8018 10248 8024 10260
rect 7607 10220 8024 10248
rect 7607 10217 7619 10220
rect 7561 10211 7619 10217
rect 8018 10208 8024 10220
rect 8076 10248 8082 10260
rect 8205 10251 8263 10257
rect 8205 10248 8217 10251
rect 8076 10220 8217 10248
rect 8076 10208 8082 10220
rect 8205 10217 8217 10220
rect 8251 10217 8263 10251
rect 8570 10248 8576 10260
rect 8531 10220 8576 10248
rect 8205 10211 8263 10217
rect 8570 10208 8576 10220
rect 8628 10248 8634 10260
rect 9677 10251 9735 10257
rect 9677 10248 9689 10251
rect 8628 10220 9689 10248
rect 8628 10208 8634 10220
rect 9677 10217 9689 10220
rect 9723 10217 9735 10251
rect 10686 10248 10692 10260
rect 10647 10220 10692 10248
rect 9677 10211 9735 10217
rect 10686 10208 10692 10220
rect 10744 10208 10750 10260
rect 10870 10208 10876 10260
rect 10928 10248 10934 10260
rect 10928 10220 11928 10248
rect 10928 10208 10934 10220
rect 2869 10183 2927 10189
rect 2869 10149 2881 10183
rect 2915 10180 2927 10183
rect 3510 10180 3516 10192
rect 2915 10152 3516 10180
rect 2915 10149 2927 10152
rect 2869 10143 2927 10149
rect 3510 10140 3516 10152
rect 3568 10140 3574 10192
rect 3697 10183 3755 10189
rect 3697 10149 3709 10183
rect 3743 10180 3755 10183
rect 4430 10180 4436 10192
rect 3743 10152 4436 10180
rect 3743 10149 3755 10152
rect 3697 10143 3755 10149
rect 4430 10140 4436 10152
rect 4488 10140 4494 10192
rect 5997 10183 6055 10189
rect 5997 10149 6009 10183
rect 6043 10180 6055 10183
rect 8110 10180 8116 10192
rect 6043 10152 8116 10180
rect 6043 10149 6055 10152
rect 5997 10143 6055 10149
rect 8110 10140 8116 10152
rect 8168 10140 8174 10192
rect 9214 10180 9220 10192
rect 9175 10152 9220 10180
rect 9214 10140 9220 10152
rect 9272 10140 9278 10192
rect 10137 10183 10195 10189
rect 10137 10149 10149 10183
rect 10183 10180 10195 10183
rect 10778 10180 10784 10192
rect 10183 10152 10784 10180
rect 10183 10149 10195 10152
rect 10137 10143 10195 10149
rect 10778 10140 10784 10152
rect 10836 10180 10842 10192
rect 11054 10180 11060 10192
rect 10836 10152 11060 10180
rect 10836 10140 10842 10152
rect 11054 10140 11060 10152
rect 11112 10140 11118 10192
rect 11330 10140 11336 10192
rect 11388 10180 11394 10192
rect 11762 10183 11820 10189
rect 11762 10180 11774 10183
rect 11388 10152 11774 10180
rect 11388 10140 11394 10152
rect 11762 10149 11774 10152
rect 11808 10149 11820 10183
rect 11900 10180 11928 10220
rect 12894 10208 12900 10260
rect 12952 10248 12958 10260
rect 13817 10251 13875 10257
rect 13817 10248 13829 10251
rect 12952 10220 13829 10248
rect 12952 10208 12958 10220
rect 13817 10217 13829 10220
rect 13863 10248 13875 10251
rect 13998 10248 14004 10260
rect 13863 10220 14004 10248
rect 13863 10217 13875 10220
rect 13817 10211 13875 10217
rect 13998 10208 14004 10220
rect 14056 10208 14062 10260
rect 14277 10251 14335 10257
rect 14277 10217 14289 10251
rect 14323 10248 14335 10251
rect 15378 10248 15384 10260
rect 14323 10220 15384 10248
rect 14323 10217 14335 10220
rect 14277 10211 14335 10217
rect 15378 10208 15384 10220
rect 15436 10208 15442 10260
rect 16942 10208 16948 10260
rect 17000 10248 17006 10260
rect 17681 10251 17739 10257
rect 17681 10248 17693 10251
rect 17000 10220 17693 10248
rect 17000 10208 17006 10220
rect 17681 10217 17693 10220
rect 17727 10217 17739 10251
rect 17681 10211 17739 10217
rect 14642 10180 14648 10192
rect 11900 10152 14648 10180
rect 11762 10143 11820 10149
rect 14642 10140 14648 10152
rect 14700 10140 14706 10192
rect 15556 10183 15614 10189
rect 15556 10149 15568 10183
rect 15602 10180 15614 10183
rect 16298 10180 16304 10192
rect 15602 10152 16304 10180
rect 15602 10149 15614 10152
rect 15556 10143 15614 10149
rect 16298 10140 16304 10152
rect 16356 10180 16362 10192
rect 16482 10180 16488 10192
rect 16356 10152 16488 10180
rect 16356 10140 16362 10152
rect 16482 10140 16488 10152
rect 16540 10140 16546 10192
rect 1946 10072 1952 10124
rect 2004 10112 2010 10124
rect 2774 10112 2780 10124
rect 2004 10084 2780 10112
rect 2004 10072 2010 10084
rect 2774 10072 2780 10084
rect 2832 10112 2838 10124
rect 3528 10112 3556 10140
rect 4062 10112 4068 10124
rect 2832 10084 2925 10112
rect 3528 10084 4068 10112
rect 2832 10072 2838 10084
rect 4062 10072 4068 10084
rect 4120 10072 4126 10124
rect 4525 10115 4583 10121
rect 4525 10081 4537 10115
rect 4571 10112 4583 10115
rect 4798 10112 4804 10124
rect 4571 10084 4804 10112
rect 4571 10081 4583 10084
rect 4525 10075 4583 10081
rect 4798 10072 4804 10084
rect 4856 10072 4862 10124
rect 8941 10115 8999 10121
rect 8941 10081 8953 10115
rect 8987 10112 8999 10115
rect 9306 10112 9312 10124
rect 8987 10084 9312 10112
rect 8987 10081 8999 10084
rect 8941 10075 8999 10081
rect 9306 10072 9312 10084
rect 9364 10072 9370 10124
rect 9766 10072 9772 10124
rect 9824 10112 9830 10124
rect 10045 10115 10103 10121
rect 10045 10112 10057 10115
rect 9824 10084 10057 10112
rect 9824 10072 9830 10084
rect 10045 10081 10057 10084
rect 10091 10112 10103 10115
rect 10318 10112 10324 10124
rect 10091 10084 10324 10112
rect 10091 10081 10103 10084
rect 10045 10075 10103 10081
rect 10318 10072 10324 10084
rect 10376 10072 10382 10124
rect 11514 10112 11520 10124
rect 11475 10084 11520 10112
rect 11514 10072 11520 10084
rect 11572 10072 11578 10124
rect 12618 10072 12624 10124
rect 12676 10112 12682 10124
rect 12894 10112 12900 10124
rect 12676 10084 12900 10112
rect 12676 10072 12682 10084
rect 12894 10072 12900 10084
rect 12952 10072 12958 10124
rect 13814 10072 13820 10124
rect 13872 10112 13878 10124
rect 14093 10115 14151 10121
rect 14093 10112 14105 10115
rect 13872 10084 14105 10112
rect 13872 10072 13878 10084
rect 14093 10081 14105 10084
rect 14139 10081 14151 10115
rect 17696 10112 17724 10211
rect 18046 10208 18052 10260
rect 18104 10248 18110 10260
rect 19061 10251 19119 10257
rect 19061 10248 19073 10251
rect 18104 10220 19073 10248
rect 18104 10208 18110 10220
rect 19061 10217 19073 10220
rect 19107 10217 19119 10251
rect 19242 10248 19248 10260
rect 19203 10220 19248 10248
rect 19061 10211 19119 10217
rect 18049 10115 18107 10121
rect 18049 10112 18061 10115
rect 17696 10084 18061 10112
rect 14093 10075 14151 10081
rect 18049 10081 18061 10084
rect 18095 10081 18107 10115
rect 18049 10075 18107 10081
rect 18138 10072 18144 10124
rect 18196 10112 18202 10124
rect 19076 10112 19104 10211
rect 19242 10208 19248 10220
rect 19300 10208 19306 10260
rect 19426 10208 19432 10260
rect 19484 10248 19490 10260
rect 19613 10251 19671 10257
rect 19613 10248 19625 10251
rect 19484 10220 19625 10248
rect 19484 10208 19490 10220
rect 19613 10217 19625 10220
rect 19659 10248 19671 10251
rect 20346 10248 20352 10260
rect 19659 10220 20352 10248
rect 19659 10217 19671 10220
rect 19613 10211 19671 10217
rect 20346 10208 20352 10220
rect 20404 10208 20410 10260
rect 20530 10208 20536 10260
rect 20588 10248 20594 10260
rect 21450 10248 21456 10260
rect 20588 10220 21456 10248
rect 20588 10208 20594 10220
rect 21450 10208 21456 10220
rect 21508 10208 21514 10260
rect 21634 10208 21640 10260
rect 21692 10248 21698 10260
rect 22833 10251 22891 10257
rect 22833 10248 22845 10251
rect 21692 10220 22845 10248
rect 21692 10208 21698 10220
rect 22833 10217 22845 10220
rect 22879 10217 22891 10251
rect 22833 10211 22891 10217
rect 23106 10208 23112 10260
rect 23164 10248 23170 10260
rect 23201 10251 23259 10257
rect 23201 10248 23213 10251
rect 23164 10220 23213 10248
rect 23164 10208 23170 10220
rect 23201 10217 23213 10220
rect 23247 10217 23259 10251
rect 23201 10211 23259 10217
rect 23750 10208 23756 10260
rect 23808 10248 23814 10260
rect 23845 10251 23903 10257
rect 23845 10248 23857 10251
rect 23808 10220 23857 10248
rect 23808 10208 23814 10220
rect 23845 10217 23857 10220
rect 23891 10248 23903 10251
rect 23934 10248 23940 10260
rect 23891 10220 23940 10248
rect 23891 10217 23903 10220
rect 23845 10211 23903 10217
rect 23934 10208 23940 10220
rect 23992 10208 23998 10260
rect 24489 10251 24547 10257
rect 24489 10217 24501 10251
rect 24535 10248 24547 10251
rect 24670 10248 24676 10260
rect 24535 10220 24676 10248
rect 24535 10217 24547 10220
rect 24489 10211 24547 10217
rect 24670 10208 24676 10220
rect 24728 10208 24734 10260
rect 24762 10208 24768 10260
rect 24820 10248 24826 10260
rect 25314 10248 25320 10260
rect 24820 10220 25320 10248
rect 24820 10208 24826 10220
rect 25314 10208 25320 10220
rect 25372 10208 25378 10260
rect 25498 10248 25504 10260
rect 25459 10220 25504 10248
rect 25498 10208 25504 10220
rect 25556 10248 25562 10260
rect 25869 10251 25927 10257
rect 25869 10248 25881 10251
rect 25556 10220 25881 10248
rect 25556 10208 25562 10220
rect 25869 10217 25881 10220
rect 25915 10248 25927 10251
rect 26237 10251 26295 10257
rect 26237 10248 26249 10251
rect 25915 10220 26249 10248
rect 25915 10217 25927 10220
rect 25869 10211 25927 10217
rect 26237 10217 26249 10220
rect 26283 10248 26295 10251
rect 26418 10248 26424 10260
rect 26283 10220 26424 10248
rect 26283 10217 26295 10220
rect 26237 10211 26295 10217
rect 26418 10208 26424 10220
rect 26476 10208 26482 10260
rect 20254 10180 20260 10192
rect 20215 10152 20260 10180
rect 20254 10140 20260 10152
rect 20312 10140 20318 10192
rect 20717 10183 20775 10189
rect 20717 10149 20729 10183
rect 20763 10180 20775 10183
rect 21168 10183 21226 10189
rect 21168 10180 21180 10183
rect 20763 10152 21180 10180
rect 20763 10149 20775 10152
rect 20717 10143 20775 10149
rect 21168 10149 21180 10152
rect 21214 10180 21226 10183
rect 21910 10180 21916 10192
rect 21214 10152 21916 10180
rect 21214 10149 21226 10152
rect 21168 10143 21226 10149
rect 19242 10112 19248 10124
rect 18196 10084 18241 10112
rect 19076 10084 19248 10112
rect 18196 10072 18202 10084
rect 19242 10072 19248 10084
rect 19300 10072 19306 10124
rect 20622 10072 20628 10124
rect 20680 10112 20686 10124
rect 20732 10112 20760 10143
rect 21910 10140 21916 10152
rect 21968 10140 21974 10192
rect 20680 10084 20760 10112
rect 20680 10072 20686 10084
rect 20990 10072 20996 10124
rect 21048 10112 21054 10124
rect 21048 10084 21956 10112
rect 21048 10072 21054 10084
rect 1397 10047 1455 10053
rect 1397 10013 1409 10047
rect 1443 10044 1455 10047
rect 1443 10016 2912 10044
rect 1443 10013 1455 10016
rect 1397 10007 1455 10013
rect 1118 9936 1124 9988
rect 1176 9976 1182 9988
rect 2884 9976 2912 10016
rect 2958 10004 2964 10056
rect 3016 10044 3022 10056
rect 3053 10047 3111 10053
rect 3053 10044 3065 10047
rect 3016 10016 3065 10044
rect 3016 10004 3022 10016
rect 3053 10013 3065 10016
rect 3099 10044 3111 10047
rect 3970 10044 3976 10056
rect 3099 10016 3976 10044
rect 3099 10013 3111 10016
rect 3053 10007 3111 10013
rect 3970 10004 3976 10016
rect 4028 10004 4034 10056
rect 4706 10044 4712 10056
rect 4667 10016 4712 10044
rect 4706 10004 4712 10016
rect 4764 10004 4770 10056
rect 6270 10044 6276 10056
rect 6231 10016 6276 10044
rect 6270 10004 6276 10016
rect 6328 10004 6334 10056
rect 6733 10047 6791 10053
rect 6733 10013 6745 10047
rect 6779 10044 6791 10047
rect 7650 10044 7656 10056
rect 6779 10016 7656 10044
rect 6779 10013 6791 10016
rect 6733 10007 6791 10013
rect 7650 10004 7656 10016
rect 7708 10004 7714 10056
rect 7745 10047 7803 10053
rect 7745 10013 7757 10047
rect 7791 10013 7803 10047
rect 7745 10007 7803 10013
rect 10229 10047 10287 10053
rect 10229 10013 10241 10047
rect 10275 10013 10287 10047
rect 10229 10007 10287 10013
rect 3697 9979 3755 9985
rect 3697 9976 3709 9979
rect 1176 9948 2360 9976
rect 2884 9948 3709 9976
rect 1176 9936 1182 9948
rect 2222 9908 2228 9920
rect 2183 9880 2228 9908
rect 2222 9868 2228 9880
rect 2280 9868 2286 9920
rect 2332 9908 2360 9948
rect 3697 9945 3709 9948
rect 3743 9945 3755 9979
rect 3878 9976 3884 9988
rect 3839 9948 3884 9976
rect 3697 9939 3755 9945
rect 3878 9936 3884 9948
rect 3936 9936 3942 9988
rect 5629 9979 5687 9985
rect 5629 9945 5641 9979
rect 5675 9976 5687 9979
rect 6638 9976 6644 9988
rect 5675 9948 6644 9976
rect 5675 9945 5687 9948
rect 5629 9939 5687 9945
rect 6638 9936 6644 9948
rect 6696 9936 6702 9988
rect 7190 9976 7196 9988
rect 7151 9948 7196 9976
rect 7190 9936 7196 9948
rect 7248 9936 7254 9988
rect 7760 9976 7788 10007
rect 7300 9948 7788 9976
rect 7300 9920 7328 9948
rect 9490 9936 9496 9988
rect 9548 9976 9554 9988
rect 10244 9976 10272 10007
rect 14182 10004 14188 10056
rect 14240 10044 14246 10056
rect 15013 10047 15071 10053
rect 15013 10044 15025 10047
rect 14240 10016 15025 10044
rect 14240 10004 14246 10016
rect 15013 10013 15025 10016
rect 15059 10013 15071 10047
rect 15286 10044 15292 10056
rect 15247 10016 15292 10044
rect 15013 10007 15071 10013
rect 15286 10004 15292 10016
rect 15344 10004 15350 10056
rect 18785 10047 18843 10053
rect 18785 10013 18797 10047
rect 18831 10044 18843 10047
rect 19150 10044 19156 10056
rect 18831 10016 19156 10044
rect 18831 10013 18843 10016
rect 18785 10007 18843 10013
rect 19150 10004 19156 10016
rect 19208 10044 19214 10056
rect 19705 10047 19763 10053
rect 19705 10044 19717 10047
rect 19208 10016 19717 10044
rect 19208 10004 19214 10016
rect 19705 10013 19717 10016
rect 19751 10013 19763 10047
rect 19705 10007 19763 10013
rect 19889 10047 19947 10053
rect 19889 10013 19901 10047
rect 19935 10044 19947 10047
rect 19978 10044 19984 10056
rect 19935 10016 19984 10044
rect 19935 10013 19947 10016
rect 19889 10007 19947 10013
rect 19978 10004 19984 10016
rect 20036 10004 20042 10056
rect 20162 10004 20168 10056
rect 20220 10044 20226 10056
rect 20714 10044 20720 10056
rect 20220 10016 20720 10044
rect 20220 10004 20226 10016
rect 20714 10004 20720 10016
rect 20772 10044 20778 10056
rect 20901 10047 20959 10053
rect 20901 10044 20913 10047
rect 20772 10016 20913 10044
rect 20772 10004 20778 10016
rect 20901 10013 20913 10016
rect 20947 10013 20959 10047
rect 20901 10007 20959 10013
rect 9548 9948 10272 9976
rect 9548 9936 9554 9948
rect 12802 9936 12808 9988
rect 12860 9976 12866 9988
rect 12897 9979 12955 9985
rect 12897 9976 12909 9979
rect 12860 9948 12909 9976
rect 12860 9936 12866 9948
rect 12897 9945 12909 9948
rect 12943 9945 12955 9979
rect 21928 9976 21956 10084
rect 23382 10072 23388 10124
rect 23440 10112 23446 10124
rect 23750 10112 23756 10124
rect 23440 10084 23756 10112
rect 23440 10072 23446 10084
rect 23750 10072 23756 10084
rect 23808 10072 23814 10124
rect 24946 10112 24952 10124
rect 24907 10084 24952 10112
rect 24946 10072 24952 10084
rect 25004 10112 25010 10124
rect 25590 10112 25596 10124
rect 25004 10084 25596 10112
rect 25004 10072 25010 10084
rect 25590 10072 25596 10084
rect 25648 10072 25654 10124
rect 22462 10004 22468 10056
rect 22520 10044 22526 10056
rect 23842 10044 23848 10056
rect 22520 10016 23848 10044
rect 22520 10004 22526 10016
rect 23842 10004 23848 10016
rect 23900 10004 23906 10056
rect 23937 10047 23995 10053
rect 23937 10013 23949 10047
rect 23983 10013 23995 10047
rect 23937 10007 23995 10013
rect 23385 9979 23443 9985
rect 23385 9976 23397 9979
rect 21928 9948 23397 9976
rect 12897 9939 12955 9945
rect 23385 9945 23397 9948
rect 23431 9945 23443 9979
rect 23385 9939 23443 9945
rect 23474 9936 23480 9988
rect 23532 9976 23538 9988
rect 23952 9976 23980 10007
rect 24670 10004 24676 10056
rect 24728 10044 24734 10056
rect 24728 10016 24808 10044
rect 24728 10004 24734 10016
rect 23532 9948 23980 9976
rect 23532 9936 23538 9948
rect 24780 9920 24808 10016
rect 2866 9908 2872 9920
rect 2332 9880 2872 9908
rect 2866 9868 2872 9880
rect 2924 9868 2930 9920
rect 3510 9908 3516 9920
rect 3471 9880 3516 9908
rect 3510 9868 3516 9880
rect 3568 9868 3574 9920
rect 4614 9868 4620 9920
rect 4672 9908 4678 9920
rect 5169 9911 5227 9917
rect 5169 9908 5181 9911
rect 4672 9880 5181 9908
rect 4672 9868 4678 9880
rect 5169 9877 5181 9880
rect 5215 9877 5227 9911
rect 5169 9871 5227 9877
rect 7101 9911 7159 9917
rect 7101 9877 7113 9911
rect 7147 9908 7159 9911
rect 7282 9908 7288 9920
rect 7147 9880 7288 9908
rect 7147 9877 7159 9880
rect 7101 9871 7159 9877
rect 7282 9868 7288 9880
rect 7340 9868 7346 9920
rect 8662 9868 8668 9920
rect 8720 9908 8726 9920
rect 8757 9911 8815 9917
rect 8757 9908 8769 9911
rect 8720 9880 8769 9908
rect 8720 9868 8726 9880
rect 8757 9877 8769 9880
rect 8803 9908 8815 9911
rect 11057 9911 11115 9917
rect 11057 9908 11069 9911
rect 8803 9880 11069 9908
rect 8803 9877 8815 9880
rect 8757 9871 8815 9877
rect 11057 9877 11069 9880
rect 11103 9877 11115 9911
rect 13446 9908 13452 9920
rect 13407 9880 13452 9908
rect 11057 9871 11115 9877
rect 13446 9868 13452 9880
rect 13504 9868 13510 9920
rect 14642 9908 14648 9920
rect 14603 9880 14648 9908
rect 14642 9868 14648 9880
rect 14700 9868 14706 9920
rect 16669 9911 16727 9917
rect 16669 9877 16681 9911
rect 16715 9908 16727 9911
rect 16758 9908 16764 9920
rect 16715 9880 16764 9908
rect 16715 9877 16727 9880
rect 16669 9871 16727 9877
rect 16758 9868 16764 9880
rect 16816 9868 16822 9920
rect 17218 9908 17224 9920
rect 17179 9880 17224 9908
rect 17218 9868 17224 9880
rect 17276 9868 17282 9920
rect 17310 9868 17316 9920
rect 17368 9908 17374 9920
rect 17865 9911 17923 9917
rect 17865 9908 17877 9911
rect 17368 9880 17877 9908
rect 17368 9868 17374 9880
rect 17865 9877 17877 9880
rect 17911 9877 17923 9911
rect 17865 9871 17923 9877
rect 18046 9868 18052 9920
rect 18104 9908 18110 9920
rect 18325 9911 18383 9917
rect 18325 9908 18337 9911
rect 18104 9880 18337 9908
rect 18104 9868 18110 9880
rect 18325 9877 18337 9880
rect 18371 9877 18383 9911
rect 18325 9871 18383 9877
rect 22002 9868 22008 9920
rect 22060 9908 22066 9920
rect 22281 9911 22339 9917
rect 22281 9908 22293 9911
rect 22060 9880 22293 9908
rect 22060 9868 22066 9880
rect 22281 9877 22293 9880
rect 22327 9877 22339 9911
rect 22281 9871 22339 9877
rect 24762 9868 24768 9920
rect 24820 9868 24826 9920
rect 24946 9868 24952 9920
rect 25004 9908 25010 9920
rect 25133 9911 25191 9917
rect 25133 9908 25145 9911
rect 25004 9880 25145 9908
rect 25004 9868 25010 9880
rect 25133 9877 25145 9880
rect 25179 9877 25191 9911
rect 25133 9871 25191 9877
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 2130 9664 2136 9716
rect 2188 9704 2194 9716
rect 2498 9704 2504 9716
rect 2188 9676 2504 9704
rect 2188 9664 2194 9676
rect 2498 9664 2504 9676
rect 2556 9664 2562 9716
rect 4430 9704 4436 9716
rect 4391 9676 4436 9704
rect 4430 9664 4436 9676
rect 4488 9664 4494 9716
rect 6362 9704 6368 9716
rect 5460 9676 6368 9704
rect 1946 9636 1952 9648
rect 1907 9608 1952 9636
rect 1946 9596 1952 9608
rect 2004 9596 2010 9648
rect 5169 9639 5227 9645
rect 5169 9605 5181 9639
rect 5215 9636 5227 9639
rect 5460 9636 5488 9676
rect 6362 9664 6368 9676
rect 6420 9664 6426 9716
rect 7098 9704 7104 9716
rect 6472 9676 7104 9704
rect 6270 9636 6276 9648
rect 5215 9608 5488 9636
rect 6231 9608 6276 9636
rect 5215 9605 5227 9608
rect 5169 9599 5227 9605
rect 6270 9596 6276 9608
rect 6328 9596 6334 9648
rect 1673 9571 1731 9577
rect 1673 9537 1685 9571
rect 1719 9568 1731 9571
rect 1719 9540 2268 9568
rect 1719 9537 1731 9540
rect 1673 9531 1731 9537
rect 1302 9460 1308 9512
rect 1360 9500 1366 9512
rect 2133 9503 2191 9509
rect 2133 9500 2145 9503
rect 1360 9472 2145 9500
rect 1360 9460 1366 9472
rect 2133 9469 2145 9472
rect 2179 9469 2191 9503
rect 2240 9500 2268 9540
rect 4614 9528 4620 9580
rect 4672 9568 4678 9580
rect 5721 9571 5779 9577
rect 5721 9568 5733 9571
rect 4672 9540 5733 9568
rect 4672 9528 4678 9540
rect 5721 9537 5733 9540
rect 5767 9568 5779 9571
rect 6472 9568 6500 9676
rect 7098 9664 7104 9676
rect 7156 9664 7162 9716
rect 11330 9664 11336 9716
rect 11388 9704 11394 9716
rect 11517 9707 11575 9713
rect 11517 9704 11529 9707
rect 11388 9676 11529 9704
rect 11388 9664 11394 9676
rect 11517 9673 11529 9676
rect 11563 9704 11575 9707
rect 12161 9707 12219 9713
rect 12161 9704 12173 9707
rect 11563 9676 12173 9704
rect 11563 9673 11575 9676
rect 11517 9667 11575 9673
rect 12161 9673 12173 9676
rect 12207 9673 12219 9707
rect 12161 9667 12219 9673
rect 5767 9540 6500 9568
rect 8113 9571 8171 9577
rect 5767 9537 5779 9540
rect 5721 9531 5779 9537
rect 8113 9537 8125 9571
rect 8159 9568 8171 9571
rect 8478 9568 8484 9580
rect 8159 9540 8484 9568
rect 8159 9537 8171 9540
rect 8113 9531 8171 9537
rect 8478 9528 8484 9540
rect 8536 9528 8542 9580
rect 12176 9568 12204 9667
rect 12802 9664 12808 9716
rect 12860 9704 12866 9716
rect 13449 9707 13507 9713
rect 13449 9704 13461 9707
rect 12860 9676 13461 9704
rect 12860 9664 12866 9676
rect 13449 9673 13461 9676
rect 13495 9673 13507 9707
rect 13814 9704 13820 9716
rect 13775 9676 13820 9704
rect 13449 9667 13507 9673
rect 13814 9664 13820 9676
rect 13872 9664 13878 9716
rect 13998 9704 14004 9716
rect 13959 9676 14004 9704
rect 13998 9664 14004 9676
rect 14056 9664 14062 9716
rect 14458 9664 14464 9716
rect 14516 9704 14522 9716
rect 14516 9676 14964 9704
rect 14516 9664 14522 9676
rect 14936 9648 14964 9676
rect 15654 9664 15660 9716
rect 15712 9704 15718 9716
rect 15838 9704 15844 9716
rect 15712 9676 15844 9704
rect 15712 9664 15718 9676
rect 15838 9664 15844 9676
rect 15896 9664 15902 9716
rect 16482 9664 16488 9716
rect 16540 9704 16546 9716
rect 16850 9704 16856 9716
rect 16540 9676 16856 9704
rect 16540 9664 16546 9676
rect 16850 9664 16856 9676
rect 16908 9664 16914 9716
rect 18138 9704 18144 9716
rect 17880 9676 18144 9704
rect 12437 9639 12495 9645
rect 12437 9605 12449 9639
rect 12483 9636 12495 9639
rect 13722 9636 13728 9648
rect 12483 9608 13728 9636
rect 12483 9605 12495 9608
rect 12437 9599 12495 9605
rect 13722 9596 13728 9608
rect 13780 9636 13786 9648
rect 13780 9608 14504 9636
rect 13780 9596 13786 9608
rect 13078 9568 13084 9580
rect 12176 9540 13084 9568
rect 13078 9528 13084 9540
rect 13136 9528 13142 9580
rect 14476 9577 14504 9608
rect 14918 9596 14924 9648
rect 14976 9596 14982 9648
rect 15562 9636 15568 9648
rect 15523 9608 15568 9636
rect 15562 9596 15568 9608
rect 15620 9596 15626 9648
rect 16298 9636 16304 9648
rect 15856 9608 16304 9636
rect 14461 9571 14519 9577
rect 14461 9537 14473 9571
rect 14507 9537 14519 9571
rect 14461 9531 14519 9537
rect 14550 9528 14556 9580
rect 14608 9568 14614 9580
rect 15381 9571 15439 9577
rect 14608 9540 14653 9568
rect 14608 9528 14614 9540
rect 15381 9537 15393 9571
rect 15427 9568 15439 9571
rect 15856 9568 15884 9608
rect 16298 9596 16304 9608
rect 16356 9596 16362 9648
rect 16666 9596 16672 9648
rect 16724 9636 16730 9648
rect 17880 9645 17908 9676
rect 18138 9664 18144 9676
rect 18196 9664 18202 9716
rect 19150 9704 19156 9716
rect 19111 9676 19156 9704
rect 19150 9664 19156 9676
rect 19208 9664 19214 9716
rect 19242 9664 19248 9716
rect 19300 9664 19306 9716
rect 22094 9664 22100 9716
rect 22152 9704 22158 9716
rect 24026 9704 24032 9716
rect 22152 9676 22197 9704
rect 23676 9676 24032 9704
rect 22152 9664 22158 9676
rect 17865 9639 17923 9645
rect 17865 9636 17877 9639
rect 16724 9608 17877 9636
rect 16724 9596 16730 9608
rect 17865 9605 17877 9608
rect 17911 9605 17923 9639
rect 17865 9599 17923 9605
rect 18322 9596 18328 9648
rect 18380 9636 18386 9648
rect 18969 9639 19027 9645
rect 18969 9636 18981 9639
rect 18380 9608 18981 9636
rect 18380 9596 18386 9608
rect 18969 9605 18981 9608
rect 19015 9605 19027 9639
rect 19260 9636 19288 9664
rect 20257 9639 20315 9645
rect 19260 9608 19656 9636
rect 18969 9599 19027 9605
rect 15427 9540 15884 9568
rect 15427 9537 15439 9540
rect 15381 9531 15439 9537
rect 15930 9528 15936 9580
rect 15988 9568 15994 9580
rect 16117 9571 16175 9577
rect 16117 9568 16129 9571
rect 15988 9540 16129 9568
rect 15988 9528 15994 9540
rect 16117 9537 16129 9540
rect 16163 9568 16175 9571
rect 16577 9571 16635 9577
rect 16577 9568 16589 9571
rect 16163 9540 16589 9568
rect 16163 9537 16175 9540
rect 16117 9531 16175 9537
rect 16577 9537 16589 9540
rect 16623 9537 16635 9571
rect 16577 9531 16635 9537
rect 2958 9500 2964 9512
rect 2240 9472 2964 9500
rect 2133 9463 2191 9469
rect 2958 9460 2964 9472
rect 3016 9460 3022 9512
rect 5626 9500 5632 9512
rect 5587 9472 5632 9500
rect 5626 9460 5632 9472
rect 5684 9460 5690 9512
rect 7377 9503 7435 9509
rect 7377 9469 7389 9503
rect 7423 9500 7435 9503
rect 7837 9503 7895 9509
rect 7837 9500 7849 9503
rect 7423 9472 7849 9500
rect 7423 9469 7435 9472
rect 7377 9463 7435 9469
rect 7837 9469 7849 9472
rect 7883 9500 7895 9503
rect 7926 9500 7932 9512
rect 7883 9472 7932 9500
rect 7883 9469 7895 9472
rect 7837 9463 7895 9469
rect 7926 9460 7932 9472
rect 7984 9460 7990 9512
rect 8938 9500 8944 9512
rect 8899 9472 8944 9500
rect 8938 9460 8944 9472
rect 8996 9460 9002 9512
rect 9033 9503 9091 9509
rect 9033 9469 9045 9503
rect 9079 9500 9091 9503
rect 9300 9503 9358 9509
rect 9079 9472 9260 9500
rect 9079 9469 9091 9472
rect 9033 9463 9091 9469
rect 9232 9444 9260 9472
rect 9300 9469 9312 9503
rect 9346 9500 9358 9503
rect 9582 9500 9588 9512
rect 9346 9472 9588 9500
rect 9346 9469 9358 9472
rect 9300 9463 9358 9469
rect 9582 9460 9588 9472
rect 9640 9460 9646 9512
rect 12434 9460 12440 9512
rect 12492 9500 12498 9512
rect 12805 9503 12863 9509
rect 12805 9500 12817 9503
rect 12492 9472 12817 9500
rect 12492 9460 12498 9472
rect 12805 9469 12817 9472
rect 12851 9500 12863 9503
rect 13446 9500 13452 9512
rect 12851 9472 13452 9500
rect 12851 9469 12863 9472
rect 12805 9463 12863 9469
rect 13446 9460 13452 9472
rect 13504 9460 13510 9512
rect 15838 9460 15844 9512
rect 15896 9500 15902 9512
rect 16025 9503 16083 9509
rect 16025 9500 16037 9503
rect 15896 9472 16037 9500
rect 15896 9460 15902 9472
rect 16025 9469 16037 9472
rect 16071 9500 16083 9503
rect 16945 9503 17003 9509
rect 16945 9500 16957 9503
rect 16071 9472 16957 9500
rect 16071 9469 16083 9472
rect 16025 9463 16083 9469
rect 16945 9469 16957 9472
rect 16991 9469 17003 9503
rect 16945 9463 17003 9469
rect 17310 9460 17316 9512
rect 17368 9509 17374 9512
rect 17368 9500 17379 9509
rect 18049 9503 18107 9509
rect 17368 9472 17413 9500
rect 17368 9463 17379 9472
rect 18049 9469 18061 9503
rect 18095 9500 18107 9503
rect 18230 9500 18236 9512
rect 18095 9472 18236 9500
rect 18095 9469 18107 9472
rect 18049 9463 18107 9469
rect 17368 9460 17374 9463
rect 18230 9460 18236 9472
rect 18288 9500 18294 9512
rect 18601 9503 18659 9509
rect 18601 9500 18613 9503
rect 18288 9472 18613 9500
rect 18288 9460 18294 9472
rect 18601 9469 18613 9472
rect 18647 9469 18659 9503
rect 18984 9500 19012 9599
rect 19628 9577 19656 9608
rect 20257 9605 20269 9639
rect 20303 9636 20315 9639
rect 20622 9636 20628 9648
rect 20303 9608 20628 9636
rect 20303 9605 20315 9608
rect 20257 9599 20315 9605
rect 19613 9571 19671 9577
rect 19613 9537 19625 9571
rect 19659 9537 19671 9571
rect 19613 9531 19671 9537
rect 19797 9571 19855 9577
rect 19797 9537 19809 9571
rect 19843 9568 19855 9571
rect 20272 9568 20300 9599
rect 20622 9596 20628 9608
rect 20680 9596 20686 9648
rect 23109 9639 23167 9645
rect 23109 9605 23121 9639
rect 23155 9636 23167 9639
rect 23382 9636 23388 9648
rect 23155 9608 23388 9636
rect 23155 9605 23167 9608
rect 23109 9599 23167 9605
rect 23382 9596 23388 9608
rect 23440 9596 23446 9648
rect 19843 9540 20300 9568
rect 23676 9568 23704 9676
rect 24026 9664 24032 9676
rect 24084 9664 24090 9716
rect 25590 9704 25596 9716
rect 25551 9676 25596 9704
rect 25590 9664 25596 9676
rect 25648 9664 25654 9716
rect 24854 9596 24860 9648
rect 24912 9636 24918 9648
rect 25041 9639 25099 9645
rect 25041 9636 25053 9639
rect 24912 9608 25053 9636
rect 24912 9596 24918 9608
rect 25041 9605 25053 9608
rect 25087 9605 25099 9639
rect 26418 9636 26424 9648
rect 26379 9608 26424 9636
rect 25041 9599 25099 9605
rect 26418 9596 26424 9608
rect 26476 9596 26482 9648
rect 23676 9540 23796 9568
rect 19843 9537 19855 9540
rect 19797 9531 19855 9537
rect 19521 9503 19579 9509
rect 19521 9500 19533 9503
rect 18984 9472 19533 9500
rect 18601 9463 18659 9469
rect 19521 9469 19533 9472
rect 19567 9469 19579 9503
rect 20714 9500 20720 9512
rect 20675 9472 20720 9500
rect 19521 9463 19579 9469
rect 20714 9460 20720 9472
rect 20772 9460 20778 9512
rect 22646 9460 22652 9512
rect 22704 9500 22710 9512
rect 22741 9503 22799 9509
rect 22741 9500 22753 9503
rect 22704 9472 22753 9500
rect 22704 9460 22710 9472
rect 22741 9469 22753 9472
rect 22787 9500 22799 9503
rect 23106 9500 23112 9512
rect 22787 9472 23112 9500
rect 22787 9469 22799 9472
rect 22741 9463 22799 9469
rect 23106 9460 23112 9472
rect 23164 9460 23170 9512
rect 23661 9503 23719 9509
rect 23661 9500 23673 9503
rect 23308 9472 23673 9500
rect 2314 9392 2320 9444
rect 2372 9441 2378 9444
rect 2372 9435 2436 9441
rect 2372 9401 2390 9435
rect 2424 9401 2436 9435
rect 2372 9395 2436 9401
rect 2372 9392 2378 9395
rect 6086 9392 6092 9444
rect 6144 9432 6150 9444
rect 6641 9435 6699 9441
rect 6641 9432 6653 9435
rect 6144 9404 6653 9432
rect 6144 9392 6150 9404
rect 6641 9401 6653 9404
rect 6687 9432 6699 9435
rect 6687 9404 7604 9432
rect 6687 9401 6699 9404
rect 6641 9395 6699 9401
rect 7576 9376 7604 9404
rect 9214 9392 9220 9444
rect 9272 9392 9278 9444
rect 15010 9392 15016 9444
rect 15068 9432 15074 9444
rect 15286 9432 15292 9444
rect 15068 9404 15292 9432
rect 15068 9392 15074 9404
rect 15286 9392 15292 9404
rect 15344 9432 15350 9444
rect 15344 9404 17172 9432
rect 15344 9392 15350 9404
rect 3513 9367 3571 9373
rect 3513 9333 3525 9367
rect 3559 9364 3571 9367
rect 3602 9364 3608 9376
rect 3559 9336 3608 9364
rect 3559 9333 3571 9336
rect 3513 9327 3571 9333
rect 3602 9324 3608 9336
rect 3660 9324 3666 9376
rect 4157 9367 4215 9373
rect 4157 9333 4169 9367
rect 4203 9364 4215 9367
rect 4798 9364 4804 9376
rect 4203 9336 4804 9364
rect 4203 9333 4215 9336
rect 4157 9327 4215 9333
rect 4798 9324 4804 9336
rect 4856 9324 4862 9376
rect 5077 9367 5135 9373
rect 5077 9333 5089 9367
rect 5123 9364 5135 9367
rect 5534 9364 5540 9376
rect 5123 9336 5540 9364
rect 5123 9333 5135 9336
rect 5077 9327 5135 9333
rect 5534 9324 5540 9336
rect 5592 9324 5598 9376
rect 7466 9364 7472 9376
rect 7427 9336 7472 9364
rect 7466 9324 7472 9336
rect 7524 9324 7530 9376
rect 7558 9324 7564 9376
rect 7616 9364 7622 9376
rect 7929 9367 7987 9373
rect 7929 9364 7941 9367
rect 7616 9336 7941 9364
rect 7616 9324 7622 9336
rect 7929 9333 7941 9336
rect 7975 9333 7987 9367
rect 8478 9364 8484 9376
rect 8439 9336 8484 9364
rect 7929 9327 7987 9333
rect 8478 9324 8484 9336
rect 8536 9324 8542 9376
rect 8570 9324 8576 9376
rect 8628 9364 8634 9376
rect 8938 9364 8944 9376
rect 8628 9336 8944 9364
rect 8628 9324 8634 9336
rect 8938 9324 8944 9336
rect 8996 9324 9002 9376
rect 9398 9324 9404 9376
rect 9456 9364 9462 9376
rect 10413 9367 10471 9373
rect 10413 9364 10425 9367
rect 9456 9336 10425 9364
rect 9456 9324 9462 9336
rect 10413 9333 10425 9336
rect 10459 9364 10471 9367
rect 10686 9364 10692 9376
rect 10459 9336 10692 9364
rect 10459 9333 10471 9336
rect 10413 9327 10471 9333
rect 10686 9324 10692 9336
rect 10744 9324 10750 9376
rect 11054 9364 11060 9376
rect 10967 9336 11060 9364
rect 11054 9324 11060 9336
rect 11112 9364 11118 9376
rect 12066 9364 12072 9376
rect 11112 9336 12072 9364
rect 11112 9324 11118 9336
rect 12066 9324 12072 9336
rect 12124 9324 12130 9376
rect 12894 9364 12900 9376
rect 12855 9336 12900 9364
rect 12894 9324 12900 9336
rect 12952 9324 12958 9376
rect 13814 9324 13820 9376
rect 13872 9364 13878 9376
rect 14369 9367 14427 9373
rect 14369 9364 14381 9367
rect 13872 9336 14381 9364
rect 13872 9324 13878 9336
rect 14369 9333 14381 9336
rect 14415 9364 14427 9367
rect 14642 9364 14648 9376
rect 14415 9336 14648 9364
rect 14415 9333 14427 9336
rect 14369 9327 14427 9333
rect 14642 9324 14648 9336
rect 14700 9324 14706 9376
rect 15194 9324 15200 9376
rect 15252 9364 15258 9376
rect 17144 9373 17172 9404
rect 17862 9392 17868 9444
rect 17920 9432 17926 9444
rect 19426 9432 19432 9444
rect 17920 9404 19432 9432
rect 17920 9392 17926 9404
rect 19426 9392 19432 9404
rect 19484 9392 19490 9444
rect 19978 9392 19984 9444
rect 20036 9432 20042 9444
rect 20962 9435 21020 9441
rect 20962 9432 20974 9435
rect 20036 9404 20974 9432
rect 20036 9392 20042 9404
rect 20962 9401 20974 9404
rect 21008 9432 21020 9435
rect 22002 9432 22008 9444
rect 21008 9404 22008 9432
rect 21008 9401 21020 9404
rect 20962 9395 21020 9401
rect 22002 9392 22008 9404
rect 22060 9392 22066 9444
rect 22554 9392 22560 9444
rect 22612 9432 22618 9444
rect 22922 9432 22928 9444
rect 22612 9404 22928 9432
rect 22612 9392 22618 9404
rect 22922 9392 22928 9404
rect 22980 9392 22986 9444
rect 15933 9367 15991 9373
rect 15933 9364 15945 9367
rect 15252 9336 15945 9364
rect 15252 9324 15258 9336
rect 15933 9333 15945 9336
rect 15979 9333 15991 9367
rect 15933 9327 15991 9333
rect 17129 9367 17187 9373
rect 17129 9333 17141 9367
rect 17175 9364 17187 9367
rect 17494 9364 17500 9376
rect 17175 9336 17500 9364
rect 17175 9333 17187 9336
rect 17129 9327 17187 9333
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 18138 9324 18144 9376
rect 18196 9364 18202 9376
rect 18233 9367 18291 9373
rect 18233 9364 18245 9367
rect 18196 9336 18245 9364
rect 18196 9324 18202 9336
rect 18233 9333 18245 9336
rect 18279 9333 18291 9367
rect 18233 9327 18291 9333
rect 20806 9324 20812 9376
rect 20864 9364 20870 9376
rect 23308 9364 23336 9472
rect 23661 9469 23673 9472
rect 23707 9500 23719 9503
rect 23768 9500 23796 9540
rect 25590 9528 25596 9580
rect 25648 9568 25654 9580
rect 25958 9568 25964 9580
rect 25648 9540 25964 9568
rect 25648 9528 25654 9540
rect 25958 9528 25964 9540
rect 26016 9528 26022 9580
rect 23707 9472 23796 9500
rect 23928 9503 23986 9509
rect 23707 9469 23719 9472
rect 23661 9463 23719 9469
rect 23928 9469 23940 9503
rect 23974 9500 23986 9503
rect 24762 9500 24768 9512
rect 23974 9472 24768 9500
rect 23974 9469 23986 9472
rect 23928 9463 23986 9469
rect 24762 9460 24768 9472
rect 24820 9460 24826 9512
rect 23477 9435 23535 9441
rect 23477 9401 23489 9435
rect 23523 9432 23535 9435
rect 25774 9432 25780 9444
rect 23523 9404 25780 9432
rect 23523 9401 23535 9404
rect 23477 9395 23535 9401
rect 23952 9376 23980 9404
rect 25774 9392 25780 9404
rect 25832 9392 25838 9444
rect 20864 9336 23336 9364
rect 20864 9324 20870 9336
rect 23934 9324 23940 9376
rect 23992 9324 23998 9376
rect 25314 9324 25320 9376
rect 25372 9364 25378 9376
rect 25961 9367 26019 9373
rect 25961 9364 25973 9367
rect 25372 9336 25973 9364
rect 25372 9324 25378 9336
rect 25961 9333 25973 9336
rect 26007 9333 26019 9367
rect 25961 9327 26019 9333
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1397 9163 1455 9169
rect 1397 9129 1409 9163
rect 1443 9160 1455 9163
rect 1854 9160 1860 9172
rect 1443 9132 1860 9160
rect 1443 9129 1455 9132
rect 1397 9123 1455 9129
rect 1854 9120 1860 9132
rect 1912 9120 1918 9172
rect 2225 9163 2283 9169
rect 2225 9129 2237 9163
rect 2271 9160 2283 9163
rect 2314 9160 2320 9172
rect 2271 9132 2320 9160
rect 2271 9129 2283 9132
rect 2225 9123 2283 9129
rect 2314 9120 2320 9132
rect 2372 9120 2378 9172
rect 2869 9163 2927 9169
rect 2869 9129 2881 9163
rect 2915 9160 2927 9163
rect 3878 9160 3884 9172
rect 2915 9132 3884 9160
rect 2915 9129 2927 9132
rect 2869 9123 2927 9129
rect 3878 9120 3884 9132
rect 3936 9120 3942 9172
rect 4062 9160 4068 9172
rect 4023 9132 4068 9160
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 4154 9120 4160 9172
rect 4212 9160 4218 9172
rect 4706 9160 4712 9172
rect 4212 9132 4712 9160
rect 4212 9120 4218 9132
rect 4706 9120 4712 9132
rect 4764 9120 4770 9172
rect 5261 9163 5319 9169
rect 5261 9129 5273 9163
rect 5307 9160 5319 9163
rect 5626 9160 5632 9172
rect 5307 9132 5632 9160
rect 5307 9129 5319 9132
rect 5261 9123 5319 9129
rect 5626 9120 5632 9132
rect 5684 9120 5690 9172
rect 9125 9163 9183 9169
rect 9125 9129 9137 9163
rect 9171 9160 9183 9163
rect 9398 9160 9404 9172
rect 9171 9132 9404 9160
rect 9171 9129 9183 9132
rect 9125 9123 9183 9129
rect 9398 9120 9404 9132
rect 9456 9160 9462 9172
rect 9582 9160 9588 9172
rect 9456 9132 9588 9160
rect 9456 9120 9462 9132
rect 9582 9120 9588 9132
rect 9640 9120 9646 9172
rect 9950 9120 9956 9172
rect 10008 9160 10014 9172
rect 10045 9163 10103 9169
rect 10045 9160 10057 9163
rect 10008 9132 10057 9160
rect 10008 9120 10014 9132
rect 10045 9129 10057 9132
rect 10091 9129 10103 9163
rect 10045 9123 10103 9129
rect 10873 9163 10931 9169
rect 10873 9129 10885 9163
rect 10919 9160 10931 9163
rect 11238 9160 11244 9172
rect 10919 9132 11244 9160
rect 10919 9129 10931 9132
rect 10873 9123 10931 9129
rect 3326 9052 3332 9104
rect 3384 9092 3390 9104
rect 6362 9101 6368 9104
rect 4433 9095 4491 9101
rect 4433 9092 4445 9095
rect 3384 9064 4445 9092
rect 3384 9052 3390 9064
rect 4433 9061 4445 9064
rect 4479 9061 4491 9095
rect 6356 9092 6368 9101
rect 6275 9064 6368 9092
rect 4433 9055 4491 9061
rect 6356 9055 6368 9064
rect 6420 9092 6426 9104
rect 9306 9092 9312 9104
rect 6420 9064 9312 9092
rect 6362 9052 6368 9055
rect 6420 9052 6426 9064
rect 9306 9052 9312 9064
rect 9364 9052 9370 9104
rect 9490 9092 9496 9104
rect 9451 9064 9496 9092
rect 9490 9052 9496 9064
rect 9548 9052 9554 9104
rect 10060 9092 10088 9123
rect 11238 9120 11244 9132
rect 11296 9160 11302 9172
rect 11790 9160 11796 9172
rect 11296 9132 11796 9160
rect 11296 9120 11302 9132
rect 11790 9120 11796 9132
rect 11848 9120 11854 9172
rect 13722 9120 13728 9172
rect 13780 9160 13786 9172
rect 14645 9163 14703 9169
rect 14645 9160 14657 9163
rect 13780 9132 14657 9160
rect 13780 9120 13786 9132
rect 14645 9129 14657 9132
rect 14691 9129 14703 9163
rect 14645 9123 14703 9129
rect 14918 9120 14924 9172
rect 14976 9160 14982 9172
rect 15838 9160 15844 9172
rect 14976 9132 15844 9160
rect 14976 9120 14982 9132
rect 15838 9120 15844 9132
rect 15896 9120 15902 9172
rect 19978 9160 19984 9172
rect 17880 9132 19104 9160
rect 19939 9132 19984 9160
rect 11149 9095 11207 9101
rect 11149 9092 11161 9095
rect 10060 9064 11161 9092
rect 11149 9061 11161 9064
rect 11195 9061 11207 9095
rect 11149 9055 11207 9061
rect 14734 9052 14740 9104
rect 14792 9092 14798 9104
rect 16298 9092 16304 9104
rect 14792 9064 16304 9092
rect 14792 9052 14798 9064
rect 16298 9052 16304 9064
rect 16356 9052 16362 9104
rect 17310 9092 17316 9104
rect 17223 9064 17316 9092
rect 17310 9052 17316 9064
rect 17368 9092 17374 9104
rect 17880 9092 17908 9132
rect 17368 9064 17908 9092
rect 18224 9095 18282 9101
rect 17368 9052 17374 9064
rect 18224 9061 18236 9095
rect 18270 9092 18282 9095
rect 18966 9092 18972 9104
rect 18270 9064 18972 9092
rect 18270 9061 18282 9064
rect 18224 9055 18282 9061
rect 18966 9052 18972 9064
rect 19024 9052 19030 9104
rect 19076 9092 19104 9132
rect 19978 9120 19984 9132
rect 20036 9160 20042 9172
rect 20257 9163 20315 9169
rect 20257 9160 20269 9163
rect 20036 9132 20269 9160
rect 20036 9120 20042 9132
rect 20257 9129 20269 9132
rect 20303 9129 20315 9163
rect 21358 9160 21364 9172
rect 21319 9132 21364 9160
rect 20257 9123 20315 9129
rect 21358 9120 21364 9132
rect 21416 9120 21422 9172
rect 22925 9163 22983 9169
rect 22925 9129 22937 9163
rect 22971 9160 22983 9163
rect 23014 9160 23020 9172
rect 22971 9132 23020 9160
rect 22971 9129 22983 9132
rect 22925 9123 22983 9129
rect 23014 9120 23020 9132
rect 23072 9120 23078 9172
rect 23474 9160 23480 9172
rect 23435 9132 23480 9160
rect 23474 9120 23480 9132
rect 23532 9120 23538 9172
rect 24118 9120 24124 9172
rect 24176 9160 24182 9172
rect 24489 9163 24547 9169
rect 24489 9160 24501 9163
rect 24176 9132 24501 9160
rect 24176 9120 24182 9132
rect 24489 9129 24501 9132
rect 24535 9129 24547 9163
rect 24489 9123 24547 9129
rect 25314 9120 25320 9172
rect 25372 9160 25378 9172
rect 25409 9163 25467 9169
rect 25409 9160 25421 9163
rect 25372 9132 25421 9160
rect 25372 9120 25378 9132
rect 25409 9129 25421 9132
rect 25455 9160 25467 9163
rect 25777 9163 25835 9169
rect 25777 9160 25789 9163
rect 25455 9132 25789 9160
rect 25455 9129 25467 9132
rect 25409 9123 25467 9129
rect 25777 9129 25789 9132
rect 25823 9160 25835 9163
rect 26142 9160 26148 9172
rect 25823 9132 26148 9160
rect 25823 9129 25835 9132
rect 25777 9123 25835 9129
rect 26142 9120 26148 9132
rect 26200 9120 26206 9172
rect 26237 9163 26295 9169
rect 26237 9129 26249 9163
rect 26283 9160 26295 9163
rect 26418 9160 26424 9172
rect 26283 9132 26424 9160
rect 26283 9129 26295 9132
rect 26237 9123 26295 9129
rect 26418 9120 26424 9132
rect 26476 9120 26482 9172
rect 22281 9095 22339 9101
rect 22281 9092 22293 9095
rect 19076 9064 22293 9092
rect 2774 8984 2780 9036
rect 2832 9024 2838 9036
rect 3881 9027 3939 9033
rect 2832 8996 2877 9024
rect 2832 8984 2838 8996
rect 3881 8993 3893 9027
rect 3927 9024 3939 9027
rect 3970 9024 3976 9036
rect 3927 8996 3976 9024
rect 3927 8993 3939 8996
rect 3881 8987 3939 8993
rect 3970 8984 3976 8996
rect 4028 8984 4034 9036
rect 5074 9024 5080 9036
rect 4540 8996 5080 9024
rect 2958 8956 2964 8968
rect 2919 8928 2964 8956
rect 2958 8916 2964 8928
rect 3016 8916 3022 8968
rect 4154 8916 4160 8968
rect 4212 8956 4218 8968
rect 4540 8965 4568 8996
rect 5074 8984 5080 8996
rect 5132 8984 5138 9036
rect 5997 9027 6055 9033
rect 5997 8993 6009 9027
rect 6043 9024 6055 9027
rect 6178 9024 6184 9036
rect 6043 8996 6184 9024
rect 6043 8993 6055 8996
rect 5997 8987 6055 8993
rect 6178 8984 6184 8996
rect 6236 8984 6242 9036
rect 8113 9027 8171 9033
rect 8113 8993 8125 9027
rect 8159 9024 8171 9027
rect 8478 9024 8484 9036
rect 8159 8996 8484 9024
rect 8159 8993 8171 8996
rect 8113 8987 8171 8993
rect 8478 8984 8484 8996
rect 8536 8984 8542 9036
rect 11330 8984 11336 9036
rect 11388 9024 11394 9036
rect 11773 9027 11831 9033
rect 11773 9024 11785 9027
rect 11388 8996 11785 9024
rect 11388 8984 11394 8996
rect 11773 8993 11785 8996
rect 11819 8993 11831 9027
rect 11773 8987 11831 8993
rect 13906 8984 13912 9036
rect 13964 9024 13970 9036
rect 15562 9033 15568 9036
rect 14093 9027 14151 9033
rect 14093 9024 14105 9027
rect 13964 8996 14105 9024
rect 13964 8984 13970 8996
rect 14093 8993 14105 8996
rect 14139 8993 14151 9027
rect 15556 9024 15568 9033
rect 15523 8996 15568 9024
rect 14093 8987 14151 8993
rect 15556 8987 15568 8996
rect 15562 8984 15568 8987
rect 15620 8984 15626 9036
rect 17494 8984 17500 9036
rect 17552 9024 17558 9036
rect 20640 9033 20668 9064
rect 22281 9061 22293 9064
rect 22327 9061 22339 9095
rect 22281 9055 22339 9061
rect 23290 9052 23296 9104
rect 23348 9092 23354 9104
rect 23845 9095 23903 9101
rect 23845 9092 23857 9095
rect 23348 9064 23857 9092
rect 23348 9052 23354 9064
rect 23845 9061 23857 9064
rect 23891 9061 23903 9095
rect 23845 9055 23903 9061
rect 17957 9027 18015 9033
rect 17957 9024 17969 9027
rect 17552 8996 17969 9024
rect 17552 8984 17558 8996
rect 17957 8993 17969 8996
rect 18003 8993 18015 9027
rect 17957 8987 18015 8993
rect 20625 9027 20683 9033
rect 20625 8993 20637 9027
rect 20671 8993 20683 9027
rect 20625 8987 20683 8993
rect 21269 9027 21327 9033
rect 21269 8993 21281 9027
rect 21315 8993 21327 9027
rect 22830 9024 22836 9036
rect 22791 8996 22836 9024
rect 21269 8987 21327 8993
rect 4525 8959 4583 8965
rect 4525 8956 4537 8959
rect 4212 8928 4537 8956
rect 4212 8916 4218 8928
rect 4525 8925 4537 8928
rect 4571 8925 4583 8959
rect 4525 8919 4583 8925
rect 4614 8916 4620 8968
rect 4672 8956 4678 8968
rect 6089 8959 6147 8965
rect 6089 8956 6101 8959
rect 4672 8928 4765 8956
rect 5828 8928 6101 8956
rect 4672 8916 4678 8928
rect 1578 8848 1584 8900
rect 1636 8888 1642 8900
rect 2409 8891 2467 8897
rect 2409 8888 2421 8891
rect 1636 8860 2421 8888
rect 1636 8848 1642 8860
rect 2409 8857 2421 8860
rect 2455 8857 2467 8891
rect 2409 8851 2467 8857
rect 3602 8848 3608 8900
rect 3660 8888 3666 8900
rect 4632 8888 4660 8916
rect 5626 8888 5632 8900
rect 3660 8860 4660 8888
rect 5587 8860 5632 8888
rect 3660 8848 3666 8860
rect 5626 8848 5632 8860
rect 5684 8848 5690 8900
rect 3142 8780 3148 8832
rect 3200 8820 3206 8832
rect 3421 8823 3479 8829
rect 3421 8820 3433 8823
rect 3200 8792 3433 8820
rect 3200 8780 3206 8792
rect 3421 8789 3433 8792
rect 3467 8789 3479 8823
rect 3421 8783 3479 8789
rect 4246 8780 4252 8832
rect 4304 8820 4310 8832
rect 4614 8820 4620 8832
rect 4304 8792 4620 8820
rect 4304 8780 4310 8792
rect 4614 8780 4620 8792
rect 4672 8820 4678 8832
rect 5828 8829 5856 8928
rect 6089 8925 6101 8928
rect 6135 8925 6147 8959
rect 8570 8956 8576 8968
rect 8531 8928 8576 8956
rect 6089 8919 6147 8925
rect 8570 8916 8576 8928
rect 8628 8916 8634 8968
rect 9766 8916 9772 8968
rect 9824 8956 9830 8968
rect 10137 8959 10195 8965
rect 10137 8956 10149 8959
rect 9824 8928 10149 8956
rect 9824 8916 9830 8928
rect 10137 8925 10149 8928
rect 10183 8925 10195 8959
rect 10137 8919 10195 8925
rect 10226 8916 10232 8968
rect 10284 8956 10290 8968
rect 11514 8956 11520 8968
rect 10284 8928 10329 8956
rect 11475 8928 11520 8956
rect 10284 8916 10290 8928
rect 11514 8916 11520 8928
rect 11572 8916 11578 8968
rect 12894 8916 12900 8968
rect 12952 8956 12958 8968
rect 13449 8959 13507 8965
rect 13449 8956 13461 8959
rect 12952 8928 13461 8956
rect 12952 8916 12958 8928
rect 13449 8925 13461 8928
rect 13495 8925 13507 8959
rect 13449 8919 13507 8925
rect 14182 8916 14188 8968
rect 14240 8916 14246 8968
rect 14274 8916 14280 8968
rect 14332 8956 14338 8968
rect 15013 8959 15071 8965
rect 15013 8956 15025 8959
rect 14332 8928 15025 8956
rect 14332 8916 14338 8928
rect 15013 8925 15025 8928
rect 15059 8956 15071 8959
rect 15194 8956 15200 8968
rect 15059 8928 15200 8956
rect 15059 8925 15071 8928
rect 15013 8919 15071 8925
rect 15194 8916 15200 8928
rect 15252 8916 15258 8968
rect 15289 8959 15347 8965
rect 15289 8925 15301 8959
rect 15335 8925 15347 8959
rect 15289 8919 15347 8925
rect 9674 8888 9680 8900
rect 9635 8860 9680 8888
rect 9674 8848 9680 8860
rect 9732 8848 9738 8900
rect 13909 8891 13967 8897
rect 13909 8857 13921 8891
rect 13955 8888 13967 8891
rect 14200 8888 14228 8916
rect 14458 8888 14464 8900
rect 13955 8860 14464 8888
rect 13955 8857 13967 8860
rect 13909 8851 13967 8857
rect 14458 8848 14464 8860
rect 14516 8848 14522 8900
rect 14918 8848 14924 8900
rect 14976 8888 14982 8900
rect 15304 8888 15332 8919
rect 17310 8916 17316 8968
rect 17368 8956 17374 8968
rect 17512 8956 17540 8984
rect 17862 8956 17868 8968
rect 17368 8928 17540 8956
rect 17823 8928 17868 8956
rect 17368 8916 17374 8928
rect 17862 8916 17868 8928
rect 17920 8916 17926 8968
rect 19518 8916 19524 8968
rect 19576 8956 19582 8968
rect 21284 8956 21312 8987
rect 22830 8984 22836 8996
rect 22888 8984 22894 9036
rect 24394 9024 24400 9036
rect 24355 8996 24400 9024
rect 24394 8984 24400 8996
rect 24452 9024 24458 9036
rect 24854 9024 24860 9036
rect 24452 8996 24860 9024
rect 24452 8984 24458 8996
rect 24854 8984 24860 8996
rect 24912 8984 24918 9036
rect 21450 8956 21456 8968
rect 19576 8928 21312 8956
rect 21411 8928 21456 8956
rect 19576 8916 19582 8928
rect 21450 8916 21456 8928
rect 21508 8956 21514 8968
rect 21913 8959 21971 8965
rect 21913 8956 21925 8959
rect 21508 8928 21925 8956
rect 21508 8916 21514 8928
rect 21913 8925 21925 8928
rect 21959 8925 21971 8959
rect 21913 8919 21971 8925
rect 22922 8916 22928 8968
rect 22980 8956 22986 8968
rect 23017 8959 23075 8965
rect 23017 8956 23029 8959
rect 22980 8928 23029 8956
rect 22980 8916 22986 8928
rect 23017 8925 23029 8928
rect 23063 8925 23075 8959
rect 23017 8919 23075 8925
rect 24581 8959 24639 8965
rect 24581 8925 24593 8959
rect 24627 8925 24639 8959
rect 24581 8919 24639 8925
rect 14976 8860 15332 8888
rect 20441 8891 20499 8897
rect 14976 8848 14982 8860
rect 20441 8857 20453 8891
rect 20487 8888 20499 8891
rect 20806 8888 20812 8900
rect 20487 8860 20812 8888
rect 20487 8857 20499 8860
rect 20441 8851 20499 8857
rect 20806 8848 20812 8860
rect 20864 8848 20870 8900
rect 23032 8888 23060 8919
rect 24596 8888 24624 8919
rect 24946 8888 24952 8900
rect 23032 8860 24952 8888
rect 24946 8848 24952 8860
rect 25004 8848 25010 8900
rect 5813 8823 5871 8829
rect 5813 8820 5825 8823
rect 4672 8792 5825 8820
rect 4672 8780 4678 8792
rect 5813 8789 5825 8792
rect 5859 8789 5871 8823
rect 5813 8783 5871 8789
rect 7282 8780 7288 8832
rect 7340 8820 7346 8832
rect 7469 8823 7527 8829
rect 7469 8820 7481 8823
rect 7340 8792 7481 8820
rect 7340 8780 7346 8792
rect 7469 8789 7481 8792
rect 7515 8789 7527 8823
rect 7469 8783 7527 8789
rect 8202 8780 8208 8832
rect 8260 8820 8266 8832
rect 8389 8823 8447 8829
rect 8389 8820 8401 8823
rect 8260 8792 8401 8820
rect 8260 8780 8266 8792
rect 8389 8789 8401 8792
rect 8435 8789 8447 8823
rect 8389 8783 8447 8789
rect 12897 8823 12955 8829
rect 12897 8789 12909 8823
rect 12943 8820 12955 8823
rect 13078 8820 13084 8832
rect 12943 8792 13084 8820
rect 12943 8789 12955 8792
rect 12897 8783 12955 8789
rect 13078 8780 13084 8792
rect 13136 8820 13142 8832
rect 13722 8820 13728 8832
rect 13136 8792 13728 8820
rect 13136 8780 13142 8792
rect 13722 8780 13728 8792
rect 13780 8780 13786 8832
rect 14182 8780 14188 8832
rect 14240 8820 14246 8832
rect 14277 8823 14335 8829
rect 14277 8820 14289 8823
rect 14240 8792 14289 8820
rect 14240 8780 14246 8792
rect 14277 8789 14289 8792
rect 14323 8789 14335 8823
rect 14277 8783 14335 8789
rect 16298 8780 16304 8832
rect 16356 8820 16362 8832
rect 16669 8823 16727 8829
rect 16669 8820 16681 8823
rect 16356 8792 16681 8820
rect 16356 8780 16362 8792
rect 16669 8789 16681 8792
rect 16715 8820 16727 8823
rect 17862 8820 17868 8832
rect 16715 8792 17868 8820
rect 16715 8789 16727 8792
rect 16669 8783 16727 8789
rect 17862 8780 17868 8792
rect 17920 8780 17926 8832
rect 18230 8780 18236 8832
rect 18288 8820 18294 8832
rect 19337 8823 19395 8829
rect 19337 8820 19349 8823
rect 18288 8792 19349 8820
rect 18288 8780 18294 8792
rect 19337 8789 19349 8792
rect 19383 8789 19395 8823
rect 20898 8820 20904 8832
rect 20859 8792 20904 8820
rect 19337 8783 19395 8789
rect 20898 8780 20904 8792
rect 20956 8780 20962 8832
rect 22462 8820 22468 8832
rect 22423 8792 22468 8820
rect 22462 8780 22468 8792
rect 22520 8780 22526 8832
rect 23934 8780 23940 8832
rect 23992 8820 23998 8832
rect 24029 8823 24087 8829
rect 24029 8820 24041 8823
rect 23992 8792 24041 8820
rect 23992 8780 23998 8792
rect 24029 8789 24041 8792
rect 24075 8789 24087 8823
rect 24029 8783 24087 8789
rect 24118 8780 24124 8832
rect 24176 8820 24182 8832
rect 25041 8823 25099 8829
rect 25041 8820 25053 8823
rect 24176 8792 25053 8820
rect 24176 8780 24182 8792
rect 25041 8789 25053 8792
rect 25087 8789 25099 8823
rect 25041 8783 25099 8789
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 2682 8616 2688 8628
rect 2643 8588 2688 8616
rect 2682 8576 2688 8588
rect 2740 8576 2746 8628
rect 4890 8616 4896 8628
rect 2976 8588 4896 8616
rect 2976 8560 3004 8588
rect 4890 8576 4896 8588
rect 4948 8616 4954 8628
rect 5629 8619 5687 8625
rect 5629 8616 5641 8619
rect 4948 8588 5641 8616
rect 4948 8576 4954 8588
rect 5629 8585 5641 8588
rect 5675 8585 5687 8619
rect 5629 8579 5687 8585
rect 6273 8619 6331 8625
rect 6273 8585 6285 8619
rect 6319 8616 6331 8619
rect 6362 8616 6368 8628
rect 6319 8588 6368 8616
rect 6319 8585 6331 8588
rect 6273 8579 6331 8585
rect 6362 8576 6368 8588
rect 6420 8576 6426 8628
rect 7282 8576 7288 8628
rect 7340 8616 7346 8628
rect 9309 8619 9367 8625
rect 9309 8616 9321 8619
rect 7340 8588 9321 8616
rect 7340 8576 7346 8588
rect 9309 8585 9321 8588
rect 9355 8616 9367 8619
rect 10226 8616 10232 8628
rect 9355 8588 10232 8616
rect 9355 8585 9367 8588
rect 9309 8579 9367 8585
rect 10226 8576 10232 8588
rect 10284 8576 10290 8628
rect 11790 8616 11796 8628
rect 11751 8588 11796 8616
rect 11790 8576 11796 8588
rect 11848 8576 11854 8628
rect 12437 8619 12495 8625
rect 12437 8585 12449 8619
rect 12483 8616 12495 8619
rect 12894 8616 12900 8628
rect 12483 8588 12900 8616
rect 12483 8585 12495 8588
rect 12437 8579 12495 8585
rect 12894 8576 12900 8588
rect 12952 8576 12958 8628
rect 13906 8616 13912 8628
rect 13867 8588 13912 8616
rect 13906 8576 13912 8588
rect 13964 8576 13970 8628
rect 15378 8616 15384 8628
rect 15339 8588 15384 8616
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 17310 8576 17316 8628
rect 17368 8576 17374 8628
rect 17494 8576 17500 8628
rect 17552 8616 17558 8628
rect 17865 8619 17923 8625
rect 17865 8616 17877 8619
rect 17552 8588 17877 8616
rect 17552 8576 17558 8588
rect 17865 8585 17877 8588
rect 17911 8616 17923 8619
rect 18966 8616 18972 8628
rect 17911 8588 18972 8616
rect 17911 8585 17923 8588
rect 17865 8579 17923 8585
rect 18966 8576 18972 8588
rect 19024 8576 19030 8628
rect 19518 8576 19524 8628
rect 19576 8616 19582 8628
rect 19981 8619 20039 8625
rect 19981 8616 19993 8619
rect 19576 8588 19993 8616
rect 19576 8576 19582 8588
rect 19981 8585 19993 8588
rect 20027 8585 20039 8619
rect 20438 8616 20444 8628
rect 20399 8588 20444 8616
rect 19981 8579 20039 8585
rect 20438 8576 20444 8588
rect 20496 8576 20502 8628
rect 21358 8576 21364 8628
rect 21416 8616 21422 8628
rect 21545 8619 21603 8625
rect 21545 8616 21557 8619
rect 21416 8588 21557 8616
rect 21416 8576 21422 8588
rect 21545 8585 21557 8588
rect 21591 8585 21603 8619
rect 21545 8579 21603 8585
rect 22373 8619 22431 8625
rect 22373 8585 22385 8619
rect 22419 8616 22431 8619
rect 23014 8616 23020 8628
rect 22419 8588 23020 8616
rect 22419 8585 22431 8588
rect 22373 8579 22431 8585
rect 23014 8576 23020 8588
rect 23072 8576 23078 8628
rect 23658 8616 23664 8628
rect 23619 8588 23664 8616
rect 23658 8576 23664 8588
rect 23716 8576 23722 8628
rect 24765 8619 24823 8625
rect 24765 8585 24777 8619
rect 24811 8616 24823 8619
rect 24854 8616 24860 8628
rect 24811 8588 24860 8616
rect 24811 8585 24823 8588
rect 24765 8579 24823 8585
rect 24854 8576 24860 8588
rect 24912 8576 24918 8628
rect 24946 8576 24952 8628
rect 25004 8616 25010 8628
rect 25041 8619 25099 8625
rect 25041 8616 25053 8619
rect 25004 8588 25053 8616
rect 25004 8576 25010 8588
rect 25041 8585 25053 8588
rect 25087 8585 25099 8619
rect 26142 8616 26148 8628
rect 26103 8588 26148 8616
rect 25041 8579 25099 8585
rect 26142 8576 26148 8588
rect 26200 8576 26206 8628
rect 2225 8551 2283 8557
rect 2225 8517 2237 8551
rect 2271 8548 2283 8551
rect 2958 8548 2964 8560
rect 2271 8520 2964 8548
rect 2271 8517 2283 8520
rect 2225 8511 2283 8517
rect 2958 8508 2964 8520
rect 3016 8508 3022 8560
rect 7009 8551 7067 8557
rect 7009 8517 7021 8551
rect 7055 8548 7067 8551
rect 7190 8548 7196 8560
rect 7055 8520 7196 8548
rect 7055 8517 7067 8520
rect 7009 8511 7067 8517
rect 7190 8508 7196 8520
rect 7248 8508 7254 8560
rect 12253 8551 12311 8557
rect 12253 8517 12265 8551
rect 12299 8548 12311 8551
rect 12802 8548 12808 8560
rect 12299 8520 12808 8548
rect 12299 8517 12311 8520
rect 12253 8511 12311 8517
rect 12802 8508 12808 8520
rect 12860 8508 12866 8560
rect 13924 8548 13952 8576
rect 12912 8520 13952 8548
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8480 1731 8483
rect 2406 8480 2412 8492
rect 1719 8452 2412 8480
rect 1719 8449 1731 8452
rect 1673 8443 1731 8449
rect 2406 8440 2412 8452
rect 2464 8440 2470 8492
rect 2866 8440 2872 8492
rect 2924 8480 2930 8492
rect 3237 8483 3295 8489
rect 3237 8480 3249 8483
rect 2924 8452 3249 8480
rect 2924 8440 2930 8452
rect 3237 8449 3249 8452
rect 3283 8449 3295 8483
rect 3237 8443 3295 8449
rect 3970 8440 3976 8492
rect 4028 8480 4034 8492
rect 8478 8480 8484 8492
rect 4028 8452 4384 8480
rect 4028 8440 4034 8452
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 1578 8412 1584 8424
rect 1443 8384 1584 8412
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 1578 8372 1584 8384
rect 1636 8412 1642 8424
rect 2222 8412 2228 8424
rect 1636 8384 2228 8412
rect 1636 8372 1642 8384
rect 2222 8372 2228 8384
rect 2280 8372 2286 8424
rect 3053 8415 3111 8421
rect 3053 8381 3065 8415
rect 3099 8412 3111 8415
rect 3510 8412 3516 8424
rect 3099 8384 3516 8412
rect 3099 8381 3111 8384
rect 3053 8375 3111 8381
rect 3510 8372 3516 8384
rect 3568 8412 3574 8424
rect 4062 8412 4068 8424
rect 3568 8384 4068 8412
rect 3568 8372 3574 8384
rect 4062 8372 4068 8384
rect 4120 8372 4126 8424
rect 4249 8415 4307 8421
rect 4249 8381 4261 8415
rect 4295 8381 4307 8415
rect 4356 8412 4384 8452
rect 5276 8452 7880 8480
rect 8439 8452 8484 8480
rect 5276 8412 5304 8452
rect 4356 8384 5304 8412
rect 6825 8415 6883 8421
rect 4249 8375 4307 8381
rect 6825 8381 6837 8415
rect 6871 8381 6883 8415
rect 6825 8375 6883 8381
rect 1946 8304 1952 8356
rect 2004 8344 2010 8356
rect 2004 8316 2268 8344
rect 2004 8304 2010 8316
rect 2240 8288 2268 8316
rect 2958 8304 2964 8356
rect 3016 8344 3022 8356
rect 3234 8344 3240 8356
rect 3016 8316 3240 8344
rect 3016 8304 3022 8316
rect 3234 8304 3240 8316
rect 3292 8304 3298 8356
rect 4154 8344 4160 8356
rect 4115 8316 4160 8344
rect 4154 8304 4160 8316
rect 4212 8304 4218 8356
rect 4264 8344 4292 8375
rect 4264 8316 4375 8344
rect 2222 8236 2228 8288
rect 2280 8236 2286 8288
rect 2593 8279 2651 8285
rect 2593 8245 2605 8279
rect 2639 8276 2651 8279
rect 2866 8276 2872 8288
rect 2639 8248 2872 8276
rect 2639 8245 2651 8248
rect 2593 8239 2651 8245
rect 2866 8236 2872 8248
rect 2924 8236 2930 8288
rect 3142 8276 3148 8288
rect 3103 8248 3148 8276
rect 3142 8236 3148 8248
rect 3200 8236 3206 8288
rect 3326 8236 3332 8288
rect 3384 8276 3390 8288
rect 3694 8276 3700 8288
rect 3384 8248 3700 8276
rect 3384 8236 3390 8248
rect 3694 8236 3700 8248
rect 3752 8236 3758 8288
rect 4347 8276 4375 8316
rect 4430 8304 4436 8356
rect 4488 8353 4494 8356
rect 4488 8347 4552 8353
rect 4488 8313 4506 8347
rect 4540 8313 4552 8347
rect 6638 8344 6644 8356
rect 6599 8316 6644 8344
rect 4488 8307 4552 8313
rect 4488 8304 4494 8307
rect 6638 8304 6644 8316
rect 6696 8344 6702 8356
rect 6840 8344 6868 8375
rect 7098 8372 7104 8424
rect 7156 8412 7162 8424
rect 7852 8421 7880 8452
rect 8478 8440 8484 8452
rect 8536 8440 8542 8492
rect 10321 8483 10379 8489
rect 10321 8449 10333 8483
rect 10367 8480 10379 8483
rect 11330 8480 11336 8492
rect 10367 8452 11336 8480
rect 10367 8449 10379 8452
rect 10321 8443 10379 8449
rect 11330 8440 11336 8452
rect 11388 8440 11394 8492
rect 12912 8489 12940 8520
rect 15194 8508 15200 8560
rect 15252 8548 15258 8560
rect 16574 8548 16580 8560
rect 15252 8520 16580 8548
rect 15252 8508 15258 8520
rect 16574 8508 16580 8520
rect 16632 8508 16638 8560
rect 17328 8548 17356 8576
rect 17328 8520 18092 8548
rect 12897 8483 12955 8489
rect 12897 8449 12909 8483
rect 12943 8449 12955 8483
rect 13078 8480 13084 8492
rect 13039 8452 13084 8480
rect 12897 8443 12955 8449
rect 7377 8415 7435 8421
rect 7377 8412 7389 8415
rect 7156 8384 7389 8412
rect 7156 8372 7162 8384
rect 7377 8381 7389 8384
rect 7423 8381 7435 8415
rect 7377 8375 7435 8381
rect 7837 8415 7895 8421
rect 7837 8381 7849 8415
rect 7883 8412 7895 8415
rect 8389 8415 8447 8421
rect 8389 8412 8401 8415
rect 7883 8384 8401 8412
rect 7883 8381 7895 8384
rect 7837 8375 7895 8381
rect 8389 8381 8401 8384
rect 8435 8412 8447 8415
rect 8846 8412 8852 8424
rect 8435 8384 8852 8412
rect 8435 8381 8447 8384
rect 8389 8375 8447 8381
rect 6696 8316 6868 8344
rect 7392 8344 7420 8375
rect 8846 8372 8852 8384
rect 8904 8372 8910 8424
rect 9033 8415 9091 8421
rect 9033 8381 9045 8415
rect 9079 8412 9091 8415
rect 9493 8415 9551 8421
rect 9493 8412 9505 8415
rect 9079 8384 9505 8412
rect 9079 8381 9091 8384
rect 9033 8375 9091 8381
rect 9493 8381 9505 8384
rect 9539 8412 9551 8415
rect 9582 8412 9588 8424
rect 9539 8384 9588 8412
rect 9539 8381 9551 8384
rect 9493 8375 9551 8381
rect 9582 8372 9588 8384
rect 9640 8372 9646 8424
rect 11238 8412 11244 8424
rect 11199 8384 11244 8412
rect 11238 8372 11244 8384
rect 11296 8372 11302 8424
rect 11790 8372 11796 8424
rect 11848 8412 11854 8424
rect 12912 8412 12940 8443
rect 13078 8440 13084 8452
rect 13136 8440 13142 8492
rect 15010 8440 15016 8492
rect 15068 8440 15074 8492
rect 15562 8440 15568 8492
rect 15620 8480 15626 8492
rect 16025 8483 16083 8489
rect 16025 8480 16037 8483
rect 15620 8452 16037 8480
rect 15620 8440 15626 8452
rect 16025 8449 16037 8452
rect 16071 8480 16083 8483
rect 16758 8480 16764 8492
rect 16071 8452 16764 8480
rect 16071 8449 16083 8452
rect 16025 8443 16083 8449
rect 16758 8440 16764 8452
rect 16816 8480 16822 8492
rect 17310 8480 17316 8492
rect 16816 8452 17316 8480
rect 16816 8440 16822 8452
rect 17310 8440 17316 8452
rect 17368 8440 17374 8492
rect 18064 8489 18092 8520
rect 19334 8508 19340 8560
rect 19392 8548 19398 8560
rect 20533 8551 20591 8557
rect 20533 8548 20545 8551
rect 19392 8520 20545 8548
rect 19392 8508 19398 8520
rect 20533 8517 20545 8520
rect 20579 8517 20591 8551
rect 20533 8511 20591 8517
rect 23290 8508 23296 8560
rect 23348 8548 23354 8560
rect 23348 8520 24256 8548
rect 23348 8508 23354 8520
rect 18049 8483 18107 8489
rect 18049 8449 18061 8483
rect 18095 8449 18107 8483
rect 18049 8443 18107 8449
rect 21177 8483 21235 8489
rect 21177 8449 21189 8483
rect 21223 8480 21235 8483
rect 21450 8480 21456 8492
rect 21223 8452 21456 8480
rect 21223 8449 21235 8452
rect 21177 8443 21235 8449
rect 11848 8384 12940 8412
rect 11848 8372 11854 8384
rect 13446 8372 13452 8424
rect 13504 8412 13510 8424
rect 13630 8412 13636 8424
rect 13504 8384 13636 8412
rect 13504 8372 13510 8384
rect 13630 8372 13636 8384
rect 13688 8372 13694 8424
rect 13906 8372 13912 8424
rect 13964 8412 13970 8424
rect 14001 8415 14059 8421
rect 14001 8412 14013 8415
rect 13964 8384 14013 8412
rect 13964 8372 13970 8384
rect 14001 8381 14013 8384
rect 14047 8381 14059 8415
rect 14268 8415 14326 8421
rect 14268 8412 14280 8415
rect 14001 8375 14059 8381
rect 14200 8384 14280 8412
rect 8297 8347 8355 8353
rect 8297 8344 8309 8347
rect 7392 8316 8309 8344
rect 6696 8304 6702 8316
rect 8297 8313 8309 8316
rect 8343 8344 8355 8347
rect 9122 8344 9128 8356
rect 8343 8316 9128 8344
rect 8343 8313 8355 8316
rect 8297 8307 8355 8313
rect 9122 8304 9128 8316
rect 9180 8304 9186 8356
rect 9766 8344 9772 8356
rect 9727 8316 9772 8344
rect 9766 8304 9772 8316
rect 9824 8304 9830 8356
rect 10594 8344 10600 8356
rect 10555 8316 10600 8344
rect 10594 8304 10600 8316
rect 10652 8344 10658 8356
rect 11149 8347 11207 8353
rect 11149 8344 11161 8347
rect 10652 8316 11161 8344
rect 10652 8304 10658 8316
rect 11149 8313 11161 8316
rect 11195 8344 11207 8347
rect 11882 8344 11888 8356
rect 11195 8316 11888 8344
rect 11195 8313 11207 8316
rect 11149 8307 11207 8313
rect 11882 8304 11888 8316
rect 11940 8304 11946 8356
rect 12802 8344 12808 8356
rect 12763 8316 12808 8344
rect 12802 8304 12808 8316
rect 12860 8304 12866 8356
rect 13541 8347 13599 8353
rect 13541 8313 13553 8347
rect 13587 8344 13599 8347
rect 14200 8344 14228 8384
rect 14268 8381 14280 8384
rect 14314 8412 14326 8415
rect 15028 8412 15056 8440
rect 14314 8384 15056 8412
rect 16393 8415 16451 8421
rect 14314 8381 14326 8384
rect 14268 8375 14326 8381
rect 16393 8381 16405 8415
rect 16439 8412 16451 8415
rect 16516 8415 16574 8421
rect 16516 8412 16528 8415
rect 16439 8384 16528 8412
rect 16439 8381 16451 8384
rect 16393 8375 16451 8381
rect 16516 8381 16528 8384
rect 16562 8412 16574 8415
rect 17678 8412 17684 8424
rect 16562 8384 17684 8412
rect 16562 8381 16574 8384
rect 16516 8375 16574 8381
rect 17678 8372 17684 8384
rect 17736 8372 17742 8424
rect 18064 8412 18092 8443
rect 21450 8440 21456 8452
rect 21508 8440 21514 8492
rect 22370 8440 22376 8492
rect 22428 8480 22434 8492
rect 22646 8480 22652 8492
rect 22428 8452 22652 8480
rect 22428 8440 22434 8452
rect 22646 8440 22652 8452
rect 22704 8440 22710 8492
rect 24118 8480 24124 8492
rect 24079 8452 24124 8480
rect 24118 8440 24124 8452
rect 24176 8440 24182 8492
rect 24228 8489 24256 8520
rect 24213 8483 24271 8489
rect 24213 8449 24225 8483
rect 24259 8480 24271 8483
rect 24854 8480 24860 8492
rect 24259 8452 24860 8480
rect 24259 8449 24271 8452
rect 24213 8443 24271 8449
rect 24854 8440 24860 8452
rect 24912 8440 24918 8492
rect 19610 8412 19616 8424
rect 18064 8384 19616 8412
rect 19610 8372 19616 8384
rect 19668 8372 19674 8424
rect 20714 8372 20720 8424
rect 20772 8412 20778 8424
rect 21913 8415 21971 8421
rect 21913 8412 21925 8415
rect 20772 8384 21925 8412
rect 20772 8372 20778 8384
rect 21913 8381 21925 8384
rect 21959 8412 21971 8415
rect 22465 8415 22523 8421
rect 22465 8412 22477 8415
rect 21959 8384 22477 8412
rect 21959 8381 21971 8384
rect 21913 8375 21971 8381
rect 22465 8381 22477 8384
rect 22511 8412 22523 8415
rect 23658 8412 23664 8424
rect 22511 8384 23664 8412
rect 22511 8381 22523 8384
rect 22465 8375 22523 8381
rect 23658 8372 23664 8384
rect 23716 8372 23722 8424
rect 25222 8412 25228 8424
rect 25183 8384 25228 8412
rect 25222 8372 25228 8384
rect 25280 8412 25286 8424
rect 25777 8415 25835 8421
rect 25777 8412 25789 8415
rect 25280 8384 25789 8412
rect 25280 8372 25286 8384
rect 25777 8381 25789 8384
rect 25823 8381 25835 8415
rect 25777 8375 25835 8381
rect 13587 8316 14228 8344
rect 13587 8313 13599 8316
rect 13541 8307 13599 8313
rect 14458 8304 14464 8356
rect 14516 8344 14522 8356
rect 15010 8344 15016 8356
rect 14516 8316 15016 8344
rect 14516 8304 14522 8316
rect 15010 8304 15016 8316
rect 15068 8304 15074 8356
rect 16758 8344 16764 8356
rect 16719 8316 16764 8344
rect 16758 8304 16764 8316
rect 16816 8304 16822 8356
rect 17497 8347 17555 8353
rect 17497 8313 17509 8347
rect 17543 8344 17555 8347
rect 18230 8344 18236 8356
rect 17543 8316 18236 8344
rect 17543 8313 17555 8316
rect 17497 8307 17555 8313
rect 18230 8304 18236 8316
rect 18288 8353 18294 8356
rect 18288 8347 18352 8353
rect 18288 8313 18306 8347
rect 18340 8313 18352 8347
rect 20438 8344 20444 8356
rect 18288 8307 18352 8313
rect 18432 8316 20444 8344
rect 18288 8304 18294 8307
rect 4614 8276 4620 8288
rect 4347 8248 4620 8276
rect 4614 8236 4620 8248
rect 4672 8236 4678 8288
rect 7929 8279 7987 8285
rect 7929 8245 7941 8279
rect 7975 8276 7987 8279
rect 8018 8276 8024 8288
rect 7975 8248 8024 8276
rect 7975 8245 7987 8248
rect 7929 8239 7987 8245
rect 8018 8236 8024 8248
rect 8076 8236 8082 8288
rect 10781 8279 10839 8285
rect 10781 8245 10793 8279
rect 10827 8276 10839 8279
rect 11054 8276 11060 8288
rect 10827 8248 11060 8276
rect 10827 8245 10839 8248
rect 10781 8239 10839 8245
rect 11054 8236 11060 8248
rect 11112 8236 11118 8288
rect 12894 8236 12900 8288
rect 12952 8276 12958 8288
rect 18432 8276 18460 8316
rect 20438 8304 20444 8316
rect 20496 8304 20502 8356
rect 20901 8347 20959 8353
rect 20901 8344 20913 8347
rect 20640 8316 20913 8344
rect 12952 8248 18460 8276
rect 12952 8236 12958 8248
rect 19334 8236 19340 8288
rect 19392 8276 19398 8288
rect 19429 8279 19487 8285
rect 19429 8276 19441 8279
rect 19392 8248 19441 8276
rect 19392 8236 19398 8248
rect 19429 8245 19441 8248
rect 19475 8245 19487 8279
rect 19429 8239 19487 8245
rect 20530 8236 20536 8288
rect 20588 8276 20594 8288
rect 20640 8276 20668 8316
rect 20901 8313 20913 8316
rect 20947 8313 20959 8347
rect 20901 8307 20959 8313
rect 22830 8304 22836 8356
rect 22888 8344 22894 8356
rect 23017 8347 23075 8353
rect 23017 8344 23029 8347
rect 22888 8316 23029 8344
rect 22888 8304 22894 8316
rect 23017 8313 23029 8316
rect 23063 8313 23075 8347
rect 23017 8307 23075 8313
rect 20588 8248 20668 8276
rect 20588 8236 20594 8248
rect 20714 8236 20720 8288
rect 20772 8276 20778 8288
rect 20993 8279 21051 8285
rect 20993 8276 21005 8279
rect 20772 8248 21005 8276
rect 20772 8236 20778 8248
rect 20993 8245 21005 8248
rect 21039 8245 21051 8279
rect 22646 8276 22652 8288
rect 22607 8248 22652 8276
rect 20993 8239 21051 8245
rect 22646 8236 22652 8248
rect 22704 8236 22710 8288
rect 23382 8276 23388 8288
rect 23343 8248 23388 8276
rect 23382 8236 23388 8248
rect 23440 8276 23446 8288
rect 24029 8279 24087 8285
rect 24029 8276 24041 8279
rect 23440 8248 24041 8276
rect 23440 8236 23446 8248
rect 24029 8245 24041 8248
rect 24075 8245 24087 8279
rect 25406 8276 25412 8288
rect 25367 8248 25412 8276
rect 24029 8239 24087 8245
rect 25406 8236 25412 8248
rect 25464 8236 25470 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1394 8032 1400 8084
rect 1452 8072 1458 8084
rect 1670 8072 1676 8084
rect 1452 8044 1676 8072
rect 1452 8032 1458 8044
rect 1670 8032 1676 8044
rect 1728 8032 1734 8084
rect 2314 8032 2320 8084
rect 2372 8072 2378 8084
rect 2777 8075 2835 8081
rect 2777 8072 2789 8075
rect 2372 8044 2789 8072
rect 2372 8032 2378 8044
rect 2777 8041 2789 8044
rect 2823 8041 2835 8075
rect 2777 8035 2835 8041
rect 3602 8032 3608 8084
rect 3660 8072 3666 8084
rect 3789 8075 3847 8081
rect 3789 8072 3801 8075
rect 3660 8044 3801 8072
rect 3660 8032 3666 8044
rect 3789 8041 3801 8044
rect 3835 8041 3847 8075
rect 3789 8035 3847 8041
rect 4341 8075 4399 8081
rect 4341 8041 4353 8075
rect 4387 8072 4399 8075
rect 4430 8072 4436 8084
rect 4387 8044 4436 8072
rect 4387 8041 4399 8044
rect 4341 8035 4399 8041
rect 4430 8032 4436 8044
rect 4488 8032 4494 8084
rect 5077 8075 5135 8081
rect 5077 8041 5089 8075
rect 5123 8072 5135 8075
rect 5442 8072 5448 8084
rect 5123 8044 5448 8072
rect 5123 8041 5135 8044
rect 5077 8035 5135 8041
rect 5442 8032 5448 8044
rect 5500 8032 5506 8084
rect 5534 8032 5540 8084
rect 5592 8072 5598 8084
rect 5810 8072 5816 8084
rect 5592 8044 5816 8072
rect 5592 8032 5598 8044
rect 5810 8032 5816 8044
rect 5868 8032 5874 8084
rect 8386 8072 8392 8084
rect 8347 8044 8392 8072
rect 8386 8032 8392 8044
rect 8444 8032 8450 8084
rect 9306 8032 9312 8084
rect 9364 8072 9370 8084
rect 9401 8075 9459 8081
rect 9401 8072 9413 8075
rect 9364 8044 9413 8072
rect 9364 8032 9370 8044
rect 9401 8041 9413 8044
rect 9447 8041 9459 8075
rect 9401 8035 9459 8041
rect 10505 8075 10563 8081
rect 10505 8041 10517 8075
rect 10551 8072 10563 8075
rect 10686 8072 10692 8084
rect 10551 8044 10692 8072
rect 10551 8041 10563 8044
rect 10505 8035 10563 8041
rect 10686 8032 10692 8044
rect 10744 8032 10750 8084
rect 11330 8072 11336 8084
rect 11291 8044 11336 8072
rect 11330 8032 11336 8044
rect 11388 8072 11394 8084
rect 11701 8075 11759 8081
rect 11701 8072 11713 8075
rect 11388 8044 11713 8072
rect 11388 8032 11394 8044
rect 11701 8041 11713 8044
rect 11747 8041 11759 8075
rect 11701 8035 11759 8041
rect 11885 8075 11943 8081
rect 11885 8041 11897 8075
rect 11931 8072 11943 8075
rect 12342 8072 12348 8084
rect 11931 8044 12348 8072
rect 11931 8041 11943 8044
rect 11885 8035 11943 8041
rect 4706 7964 4712 8016
rect 4764 8004 4770 8016
rect 11716 8004 11744 8035
rect 12342 8032 12348 8044
rect 12400 8032 12406 8084
rect 13078 8072 13084 8084
rect 12452 8044 13084 8072
rect 12452 8004 12480 8044
rect 13078 8032 13084 8044
rect 13136 8072 13142 8084
rect 13265 8075 13323 8081
rect 13265 8072 13277 8075
rect 13136 8044 13277 8072
rect 13136 8032 13142 8044
rect 13265 8041 13277 8044
rect 13311 8041 13323 8075
rect 13265 8035 13323 8041
rect 13449 8075 13507 8081
rect 13449 8041 13461 8075
rect 13495 8072 13507 8075
rect 13814 8072 13820 8084
rect 13495 8044 13820 8072
rect 13495 8041 13507 8044
rect 13449 8035 13507 8041
rect 13814 8032 13820 8044
rect 13872 8032 13878 8084
rect 14458 8072 14464 8084
rect 13924 8044 14464 8072
rect 4764 7976 6500 8004
rect 11716 7976 12480 8004
rect 4764 7964 4770 7976
rect 1664 7939 1722 7945
rect 1664 7905 1676 7939
rect 1710 7936 1722 7939
rect 2866 7936 2872 7948
rect 1710 7908 2872 7936
rect 1710 7905 1722 7908
rect 1664 7899 1722 7905
rect 2866 7896 2872 7908
rect 2924 7896 2930 7948
rect 4522 7896 4528 7948
rect 4580 7936 4586 7948
rect 5169 7939 5227 7945
rect 5169 7936 5181 7939
rect 4580 7908 5181 7936
rect 4580 7896 4586 7908
rect 5169 7905 5181 7908
rect 5215 7936 5227 7939
rect 5258 7936 5264 7948
rect 5215 7908 5264 7936
rect 5215 7905 5227 7908
rect 5169 7899 5227 7905
rect 5258 7896 5264 7908
rect 5316 7896 5322 7948
rect 6472 7936 6500 7976
rect 6733 7939 6791 7945
rect 6733 7936 6745 7939
rect 6472 7908 6745 7936
rect 6472 7880 6500 7908
rect 6733 7905 6745 7908
rect 6779 7905 6791 7939
rect 6733 7899 6791 7905
rect 7282 7896 7288 7948
rect 7340 7936 7346 7948
rect 8297 7939 8355 7945
rect 8297 7936 8309 7939
rect 7340 7908 8309 7936
rect 7340 7896 7346 7908
rect 8297 7905 8309 7908
rect 8343 7905 8355 7939
rect 12250 7936 12256 7948
rect 12211 7908 12256 7936
rect 8297 7899 8355 7905
rect 12250 7896 12256 7908
rect 12308 7896 12314 7948
rect 1394 7868 1400 7880
rect 1355 7840 1400 7868
rect 1394 7828 1400 7840
rect 1452 7828 1458 7880
rect 5350 7868 5356 7880
rect 5311 7840 5356 7868
rect 5350 7828 5356 7840
rect 5408 7828 5414 7880
rect 6454 7828 6460 7880
rect 6512 7828 6518 7880
rect 6822 7868 6828 7880
rect 6783 7840 6828 7868
rect 6822 7828 6828 7840
rect 6880 7828 6886 7880
rect 7009 7871 7067 7877
rect 7009 7837 7021 7871
rect 7055 7868 7067 7871
rect 7098 7868 7104 7880
rect 7055 7840 7104 7868
rect 7055 7837 7067 7840
rect 7009 7831 7067 7837
rect 7098 7828 7104 7840
rect 7156 7828 7162 7880
rect 8478 7868 8484 7880
rect 8439 7840 8484 7868
rect 8478 7828 8484 7840
rect 8536 7828 8542 7880
rect 10597 7871 10655 7877
rect 10597 7837 10609 7871
rect 10643 7837 10655 7871
rect 10597 7831 10655 7837
rect 10781 7871 10839 7877
rect 10781 7837 10793 7871
rect 10827 7868 10839 7871
rect 11054 7868 11060 7880
rect 10827 7840 11060 7868
rect 10827 7837 10839 7840
rect 10781 7831 10839 7837
rect 5074 7760 5080 7812
rect 5132 7800 5138 7812
rect 5368 7800 5396 7828
rect 5132 7772 5396 7800
rect 7653 7803 7711 7809
rect 5132 7760 5138 7772
rect 7653 7769 7665 7803
rect 7699 7800 7711 7803
rect 8110 7800 8116 7812
rect 7699 7772 8116 7800
rect 7699 7769 7711 7772
rect 7653 7763 7711 7769
rect 8110 7760 8116 7772
rect 8168 7760 8174 7812
rect 9766 7760 9772 7812
rect 9824 7800 9830 7812
rect 10612 7800 10640 7831
rect 11054 7828 11060 7840
rect 11112 7828 11118 7880
rect 12342 7868 12348 7880
rect 12303 7840 12348 7868
rect 12342 7828 12348 7840
rect 12400 7828 12406 7880
rect 12452 7877 12480 7976
rect 12989 8007 13047 8013
rect 12989 7973 13001 8007
rect 13035 8004 13047 8007
rect 13170 8004 13176 8016
rect 13035 7976 13176 8004
rect 13035 7973 13047 7976
rect 12989 7967 13047 7973
rect 13170 7964 13176 7976
rect 13228 7964 13234 8016
rect 13924 8004 13952 8044
rect 14458 8032 14464 8044
rect 14516 8032 14522 8084
rect 15286 8072 15292 8084
rect 15247 8044 15292 8072
rect 15286 8032 15292 8044
rect 15344 8032 15350 8084
rect 16298 8032 16304 8084
rect 16356 8072 16362 8084
rect 17681 8075 17739 8081
rect 17681 8072 17693 8075
rect 16356 8044 17693 8072
rect 16356 8032 16362 8044
rect 17681 8041 17693 8044
rect 17727 8072 17739 8075
rect 17770 8072 17776 8084
rect 17727 8044 17776 8072
rect 17727 8041 17739 8044
rect 17681 8035 17739 8041
rect 17770 8032 17776 8044
rect 17828 8032 17834 8084
rect 18782 8072 18788 8084
rect 18743 8044 18788 8072
rect 18782 8032 18788 8044
rect 18840 8032 18846 8084
rect 18966 8032 18972 8084
rect 19024 8072 19030 8084
rect 20257 8075 20315 8081
rect 20257 8072 20269 8075
rect 19024 8044 20269 8072
rect 19024 8032 19030 8044
rect 20257 8041 20269 8044
rect 20303 8072 20315 8075
rect 21450 8072 21456 8084
rect 20303 8044 21456 8072
rect 20303 8041 20315 8044
rect 20257 8035 20315 8041
rect 21450 8032 21456 8044
rect 21508 8032 21514 8084
rect 22922 8072 22928 8084
rect 22883 8044 22928 8072
rect 22922 8032 22928 8044
rect 22980 8032 22986 8084
rect 23290 8072 23296 8084
rect 23251 8044 23296 8072
rect 23290 8032 23296 8044
rect 23348 8032 23354 8084
rect 24026 8072 24032 8084
rect 23987 8044 24032 8072
rect 24026 8032 24032 8044
rect 24084 8032 24090 8084
rect 24210 8032 24216 8084
rect 24268 8072 24274 8084
rect 24489 8075 24547 8081
rect 24489 8072 24501 8075
rect 24268 8044 24501 8072
rect 24268 8032 24274 8044
rect 24489 8041 24501 8044
rect 24535 8041 24547 8075
rect 24489 8035 24547 8041
rect 25961 8075 26019 8081
rect 25961 8041 25973 8075
rect 26007 8072 26019 8075
rect 26142 8072 26148 8084
rect 26007 8044 26148 8072
rect 26007 8041 26019 8044
rect 25961 8035 26019 8041
rect 26142 8032 26148 8044
rect 26200 8032 26206 8084
rect 26329 8075 26387 8081
rect 26329 8041 26341 8075
rect 26375 8072 26387 8075
rect 26418 8072 26424 8084
rect 26375 8044 26424 8072
rect 26375 8041 26387 8044
rect 26329 8035 26387 8041
rect 26418 8032 26424 8044
rect 26476 8032 26482 8084
rect 13832 7976 13952 8004
rect 13630 7896 13636 7948
rect 13688 7936 13694 7948
rect 13832 7945 13860 7976
rect 14090 7964 14096 8016
rect 14148 7964 14154 8016
rect 14921 8007 14979 8013
rect 14921 7973 14933 8007
rect 14967 8004 14979 8007
rect 15010 8004 15016 8016
rect 14967 7976 15016 8004
rect 14967 7973 14979 7976
rect 14921 7967 14979 7973
rect 15010 7964 15016 7976
rect 15068 8004 15074 8016
rect 15841 8007 15899 8013
rect 15841 8004 15853 8007
rect 15068 7976 15853 8004
rect 15068 7964 15074 7976
rect 15841 7973 15853 7976
rect 15887 8004 15899 8007
rect 16209 8007 16267 8013
rect 16209 8004 16221 8007
rect 15887 7976 16221 8004
rect 15887 7973 15899 7976
rect 15841 7967 15899 7973
rect 16209 7973 16221 7976
rect 16255 8004 16267 8007
rect 16390 8004 16396 8016
rect 16255 7976 16396 8004
rect 16255 7973 16267 7976
rect 16209 7967 16267 7973
rect 16390 7964 16396 7976
rect 16448 7964 16454 8016
rect 18322 8004 18328 8016
rect 18283 7976 18328 8004
rect 18322 7964 18328 7976
rect 18380 7964 18386 8016
rect 20070 7964 20076 8016
rect 20128 8004 20134 8016
rect 21168 8007 21226 8013
rect 21168 8004 21180 8007
rect 20128 7976 21180 8004
rect 20128 7964 20134 7976
rect 21168 7973 21180 7976
rect 21214 8004 21226 8007
rect 22002 8004 22008 8016
rect 21214 7976 22008 8004
rect 21214 7973 21226 7976
rect 21168 7967 21226 7973
rect 22002 7964 22008 7976
rect 22060 7964 22066 8016
rect 13817 7939 13875 7945
rect 13817 7936 13829 7939
rect 13688 7908 13829 7936
rect 13688 7896 13694 7908
rect 13817 7905 13829 7908
rect 13863 7905 13875 7939
rect 13817 7899 13875 7905
rect 13906 7896 13912 7948
rect 13964 7936 13970 7948
rect 14108 7936 14136 7964
rect 13964 7908 14009 7936
rect 14108 7908 14228 7936
rect 13964 7896 13970 7908
rect 12437 7871 12495 7877
rect 12437 7837 12449 7871
rect 12483 7837 12495 7871
rect 12437 7831 12495 7837
rect 13722 7828 13728 7880
rect 13780 7868 13786 7880
rect 14090 7868 14096 7880
rect 13780 7840 14096 7868
rect 13780 7828 13786 7840
rect 14090 7828 14096 7840
rect 14148 7828 14154 7880
rect 13078 7800 13084 7812
rect 9824 7772 13084 7800
rect 9824 7760 9830 7772
rect 13078 7760 13084 7772
rect 13136 7760 13142 7812
rect 13814 7760 13820 7812
rect 13872 7800 13878 7812
rect 14200 7800 14228 7908
rect 15562 7896 15568 7948
rect 15620 7936 15626 7948
rect 16557 7939 16615 7945
rect 16557 7936 16569 7939
rect 15620 7908 16569 7936
rect 15620 7896 15626 7908
rect 16557 7905 16569 7908
rect 16603 7936 16615 7939
rect 16603 7908 18828 7936
rect 16603 7905 16615 7908
rect 16557 7899 16615 7905
rect 14918 7828 14924 7880
rect 14976 7868 14982 7880
rect 16301 7871 16359 7877
rect 16301 7868 16313 7871
rect 14976 7840 16313 7868
rect 14976 7828 14982 7840
rect 16301 7837 16313 7840
rect 16347 7837 16359 7871
rect 16301 7831 16359 7837
rect 17678 7828 17684 7880
rect 17736 7868 17742 7880
rect 18414 7868 18420 7880
rect 17736 7840 18420 7868
rect 17736 7828 17742 7840
rect 18414 7828 18420 7840
rect 18472 7828 18478 7880
rect 15654 7800 15660 7812
rect 13872 7772 14228 7800
rect 14283 7772 15660 7800
rect 13872 7760 13878 7772
rect 3326 7732 3332 7744
rect 3287 7704 3332 7732
rect 3326 7692 3332 7704
rect 3384 7692 3390 7744
rect 4430 7692 4436 7744
rect 4488 7732 4494 7744
rect 4709 7735 4767 7741
rect 4709 7732 4721 7735
rect 4488 7704 4721 7732
rect 4488 7692 4494 7704
rect 4709 7701 4721 7704
rect 4755 7701 4767 7735
rect 6086 7732 6092 7744
rect 6047 7704 6092 7732
rect 4709 7695 4767 7701
rect 6086 7692 6092 7704
rect 6144 7692 6150 7744
rect 6365 7735 6423 7741
rect 6365 7701 6377 7735
rect 6411 7732 6423 7735
rect 6914 7732 6920 7744
rect 6411 7704 6920 7732
rect 6411 7701 6423 7704
rect 6365 7695 6423 7701
rect 6914 7692 6920 7704
rect 6972 7692 6978 7744
rect 7926 7732 7932 7744
rect 7839 7704 7932 7732
rect 7926 7692 7932 7704
rect 7984 7732 7990 7744
rect 8941 7735 8999 7741
rect 8941 7732 8953 7735
rect 7984 7704 8953 7732
rect 7984 7692 7990 7704
rect 8941 7701 8953 7704
rect 8987 7701 8999 7735
rect 9950 7732 9956 7744
rect 9911 7704 9956 7732
rect 8941 7695 8999 7701
rect 9950 7692 9956 7704
rect 10008 7692 10014 7744
rect 10042 7692 10048 7744
rect 10100 7732 10106 7744
rect 10137 7735 10195 7741
rect 10137 7732 10149 7735
rect 10100 7704 10149 7732
rect 10100 7692 10106 7704
rect 10137 7701 10149 7704
rect 10183 7701 10195 7735
rect 10137 7695 10195 7701
rect 11882 7692 11888 7744
rect 11940 7732 11946 7744
rect 14283 7732 14311 7772
rect 15654 7760 15660 7772
rect 15712 7760 15718 7812
rect 18800 7800 18828 7908
rect 18874 7896 18880 7948
rect 18932 7936 18938 7948
rect 19153 7939 19211 7945
rect 19153 7936 19165 7939
rect 18932 7908 19165 7936
rect 18932 7896 18938 7908
rect 19153 7905 19165 7908
rect 19199 7936 19211 7939
rect 19797 7939 19855 7945
rect 19797 7936 19809 7939
rect 19199 7908 19809 7936
rect 19199 7905 19211 7908
rect 19153 7899 19211 7905
rect 19797 7905 19809 7908
rect 19843 7905 19855 7939
rect 23382 7936 23388 7948
rect 23343 7908 23388 7936
rect 19797 7899 19855 7905
rect 23382 7896 23388 7908
rect 23440 7896 23446 7948
rect 23566 7896 23572 7948
rect 23624 7936 23630 7948
rect 23750 7936 23756 7948
rect 23624 7908 23756 7936
rect 23624 7896 23630 7908
rect 23750 7896 23756 7908
rect 23808 7896 23814 7948
rect 24857 7939 24915 7945
rect 24857 7905 24869 7939
rect 24903 7936 24915 7939
rect 25222 7936 25228 7948
rect 24903 7908 25228 7936
rect 24903 7905 24915 7908
rect 24857 7899 24915 7905
rect 25222 7896 25228 7908
rect 25280 7896 25286 7948
rect 19242 7868 19248 7880
rect 19203 7840 19248 7868
rect 19242 7828 19248 7840
rect 19300 7828 19306 7880
rect 19334 7828 19340 7880
rect 19392 7868 19398 7880
rect 19392 7840 19437 7868
rect 19392 7828 19398 7840
rect 20806 7828 20812 7880
rect 20864 7868 20870 7880
rect 20901 7871 20959 7877
rect 20901 7868 20913 7871
rect 20864 7840 20913 7868
rect 20864 7828 20870 7840
rect 20901 7837 20913 7840
rect 20947 7837 20959 7871
rect 24946 7868 24952 7880
rect 24907 7840 24952 7868
rect 20901 7831 20959 7837
rect 24946 7828 24952 7840
rect 25004 7828 25010 7880
rect 25041 7871 25099 7877
rect 25041 7837 25053 7871
rect 25087 7837 25099 7871
rect 25041 7831 25099 7837
rect 19352 7800 19380 7828
rect 18800 7772 19380 7800
rect 24854 7760 24860 7812
rect 24912 7800 24918 7812
rect 25056 7800 25084 7831
rect 24912 7772 25084 7800
rect 24912 7760 24918 7772
rect 14458 7732 14464 7744
rect 11940 7704 14311 7732
rect 14419 7704 14464 7732
rect 11940 7692 11946 7704
rect 14458 7692 14464 7704
rect 14516 7692 14522 7744
rect 18598 7732 18604 7744
rect 18559 7704 18604 7732
rect 18598 7692 18604 7704
rect 18656 7692 18662 7744
rect 20530 7732 20536 7744
rect 20491 7704 20536 7732
rect 20530 7692 20536 7704
rect 20588 7692 20594 7744
rect 22281 7735 22339 7741
rect 22281 7701 22293 7735
rect 22327 7732 22339 7735
rect 23290 7732 23296 7744
rect 22327 7704 23296 7732
rect 22327 7701 22339 7704
rect 22281 7695 22339 7701
rect 23290 7692 23296 7704
rect 23348 7692 23354 7744
rect 23569 7735 23627 7741
rect 23569 7701 23581 7735
rect 23615 7732 23627 7735
rect 25314 7732 25320 7744
rect 23615 7704 25320 7732
rect 23615 7701 23627 7704
rect 23569 7695 23627 7701
rect 25314 7692 25320 7704
rect 25372 7692 25378 7744
rect 25498 7732 25504 7744
rect 25459 7704 25504 7732
rect 25498 7692 25504 7704
rect 25556 7692 25562 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1489 7531 1547 7537
rect 1489 7497 1501 7531
rect 1535 7528 1547 7531
rect 1578 7528 1584 7540
rect 1535 7500 1584 7528
rect 1535 7497 1547 7500
rect 1489 7491 1547 7497
rect 1578 7488 1584 7500
rect 1636 7488 1642 7540
rect 2314 7488 2320 7540
rect 2372 7528 2378 7540
rect 2501 7531 2559 7537
rect 2501 7528 2513 7531
rect 2372 7500 2513 7528
rect 2372 7488 2378 7500
rect 2501 7497 2513 7500
rect 2547 7497 2559 7531
rect 2501 7491 2559 7497
rect 3142 7488 3148 7540
rect 3200 7528 3206 7540
rect 3973 7531 4031 7537
rect 3973 7528 3985 7531
rect 3200 7500 3985 7528
rect 3200 7488 3206 7500
rect 3973 7497 3985 7500
rect 4019 7497 4031 7531
rect 5442 7528 5448 7540
rect 5403 7500 5448 7528
rect 3973 7491 4031 7497
rect 5442 7488 5448 7500
rect 5500 7488 5506 7540
rect 8386 7488 8392 7540
rect 8444 7528 8450 7540
rect 8573 7531 8631 7537
rect 8573 7528 8585 7531
rect 8444 7500 8585 7528
rect 8444 7488 8450 7500
rect 8573 7497 8585 7500
rect 8619 7497 8631 7531
rect 9766 7528 9772 7540
rect 9727 7500 9772 7528
rect 8573 7491 8631 7497
rect 9766 7488 9772 7500
rect 9824 7488 9830 7540
rect 11241 7531 11299 7537
rect 11241 7497 11253 7531
rect 11287 7528 11299 7531
rect 11330 7528 11336 7540
rect 11287 7500 11336 7528
rect 11287 7497 11299 7500
rect 11241 7491 11299 7497
rect 11330 7488 11336 7500
rect 11388 7488 11394 7540
rect 11885 7531 11943 7537
rect 11885 7497 11897 7531
rect 11931 7528 11943 7531
rect 12342 7528 12348 7540
rect 11931 7500 12348 7528
rect 11931 7497 11943 7500
rect 11885 7491 11943 7497
rect 12342 7488 12348 7500
rect 12400 7488 12406 7540
rect 12618 7488 12624 7540
rect 12676 7528 12682 7540
rect 13541 7531 13599 7537
rect 13541 7528 13553 7531
rect 12676 7500 13553 7528
rect 12676 7488 12682 7500
rect 13541 7497 13553 7500
rect 13587 7528 13599 7531
rect 13630 7528 13636 7540
rect 13587 7500 13636 7528
rect 13587 7497 13599 7500
rect 13541 7491 13599 7497
rect 13630 7488 13636 7500
rect 13688 7488 13694 7540
rect 13906 7488 13912 7540
rect 13964 7528 13970 7540
rect 15013 7531 15071 7537
rect 15013 7528 15025 7531
rect 13964 7500 15025 7528
rect 13964 7488 13970 7500
rect 15013 7497 15025 7500
rect 15059 7497 15071 7531
rect 15562 7528 15568 7540
rect 15523 7500 15568 7528
rect 15013 7491 15071 7497
rect 15562 7488 15568 7500
rect 15620 7488 15626 7540
rect 15838 7528 15844 7540
rect 15799 7500 15844 7528
rect 15838 7488 15844 7500
rect 15896 7488 15902 7540
rect 17494 7528 17500 7540
rect 17455 7500 17500 7528
rect 17494 7488 17500 7500
rect 17552 7488 17558 7540
rect 17770 7488 17776 7540
rect 17828 7528 17834 7540
rect 18966 7528 18972 7540
rect 17828 7500 18972 7528
rect 17828 7488 17834 7500
rect 18966 7488 18972 7500
rect 19024 7488 19030 7540
rect 19334 7488 19340 7540
rect 19392 7528 19398 7540
rect 20070 7528 20076 7540
rect 19392 7500 19437 7528
rect 20031 7500 20076 7528
rect 19392 7488 19398 7500
rect 20070 7488 20076 7500
rect 20128 7488 20134 7540
rect 23382 7528 23388 7540
rect 23343 7500 23388 7528
rect 23382 7488 23388 7500
rect 23440 7488 23446 7540
rect 23934 7528 23940 7540
rect 23895 7500 23940 7528
rect 23934 7488 23940 7500
rect 23992 7488 23998 7540
rect 26418 7528 26424 7540
rect 26379 7500 26424 7528
rect 26418 7488 26424 7500
rect 26476 7488 26482 7540
rect 2133 7395 2191 7401
rect 2133 7361 2145 7395
rect 2179 7392 2191 7395
rect 2332 7392 2360 7488
rect 7006 7420 7012 7472
rect 7064 7460 7070 7472
rect 7561 7463 7619 7469
rect 7561 7460 7573 7463
rect 7064 7432 7573 7460
rect 7064 7420 7070 7432
rect 7561 7429 7573 7432
rect 7607 7429 7619 7463
rect 12158 7460 12164 7472
rect 12119 7432 12164 7460
rect 7561 7423 7619 7429
rect 12158 7420 12164 7432
rect 12216 7460 12222 7472
rect 12894 7460 12900 7472
rect 12216 7432 12900 7460
rect 12216 7420 12222 7432
rect 12894 7420 12900 7432
rect 12952 7420 12958 7472
rect 13814 7420 13820 7472
rect 13872 7460 13878 7472
rect 13872 7432 14596 7460
rect 13872 7420 13878 7432
rect 4430 7392 4436 7404
rect 2179 7364 2360 7392
rect 4391 7364 4436 7392
rect 2179 7361 2191 7364
rect 2133 7355 2191 7361
rect 4430 7352 4436 7364
rect 4488 7352 4494 7404
rect 4525 7395 4583 7401
rect 4525 7361 4537 7395
rect 4571 7361 4583 7395
rect 8018 7392 8024 7404
rect 7979 7364 8024 7392
rect 4525 7355 4583 7361
rect 3326 7324 3332 7336
rect 1872 7296 3332 7324
rect 1872 7200 1900 7296
rect 3326 7284 3332 7296
rect 3384 7284 3390 7336
rect 3513 7327 3571 7333
rect 3513 7293 3525 7327
rect 3559 7324 3571 7327
rect 3602 7324 3608 7336
rect 3559 7296 3608 7324
rect 3559 7293 3571 7296
rect 3513 7287 3571 7293
rect 3602 7284 3608 7296
rect 3660 7324 3666 7336
rect 4540 7324 4568 7355
rect 8018 7352 8024 7364
rect 8076 7352 8082 7404
rect 8110 7352 8116 7404
rect 8168 7392 8174 7404
rect 8168 7364 8213 7392
rect 8168 7352 8174 7364
rect 12710 7352 12716 7404
rect 12768 7392 12774 7404
rect 13081 7395 13139 7401
rect 13081 7392 13093 7395
rect 12768 7364 13093 7392
rect 12768 7352 12774 7364
rect 13081 7361 13093 7364
rect 13127 7392 13139 7395
rect 13170 7392 13176 7404
rect 13127 7364 13176 7392
rect 13127 7361 13139 7364
rect 13081 7355 13139 7361
rect 13170 7352 13176 7364
rect 13228 7352 13234 7404
rect 13906 7352 13912 7404
rect 13964 7392 13970 7404
rect 14274 7392 14280 7404
rect 13964 7364 14280 7392
rect 13964 7352 13970 7364
rect 14274 7352 14280 7364
rect 14332 7352 14338 7404
rect 14458 7392 14464 7404
rect 14419 7364 14464 7392
rect 14458 7352 14464 7364
rect 14516 7352 14522 7404
rect 14568 7401 14596 7432
rect 14553 7395 14611 7401
rect 14553 7361 14565 7395
rect 14599 7361 14611 7395
rect 14553 7355 14611 7361
rect 17037 7395 17095 7401
rect 17037 7361 17049 7395
rect 17083 7392 17095 7395
rect 17512 7392 17540 7488
rect 18233 7463 18291 7469
rect 18233 7429 18245 7463
rect 18279 7460 18291 7463
rect 19242 7460 19248 7472
rect 18279 7432 19248 7460
rect 18279 7429 18291 7432
rect 18233 7423 18291 7429
rect 19242 7420 19248 7432
rect 19300 7420 19306 7472
rect 21637 7463 21695 7469
rect 21637 7429 21649 7463
rect 21683 7460 21695 7463
rect 22922 7460 22928 7472
rect 21683 7432 22928 7460
rect 21683 7429 21695 7432
rect 21637 7423 21695 7429
rect 17083 7364 17540 7392
rect 17865 7395 17923 7401
rect 17083 7361 17095 7364
rect 17037 7355 17095 7361
rect 17865 7361 17877 7395
rect 17911 7392 17923 7395
rect 18877 7395 18935 7401
rect 18877 7392 18889 7395
rect 17911 7364 18889 7392
rect 17911 7361 17923 7364
rect 17865 7355 17923 7361
rect 18248 7336 18276 7364
rect 18800 7336 18828 7364
rect 18877 7361 18889 7364
rect 18923 7361 18935 7395
rect 18877 7355 18935 7361
rect 20254 7352 20260 7404
rect 20312 7392 20318 7404
rect 20717 7395 20775 7401
rect 20717 7392 20729 7395
rect 20312 7364 20729 7392
rect 20312 7352 20318 7364
rect 20717 7361 20729 7364
rect 20763 7361 20775 7395
rect 20717 7355 20775 7361
rect 21450 7352 21456 7404
rect 21508 7392 21514 7404
rect 21910 7392 21916 7404
rect 21508 7364 21916 7392
rect 21508 7352 21514 7364
rect 21910 7352 21916 7364
rect 21968 7392 21974 7404
rect 22204 7401 22232 7432
rect 22922 7420 22928 7432
rect 22980 7420 22986 7472
rect 24949 7463 25007 7469
rect 24949 7460 24961 7463
rect 24136 7432 24961 7460
rect 22189 7395 22247 7401
rect 21968 7364 22140 7392
rect 21968 7352 21974 7364
rect 3660 7296 4568 7324
rect 3660 7284 3666 7296
rect 5534 7284 5540 7336
rect 5592 7324 5598 7336
rect 5629 7327 5687 7333
rect 5629 7324 5641 7327
rect 5592 7296 5641 7324
rect 5592 7284 5598 7296
rect 5629 7293 5641 7296
rect 5675 7293 5687 7327
rect 7926 7324 7932 7336
rect 7887 7296 7932 7324
rect 5629 7287 5687 7293
rect 7926 7284 7932 7296
rect 7984 7284 7990 7336
rect 8662 7284 8668 7336
rect 8720 7324 8726 7336
rect 9309 7327 9367 7333
rect 9309 7324 9321 7327
rect 8720 7296 9321 7324
rect 8720 7284 8726 7296
rect 9309 7293 9321 7296
rect 9355 7293 9367 7327
rect 9309 7287 9367 7293
rect 9582 7284 9588 7336
rect 9640 7324 9646 7336
rect 9861 7327 9919 7333
rect 9861 7324 9873 7327
rect 9640 7296 9873 7324
rect 9640 7284 9646 7296
rect 9861 7293 9873 7296
rect 9907 7293 9919 7327
rect 9861 7287 9919 7293
rect 9950 7284 9956 7336
rect 10008 7324 10014 7336
rect 10117 7327 10175 7333
rect 10117 7324 10129 7327
rect 10008 7296 10129 7324
rect 10008 7284 10014 7296
rect 10117 7293 10129 7296
rect 10163 7293 10175 7327
rect 10117 7287 10175 7293
rect 12434 7284 12440 7336
rect 12492 7324 12498 7336
rect 12805 7327 12863 7333
rect 12805 7324 12817 7327
rect 12492 7296 12817 7324
rect 12492 7284 12498 7296
rect 12805 7293 12817 7296
rect 12851 7293 12863 7327
rect 12805 7287 12863 7293
rect 13832 7296 14504 7324
rect 1949 7259 2007 7265
rect 1949 7225 1961 7259
rect 1995 7256 2007 7259
rect 2682 7256 2688 7268
rect 1995 7228 2688 7256
rect 1995 7225 2007 7228
rect 1949 7219 2007 7225
rect 2682 7216 2688 7228
rect 2740 7216 2746 7268
rect 3881 7259 3939 7265
rect 3881 7225 3893 7259
rect 3927 7256 3939 7259
rect 5074 7256 5080 7268
rect 3927 7228 5080 7256
rect 3927 7225 3939 7228
rect 3881 7219 3939 7225
rect 5074 7216 5080 7228
rect 5132 7216 5138 7268
rect 7098 7256 7104 7268
rect 7011 7228 7104 7256
rect 7098 7216 7104 7228
rect 7156 7256 7162 7268
rect 8386 7256 8392 7268
rect 7156 7228 8392 7256
rect 7156 7216 7162 7228
rect 8386 7216 8392 7228
rect 8444 7216 8450 7268
rect 8846 7216 8852 7268
rect 8904 7256 8910 7268
rect 9033 7259 9091 7265
rect 9033 7256 9045 7259
rect 8904 7228 9045 7256
rect 8904 7216 8910 7228
rect 9033 7225 9045 7228
rect 9079 7256 9091 7259
rect 11054 7256 11060 7268
rect 9079 7228 11060 7256
rect 9079 7225 9091 7228
rect 9033 7219 9091 7225
rect 11054 7216 11060 7228
rect 11112 7216 11118 7268
rect 11146 7216 11152 7268
rect 11204 7256 11210 7268
rect 13832 7256 13860 7296
rect 11204 7228 13860 7256
rect 13909 7259 13967 7265
rect 11204 7216 11210 7228
rect 13909 7225 13921 7259
rect 13955 7256 13967 7259
rect 14476 7256 14504 7296
rect 15838 7284 15844 7336
rect 15896 7324 15902 7336
rect 16761 7327 16819 7333
rect 16761 7324 16773 7327
rect 15896 7296 16773 7324
rect 15896 7284 15902 7296
rect 16761 7293 16773 7296
rect 16807 7324 16819 7327
rect 17402 7324 17408 7336
rect 16807 7296 17408 7324
rect 16807 7293 16819 7296
rect 16761 7287 16819 7293
rect 17402 7284 17408 7296
rect 17460 7284 17466 7336
rect 18230 7284 18236 7336
rect 18288 7284 18294 7336
rect 18782 7284 18788 7336
rect 18840 7284 18846 7336
rect 19889 7327 19947 7333
rect 19889 7293 19901 7327
rect 19935 7324 19947 7327
rect 20625 7327 20683 7333
rect 20625 7324 20637 7327
rect 19935 7296 20637 7324
rect 19935 7293 19947 7296
rect 19889 7287 19947 7293
rect 20625 7293 20637 7296
rect 20671 7293 20683 7327
rect 20625 7287 20683 7293
rect 21269 7327 21327 7333
rect 21269 7293 21281 7327
rect 21315 7324 21327 7327
rect 22002 7324 22008 7336
rect 21315 7296 22008 7324
rect 21315 7293 21327 7296
rect 21269 7287 21327 7293
rect 22002 7284 22008 7296
rect 22060 7284 22066 7336
rect 22112 7324 22140 7364
rect 22189 7361 22201 7395
rect 22235 7361 22247 7395
rect 22189 7355 22247 7361
rect 22281 7395 22339 7401
rect 22281 7361 22293 7395
rect 22327 7361 22339 7395
rect 22281 7355 22339 7361
rect 22296 7324 22324 7355
rect 22112 7296 22324 7324
rect 23750 7284 23756 7336
rect 23808 7324 23814 7336
rect 23934 7324 23940 7336
rect 23808 7296 23940 7324
rect 23808 7284 23814 7296
rect 23934 7284 23940 7296
rect 23992 7324 23998 7336
rect 24136 7324 24164 7432
rect 24949 7429 24961 7432
rect 24995 7429 25007 7463
rect 24949 7423 25007 7429
rect 24581 7395 24639 7401
rect 24581 7361 24593 7395
rect 24627 7392 24639 7395
rect 24854 7392 24860 7404
rect 24627 7364 24860 7392
rect 24627 7361 24639 7364
rect 24581 7355 24639 7361
rect 24854 7352 24860 7364
rect 24912 7392 24918 7404
rect 26053 7395 26111 7401
rect 26053 7392 26065 7395
rect 24912 7364 26065 7392
rect 24912 7352 24918 7364
rect 26053 7361 26065 7364
rect 26099 7361 26111 7395
rect 26053 7355 26111 7361
rect 24305 7327 24363 7333
rect 24305 7324 24317 7327
rect 23992 7296 24317 7324
rect 23992 7284 23998 7296
rect 24305 7293 24317 7296
rect 24351 7293 24363 7327
rect 24305 7287 24363 7293
rect 24946 7284 24952 7336
rect 25004 7284 25010 7336
rect 25498 7324 25504 7336
rect 25459 7296 25504 7324
rect 25498 7284 25504 7296
rect 25556 7284 25562 7336
rect 16209 7259 16267 7265
rect 16209 7256 16221 7259
rect 13955 7228 14412 7256
rect 14476 7228 16221 7256
rect 13955 7225 13967 7228
rect 13909 7219 13967 7225
rect 1854 7188 1860 7200
rect 1815 7160 1860 7188
rect 1854 7148 1860 7160
rect 1912 7148 1918 7200
rect 2866 7148 2872 7200
rect 2924 7188 2930 7200
rect 2961 7191 3019 7197
rect 2961 7188 2973 7191
rect 2924 7160 2973 7188
rect 2924 7148 2930 7160
rect 2961 7157 2973 7160
rect 3007 7188 3019 7191
rect 3142 7188 3148 7200
rect 3007 7160 3148 7188
rect 3007 7157 3019 7160
rect 2961 7151 3019 7157
rect 3142 7148 3148 7160
rect 3200 7148 3206 7200
rect 4246 7148 4252 7200
rect 4304 7188 4310 7200
rect 4341 7191 4399 7197
rect 4341 7188 4353 7191
rect 4304 7160 4353 7188
rect 4304 7148 4310 7160
rect 4341 7157 4353 7160
rect 4387 7157 4399 7191
rect 4341 7151 4399 7157
rect 4985 7191 5043 7197
rect 4985 7157 4997 7191
rect 5031 7188 5043 7191
rect 5258 7188 5264 7200
rect 5031 7160 5264 7188
rect 5031 7157 5043 7160
rect 4985 7151 5043 7157
rect 5258 7148 5264 7160
rect 5316 7148 5322 7200
rect 5813 7191 5871 7197
rect 5813 7157 5825 7191
rect 5859 7188 5871 7191
rect 6270 7188 6276 7200
rect 5859 7160 6276 7188
rect 5859 7157 5871 7160
rect 5813 7151 5871 7157
rect 6270 7148 6276 7160
rect 6328 7148 6334 7200
rect 6454 7188 6460 7200
rect 6415 7160 6460 7188
rect 6454 7148 6460 7160
rect 6512 7148 6518 7200
rect 7282 7148 7288 7200
rect 7340 7188 7346 7200
rect 7377 7191 7435 7197
rect 7377 7188 7389 7191
rect 7340 7160 7389 7188
rect 7340 7148 7346 7160
rect 7377 7157 7389 7160
rect 7423 7157 7435 7191
rect 7377 7151 7435 7157
rect 9125 7191 9183 7197
rect 9125 7157 9137 7191
rect 9171 7188 9183 7191
rect 9214 7188 9220 7200
rect 9171 7160 9220 7188
rect 9171 7157 9183 7160
rect 9125 7151 9183 7157
rect 9214 7148 9220 7160
rect 9272 7188 9278 7200
rect 9582 7188 9588 7200
rect 9272 7160 9588 7188
rect 9272 7148 9278 7160
rect 9582 7148 9588 7160
rect 9640 7148 9646 7200
rect 12437 7191 12495 7197
rect 12437 7157 12449 7191
rect 12483 7188 12495 7191
rect 12526 7188 12532 7200
rect 12483 7160 12532 7188
rect 12483 7157 12495 7160
rect 12437 7151 12495 7157
rect 12526 7148 12532 7160
rect 12584 7148 12590 7200
rect 12894 7188 12900 7200
rect 12855 7160 12900 7188
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 14001 7191 14059 7197
rect 14001 7157 14013 7191
rect 14047 7188 14059 7191
rect 14274 7188 14280 7200
rect 14047 7160 14280 7188
rect 14047 7157 14059 7160
rect 14001 7151 14059 7157
rect 14274 7148 14280 7160
rect 14332 7148 14338 7200
rect 14384 7197 14412 7228
rect 16209 7225 16221 7228
rect 16255 7256 16267 7259
rect 16853 7259 16911 7265
rect 16853 7256 16865 7259
rect 16255 7228 16865 7256
rect 16255 7225 16267 7228
rect 16209 7219 16267 7225
rect 16853 7225 16865 7228
rect 16899 7256 16911 7259
rect 17586 7256 17592 7268
rect 16899 7228 17592 7256
rect 16899 7225 16911 7228
rect 16853 7219 16911 7225
rect 17586 7216 17592 7228
rect 17644 7216 17650 7268
rect 18598 7256 18604 7268
rect 18511 7228 18604 7256
rect 18598 7216 18604 7228
rect 18656 7256 18662 7268
rect 18656 7228 21312 7256
rect 18656 7216 18662 7228
rect 14369 7191 14427 7197
rect 14369 7157 14381 7191
rect 14415 7188 14427 7191
rect 14458 7188 14464 7200
rect 14415 7160 14464 7188
rect 14415 7157 14427 7160
rect 14369 7151 14427 7157
rect 14458 7148 14464 7160
rect 14516 7148 14522 7200
rect 16390 7188 16396 7200
rect 16351 7160 16396 7188
rect 16390 7148 16396 7160
rect 16448 7148 16454 7200
rect 18322 7148 18328 7200
rect 18380 7188 18386 7200
rect 18693 7191 18751 7197
rect 18693 7188 18705 7191
rect 18380 7160 18705 7188
rect 18380 7148 18386 7160
rect 18693 7157 18705 7160
rect 18739 7157 18751 7191
rect 18693 7151 18751 7157
rect 19334 7148 19340 7200
rect 19392 7188 19398 7200
rect 19613 7191 19671 7197
rect 19613 7188 19625 7191
rect 19392 7160 19625 7188
rect 19392 7148 19398 7160
rect 19613 7157 19625 7160
rect 19659 7188 19671 7191
rect 19889 7191 19947 7197
rect 19889 7188 19901 7191
rect 19659 7160 19901 7188
rect 19659 7157 19671 7160
rect 19613 7151 19671 7157
rect 19889 7157 19901 7160
rect 19935 7157 19947 7191
rect 19889 7151 19947 7157
rect 20165 7191 20223 7197
rect 20165 7157 20177 7191
rect 20211 7188 20223 7191
rect 20438 7188 20444 7200
rect 20211 7160 20444 7188
rect 20211 7157 20223 7160
rect 20165 7151 20223 7157
rect 20438 7148 20444 7160
rect 20496 7148 20502 7200
rect 20533 7191 20591 7197
rect 20533 7157 20545 7191
rect 20579 7188 20591 7191
rect 20622 7188 20628 7200
rect 20579 7160 20628 7188
rect 20579 7157 20591 7160
rect 20533 7151 20591 7157
rect 20622 7148 20628 7160
rect 20680 7148 20686 7200
rect 21284 7188 21312 7228
rect 24118 7216 24124 7268
rect 24176 7256 24182 7268
rect 24964 7256 24992 7284
rect 25317 7259 25375 7265
rect 25317 7256 25329 7259
rect 24176 7228 25329 7256
rect 24176 7216 24182 7228
rect 25317 7225 25329 7228
rect 25363 7225 25375 7259
rect 25317 7219 25375 7225
rect 21729 7191 21787 7197
rect 21729 7188 21741 7191
rect 21284 7160 21741 7188
rect 21729 7157 21741 7160
rect 21775 7157 21787 7191
rect 21729 7151 21787 7157
rect 22002 7148 22008 7200
rect 22060 7188 22066 7200
rect 22097 7191 22155 7197
rect 22097 7188 22109 7191
rect 22060 7160 22109 7188
rect 22060 7148 22066 7160
rect 22097 7157 22109 7160
rect 22143 7188 22155 7191
rect 22186 7188 22192 7200
rect 22143 7160 22192 7188
rect 22143 7157 22155 7160
rect 22097 7151 22155 7157
rect 22186 7148 22192 7160
rect 22244 7148 22250 7200
rect 22278 7148 22284 7200
rect 22336 7188 22342 7200
rect 23109 7191 23167 7197
rect 23109 7188 23121 7191
rect 22336 7160 23121 7188
rect 22336 7148 22342 7160
rect 23109 7157 23121 7160
rect 23155 7188 23167 7191
rect 23750 7188 23756 7200
rect 23155 7160 23756 7188
rect 23155 7157 23167 7160
rect 23109 7151 23167 7157
rect 23750 7148 23756 7160
rect 23808 7188 23814 7200
rect 24397 7191 24455 7197
rect 24397 7188 24409 7191
rect 23808 7160 24409 7188
rect 23808 7148 23814 7160
rect 24397 7157 24409 7160
rect 24443 7157 24455 7191
rect 24397 7151 24455 7157
rect 25685 7191 25743 7197
rect 25685 7157 25697 7191
rect 25731 7188 25743 7191
rect 25958 7188 25964 7200
rect 25731 7160 25964 7188
rect 25731 7157 25743 7160
rect 25685 7151 25743 7157
rect 25958 7148 25964 7160
rect 26016 7148 26022 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 4341 6987 4399 6993
rect 4341 6953 4353 6987
rect 4387 6984 4399 6987
rect 4430 6984 4436 6996
rect 4387 6956 4436 6984
rect 4387 6953 4399 6956
rect 4341 6947 4399 6953
rect 4430 6944 4436 6956
rect 4488 6944 4494 6996
rect 7193 6987 7251 6993
rect 7193 6953 7205 6987
rect 7239 6984 7251 6987
rect 7466 6984 7472 6996
rect 7239 6956 7472 6984
rect 7239 6953 7251 6956
rect 7193 6947 7251 6953
rect 7466 6944 7472 6956
rect 7524 6984 7530 6996
rect 7653 6987 7711 6993
rect 7653 6984 7665 6987
rect 7524 6956 7665 6984
rect 7524 6944 7530 6956
rect 7653 6953 7665 6956
rect 7699 6953 7711 6987
rect 7653 6947 7711 6953
rect 10045 6987 10103 6993
rect 10045 6953 10057 6987
rect 10091 6984 10103 6987
rect 10686 6984 10692 6996
rect 10091 6956 10692 6984
rect 10091 6953 10103 6956
rect 10045 6947 10103 6953
rect 10686 6944 10692 6956
rect 10744 6944 10750 6996
rect 12161 6987 12219 6993
rect 12161 6953 12173 6987
rect 12207 6984 12219 6987
rect 12250 6984 12256 6996
rect 12207 6956 12256 6984
rect 12207 6953 12219 6956
rect 12161 6947 12219 6953
rect 12250 6944 12256 6956
rect 12308 6944 12314 6996
rect 12434 6944 12440 6996
rect 12492 6984 12498 6996
rect 13078 6984 13084 6996
rect 12492 6956 12537 6984
rect 12991 6956 13084 6984
rect 12492 6944 12498 6956
rect 13078 6944 13084 6956
rect 13136 6984 13142 6996
rect 13262 6984 13268 6996
rect 13136 6956 13268 6984
rect 13136 6944 13142 6956
rect 13262 6944 13268 6956
rect 13320 6944 13326 6996
rect 13633 6987 13691 6993
rect 13633 6953 13645 6987
rect 13679 6984 13691 6987
rect 14090 6984 14096 6996
rect 13679 6956 14096 6984
rect 13679 6953 13691 6956
rect 13633 6947 13691 6953
rect 14090 6944 14096 6956
rect 14148 6944 14154 6996
rect 16577 6987 16635 6993
rect 16577 6953 16589 6987
rect 16623 6984 16635 6987
rect 17586 6984 17592 6996
rect 16623 6956 17592 6984
rect 16623 6953 16635 6956
rect 16577 6947 16635 6953
rect 17586 6944 17592 6956
rect 17644 6944 17650 6996
rect 17865 6987 17923 6993
rect 17865 6953 17877 6987
rect 17911 6984 17923 6987
rect 18874 6984 18880 6996
rect 17911 6956 18880 6984
rect 17911 6953 17923 6956
rect 17865 6947 17923 6953
rect 18874 6944 18880 6956
rect 18932 6944 18938 6996
rect 18969 6987 19027 6993
rect 18969 6953 18981 6987
rect 19015 6984 19027 6987
rect 19242 6984 19248 6996
rect 19015 6956 19248 6984
rect 19015 6953 19027 6956
rect 18969 6947 19027 6953
rect 19242 6944 19248 6956
rect 19300 6944 19306 6996
rect 20254 6984 20260 6996
rect 20215 6956 20260 6984
rect 20254 6944 20260 6956
rect 20312 6944 20318 6996
rect 21910 6984 21916 6996
rect 21871 6956 21916 6984
rect 21910 6944 21916 6956
rect 21968 6944 21974 6996
rect 25685 6987 25743 6993
rect 25685 6953 25697 6987
rect 25731 6984 25743 6987
rect 26142 6984 26148 6996
rect 25731 6956 26148 6984
rect 25731 6953 25743 6956
rect 25685 6947 25743 6953
rect 26142 6944 26148 6956
rect 26200 6944 26206 6996
rect 8018 6876 8024 6928
rect 8076 6916 8082 6928
rect 12989 6919 13047 6925
rect 8076 6888 8248 6916
rect 8076 6876 8082 6888
rect 1394 6808 1400 6860
rect 1452 6848 1458 6860
rect 1489 6851 1547 6857
rect 1489 6848 1501 6851
rect 1452 6820 1501 6848
rect 1452 6808 1458 6820
rect 1489 6817 1501 6820
rect 1535 6848 1547 6851
rect 1578 6848 1584 6860
rect 1535 6820 1584 6848
rect 1535 6817 1547 6820
rect 1489 6811 1547 6817
rect 1578 6808 1584 6820
rect 1636 6808 1642 6860
rect 1756 6851 1814 6857
rect 1756 6817 1768 6851
rect 1802 6848 1814 6851
rect 3602 6848 3608 6860
rect 1802 6820 3608 6848
rect 1802 6817 1814 6820
rect 1756 6811 1814 6817
rect 3602 6808 3608 6820
rect 3660 6808 3666 6860
rect 4890 6808 4896 6860
rect 4948 6848 4954 6860
rect 5057 6851 5115 6857
rect 5057 6848 5069 6851
rect 4948 6820 5069 6848
rect 4948 6808 4954 6820
rect 5057 6817 5069 6820
rect 5103 6817 5115 6851
rect 5057 6811 5115 6817
rect 5534 6808 5540 6860
rect 5592 6848 5598 6860
rect 6733 6851 6791 6857
rect 6733 6848 6745 6851
rect 5592 6820 6745 6848
rect 5592 6808 5598 6820
rect 6733 6817 6745 6820
rect 6779 6848 6791 6851
rect 6822 6848 6828 6860
rect 6779 6820 6828 6848
rect 6779 6817 6791 6820
rect 6733 6811 6791 6817
rect 6822 6808 6828 6820
rect 6880 6808 6886 6860
rect 6914 6808 6920 6860
rect 6972 6848 6978 6860
rect 7745 6851 7803 6857
rect 7745 6848 7757 6851
rect 6972 6820 7757 6848
rect 6972 6808 6978 6820
rect 7745 6817 7757 6820
rect 7791 6817 7803 6851
rect 8220 6848 8248 6888
rect 12989 6885 13001 6919
rect 13035 6916 13047 6919
rect 13722 6916 13728 6928
rect 13035 6888 13728 6916
rect 13035 6885 13047 6888
rect 12989 6879 13047 6885
rect 13722 6876 13728 6888
rect 13780 6876 13786 6928
rect 13814 6876 13820 6928
rect 13872 6916 13878 6928
rect 14001 6919 14059 6925
rect 14001 6916 14013 6919
rect 13872 6888 14013 6916
rect 13872 6876 13878 6888
rect 14001 6885 14013 6888
rect 14047 6885 14059 6919
rect 14001 6879 14059 6885
rect 8665 6851 8723 6857
rect 8665 6848 8677 6851
rect 8220 6820 8677 6848
rect 7745 6811 7803 6817
rect 8665 6817 8677 6820
rect 8711 6817 8723 6851
rect 8665 6811 8723 6817
rect 9766 6808 9772 6860
rect 9824 6848 9830 6860
rect 10393 6851 10451 6857
rect 10393 6848 10405 6851
rect 9824 6820 10405 6848
rect 9824 6808 9830 6820
rect 10393 6817 10405 6820
rect 10439 6848 10451 6851
rect 11330 6848 11336 6860
rect 10439 6820 11336 6848
rect 10439 6817 10451 6820
rect 10393 6811 10451 6817
rect 11330 6808 11336 6820
rect 11388 6808 11394 6860
rect 14016 6848 14044 6879
rect 14642 6876 14648 6928
rect 14700 6916 14706 6928
rect 14826 6916 14832 6928
rect 14700 6888 14832 6916
rect 14700 6876 14706 6888
rect 14826 6876 14832 6888
rect 14884 6876 14890 6928
rect 16390 6876 16396 6928
rect 16448 6916 16454 6928
rect 17405 6919 17463 6925
rect 16448 6888 16712 6916
rect 16448 6876 16454 6888
rect 15838 6848 15844 6860
rect 14016 6820 15844 6848
rect 15838 6808 15844 6820
rect 15896 6808 15902 6860
rect 16117 6851 16175 6857
rect 16117 6817 16129 6851
rect 16163 6848 16175 6851
rect 16206 6848 16212 6860
rect 16163 6820 16212 6848
rect 16163 6817 16175 6820
rect 16117 6811 16175 6817
rect 16206 6808 16212 6820
rect 16264 6808 16270 6860
rect 16684 6848 16712 6888
rect 17405 6885 17417 6919
rect 17451 6916 17463 6919
rect 18233 6919 18291 6925
rect 18233 6916 18245 6919
rect 17451 6888 18245 6916
rect 17451 6885 17463 6888
rect 17405 6879 17463 6885
rect 18233 6885 18245 6888
rect 18279 6916 18291 6919
rect 19150 6916 19156 6928
rect 18279 6888 19156 6916
rect 18279 6885 18291 6888
rect 18233 6879 18291 6885
rect 19150 6876 19156 6888
rect 19208 6876 19214 6928
rect 23106 6876 23112 6928
rect 23164 6916 23170 6928
rect 23560 6919 23618 6925
rect 23560 6916 23572 6919
rect 23164 6888 23572 6916
rect 23164 6876 23170 6888
rect 23560 6885 23572 6888
rect 23606 6916 23618 6919
rect 24854 6916 24860 6928
rect 23606 6888 24860 6916
rect 23606 6885 23618 6888
rect 23560 6879 23618 6885
rect 24854 6876 24860 6888
rect 24912 6916 24918 6928
rect 25038 6916 25044 6928
rect 24912 6888 25044 6916
rect 24912 6876 24918 6888
rect 25038 6876 25044 6888
rect 25096 6876 25102 6928
rect 17681 6851 17739 6857
rect 17681 6848 17693 6851
rect 16684 6820 17693 6848
rect 17681 6817 17693 6820
rect 17727 6817 17739 6851
rect 19426 6848 19432 6860
rect 19387 6820 19432 6848
rect 17681 6811 17739 6817
rect 4614 6740 4620 6792
rect 4672 6780 4678 6792
rect 4801 6783 4859 6789
rect 4801 6780 4813 6783
rect 4672 6752 4813 6780
rect 4672 6740 4678 6752
rect 4801 6749 4813 6752
rect 4847 6749 4859 6783
rect 4801 6743 4859 6749
rect 2869 6647 2927 6653
rect 2869 6613 2881 6647
rect 2915 6644 2927 6647
rect 3142 6644 3148 6656
rect 2915 6616 3148 6644
rect 2915 6613 2927 6616
rect 2869 6607 2927 6613
rect 3142 6604 3148 6616
rect 3200 6604 3206 6656
rect 3418 6644 3424 6656
rect 3379 6616 3424 6644
rect 3418 6604 3424 6616
rect 3476 6604 3482 6656
rect 3878 6644 3884 6656
rect 3839 6616 3884 6644
rect 3878 6604 3884 6616
rect 3936 6604 3942 6656
rect 4246 6604 4252 6656
rect 4304 6644 4310 6656
rect 4617 6647 4675 6653
rect 4617 6644 4629 6647
rect 4304 6616 4629 6644
rect 4304 6604 4310 6616
rect 4617 6613 4629 6616
rect 4663 6613 4675 6647
rect 4816 6644 4844 6743
rect 7466 6740 7472 6792
rect 7524 6780 7530 6792
rect 7837 6783 7895 6789
rect 7837 6780 7849 6783
rect 7524 6752 7849 6780
rect 7524 6740 7530 6752
rect 7837 6749 7849 6752
rect 7883 6780 7895 6783
rect 8110 6780 8116 6792
rect 7883 6752 8116 6780
rect 7883 6749 7895 6752
rect 7837 6743 7895 6749
rect 8110 6740 8116 6752
rect 8168 6740 8174 6792
rect 9582 6740 9588 6792
rect 9640 6780 9646 6792
rect 10137 6783 10195 6789
rect 10137 6780 10149 6783
rect 9640 6752 10149 6780
rect 9640 6740 9646 6752
rect 10137 6749 10149 6752
rect 10183 6749 10195 6783
rect 10137 6743 10195 6749
rect 7285 6715 7343 6721
rect 7285 6681 7297 6715
rect 7331 6712 7343 6715
rect 7926 6712 7932 6724
rect 7331 6684 7932 6712
rect 7331 6681 7343 6684
rect 7285 6675 7343 6681
rect 7926 6672 7932 6684
rect 7984 6712 7990 6724
rect 9033 6715 9091 6721
rect 9033 6712 9045 6715
rect 7984 6684 9045 6712
rect 7984 6672 7990 6684
rect 9033 6681 9045 6684
rect 9079 6681 9091 6715
rect 9033 6675 9091 6681
rect 5534 6644 5540 6656
rect 4816 6616 5540 6644
rect 4617 6607 4675 6613
rect 5534 6604 5540 6616
rect 5592 6604 5598 6656
rect 6086 6604 6092 6656
rect 6144 6644 6150 6656
rect 6181 6647 6239 6653
rect 6181 6644 6193 6647
rect 6144 6616 6193 6644
rect 6144 6604 6150 6616
rect 6181 6613 6193 6616
rect 6227 6613 6239 6647
rect 8386 6644 8392 6656
rect 8299 6616 8392 6644
rect 6181 6607 6239 6613
rect 8386 6604 8392 6616
rect 8444 6644 8450 6656
rect 9214 6644 9220 6656
rect 8444 6616 9220 6644
rect 8444 6604 8450 6616
rect 9214 6604 9220 6616
rect 9272 6604 9278 6656
rect 9306 6604 9312 6656
rect 9364 6644 9370 6656
rect 9401 6647 9459 6653
rect 9401 6644 9413 6647
rect 9364 6616 9413 6644
rect 9364 6604 9370 6616
rect 9401 6613 9413 6616
rect 9447 6613 9459 6647
rect 10152 6644 10180 6743
rect 13170 6740 13176 6792
rect 13228 6780 13234 6792
rect 13228 6752 13273 6780
rect 13228 6740 13234 6752
rect 14090 6740 14096 6792
rect 14148 6780 14154 6792
rect 14185 6783 14243 6789
rect 14185 6780 14197 6783
rect 14148 6752 14197 6780
rect 14148 6740 14154 6752
rect 14185 6749 14197 6752
rect 14231 6749 14243 6783
rect 15470 6780 15476 6792
rect 15431 6752 15476 6780
rect 14185 6743 14243 6749
rect 15470 6740 15476 6752
rect 15528 6740 15534 6792
rect 16224 6780 16252 6808
rect 16666 6780 16672 6792
rect 16224 6752 16528 6780
rect 16627 6752 16672 6780
rect 16114 6672 16120 6724
rect 16172 6712 16178 6724
rect 16209 6715 16267 6721
rect 16209 6712 16221 6715
rect 16172 6684 16221 6712
rect 16172 6672 16178 6684
rect 16209 6681 16221 6684
rect 16255 6681 16267 6715
rect 16500 6712 16528 6752
rect 16666 6740 16672 6752
rect 16724 6740 16730 6792
rect 16761 6783 16819 6789
rect 16761 6749 16773 6783
rect 16807 6749 16819 6783
rect 17696 6780 17724 6811
rect 19426 6808 19432 6820
rect 19484 6808 19490 6860
rect 21266 6848 21272 6860
rect 21227 6820 21272 6848
rect 21266 6808 21272 6820
rect 21324 6808 21330 6860
rect 23017 6851 23075 6857
rect 23017 6848 23029 6851
rect 21376 6820 23029 6848
rect 18325 6783 18383 6789
rect 18325 6780 18337 6783
rect 17696 6752 18337 6780
rect 16761 6743 16819 6749
rect 18325 6749 18337 6752
rect 18371 6749 18383 6783
rect 18325 6743 18383 6749
rect 18509 6783 18567 6789
rect 18509 6749 18521 6783
rect 18555 6780 18567 6783
rect 18598 6780 18604 6792
rect 18555 6752 18604 6780
rect 18555 6749 18567 6752
rect 18509 6743 18567 6749
rect 16776 6712 16804 6743
rect 18598 6740 18604 6752
rect 18656 6780 18662 6792
rect 18782 6780 18788 6792
rect 18656 6752 18788 6780
rect 18656 6740 18662 6752
rect 18782 6740 18788 6752
rect 18840 6740 18846 6792
rect 19610 6780 19616 6792
rect 19571 6752 19616 6780
rect 19610 6740 19616 6752
rect 19668 6740 19674 6792
rect 20714 6740 20720 6792
rect 20772 6780 20778 6792
rect 21376 6789 21404 6820
rect 23017 6817 23029 6820
rect 23063 6817 23075 6851
rect 23017 6811 23075 6817
rect 21361 6783 21419 6789
rect 21361 6780 21373 6783
rect 20772 6752 21373 6780
rect 20772 6740 20778 6752
rect 21361 6749 21373 6752
rect 21407 6749 21419 6783
rect 21361 6743 21419 6749
rect 21545 6783 21603 6789
rect 21545 6749 21557 6783
rect 21591 6780 21603 6783
rect 21818 6780 21824 6792
rect 21591 6752 21824 6780
rect 21591 6749 21603 6752
rect 21545 6743 21603 6749
rect 21818 6740 21824 6752
rect 21876 6740 21882 6792
rect 23290 6780 23296 6792
rect 23251 6752 23296 6780
rect 23290 6740 23296 6752
rect 23348 6740 23354 6792
rect 16500 6684 16804 6712
rect 16209 6675 16267 6681
rect 16850 6672 16856 6724
rect 16908 6672 16914 6724
rect 19337 6715 19395 6721
rect 19337 6681 19349 6715
rect 19383 6712 19395 6715
rect 20438 6712 20444 6724
rect 19383 6684 20444 6712
rect 19383 6681 19395 6684
rect 19337 6675 19395 6681
rect 20438 6672 20444 6684
rect 20496 6672 20502 6724
rect 20901 6715 20959 6721
rect 20901 6681 20913 6715
rect 20947 6712 20959 6715
rect 20990 6712 20996 6724
rect 20947 6684 20996 6712
rect 20947 6681 20959 6684
rect 20901 6675 20959 6681
rect 20990 6672 20996 6684
rect 21048 6672 21054 6724
rect 21726 6672 21732 6724
rect 21784 6712 21790 6724
rect 22649 6715 22707 6721
rect 22649 6712 22661 6715
rect 21784 6684 22661 6712
rect 21784 6672 21790 6684
rect 22649 6681 22661 6684
rect 22695 6681 22707 6715
rect 22649 6675 22707 6681
rect 24673 6715 24731 6721
rect 24673 6681 24685 6715
rect 24719 6712 24731 6715
rect 24762 6712 24768 6724
rect 24719 6684 24768 6712
rect 24719 6681 24731 6684
rect 24673 6675 24731 6681
rect 24762 6672 24768 6684
rect 24820 6672 24826 6724
rect 25222 6672 25228 6724
rect 25280 6712 25286 6724
rect 25317 6715 25375 6721
rect 25317 6712 25329 6715
rect 25280 6684 25329 6712
rect 25280 6672 25286 6684
rect 25317 6681 25329 6684
rect 25363 6712 25375 6715
rect 25866 6712 25872 6724
rect 25363 6684 25872 6712
rect 25363 6681 25375 6684
rect 25317 6675 25375 6681
rect 25866 6672 25872 6684
rect 25924 6672 25930 6724
rect 10410 6644 10416 6656
rect 10152 6616 10416 6644
rect 9401 6607 9459 6613
rect 10410 6604 10416 6616
rect 10468 6604 10474 6656
rect 11054 6604 11060 6656
rect 11112 6644 11118 6656
rect 11517 6647 11575 6653
rect 11517 6644 11529 6647
rect 11112 6616 11529 6644
rect 11112 6604 11118 6616
rect 11517 6613 11529 6616
rect 11563 6613 11575 6647
rect 11517 6607 11575 6613
rect 12621 6647 12679 6653
rect 12621 6613 12633 6647
rect 12667 6644 12679 6647
rect 12894 6644 12900 6656
rect 12667 6616 12900 6644
rect 12667 6613 12679 6616
rect 12621 6607 12679 6613
rect 12894 6604 12900 6616
rect 12952 6644 12958 6656
rect 14645 6647 14703 6653
rect 14645 6644 14657 6647
rect 12952 6616 14657 6644
rect 12952 6604 12958 6616
rect 14645 6613 14657 6616
rect 14691 6613 14703 6647
rect 14645 6607 14703 6613
rect 14826 6604 14832 6656
rect 14884 6644 14890 6656
rect 15013 6647 15071 6653
rect 15013 6644 15025 6647
rect 14884 6616 15025 6644
rect 14884 6604 14890 6616
rect 15013 6613 15025 6616
rect 15059 6613 15071 6647
rect 15013 6607 15071 6613
rect 16390 6604 16396 6656
rect 16448 6644 16454 6656
rect 16868 6644 16896 6672
rect 20622 6644 20628 6656
rect 16448 6616 16896 6644
rect 20583 6616 20628 6644
rect 16448 6604 16454 6616
rect 20622 6604 20628 6616
rect 20680 6604 20686 6656
rect 21358 6604 21364 6656
rect 21416 6644 21422 6656
rect 22281 6647 22339 6653
rect 22281 6644 22293 6647
rect 21416 6616 22293 6644
rect 21416 6604 21422 6616
rect 22281 6613 22293 6616
rect 22327 6613 22339 6647
rect 22281 6607 22339 6613
rect 24854 6604 24860 6656
rect 24912 6644 24918 6656
rect 25961 6647 26019 6653
rect 25961 6644 25973 6647
rect 24912 6616 25973 6644
rect 24912 6604 24918 6616
rect 25961 6613 25973 6616
rect 26007 6613 26019 6647
rect 25961 6607 26019 6613
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 3602 6400 3608 6452
rect 3660 6440 3666 6452
rect 3789 6443 3847 6449
rect 3789 6440 3801 6443
rect 3660 6412 3801 6440
rect 3660 6400 3666 6412
rect 3789 6409 3801 6412
rect 3835 6409 3847 6443
rect 3789 6403 3847 6409
rect 1578 6264 1584 6316
rect 1636 6304 1642 6316
rect 3804 6304 3832 6403
rect 4062 6400 4068 6452
rect 4120 6440 4126 6452
rect 4893 6443 4951 6449
rect 4893 6440 4905 6443
rect 4120 6412 4905 6440
rect 4120 6400 4126 6412
rect 4893 6409 4905 6412
rect 4939 6409 4951 6443
rect 9766 6440 9772 6452
rect 9727 6412 9772 6440
rect 4893 6403 4951 6409
rect 9766 6400 9772 6412
rect 9824 6400 9830 6452
rect 13814 6400 13820 6452
rect 13872 6440 13878 6452
rect 14737 6443 14795 6449
rect 14737 6440 14749 6443
rect 13872 6412 14749 6440
rect 13872 6400 13878 6412
rect 14737 6409 14749 6412
rect 14783 6409 14795 6443
rect 14737 6403 14795 6409
rect 16942 6400 16948 6452
rect 17000 6440 17006 6452
rect 17405 6443 17463 6449
rect 17405 6440 17417 6443
rect 17000 6412 17417 6440
rect 17000 6400 17006 6412
rect 17405 6409 17417 6412
rect 17451 6409 17463 6443
rect 17770 6440 17776 6452
rect 17731 6412 17776 6440
rect 17405 6403 17463 6409
rect 4430 6332 4436 6384
rect 4488 6372 4494 6384
rect 6454 6372 6460 6384
rect 4488 6344 6460 6372
rect 4488 6332 4494 6344
rect 6454 6332 6460 6344
rect 6512 6332 6518 6384
rect 17420 6372 17448 6403
rect 17770 6400 17776 6412
rect 17828 6440 17834 6452
rect 17828 6412 18552 6440
rect 17828 6400 17834 6412
rect 18322 6372 18328 6384
rect 17420 6344 18328 6372
rect 18322 6332 18328 6344
rect 18380 6332 18386 6384
rect 4801 6307 4859 6313
rect 4801 6304 4813 6307
rect 1636 6276 2452 6304
rect 3804 6276 4813 6304
rect 1636 6264 1642 6276
rect 1762 6196 1768 6248
rect 1820 6236 1826 6248
rect 2130 6236 2136 6248
rect 1820 6208 2136 6236
rect 1820 6196 1826 6208
rect 2130 6196 2136 6208
rect 2188 6196 2194 6248
rect 2424 6245 2452 6276
rect 4801 6273 4813 6276
rect 4847 6304 4859 6307
rect 5445 6307 5503 6313
rect 5445 6304 5457 6307
rect 4847 6276 5457 6304
rect 4847 6273 4859 6276
rect 4801 6267 4859 6273
rect 5445 6273 5457 6276
rect 5491 6273 5503 6307
rect 5445 6267 5503 6273
rect 15197 6307 15255 6313
rect 15197 6273 15209 6307
rect 15243 6304 15255 6307
rect 15243 6276 15424 6304
rect 15243 6273 15255 6276
rect 15197 6267 15255 6273
rect 2409 6239 2467 6245
rect 2409 6205 2421 6239
rect 2455 6236 2467 6239
rect 4433 6239 4491 6245
rect 2455 6208 4384 6236
rect 2455 6205 2467 6208
rect 2409 6199 2467 6205
rect 2682 6177 2688 6180
rect 2317 6171 2375 6177
rect 2317 6137 2329 6171
rect 2363 6168 2375 6171
rect 2654 6171 2688 6177
rect 2654 6168 2666 6171
rect 2363 6140 2666 6168
rect 2363 6137 2375 6140
rect 2317 6131 2375 6137
rect 2654 6137 2666 6140
rect 2654 6131 2688 6137
rect 2682 6128 2688 6131
rect 2740 6128 2746 6180
rect 4356 6168 4384 6208
rect 4433 6205 4445 6239
rect 4479 6236 4491 6239
rect 4890 6236 4896 6248
rect 4479 6208 4896 6236
rect 4479 6205 4491 6208
rect 4433 6199 4491 6205
rect 4890 6196 4896 6208
rect 4948 6196 4954 6248
rect 5258 6236 5264 6248
rect 5219 6208 5264 6236
rect 5258 6196 5264 6208
rect 5316 6196 5322 6248
rect 5534 6196 5540 6248
rect 5592 6236 5598 6248
rect 7377 6239 7435 6245
rect 7377 6236 7389 6239
rect 5592 6208 7389 6236
rect 5592 6196 5598 6208
rect 7377 6205 7389 6208
rect 7423 6236 7435 6239
rect 8110 6236 8116 6248
rect 7423 6208 8116 6236
rect 7423 6205 7435 6208
rect 7377 6199 7435 6205
rect 8110 6196 8116 6208
rect 8168 6196 8174 6248
rect 9861 6239 9919 6245
rect 9861 6205 9873 6239
rect 9907 6236 9919 6239
rect 10410 6236 10416 6248
rect 9907 6208 10416 6236
rect 9907 6205 9919 6208
rect 9861 6199 9919 6205
rect 10410 6196 10416 6208
rect 10468 6236 10474 6248
rect 11514 6236 11520 6248
rect 10468 6208 11520 6236
rect 10468 6196 10474 6208
rect 11514 6196 11520 6208
rect 11572 6236 11578 6248
rect 11974 6236 11980 6248
rect 11572 6208 11980 6236
rect 11572 6196 11578 6208
rect 11974 6196 11980 6208
rect 12032 6236 12038 6248
rect 12437 6239 12495 6245
rect 12437 6236 12449 6239
rect 12032 6208 12449 6236
rect 12032 6196 12038 6208
rect 12437 6205 12449 6208
rect 12483 6205 12495 6239
rect 12704 6239 12762 6245
rect 12704 6236 12716 6239
rect 12437 6199 12495 6205
rect 12636 6208 12716 6236
rect 5552 6168 5580 6196
rect 4356 6140 5580 6168
rect 6273 6171 6331 6177
rect 6273 6137 6285 6171
rect 6319 6168 6331 6171
rect 7098 6168 7104 6180
rect 6319 6140 7104 6168
rect 6319 6137 6331 6140
rect 6273 6131 6331 6137
rect 7098 6128 7104 6140
rect 7156 6128 7162 6180
rect 7622 6171 7680 6177
rect 7622 6168 7634 6171
rect 7484 6140 7634 6168
rect 7484 6112 7512 6140
rect 7622 6137 7634 6140
rect 7668 6137 7680 6171
rect 9401 6171 9459 6177
rect 9401 6168 9413 6171
rect 7622 6131 7680 6137
rect 8772 6140 9413 6168
rect 1397 6103 1455 6109
rect 1397 6069 1409 6103
rect 1443 6100 1455 6103
rect 1762 6100 1768 6112
rect 1443 6072 1768 6100
rect 1443 6069 1455 6072
rect 1397 6063 1455 6069
rect 1762 6060 1768 6072
rect 1820 6100 1826 6112
rect 1857 6103 1915 6109
rect 1857 6100 1869 6103
rect 1820 6072 1869 6100
rect 1820 6060 1826 6072
rect 1857 6069 1869 6072
rect 1903 6069 1915 6103
rect 1857 6063 1915 6069
rect 5350 6060 5356 6112
rect 5408 6100 5414 6112
rect 6641 6103 6699 6109
rect 5408 6072 5453 6100
rect 5408 6060 5414 6072
rect 6641 6069 6653 6103
rect 6687 6100 6699 6103
rect 7285 6103 7343 6109
rect 7285 6100 7297 6103
rect 6687 6072 7297 6100
rect 6687 6069 6699 6072
rect 6641 6063 6699 6069
rect 7285 6069 7297 6072
rect 7331 6100 7343 6103
rect 7466 6100 7472 6112
rect 7331 6072 7472 6100
rect 7331 6069 7343 6072
rect 7285 6063 7343 6069
rect 7466 6060 7472 6072
rect 7524 6060 7530 6112
rect 8018 6060 8024 6112
rect 8076 6100 8082 6112
rect 8772 6109 8800 6140
rect 9401 6137 9413 6140
rect 9447 6168 9459 6171
rect 10106 6171 10164 6177
rect 10106 6168 10118 6171
rect 9447 6140 10118 6168
rect 9447 6137 9459 6140
rect 9401 6131 9459 6137
rect 10106 6137 10118 6140
rect 10152 6137 10164 6171
rect 12636 6168 12664 6208
rect 12704 6205 12716 6208
rect 12750 6236 12762 6239
rect 13170 6236 13176 6248
rect 12750 6208 13176 6236
rect 12750 6205 12762 6208
rect 12704 6199 12762 6205
rect 13170 6196 13176 6208
rect 13228 6196 13234 6248
rect 15289 6239 15347 6245
rect 15289 6205 15301 6239
rect 15335 6205 15347 6239
rect 15396 6236 15424 6276
rect 16298 6264 16304 6316
rect 16356 6264 16362 6316
rect 18524 6313 18552 6412
rect 18598 6400 18604 6452
rect 18656 6440 18662 6452
rect 19429 6443 19487 6449
rect 19429 6440 19441 6443
rect 18656 6412 19441 6440
rect 18656 6400 18662 6412
rect 19429 6409 19441 6412
rect 19475 6409 19487 6443
rect 19429 6403 19487 6409
rect 20349 6443 20407 6449
rect 20349 6409 20361 6443
rect 20395 6440 20407 6443
rect 21818 6440 21824 6452
rect 20395 6412 21824 6440
rect 20395 6409 20407 6412
rect 20349 6403 20407 6409
rect 21818 6400 21824 6412
rect 21876 6400 21882 6452
rect 23106 6440 23112 6452
rect 23067 6412 23112 6440
rect 23106 6400 23112 6412
rect 23164 6400 23170 6452
rect 23382 6440 23388 6452
rect 23343 6412 23388 6440
rect 23382 6400 23388 6412
rect 23440 6400 23446 6452
rect 25038 6440 25044 6452
rect 24999 6412 25044 6440
rect 25038 6400 25044 6412
rect 25096 6400 25102 6452
rect 26053 6443 26111 6449
rect 26053 6409 26065 6443
rect 26099 6440 26111 6443
rect 26142 6440 26148 6452
rect 26099 6412 26148 6440
rect 26099 6409 26111 6412
rect 26053 6403 26111 6409
rect 26142 6400 26148 6412
rect 26200 6440 26206 6452
rect 26329 6443 26387 6449
rect 26329 6440 26341 6443
rect 26200 6412 26341 6440
rect 26200 6400 26206 6412
rect 26329 6409 26341 6412
rect 26375 6409 26387 6443
rect 26329 6403 26387 6409
rect 18509 6307 18567 6313
rect 18509 6273 18521 6307
rect 18555 6273 18567 6307
rect 18509 6267 18567 6273
rect 18693 6307 18751 6313
rect 18693 6273 18705 6307
rect 18739 6304 18751 6307
rect 18739 6276 18773 6304
rect 18739 6273 18751 6276
rect 18693 6267 18751 6273
rect 15556 6239 15614 6245
rect 15556 6236 15568 6239
rect 15396 6208 15568 6236
rect 15289 6199 15347 6205
rect 15556 6205 15568 6208
rect 15602 6236 15614 6239
rect 16316 6236 16344 6264
rect 15602 6208 16344 6236
rect 15602 6205 15614 6208
rect 15556 6199 15614 6205
rect 10106 6131 10164 6137
rect 12176 6140 12664 6168
rect 12176 6112 12204 6140
rect 15194 6128 15200 6180
rect 15252 6168 15258 6180
rect 15304 6168 15332 6199
rect 18414 6196 18420 6248
rect 18472 6236 18478 6248
rect 18708 6236 18736 6267
rect 19426 6264 19432 6316
rect 19484 6304 19490 6316
rect 19797 6307 19855 6313
rect 19797 6304 19809 6307
rect 19484 6276 19809 6304
rect 19484 6264 19490 6276
rect 19797 6273 19809 6276
rect 19843 6273 19855 6307
rect 19797 6267 19855 6273
rect 19061 6239 19119 6245
rect 19061 6236 19073 6239
rect 18472 6208 19073 6236
rect 18472 6196 18478 6208
rect 19061 6205 19073 6208
rect 19107 6205 19119 6239
rect 19061 6199 19119 6205
rect 20441 6239 20499 6245
rect 20441 6205 20453 6239
rect 20487 6236 20499 6239
rect 20530 6236 20536 6248
rect 20487 6208 20536 6236
rect 20487 6205 20499 6208
rect 20441 6199 20499 6205
rect 20530 6196 20536 6208
rect 20588 6196 20594 6248
rect 23290 6196 23296 6248
rect 23348 6236 23354 6248
rect 23661 6239 23719 6245
rect 23661 6236 23673 6239
rect 23348 6208 23673 6236
rect 23348 6196 23354 6208
rect 23661 6205 23673 6208
rect 23707 6236 23719 6239
rect 24854 6236 24860 6248
rect 23707 6208 24860 6236
rect 23707 6205 23719 6208
rect 23661 6199 23719 6205
rect 24854 6196 24860 6208
rect 24912 6196 24918 6248
rect 19334 6168 19340 6180
rect 15252 6140 15332 6168
rect 18064 6140 19340 6168
rect 15252 6128 15258 6140
rect 8757 6103 8815 6109
rect 8757 6100 8769 6103
rect 8076 6072 8769 6100
rect 8076 6060 8082 6072
rect 8757 6069 8769 6072
rect 8803 6069 8815 6103
rect 8757 6063 8815 6069
rect 9950 6060 9956 6112
rect 10008 6100 10014 6112
rect 11241 6103 11299 6109
rect 11241 6100 11253 6103
rect 10008 6072 11253 6100
rect 10008 6060 10014 6072
rect 11241 6069 11253 6072
rect 11287 6069 11299 6103
rect 11241 6063 11299 6069
rect 11885 6103 11943 6109
rect 11885 6069 11897 6103
rect 11931 6100 11943 6103
rect 12158 6100 12164 6112
rect 11931 6072 12164 6100
rect 11931 6069 11943 6072
rect 11885 6063 11943 6069
rect 12158 6060 12164 6072
rect 12216 6060 12222 6112
rect 13446 6060 13452 6112
rect 13504 6100 13510 6112
rect 13817 6103 13875 6109
rect 13817 6100 13829 6103
rect 13504 6072 13829 6100
rect 13504 6060 13510 6072
rect 13817 6069 13829 6072
rect 13863 6069 13875 6103
rect 14366 6100 14372 6112
rect 14327 6072 14372 6100
rect 13817 6063 13875 6069
rect 14366 6060 14372 6072
rect 14424 6060 14430 6112
rect 15654 6060 15660 6112
rect 15712 6100 15718 6112
rect 16206 6100 16212 6112
rect 15712 6072 16212 6100
rect 15712 6060 15718 6072
rect 16206 6060 16212 6072
rect 16264 6060 16270 6112
rect 16669 6103 16727 6109
rect 16669 6069 16681 6103
rect 16715 6100 16727 6103
rect 16942 6100 16948 6112
rect 16715 6072 16948 6100
rect 16715 6069 16727 6072
rect 16669 6063 16727 6069
rect 16942 6060 16948 6072
rect 17000 6100 17006 6112
rect 17494 6100 17500 6112
rect 17000 6072 17500 6100
rect 17000 6060 17006 6072
rect 17494 6060 17500 6072
rect 17552 6060 17558 6112
rect 18064 6109 18092 6140
rect 19334 6128 19340 6140
rect 19392 6128 19398 6180
rect 20162 6128 20168 6180
rect 20220 6168 20226 6180
rect 20686 6171 20744 6177
rect 20686 6168 20698 6171
rect 20220 6140 20698 6168
rect 20220 6128 20226 6140
rect 20686 6137 20698 6140
rect 20732 6137 20744 6171
rect 20686 6131 20744 6137
rect 23382 6128 23388 6180
rect 23440 6168 23446 6180
rect 23906 6171 23964 6177
rect 23906 6168 23918 6171
rect 23440 6140 23918 6168
rect 23440 6128 23446 6140
rect 23906 6137 23918 6140
rect 23952 6137 23964 6171
rect 23906 6131 23964 6137
rect 25038 6128 25044 6180
rect 25096 6168 25102 6180
rect 25593 6171 25651 6177
rect 25593 6168 25605 6171
rect 25096 6140 25605 6168
rect 25096 6128 25102 6140
rect 25593 6137 25605 6140
rect 25639 6137 25651 6171
rect 25593 6131 25651 6137
rect 18049 6103 18107 6109
rect 18049 6069 18061 6103
rect 18095 6069 18107 6103
rect 18049 6063 18107 6069
rect 18322 6060 18328 6112
rect 18380 6100 18386 6112
rect 18417 6103 18475 6109
rect 18417 6100 18429 6103
rect 18380 6072 18429 6100
rect 18380 6060 18386 6072
rect 18417 6069 18429 6072
rect 18463 6100 18475 6103
rect 20070 6100 20076 6112
rect 18463 6072 20076 6100
rect 18463 6069 18475 6072
rect 18417 6063 18475 6069
rect 20070 6060 20076 6072
rect 20128 6060 20134 6112
rect 22186 6060 22192 6112
rect 22244 6100 22250 6112
rect 22373 6103 22431 6109
rect 22373 6100 22385 6103
rect 22244 6072 22385 6100
rect 22244 6060 22250 6072
rect 22373 6069 22385 6072
rect 22419 6069 22431 6103
rect 22373 6063 22431 6069
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1397 5899 1455 5905
rect 1397 5865 1409 5899
rect 1443 5896 1455 5899
rect 1854 5896 1860 5908
rect 1443 5868 1860 5896
rect 1443 5865 1455 5868
rect 1397 5859 1455 5865
rect 1854 5856 1860 5868
rect 1912 5856 1918 5908
rect 3142 5856 3148 5908
rect 3200 5896 3206 5908
rect 3421 5899 3479 5905
rect 3421 5896 3433 5899
rect 3200 5868 3433 5896
rect 3200 5856 3206 5868
rect 3421 5865 3433 5868
rect 3467 5865 3479 5899
rect 4246 5896 4252 5908
rect 4207 5868 4252 5896
rect 3421 5859 3479 5865
rect 4246 5856 4252 5868
rect 4304 5856 4310 5908
rect 4706 5896 4712 5908
rect 4667 5868 4712 5896
rect 4706 5856 4712 5868
rect 4764 5856 4770 5908
rect 5074 5856 5080 5908
rect 5132 5896 5138 5908
rect 5261 5899 5319 5905
rect 5261 5896 5273 5899
rect 5132 5868 5273 5896
rect 5132 5856 5138 5868
rect 5261 5865 5273 5868
rect 5307 5865 5319 5899
rect 5261 5859 5319 5865
rect 6914 5856 6920 5908
rect 6972 5896 6978 5908
rect 7193 5899 7251 5905
rect 7193 5896 7205 5899
rect 6972 5868 7205 5896
rect 6972 5856 6978 5868
rect 7193 5865 7205 5868
rect 7239 5865 7251 5899
rect 7193 5859 7251 5865
rect 7837 5899 7895 5905
rect 7837 5865 7849 5899
rect 7883 5896 7895 5899
rect 7926 5896 7932 5908
rect 7883 5868 7932 5896
rect 7883 5865 7895 5868
rect 7837 5859 7895 5865
rect 7926 5856 7932 5868
rect 7984 5856 7990 5908
rect 9674 5896 9680 5908
rect 9635 5868 9680 5896
rect 9674 5856 9680 5868
rect 9732 5856 9738 5908
rect 11514 5896 11520 5908
rect 11475 5868 11520 5896
rect 11514 5856 11520 5868
rect 11572 5856 11578 5908
rect 11885 5899 11943 5905
rect 11885 5865 11897 5899
rect 11931 5896 11943 5899
rect 13078 5896 13084 5908
rect 11931 5868 13084 5896
rect 11931 5865 11943 5868
rect 11885 5859 11943 5865
rect 13078 5856 13084 5868
rect 13136 5856 13142 5908
rect 13262 5856 13268 5908
rect 13320 5896 13326 5908
rect 13722 5896 13728 5908
rect 13320 5868 13728 5896
rect 13320 5856 13326 5868
rect 13722 5856 13728 5868
rect 13780 5896 13786 5908
rect 14093 5899 14151 5905
rect 14093 5896 14105 5899
rect 13780 5868 14105 5896
rect 13780 5856 13786 5868
rect 14093 5865 14105 5868
rect 14139 5896 14151 5899
rect 15286 5896 15292 5908
rect 14139 5868 15292 5896
rect 14139 5865 14151 5868
rect 14093 5859 14151 5865
rect 15286 5856 15292 5868
rect 15344 5856 15350 5908
rect 15654 5896 15660 5908
rect 15615 5868 15660 5896
rect 15654 5856 15660 5868
rect 15712 5856 15718 5908
rect 15749 5899 15807 5905
rect 15749 5865 15761 5899
rect 15795 5896 15807 5899
rect 15930 5896 15936 5908
rect 15795 5868 15936 5896
rect 15795 5865 15807 5868
rect 15749 5859 15807 5865
rect 15930 5856 15936 5868
rect 15988 5856 15994 5908
rect 16666 5896 16672 5908
rect 16627 5868 16672 5896
rect 16666 5856 16672 5868
rect 16724 5856 16730 5908
rect 16850 5896 16856 5908
rect 16811 5868 16856 5896
rect 16850 5856 16856 5868
rect 16908 5856 16914 5908
rect 17678 5896 17684 5908
rect 17639 5868 17684 5896
rect 17678 5856 17684 5868
rect 17736 5856 17742 5908
rect 18230 5896 18236 5908
rect 18191 5868 18236 5896
rect 18230 5856 18236 5868
rect 18288 5856 18294 5908
rect 21177 5899 21235 5905
rect 21177 5865 21189 5899
rect 21223 5896 21235 5899
rect 21266 5896 21272 5908
rect 21223 5868 21272 5896
rect 21223 5865 21235 5868
rect 21177 5859 21235 5865
rect 21266 5856 21272 5868
rect 21324 5856 21330 5908
rect 22002 5856 22008 5908
rect 22060 5896 22066 5908
rect 22370 5896 22376 5908
rect 22060 5868 22376 5896
rect 22060 5856 22066 5868
rect 22370 5856 22376 5868
rect 22428 5856 22434 5908
rect 22925 5899 22983 5905
rect 22925 5865 22937 5899
rect 22971 5896 22983 5899
rect 23382 5896 23388 5908
rect 22971 5868 23388 5896
rect 22971 5865 22983 5868
rect 22925 5859 22983 5865
rect 23382 5856 23388 5868
rect 23440 5856 23446 5908
rect 23474 5856 23480 5908
rect 23532 5896 23538 5908
rect 23661 5899 23719 5905
rect 23661 5896 23673 5899
rect 23532 5868 23673 5896
rect 23532 5856 23538 5868
rect 23661 5865 23673 5868
rect 23707 5896 23719 5899
rect 23750 5896 23756 5908
rect 23707 5868 23756 5896
rect 23707 5865 23719 5868
rect 23661 5859 23719 5865
rect 23750 5856 23756 5868
rect 23808 5856 23814 5908
rect 24029 5899 24087 5905
rect 24029 5865 24041 5899
rect 24075 5865 24087 5899
rect 25038 5896 25044 5908
rect 24999 5868 25044 5896
rect 24029 5859 24087 5865
rect 2866 5828 2872 5840
rect 2779 5800 2872 5828
rect 2866 5788 2872 5800
rect 2924 5828 2930 5840
rect 3602 5828 3608 5840
rect 2924 5800 3608 5828
rect 2924 5788 2930 5800
rect 3602 5788 3608 5800
rect 3660 5788 3666 5840
rect 5534 5788 5540 5840
rect 5592 5828 5598 5840
rect 6181 5831 6239 5837
rect 6181 5828 6193 5831
rect 5592 5800 6193 5828
rect 5592 5788 5598 5800
rect 6181 5797 6193 5800
rect 6227 5828 6239 5831
rect 7006 5828 7012 5840
rect 6227 5800 7012 5828
rect 6227 5797 6239 5800
rect 6181 5791 6239 5797
rect 7006 5788 7012 5800
rect 7064 5788 7070 5840
rect 11146 5788 11152 5840
rect 11204 5828 11210 5840
rect 12342 5828 12348 5840
rect 11204 5800 12348 5828
rect 11204 5788 11210 5800
rect 12342 5788 12348 5800
rect 12400 5788 12406 5840
rect 15948 5828 15976 5856
rect 16574 5828 16580 5840
rect 15948 5800 16580 5828
rect 16574 5788 16580 5800
rect 16632 5788 16638 5840
rect 19242 5788 19248 5840
rect 19300 5828 19306 5840
rect 20898 5828 20904 5840
rect 19300 5800 20904 5828
rect 19300 5788 19306 5800
rect 20898 5788 20904 5800
rect 20956 5788 20962 5840
rect 21818 5837 21824 5840
rect 21812 5828 21824 5837
rect 21779 5800 21824 5828
rect 21812 5791 21824 5800
rect 21818 5788 21824 5791
rect 21876 5788 21882 5840
rect 23566 5788 23572 5840
rect 23624 5828 23630 5840
rect 24044 5828 24072 5859
rect 25038 5856 25044 5868
rect 25096 5896 25102 5908
rect 25409 5899 25467 5905
rect 25409 5896 25421 5899
rect 25096 5868 25421 5896
rect 25096 5856 25102 5868
rect 25409 5865 25421 5868
rect 25455 5865 25467 5899
rect 25409 5859 25467 5865
rect 25869 5899 25927 5905
rect 25869 5865 25881 5899
rect 25915 5896 25927 5899
rect 26142 5896 26148 5908
rect 25915 5868 26148 5896
rect 25915 5865 25927 5868
rect 25869 5859 25927 5865
rect 26142 5856 26148 5868
rect 26200 5856 26206 5908
rect 23624 5800 24072 5828
rect 23624 5788 23630 5800
rect 1394 5720 1400 5772
rect 1452 5760 1458 5772
rect 1765 5763 1823 5769
rect 1765 5760 1777 5763
rect 1452 5732 1777 5760
rect 1452 5720 1458 5732
rect 1765 5729 1777 5732
rect 1811 5729 1823 5763
rect 1765 5723 1823 5729
rect 1857 5763 1915 5769
rect 1857 5729 1869 5763
rect 1903 5760 1915 5763
rect 1946 5760 1952 5772
rect 1903 5732 1952 5760
rect 1903 5729 1915 5732
rect 1857 5723 1915 5729
rect 1946 5720 1952 5732
rect 2004 5720 2010 5772
rect 4338 5720 4344 5772
rect 4396 5760 4402 5772
rect 4617 5763 4675 5769
rect 4617 5760 4629 5763
rect 4396 5732 4629 5760
rect 4396 5720 4402 5732
rect 4617 5729 4629 5732
rect 4663 5729 4675 5763
rect 4617 5723 4675 5729
rect 6273 5763 6331 5769
rect 6273 5729 6285 5763
rect 6319 5760 6331 5763
rect 6822 5760 6828 5772
rect 6319 5732 6828 5760
rect 6319 5729 6331 5732
rect 6273 5723 6331 5729
rect 2041 5695 2099 5701
rect 2041 5661 2053 5695
rect 2087 5661 2099 5695
rect 2041 5655 2099 5661
rect 2961 5695 3019 5701
rect 2961 5661 2973 5695
rect 3007 5692 3019 5695
rect 3970 5692 3976 5704
rect 3007 5664 3976 5692
rect 3007 5661 3019 5664
rect 2961 5655 3019 5661
rect 2056 5624 2084 5655
rect 3970 5652 3976 5664
rect 4028 5652 4034 5704
rect 4062 5652 4068 5704
rect 4120 5692 4126 5704
rect 4893 5695 4951 5701
rect 4893 5692 4905 5695
rect 4120 5664 4905 5692
rect 4120 5652 4126 5664
rect 4893 5661 4905 5664
rect 4939 5692 4951 5695
rect 5074 5692 5080 5704
rect 4939 5664 5080 5692
rect 4939 5661 4951 5664
rect 4893 5655 4951 5661
rect 5074 5652 5080 5664
rect 5132 5652 5138 5704
rect 5721 5695 5779 5701
rect 5721 5661 5733 5695
rect 5767 5692 5779 5695
rect 6288 5692 6316 5723
rect 6822 5720 6828 5732
rect 6880 5720 6886 5772
rect 7282 5720 7288 5772
rect 7340 5760 7346 5772
rect 7745 5763 7803 5769
rect 7745 5760 7757 5763
rect 7340 5732 7757 5760
rect 7340 5720 7346 5732
rect 7745 5729 7757 5732
rect 7791 5729 7803 5763
rect 10042 5760 10048 5772
rect 10003 5732 10048 5760
rect 7745 5723 7803 5729
rect 10042 5720 10048 5732
rect 10100 5720 10106 5772
rect 11882 5720 11888 5772
rect 11940 5760 11946 5772
rect 12233 5763 12291 5769
rect 12233 5760 12245 5763
rect 11940 5732 12245 5760
rect 11940 5720 11946 5732
rect 12233 5729 12245 5732
rect 12279 5760 12291 5763
rect 12710 5760 12716 5772
rect 12279 5732 12716 5760
rect 12279 5729 12291 5732
rect 12233 5723 12291 5729
rect 12710 5720 12716 5732
rect 12768 5720 12774 5772
rect 13170 5720 13176 5772
rect 13228 5760 13234 5772
rect 14826 5760 14832 5772
rect 13228 5732 14832 5760
rect 13228 5720 13234 5732
rect 14826 5720 14832 5732
rect 14884 5720 14890 5772
rect 18230 5720 18236 5772
rect 18288 5760 18294 5772
rect 18325 5763 18383 5769
rect 18325 5760 18337 5763
rect 18288 5732 18337 5760
rect 18288 5720 18294 5732
rect 18325 5729 18337 5732
rect 18371 5729 18383 5763
rect 18325 5723 18383 5729
rect 19429 5763 19487 5769
rect 19429 5729 19441 5763
rect 19475 5760 19487 5763
rect 19978 5760 19984 5772
rect 19475 5732 19984 5760
rect 19475 5729 19487 5732
rect 19429 5723 19487 5729
rect 19978 5720 19984 5732
rect 20036 5720 20042 5772
rect 20530 5720 20536 5772
rect 20588 5760 20594 5772
rect 20806 5760 20812 5772
rect 20588 5732 20812 5760
rect 20588 5720 20594 5732
rect 20806 5720 20812 5732
rect 20864 5760 20870 5772
rect 21545 5763 21603 5769
rect 21545 5760 21557 5763
rect 20864 5732 21557 5760
rect 20864 5720 20870 5732
rect 21545 5729 21557 5732
rect 21591 5760 21603 5763
rect 23290 5760 23296 5772
rect 21591 5732 23296 5760
rect 21591 5729 21603 5732
rect 21545 5723 21603 5729
rect 23290 5720 23296 5732
rect 23348 5720 23354 5772
rect 23474 5720 23480 5772
rect 23532 5760 23538 5772
rect 24397 5763 24455 5769
rect 24397 5760 24409 5763
rect 23532 5732 24409 5760
rect 23532 5720 23538 5732
rect 24397 5729 24409 5732
rect 24443 5729 24455 5763
rect 24397 5723 24455 5729
rect 24489 5763 24547 5769
rect 24489 5729 24501 5763
rect 24535 5760 24547 5763
rect 24762 5760 24768 5772
rect 24535 5732 24768 5760
rect 24535 5729 24547 5732
rect 24489 5723 24547 5729
rect 24762 5720 24768 5732
rect 24820 5720 24826 5772
rect 6454 5692 6460 5704
rect 5767 5664 6316 5692
rect 6415 5664 6460 5692
rect 5767 5661 5779 5664
rect 5721 5655 5779 5661
rect 6454 5652 6460 5664
rect 6512 5652 6518 5704
rect 8018 5692 8024 5704
rect 7979 5664 8024 5692
rect 8018 5652 8024 5664
rect 8076 5652 8082 5704
rect 8849 5695 8907 5701
rect 8849 5661 8861 5695
rect 8895 5692 8907 5695
rect 10137 5695 10195 5701
rect 10137 5692 10149 5695
rect 8895 5664 10149 5692
rect 8895 5661 8907 5664
rect 8849 5655 8907 5661
rect 10137 5661 10149 5664
rect 10183 5661 10195 5695
rect 10137 5655 10195 5661
rect 10229 5695 10287 5701
rect 10229 5661 10241 5695
rect 10275 5661 10287 5695
rect 11974 5692 11980 5704
rect 11935 5664 11980 5692
rect 10229 5655 10287 5661
rect 3142 5624 3148 5636
rect 2056 5596 3148 5624
rect 3142 5584 3148 5596
rect 3200 5584 3206 5636
rect 3881 5627 3939 5633
rect 3881 5593 3893 5627
rect 3927 5624 3939 5627
rect 5350 5624 5356 5636
rect 3927 5596 5356 5624
rect 3927 5593 3939 5596
rect 3881 5587 3939 5593
rect 5350 5584 5356 5596
rect 5408 5584 5414 5636
rect 5810 5624 5816 5636
rect 5771 5596 5816 5624
rect 5810 5584 5816 5596
rect 5868 5584 5874 5636
rect 7377 5627 7435 5633
rect 7377 5593 7389 5627
rect 7423 5624 7435 5627
rect 8864 5624 8892 5655
rect 7423 5596 8892 5624
rect 7423 5593 7435 5596
rect 7377 5587 7435 5593
rect 9950 5584 9956 5636
rect 10008 5624 10014 5636
rect 10244 5624 10272 5655
rect 11974 5652 11980 5664
rect 12032 5652 12038 5704
rect 15838 5692 15844 5704
rect 15799 5664 15844 5692
rect 15838 5652 15844 5664
rect 15896 5652 15902 5704
rect 17405 5695 17463 5701
rect 17405 5661 17417 5695
rect 17451 5692 17463 5695
rect 17494 5692 17500 5704
rect 17451 5664 17500 5692
rect 17451 5661 17463 5664
rect 17405 5655 17463 5661
rect 17494 5652 17500 5664
rect 17552 5652 17558 5704
rect 18414 5692 18420 5704
rect 18375 5664 18420 5692
rect 18414 5652 18420 5664
rect 18472 5652 18478 5704
rect 19518 5652 19524 5704
rect 19576 5692 19582 5704
rect 19613 5695 19671 5701
rect 19613 5692 19625 5695
rect 19576 5664 19625 5692
rect 19576 5652 19582 5664
rect 19613 5661 19625 5664
rect 19659 5661 19671 5695
rect 24578 5692 24584 5704
rect 24539 5664 24584 5692
rect 19613 5655 19671 5661
rect 24578 5652 24584 5664
rect 24636 5652 24642 5704
rect 10008 5596 10272 5624
rect 15289 5627 15347 5633
rect 10008 5584 10014 5596
rect 15289 5593 15301 5627
rect 15335 5624 15347 5627
rect 16022 5624 16028 5636
rect 15335 5596 16028 5624
rect 15335 5593 15347 5596
rect 15289 5587 15347 5593
rect 16022 5584 16028 5596
rect 16080 5584 16086 5636
rect 17865 5627 17923 5633
rect 17865 5593 17877 5627
rect 17911 5624 17923 5627
rect 18782 5624 18788 5636
rect 17911 5596 18788 5624
rect 17911 5593 17923 5596
rect 17865 5587 17923 5593
rect 18782 5584 18788 5596
rect 18840 5624 18846 5636
rect 19337 5627 19395 5633
rect 19337 5624 19349 5627
rect 18840 5596 19349 5624
rect 18840 5584 18846 5596
rect 19337 5593 19349 5596
rect 19383 5593 19395 5627
rect 19337 5587 19395 5593
rect 19426 5584 19432 5636
rect 19484 5624 19490 5636
rect 19484 5596 20576 5624
rect 19484 5584 19490 5596
rect 2498 5556 2504 5568
rect 2411 5528 2504 5556
rect 2498 5516 2504 5528
rect 2556 5556 2562 5568
rect 2866 5556 2872 5568
rect 2556 5528 2872 5556
rect 2556 5516 2562 5528
rect 2866 5516 2872 5528
rect 2924 5516 2930 5568
rect 6917 5559 6975 5565
rect 6917 5525 6929 5559
rect 6963 5556 6975 5559
rect 7006 5556 7012 5568
rect 6963 5528 7012 5556
rect 6963 5525 6975 5528
rect 6917 5519 6975 5525
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 8478 5556 8484 5568
rect 8439 5528 8484 5556
rect 8478 5516 8484 5528
rect 8536 5516 8542 5568
rect 9214 5556 9220 5568
rect 9175 5528 9220 5556
rect 9214 5516 9220 5528
rect 9272 5516 9278 5568
rect 10042 5516 10048 5568
rect 10100 5556 10106 5568
rect 10594 5556 10600 5568
rect 10100 5528 10600 5556
rect 10100 5516 10106 5528
rect 10594 5516 10600 5528
rect 10652 5556 10658 5568
rect 10689 5559 10747 5565
rect 10689 5556 10701 5559
rect 10652 5528 10701 5556
rect 10652 5516 10658 5528
rect 10689 5525 10701 5528
rect 10735 5525 10747 5559
rect 11146 5556 11152 5568
rect 11107 5528 11152 5556
rect 10689 5519 10747 5525
rect 11146 5516 11152 5528
rect 11204 5516 11210 5568
rect 12158 5516 12164 5568
rect 12216 5556 12222 5568
rect 13357 5559 13415 5565
rect 13357 5556 13369 5559
rect 12216 5528 13369 5556
rect 12216 5516 12222 5528
rect 13357 5525 13369 5528
rect 13403 5525 13415 5559
rect 13357 5519 13415 5525
rect 14461 5559 14519 5565
rect 14461 5525 14473 5559
rect 14507 5556 14519 5559
rect 14734 5556 14740 5568
rect 14507 5528 14740 5556
rect 14507 5525 14519 5528
rect 14461 5519 14519 5525
rect 14734 5516 14740 5528
rect 14792 5516 14798 5568
rect 15105 5559 15163 5565
rect 15105 5525 15117 5559
rect 15151 5556 15163 5559
rect 15378 5556 15384 5568
rect 15151 5528 15384 5556
rect 15151 5525 15163 5528
rect 15105 5519 15163 5525
rect 15378 5516 15384 5528
rect 15436 5516 15442 5568
rect 15930 5516 15936 5568
rect 15988 5556 15994 5568
rect 16393 5559 16451 5565
rect 16393 5556 16405 5559
rect 15988 5528 16405 5556
rect 15988 5516 15994 5528
rect 16393 5525 16405 5528
rect 16439 5556 16451 5559
rect 16482 5556 16488 5568
rect 16439 5528 16488 5556
rect 16439 5525 16451 5528
rect 16393 5519 16451 5525
rect 16482 5516 16488 5528
rect 16540 5516 16546 5568
rect 18969 5559 19027 5565
rect 18969 5525 18981 5559
rect 19015 5556 19027 5559
rect 19242 5556 19248 5568
rect 19015 5528 19248 5556
rect 19015 5525 19027 5528
rect 18969 5519 19027 5525
rect 19242 5516 19248 5528
rect 19300 5516 19306 5568
rect 20162 5516 20168 5568
rect 20220 5556 20226 5568
rect 20441 5559 20499 5565
rect 20441 5556 20453 5559
rect 20220 5528 20453 5556
rect 20220 5516 20226 5528
rect 20441 5525 20453 5528
rect 20487 5525 20499 5559
rect 20548 5556 20576 5596
rect 24854 5556 24860 5568
rect 20548 5528 24860 5556
rect 20441 5519 20499 5525
rect 24854 5516 24860 5528
rect 24912 5516 24918 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 1946 5312 1952 5364
rect 2004 5352 2010 5364
rect 2961 5355 3019 5361
rect 2961 5352 2973 5355
rect 2004 5324 2973 5352
rect 2004 5312 2010 5324
rect 2961 5321 2973 5324
rect 3007 5352 3019 5355
rect 3418 5352 3424 5364
rect 3007 5324 3424 5352
rect 3007 5321 3019 5324
rect 2961 5315 3019 5321
rect 3418 5312 3424 5324
rect 3476 5312 3482 5364
rect 4338 5352 4344 5364
rect 4299 5324 4344 5352
rect 4338 5312 4344 5324
rect 4396 5312 4402 5364
rect 4706 5352 4712 5364
rect 4667 5324 4712 5352
rect 4706 5312 4712 5324
rect 4764 5312 4770 5364
rect 5074 5312 5080 5364
rect 5132 5312 5138 5364
rect 5169 5355 5227 5361
rect 5169 5321 5181 5355
rect 5215 5352 5227 5355
rect 5350 5352 5356 5364
rect 5215 5324 5356 5352
rect 5215 5321 5227 5324
rect 5169 5315 5227 5321
rect 5350 5312 5356 5324
rect 5408 5312 5414 5364
rect 6914 5312 6920 5364
rect 6972 5352 6978 5364
rect 7561 5355 7619 5361
rect 7561 5352 7573 5355
rect 6972 5324 7573 5352
rect 6972 5312 6978 5324
rect 7561 5321 7573 5324
rect 7607 5321 7619 5355
rect 7561 5315 7619 5321
rect 8202 5312 8208 5364
rect 8260 5352 8266 5364
rect 8260 5324 8616 5352
rect 8260 5312 8266 5324
rect 5092 5284 5120 5312
rect 8588 5296 8616 5324
rect 9950 5312 9956 5364
rect 10008 5352 10014 5364
rect 10137 5355 10195 5361
rect 10137 5352 10149 5355
rect 10008 5324 10149 5352
rect 10008 5312 10014 5324
rect 10137 5321 10149 5324
rect 10183 5321 10195 5355
rect 11882 5352 11888 5364
rect 11843 5324 11888 5352
rect 10137 5315 10195 5321
rect 11882 5312 11888 5324
rect 11940 5312 11946 5364
rect 12986 5312 12992 5364
rect 13044 5352 13050 5364
rect 13449 5355 13507 5361
rect 13449 5352 13461 5355
rect 13044 5324 13461 5352
rect 13044 5312 13050 5324
rect 13449 5321 13461 5324
rect 13495 5321 13507 5355
rect 13814 5352 13820 5364
rect 13775 5324 13820 5352
rect 13449 5315 13507 5321
rect 6273 5287 6331 5293
rect 5092 5256 5764 5284
rect 2041 5219 2099 5225
rect 2041 5185 2053 5219
rect 2087 5216 2099 5219
rect 2498 5216 2504 5228
rect 2087 5188 2504 5216
rect 2087 5185 2099 5188
rect 2041 5179 2099 5185
rect 2498 5176 2504 5188
rect 2556 5176 2562 5228
rect 2774 5176 2780 5228
rect 2832 5216 2838 5228
rect 3605 5219 3663 5225
rect 3605 5216 3617 5219
rect 2832 5188 3617 5216
rect 2832 5176 2838 5188
rect 3605 5185 3617 5188
rect 3651 5216 3663 5219
rect 4062 5216 4068 5228
rect 3651 5188 4068 5216
rect 3651 5185 3663 5188
rect 3605 5179 3663 5185
rect 4062 5176 4068 5188
rect 4120 5176 4126 5228
rect 5077 5219 5135 5225
rect 5077 5185 5089 5219
rect 5123 5216 5135 5219
rect 5166 5216 5172 5228
rect 5123 5188 5172 5216
rect 5123 5185 5135 5188
rect 5077 5179 5135 5185
rect 5166 5176 5172 5188
rect 5224 5216 5230 5228
rect 5736 5225 5764 5256
rect 6273 5253 6285 5287
rect 6319 5284 6331 5287
rect 6454 5284 6460 5296
rect 6319 5256 6460 5284
rect 6319 5253 6331 5256
rect 6273 5247 6331 5253
rect 6454 5244 6460 5256
rect 6512 5284 6518 5296
rect 7101 5287 7159 5293
rect 7101 5284 7113 5287
rect 6512 5256 7113 5284
rect 6512 5244 6518 5256
rect 7101 5253 7113 5256
rect 7147 5284 7159 5287
rect 8018 5284 8024 5296
rect 7147 5256 8024 5284
rect 7147 5253 7159 5256
rect 7101 5247 7159 5253
rect 8018 5244 8024 5256
rect 8076 5244 8082 5296
rect 8570 5244 8576 5296
rect 8628 5284 8634 5296
rect 10689 5287 10747 5293
rect 10689 5284 10701 5287
rect 8628 5256 10701 5284
rect 8628 5244 8634 5256
rect 10689 5253 10701 5256
rect 10735 5253 10747 5287
rect 10689 5247 10747 5253
rect 10778 5244 10784 5296
rect 10836 5284 10842 5296
rect 10962 5284 10968 5296
rect 10836 5256 10968 5284
rect 10836 5244 10842 5256
rect 10962 5244 10968 5256
rect 11020 5244 11026 5296
rect 12894 5244 12900 5296
rect 12952 5284 12958 5296
rect 13265 5287 13323 5293
rect 13265 5284 13277 5287
rect 12952 5256 13277 5284
rect 12952 5244 12958 5256
rect 13265 5253 13277 5256
rect 13311 5253 13323 5287
rect 13464 5284 13492 5315
rect 13814 5312 13820 5324
rect 13872 5312 13878 5364
rect 14001 5355 14059 5361
rect 14001 5321 14013 5355
rect 14047 5352 14059 5355
rect 14274 5352 14280 5364
rect 14047 5324 14280 5352
rect 14047 5321 14059 5324
rect 14001 5315 14059 5321
rect 14274 5312 14280 5324
rect 14332 5312 14338 5364
rect 15381 5355 15439 5361
rect 15381 5321 15393 5355
rect 15427 5352 15439 5355
rect 15654 5352 15660 5364
rect 15427 5324 15660 5352
rect 15427 5321 15439 5324
rect 15381 5315 15439 5321
rect 15654 5312 15660 5324
rect 15712 5312 15718 5364
rect 16574 5352 16580 5364
rect 16535 5324 16580 5352
rect 16574 5312 16580 5324
rect 16632 5312 16638 5364
rect 18230 5352 18236 5364
rect 18191 5324 18236 5352
rect 18230 5312 18236 5324
rect 18288 5312 18294 5364
rect 18322 5312 18328 5364
rect 18380 5352 18386 5364
rect 18601 5355 18659 5361
rect 18601 5352 18613 5355
rect 18380 5324 18613 5352
rect 18380 5312 18386 5324
rect 18601 5321 18613 5324
rect 18647 5321 18659 5355
rect 21266 5352 21272 5364
rect 21227 5324 21272 5352
rect 18601 5315 18659 5321
rect 21266 5312 21272 5324
rect 21324 5312 21330 5364
rect 22094 5312 22100 5364
rect 22152 5352 22158 5364
rect 22281 5355 22339 5361
rect 22281 5352 22293 5355
rect 22152 5324 22293 5352
rect 22152 5312 22158 5324
rect 22281 5321 22293 5324
rect 22327 5321 22339 5355
rect 22281 5315 22339 5321
rect 23109 5355 23167 5361
rect 23109 5321 23121 5355
rect 23155 5352 23167 5355
rect 23382 5352 23388 5364
rect 23155 5324 23388 5352
rect 23155 5321 23167 5324
rect 23109 5315 23167 5321
rect 23382 5312 23388 5324
rect 23440 5312 23446 5364
rect 23658 5352 23664 5364
rect 23619 5324 23664 5352
rect 23658 5312 23664 5324
rect 23716 5312 23722 5364
rect 24670 5352 24676 5364
rect 24631 5324 24676 5352
rect 24670 5312 24676 5324
rect 24728 5312 24734 5364
rect 26234 5312 26240 5364
rect 26292 5352 26298 5364
rect 26329 5355 26387 5361
rect 26329 5352 26341 5355
rect 26292 5324 26341 5352
rect 26292 5312 26298 5324
rect 26329 5321 26341 5324
rect 26375 5321 26387 5355
rect 26329 5315 26387 5321
rect 15562 5284 15568 5296
rect 13464 5256 14596 5284
rect 15523 5256 15568 5284
rect 13265 5247 13323 5253
rect 5629 5219 5687 5225
rect 5629 5216 5641 5219
rect 5224 5188 5641 5216
rect 5224 5176 5230 5188
rect 5629 5185 5641 5188
rect 5675 5185 5687 5219
rect 5629 5179 5687 5185
rect 5721 5219 5779 5225
rect 5721 5185 5733 5219
rect 5767 5185 5779 5219
rect 7466 5216 7472 5228
rect 7379 5188 7472 5216
rect 5721 5179 5779 5185
rect 7466 5176 7472 5188
rect 7524 5216 7530 5228
rect 8202 5216 8208 5228
rect 7524 5188 8208 5216
rect 7524 5176 7530 5188
rect 8202 5176 8208 5188
rect 8260 5176 8266 5228
rect 9214 5176 9220 5228
rect 9272 5216 9278 5228
rect 9677 5219 9735 5225
rect 9677 5216 9689 5219
rect 9272 5188 9689 5216
rect 9272 5176 9278 5188
rect 9677 5185 9689 5188
rect 9723 5185 9735 5219
rect 9677 5179 9735 5185
rect 10594 5176 10600 5228
rect 10652 5216 10658 5228
rect 11238 5216 11244 5228
rect 10652 5188 11244 5216
rect 10652 5176 10658 5188
rect 11238 5176 11244 5188
rect 11296 5176 11302 5228
rect 11330 5176 11336 5228
rect 11388 5216 11394 5228
rect 12161 5219 12219 5225
rect 12161 5216 12173 5219
rect 11388 5188 12173 5216
rect 11388 5176 11394 5188
rect 12161 5185 12173 5188
rect 12207 5185 12219 5219
rect 12986 5216 12992 5228
rect 12947 5188 12992 5216
rect 12161 5179 12219 5185
rect 1762 5148 1768 5160
rect 1723 5120 1768 5148
rect 1762 5108 1768 5120
rect 1820 5108 1826 5160
rect 2869 5151 2927 5157
rect 2869 5117 2881 5151
rect 2915 5148 2927 5151
rect 3142 5148 3148 5160
rect 2915 5120 3148 5148
rect 2915 5117 2927 5120
rect 2869 5111 2927 5117
rect 3142 5108 3148 5120
rect 3200 5148 3206 5160
rect 3421 5151 3479 5157
rect 3421 5148 3433 5151
rect 3200 5120 3433 5148
rect 3200 5108 3206 5120
rect 3421 5117 3433 5120
rect 3467 5148 3479 5151
rect 3786 5148 3792 5160
rect 3467 5120 3792 5148
rect 3467 5117 3479 5120
rect 3421 5111 3479 5117
rect 3786 5108 3792 5120
rect 3844 5108 3850 5160
rect 5537 5151 5595 5157
rect 5537 5117 5549 5151
rect 5583 5148 5595 5151
rect 5810 5148 5816 5160
rect 5583 5120 5816 5148
rect 5583 5117 5595 5120
rect 5537 5111 5595 5117
rect 5810 5108 5816 5120
rect 5868 5108 5874 5160
rect 7098 5108 7104 5160
rect 7156 5148 7162 5160
rect 7834 5148 7840 5160
rect 7156 5120 7840 5148
rect 7156 5108 7162 5120
rect 7834 5108 7840 5120
rect 7892 5148 7898 5160
rect 7929 5151 7987 5157
rect 7929 5148 7941 5151
rect 7892 5120 7941 5148
rect 7892 5108 7898 5120
rect 7929 5117 7941 5120
rect 7975 5117 7987 5151
rect 9122 5148 9128 5160
rect 7929 5111 7987 5117
rect 8956 5120 9128 5148
rect 3326 5080 3332 5092
rect 3287 5052 3332 5080
rect 3326 5040 3332 5052
rect 3384 5040 3390 5092
rect 6641 5083 6699 5089
rect 6641 5049 6653 5083
rect 6687 5080 6699 5083
rect 7282 5080 7288 5092
rect 6687 5052 7288 5080
rect 6687 5049 6699 5052
rect 6641 5043 6699 5049
rect 7282 5040 7288 5052
rect 7340 5040 7346 5092
rect 1394 5012 1400 5024
rect 1355 4984 1400 5012
rect 1394 4972 1400 4984
rect 1452 4972 1458 5024
rect 1670 4972 1676 5024
rect 1728 5012 1734 5024
rect 1857 5015 1915 5021
rect 1857 5012 1869 5015
rect 1728 4984 1869 5012
rect 1728 4972 1734 4984
rect 1857 4981 1869 4984
rect 1903 5012 1915 5015
rect 2406 5012 2412 5024
rect 1903 4984 2412 5012
rect 1903 4981 1915 4984
rect 1857 4975 1915 4981
rect 2406 4972 2412 4984
rect 2464 4972 2470 5024
rect 6270 4972 6276 5024
rect 6328 5012 6334 5024
rect 6822 5012 6828 5024
rect 6328 4984 6828 5012
rect 6328 4972 6334 4984
rect 6822 4972 6828 4984
rect 6880 4972 6886 5024
rect 8018 4972 8024 5024
rect 8076 5012 8082 5024
rect 8662 5012 8668 5024
rect 8076 4984 8121 5012
rect 8623 4984 8668 5012
rect 8076 4972 8082 4984
rect 8662 4972 8668 4984
rect 8720 4972 8726 5024
rect 8846 4972 8852 5024
rect 8904 5012 8910 5024
rect 8956 5021 8984 5120
rect 9122 5108 9128 5120
rect 9180 5148 9186 5160
rect 9585 5151 9643 5157
rect 9585 5148 9597 5151
rect 9180 5120 9597 5148
rect 9180 5108 9186 5120
rect 9585 5117 9597 5120
rect 9631 5117 9643 5151
rect 9585 5111 9643 5117
rect 10042 5108 10048 5160
rect 10100 5148 10106 5160
rect 10870 5148 10876 5160
rect 10100 5120 10876 5148
rect 10100 5108 10106 5120
rect 10870 5108 10876 5120
rect 10928 5108 10934 5160
rect 12176 5148 12204 5179
rect 12986 5176 12992 5188
rect 13044 5176 13050 5228
rect 13722 5176 13728 5228
rect 13780 5216 13786 5228
rect 14568 5225 14596 5256
rect 15562 5244 15568 5256
rect 15620 5244 15626 5296
rect 15838 5244 15844 5296
rect 15896 5284 15902 5296
rect 16945 5287 17003 5293
rect 16945 5284 16957 5287
rect 15896 5256 16957 5284
rect 15896 5244 15902 5256
rect 14461 5219 14519 5225
rect 14461 5216 14473 5219
rect 13780 5188 14473 5216
rect 13780 5176 13786 5188
rect 14461 5185 14473 5188
rect 14507 5185 14519 5219
rect 14461 5179 14519 5185
rect 14553 5219 14611 5225
rect 14553 5185 14565 5219
rect 14599 5185 14611 5219
rect 16022 5216 16028 5228
rect 15983 5188 16028 5216
rect 14553 5179 14611 5185
rect 16022 5176 16028 5188
rect 16080 5176 16086 5228
rect 16132 5225 16160 5256
rect 16945 5253 16957 5256
rect 16991 5284 17003 5287
rect 17313 5287 17371 5293
rect 17313 5284 17325 5287
rect 16991 5256 17325 5284
rect 16991 5253 17003 5256
rect 16945 5247 17003 5253
rect 17313 5253 17325 5256
rect 17359 5253 17371 5287
rect 17313 5247 17371 5253
rect 23477 5287 23535 5293
rect 23477 5253 23489 5287
rect 23523 5284 23535 5287
rect 23566 5284 23572 5296
rect 23523 5256 23572 5284
rect 23523 5253 23535 5256
rect 23477 5247 23535 5253
rect 23566 5244 23572 5256
rect 23624 5244 23630 5296
rect 23842 5244 23848 5296
rect 23900 5284 23906 5296
rect 24118 5284 24124 5296
rect 23900 5256 24124 5284
rect 23900 5244 23906 5256
rect 24118 5244 24124 5256
rect 24176 5244 24182 5296
rect 16117 5219 16175 5225
rect 16117 5185 16129 5219
rect 16163 5185 16175 5219
rect 21821 5219 21879 5225
rect 21821 5216 21833 5219
rect 16117 5179 16175 5185
rect 21100 5188 21833 5216
rect 12176 5120 12848 5148
rect 9490 5080 9496 5092
rect 9451 5052 9496 5080
rect 9490 5040 9496 5052
rect 9548 5040 9554 5092
rect 10597 5083 10655 5089
rect 10597 5049 10609 5083
rect 10643 5080 10655 5083
rect 11149 5083 11207 5089
rect 11149 5080 11161 5083
rect 10643 5052 11161 5080
rect 10643 5049 10655 5052
rect 10597 5043 10655 5049
rect 11149 5049 11161 5052
rect 11195 5080 11207 5083
rect 11606 5080 11612 5092
rect 11195 5052 11612 5080
rect 11195 5049 11207 5052
rect 11149 5043 11207 5049
rect 11606 5040 11612 5052
rect 11664 5040 11670 5092
rect 11882 5040 11888 5092
rect 11940 5080 11946 5092
rect 12820 5080 12848 5120
rect 13814 5108 13820 5160
rect 13872 5148 13878 5160
rect 14369 5151 14427 5157
rect 14369 5148 14381 5151
rect 13872 5120 14381 5148
rect 13872 5108 13878 5120
rect 14369 5117 14381 5120
rect 14415 5117 14427 5151
rect 14369 5111 14427 5117
rect 15378 5108 15384 5160
rect 15436 5148 15442 5160
rect 15838 5148 15844 5160
rect 15436 5120 15844 5148
rect 15436 5108 15442 5120
rect 15838 5108 15844 5120
rect 15896 5148 15902 5160
rect 15933 5151 15991 5157
rect 15933 5148 15945 5151
rect 15896 5120 15945 5148
rect 15896 5108 15902 5120
rect 15933 5117 15945 5120
rect 15979 5117 15991 5151
rect 15933 5111 15991 5117
rect 18690 5108 18696 5160
rect 18748 5148 18754 5160
rect 18785 5151 18843 5157
rect 18785 5148 18797 5151
rect 18748 5120 18797 5148
rect 18748 5108 18754 5120
rect 18785 5117 18797 5120
rect 18831 5117 18843 5151
rect 18785 5111 18843 5117
rect 12986 5080 12992 5092
rect 11940 5052 12664 5080
rect 12820 5052 12992 5080
rect 11940 5040 11946 5052
rect 8941 5015 8999 5021
rect 8941 5012 8953 5015
rect 8904 4984 8953 5012
rect 8904 4972 8910 4984
rect 8941 4981 8953 4984
rect 8987 4981 8999 5015
rect 9122 5012 9128 5024
rect 9083 4984 9128 5012
rect 8941 4975 8999 4981
rect 9122 4972 9128 4984
rect 9180 4972 9186 5024
rect 10778 4972 10784 5024
rect 10836 5012 10842 5024
rect 11054 5012 11060 5024
rect 10836 4984 11060 5012
rect 10836 4972 10842 4984
rect 11054 4972 11060 4984
rect 11112 4972 11118 5024
rect 11514 4972 11520 5024
rect 11572 5012 11578 5024
rect 12342 5012 12348 5024
rect 11572 4984 12348 5012
rect 11572 4972 11578 4984
rect 12342 4972 12348 4984
rect 12400 4972 12406 5024
rect 12434 4972 12440 5024
rect 12492 5012 12498 5024
rect 12636 5012 12664 5052
rect 12986 5040 12992 5052
rect 13044 5080 13050 5092
rect 13446 5080 13452 5092
rect 13044 5052 13452 5080
rect 13044 5040 13050 5052
rect 13446 5040 13452 5052
rect 13504 5040 13510 5092
rect 14274 5040 14280 5092
rect 14332 5080 14338 5092
rect 14642 5080 14648 5092
rect 14332 5052 14648 5080
rect 14332 5040 14338 5052
rect 14642 5040 14648 5052
rect 14700 5040 14706 5092
rect 17865 5083 17923 5089
rect 17865 5049 17877 5083
rect 17911 5080 17923 5083
rect 18322 5080 18328 5092
rect 17911 5052 18328 5080
rect 17911 5049 17923 5052
rect 17865 5043 17923 5049
rect 18322 5040 18328 5052
rect 18380 5040 18386 5092
rect 19052 5083 19110 5089
rect 19052 5049 19064 5083
rect 19098 5080 19110 5083
rect 19242 5080 19248 5092
rect 19098 5052 19248 5080
rect 19098 5049 19110 5052
rect 19052 5043 19110 5049
rect 19242 5040 19248 5052
rect 19300 5080 19306 5092
rect 19426 5080 19432 5092
rect 19300 5052 19432 5080
rect 19300 5040 19306 5052
rect 19426 5040 19432 5052
rect 19484 5040 19490 5092
rect 21100 5089 21128 5188
rect 21821 5185 21833 5188
rect 21867 5185 21879 5219
rect 21821 5179 21879 5185
rect 21637 5151 21695 5157
rect 21637 5117 21649 5151
rect 21683 5148 21695 5151
rect 21726 5148 21732 5160
rect 21683 5120 21732 5148
rect 21683 5117 21695 5120
rect 21637 5111 21695 5117
rect 21726 5108 21732 5120
rect 21784 5108 21790 5160
rect 23584 5148 23612 5244
rect 23750 5176 23756 5228
rect 23808 5216 23814 5228
rect 24213 5219 24271 5225
rect 24213 5216 24225 5219
rect 23808 5188 24225 5216
rect 23808 5176 23814 5188
rect 24213 5185 24225 5188
rect 24259 5185 24271 5219
rect 25498 5216 25504 5228
rect 25459 5188 25504 5216
rect 24213 5179 24271 5185
rect 25498 5176 25504 5188
rect 25556 5176 25562 5228
rect 23658 5148 23664 5160
rect 23571 5120 23664 5148
rect 23658 5108 23664 5120
rect 23716 5148 23722 5160
rect 24121 5151 24179 5157
rect 24121 5148 24133 5151
rect 23716 5120 24133 5148
rect 23716 5108 23722 5120
rect 24121 5117 24133 5120
rect 24167 5117 24179 5151
rect 25222 5148 25228 5160
rect 25183 5120 25228 5148
rect 24121 5111 24179 5117
rect 25222 5108 25228 5120
rect 25280 5148 25286 5160
rect 25961 5151 26019 5157
rect 25961 5148 25973 5151
rect 25280 5120 25973 5148
rect 25280 5108 25286 5120
rect 25961 5117 25973 5120
rect 26007 5117 26019 5151
rect 25961 5111 26019 5117
rect 21085 5083 21143 5089
rect 21085 5080 21097 5083
rect 20180 5052 21097 5080
rect 20180 5024 20208 5052
rect 21085 5049 21097 5052
rect 21131 5049 21143 5083
rect 21085 5043 21143 5049
rect 21818 5040 21824 5092
rect 21876 5080 21882 5092
rect 22649 5083 22707 5089
rect 22649 5080 22661 5083
rect 21876 5052 22661 5080
rect 21876 5040 21882 5052
rect 22649 5049 22661 5052
rect 22695 5049 22707 5083
rect 24026 5080 24032 5092
rect 23987 5052 24032 5080
rect 22649 5043 22707 5049
rect 24026 5040 24032 5052
rect 24084 5040 24090 5092
rect 12805 5015 12863 5021
rect 12805 5012 12817 5015
rect 12492 4984 12537 5012
rect 12636 4984 12817 5012
rect 12492 4972 12498 4984
rect 12805 4981 12817 4984
rect 12851 4981 12863 5015
rect 12805 4975 12863 4981
rect 12897 5015 12955 5021
rect 12897 4981 12909 5015
rect 12943 5012 12955 5015
rect 13265 5015 13323 5021
rect 13265 5012 13277 5015
rect 12943 4984 13277 5012
rect 12943 4981 12955 4984
rect 12897 4975 12955 4981
rect 13265 4981 13277 4984
rect 13311 4981 13323 5015
rect 20162 5012 20168 5024
rect 20123 4984 20168 5012
rect 13265 4975 13323 4981
rect 20162 4972 20168 4984
rect 20220 4972 20226 5024
rect 20714 5012 20720 5024
rect 20675 4984 20720 5012
rect 20714 4972 20720 4984
rect 20772 4972 20778 5024
rect 21450 4972 21456 5024
rect 21508 5012 21514 5024
rect 21729 5015 21787 5021
rect 21729 5012 21741 5015
rect 21508 4984 21741 5012
rect 21508 4972 21514 4984
rect 21729 4981 21741 4984
rect 21775 4981 21787 5015
rect 21729 4975 21787 4981
rect 24854 4972 24860 5024
rect 24912 5012 24918 5024
rect 25041 5015 25099 5021
rect 25041 5012 25053 5015
rect 24912 4984 25053 5012
rect 24912 4972 24918 4984
rect 25041 4981 25053 4984
rect 25087 4981 25099 5015
rect 25041 4975 25099 4981
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1489 4811 1547 4817
rect 1489 4777 1501 4811
rect 1535 4808 1547 4811
rect 1762 4808 1768 4820
rect 1535 4780 1768 4808
rect 1535 4777 1547 4780
rect 1489 4771 1547 4777
rect 1762 4768 1768 4780
rect 1820 4768 1826 4820
rect 1946 4808 1952 4820
rect 1907 4780 1952 4808
rect 1946 4768 1952 4780
rect 2004 4768 2010 4820
rect 2498 4808 2504 4820
rect 2459 4780 2504 4808
rect 2498 4768 2504 4780
rect 2556 4768 2562 4820
rect 3234 4768 3240 4820
rect 3292 4808 3298 4820
rect 4065 4811 4123 4817
rect 4065 4808 4077 4811
rect 3292 4780 4077 4808
rect 3292 4768 3298 4780
rect 4065 4777 4077 4780
rect 4111 4777 4123 4811
rect 4430 4808 4436 4820
rect 4391 4780 4436 4808
rect 4065 4771 4123 4777
rect 4430 4768 4436 4780
rect 4488 4768 4494 4820
rect 5534 4808 5540 4820
rect 5495 4780 5540 4808
rect 5534 4768 5540 4780
rect 5592 4768 5598 4820
rect 5721 4811 5779 4817
rect 5721 4777 5733 4811
rect 5767 4808 5779 4811
rect 7006 4808 7012 4820
rect 5767 4780 7012 4808
rect 5767 4777 5779 4780
rect 5721 4771 5779 4777
rect 7006 4768 7012 4780
rect 7064 4768 7070 4820
rect 7282 4808 7288 4820
rect 7243 4780 7288 4808
rect 7282 4768 7288 4780
rect 7340 4768 7346 4820
rect 7745 4811 7803 4817
rect 7745 4777 7757 4811
rect 7791 4808 7803 4811
rect 9122 4808 9128 4820
rect 7791 4780 9128 4808
rect 7791 4777 7803 4780
rect 7745 4771 7803 4777
rect 1857 4743 1915 4749
rect 1857 4709 1869 4743
rect 1903 4740 1915 4743
rect 2590 4740 2596 4752
rect 1903 4712 2596 4740
rect 1903 4709 1915 4712
rect 1857 4703 1915 4709
rect 2590 4700 2596 4712
rect 2648 4700 2654 4752
rect 2774 4700 2780 4752
rect 2832 4740 2838 4752
rect 3053 4743 3111 4749
rect 3053 4740 3065 4743
rect 2832 4712 3065 4740
rect 2832 4700 2838 4712
rect 3053 4709 3065 4712
rect 3099 4740 3111 4743
rect 3326 4740 3332 4752
rect 3099 4712 3332 4740
rect 3099 4709 3111 4712
rect 3053 4703 3111 4709
rect 3326 4700 3332 4712
rect 3384 4700 3390 4752
rect 5261 4743 5319 4749
rect 5261 4709 5273 4743
rect 5307 4740 5319 4743
rect 5810 4740 5816 4752
rect 5307 4712 5816 4740
rect 5307 4709 5319 4712
rect 5261 4703 5319 4709
rect 5810 4700 5816 4712
rect 5868 4700 5874 4752
rect 5994 4700 6000 4752
rect 6052 4740 6058 4752
rect 6181 4743 6239 4749
rect 6181 4740 6193 4743
rect 6052 4712 6193 4740
rect 6052 4700 6058 4712
rect 6181 4709 6193 4712
rect 6227 4709 6239 4743
rect 6181 4703 6239 4709
rect 6825 4743 6883 4749
rect 6825 4709 6837 4743
rect 6871 4740 6883 4743
rect 7760 4740 7788 4771
rect 9122 4768 9128 4780
rect 9180 4768 9186 4820
rect 9217 4811 9275 4817
rect 9217 4777 9229 4811
rect 9263 4808 9275 4811
rect 9490 4808 9496 4820
rect 9263 4780 9496 4808
rect 9263 4777 9275 4780
rect 9217 4771 9275 4777
rect 8386 4740 8392 4752
rect 6871 4712 7788 4740
rect 8347 4712 8392 4740
rect 6871 4709 6883 4712
rect 6825 4703 6883 4709
rect 8386 4700 8392 4712
rect 8444 4700 8450 4752
rect 8478 4700 8484 4752
rect 8536 4740 8542 4752
rect 9232 4740 9260 4771
rect 9490 4768 9496 4780
rect 9548 4768 9554 4820
rect 9677 4811 9735 4817
rect 9677 4777 9689 4811
rect 9723 4808 9735 4811
rect 9766 4808 9772 4820
rect 9723 4780 9772 4808
rect 9723 4777 9735 4780
rect 9677 4771 9735 4777
rect 9766 4768 9772 4780
rect 9824 4768 9830 4820
rect 10137 4811 10195 4817
rect 10137 4777 10149 4811
rect 10183 4808 10195 4811
rect 10686 4808 10692 4820
rect 10183 4780 10692 4808
rect 10183 4777 10195 4780
rect 10137 4771 10195 4777
rect 10686 4768 10692 4780
rect 10744 4768 10750 4820
rect 12342 4808 12348 4820
rect 12303 4780 12348 4808
rect 12342 4768 12348 4780
rect 12400 4768 12406 4820
rect 12710 4768 12716 4820
rect 12768 4808 12774 4820
rect 13265 4811 13323 4817
rect 13265 4808 13277 4811
rect 12768 4780 13277 4808
rect 12768 4768 12774 4780
rect 13265 4777 13277 4780
rect 13311 4777 13323 4811
rect 13265 4771 13323 4777
rect 13449 4811 13507 4817
rect 13449 4777 13461 4811
rect 13495 4808 13507 4811
rect 13630 4808 13636 4820
rect 13495 4780 13636 4808
rect 13495 4777 13507 4780
rect 13449 4771 13507 4777
rect 8536 4712 9260 4740
rect 10045 4743 10103 4749
rect 8536 4700 8542 4712
rect 10045 4709 10057 4743
rect 10091 4740 10103 4743
rect 10962 4740 10968 4752
rect 10091 4712 10968 4740
rect 10091 4709 10103 4712
rect 10045 4703 10103 4709
rect 10962 4700 10968 4712
rect 11020 4700 11026 4752
rect 11238 4700 11244 4752
rect 11296 4740 11302 4752
rect 12894 4740 12900 4752
rect 11296 4712 12900 4740
rect 11296 4700 11302 4712
rect 12894 4700 12900 4712
rect 12952 4700 12958 4752
rect 3421 4675 3479 4681
rect 3421 4641 3433 4675
rect 3467 4672 3479 4675
rect 3881 4675 3939 4681
rect 3881 4672 3893 4675
rect 3467 4644 3893 4672
rect 3467 4641 3479 4644
rect 3421 4635 3479 4641
rect 3881 4641 3893 4644
rect 3927 4672 3939 4675
rect 4062 4672 4068 4684
rect 3927 4644 4068 4672
rect 3927 4641 3939 4644
rect 3881 4635 3939 4641
rect 4062 4632 4068 4644
rect 4120 4632 4126 4684
rect 6089 4675 6147 4681
rect 6089 4641 6101 4675
rect 6135 4672 6147 4675
rect 6362 4672 6368 4684
rect 6135 4644 6368 4672
rect 6135 4641 6147 4644
rect 6089 4635 6147 4641
rect 6362 4632 6368 4644
rect 6420 4632 6426 4684
rect 7006 4632 7012 4684
rect 7064 4672 7070 4684
rect 7653 4675 7711 4681
rect 7653 4672 7665 4675
rect 7064 4644 7665 4672
rect 7064 4632 7070 4644
rect 7653 4641 7665 4644
rect 7699 4641 7711 4675
rect 11330 4672 11336 4684
rect 11291 4644 11336 4672
rect 7653 4635 7711 4641
rect 11330 4632 11336 4644
rect 11388 4632 11394 4684
rect 12253 4675 12311 4681
rect 12253 4672 12265 4675
rect 11900 4644 12265 4672
rect 2133 4607 2191 4613
rect 2133 4573 2145 4607
rect 2179 4604 2191 4607
rect 2498 4604 2504 4616
rect 2179 4576 2504 4604
rect 2179 4573 2191 4576
rect 2133 4567 2191 4573
rect 2498 4564 2504 4576
rect 2556 4564 2562 4616
rect 4522 4604 4528 4616
rect 4483 4576 4528 4604
rect 4522 4564 4528 4576
rect 4580 4564 4586 4616
rect 4706 4564 4712 4616
rect 4764 4604 4770 4616
rect 5442 4604 5448 4616
rect 4764 4576 5448 4604
rect 4764 4564 4770 4576
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 6270 4604 6276 4616
rect 6231 4576 6276 4604
rect 6270 4564 6276 4576
rect 6328 4564 6334 4616
rect 7193 4607 7251 4613
rect 7193 4573 7205 4607
rect 7239 4604 7251 4607
rect 7929 4607 7987 4613
rect 7929 4604 7941 4607
rect 7239 4576 7941 4604
rect 7239 4573 7251 4576
rect 7193 4567 7251 4573
rect 7929 4573 7941 4576
rect 7975 4604 7987 4607
rect 8202 4604 8208 4616
rect 7975 4576 8208 4604
rect 7975 4573 7987 4576
rect 7929 4567 7987 4573
rect 8202 4564 8208 4576
rect 8260 4564 8266 4616
rect 8849 4607 8907 4613
rect 8849 4573 8861 4607
rect 8895 4604 8907 4607
rect 9398 4604 9404 4616
rect 8895 4576 9404 4604
rect 8895 4573 8907 4576
rect 8849 4567 8907 4573
rect 9398 4564 9404 4576
rect 9456 4604 9462 4616
rect 10229 4607 10287 4613
rect 10229 4604 10241 4607
rect 9456 4576 10241 4604
rect 9456 4564 9462 4576
rect 10229 4573 10241 4576
rect 10275 4573 10287 4607
rect 10229 4567 10287 4573
rect 11146 4564 11152 4616
rect 11204 4604 11210 4616
rect 11900 4604 11928 4644
rect 12253 4641 12265 4644
rect 12299 4641 12311 4675
rect 12253 4635 12311 4641
rect 11204 4576 11928 4604
rect 11204 4564 11210 4576
rect 12158 4564 12164 4616
rect 12216 4604 12222 4616
rect 12437 4607 12495 4613
rect 12437 4604 12449 4607
rect 12216 4576 12449 4604
rect 12216 4564 12222 4576
rect 12437 4573 12449 4576
rect 12483 4573 12495 4607
rect 13280 4604 13308 4771
rect 13630 4768 13636 4780
rect 13688 4768 13694 4820
rect 13909 4811 13967 4817
rect 13909 4777 13921 4811
rect 13955 4808 13967 4811
rect 13998 4808 14004 4820
rect 13955 4780 14004 4808
rect 13955 4777 13967 4780
rect 13909 4771 13967 4777
rect 13998 4768 14004 4780
rect 14056 4768 14062 4820
rect 15105 4811 15163 4817
rect 15105 4777 15117 4811
rect 15151 4808 15163 4811
rect 16022 4808 16028 4820
rect 15151 4780 16028 4808
rect 15151 4777 15163 4780
rect 15105 4771 15163 4777
rect 16022 4768 16028 4780
rect 16080 4768 16086 4820
rect 19426 4808 19432 4820
rect 19339 4780 19432 4808
rect 19426 4768 19432 4780
rect 19484 4808 19490 4820
rect 20254 4808 20260 4820
rect 19484 4780 20260 4808
rect 19484 4768 19490 4780
rect 20254 4768 20260 4780
rect 20312 4808 20318 4820
rect 20625 4811 20683 4817
rect 20625 4808 20637 4811
rect 20312 4780 20637 4808
rect 20312 4768 20318 4780
rect 20625 4777 20637 4780
rect 20671 4777 20683 4811
rect 20625 4771 20683 4777
rect 20901 4811 20959 4817
rect 20901 4777 20913 4811
rect 20947 4808 20959 4811
rect 21726 4808 21732 4820
rect 20947 4780 21732 4808
rect 20947 4777 20959 4780
rect 20901 4771 20959 4777
rect 15286 4700 15292 4752
rect 15344 4740 15350 4752
rect 18690 4740 18696 4752
rect 15344 4712 18696 4740
rect 15344 4700 15350 4712
rect 13814 4672 13820 4684
rect 13775 4644 13820 4672
rect 13814 4632 13820 4644
rect 13872 4632 13878 4684
rect 15556 4675 15614 4681
rect 15556 4641 15568 4675
rect 15602 4672 15614 4675
rect 16482 4672 16488 4684
rect 15602 4644 16488 4672
rect 15602 4641 15614 4644
rect 15556 4635 15614 4641
rect 16482 4632 16488 4644
rect 16540 4632 16546 4684
rect 18064 4681 18092 4712
rect 18690 4700 18696 4712
rect 18748 4700 18754 4752
rect 20640 4740 20668 4771
rect 21726 4768 21732 4780
rect 21784 4768 21790 4820
rect 22278 4768 22284 4820
rect 22336 4808 22342 4820
rect 22336 4780 23336 4808
rect 22336 4768 22342 4780
rect 20640 4712 21496 4740
rect 18322 4681 18328 4684
rect 18049 4675 18107 4681
rect 18049 4641 18061 4675
rect 18095 4641 18107 4675
rect 18316 4672 18328 4681
rect 18283 4644 18328 4672
rect 18049 4635 18107 4641
rect 18316 4635 18328 4644
rect 18322 4632 18328 4635
rect 18380 4632 18386 4684
rect 21266 4672 21272 4684
rect 21227 4644 21272 4672
rect 21266 4632 21272 4644
rect 21324 4632 21330 4684
rect 21468 4616 21496 4712
rect 22554 4700 22560 4752
rect 22612 4740 22618 4752
rect 22833 4743 22891 4749
rect 22833 4740 22845 4743
rect 22612 4712 22845 4740
rect 22612 4700 22618 4712
rect 22833 4709 22845 4712
rect 22879 4709 22891 4743
rect 23308 4740 23336 4780
rect 23382 4768 23388 4820
rect 23440 4808 23446 4820
rect 23753 4811 23811 4817
rect 23753 4808 23765 4811
rect 23440 4780 23765 4808
rect 23440 4768 23446 4780
rect 23753 4777 23765 4780
rect 23799 4808 23811 4811
rect 24118 4808 24124 4820
rect 23799 4780 24124 4808
rect 23799 4777 23811 4780
rect 23753 4771 23811 4777
rect 24118 4768 24124 4780
rect 24176 4768 24182 4820
rect 24489 4811 24547 4817
rect 24489 4777 24501 4811
rect 24535 4808 24547 4811
rect 24854 4808 24860 4820
rect 24535 4780 24860 4808
rect 24535 4777 24547 4780
rect 24489 4771 24547 4777
rect 24854 4768 24860 4780
rect 24912 4808 24918 4820
rect 25590 4808 25596 4820
rect 24912 4780 25596 4808
rect 24912 4768 24918 4780
rect 25590 4768 25596 4780
rect 25648 4768 25654 4820
rect 26234 4768 26240 4820
rect 26292 4808 26298 4820
rect 26292 4780 26337 4808
rect 26292 4768 26298 4780
rect 25409 4743 25467 4749
rect 25409 4740 25421 4743
rect 23308 4712 25421 4740
rect 22833 4703 22891 4709
rect 25409 4709 25421 4712
rect 25455 4740 25467 4743
rect 26326 4740 26332 4752
rect 25455 4712 26332 4740
rect 25455 4709 25467 4712
rect 25409 4703 25467 4709
rect 26326 4700 26332 4712
rect 26384 4700 26390 4752
rect 23934 4632 23940 4684
rect 23992 4672 23998 4684
rect 24397 4675 24455 4681
rect 24397 4672 24409 4675
rect 23992 4644 24409 4672
rect 23992 4632 23998 4644
rect 24397 4641 24409 4644
rect 24443 4641 24455 4675
rect 24397 4635 24455 4641
rect 25038 4632 25044 4684
rect 25096 4672 25102 4684
rect 25774 4672 25780 4684
rect 25096 4644 25780 4672
rect 25096 4632 25102 4644
rect 25774 4632 25780 4644
rect 25832 4632 25838 4684
rect 14001 4607 14059 4613
rect 14001 4604 14013 4607
rect 13280 4576 14013 4604
rect 12437 4567 12495 4573
rect 14001 4573 14013 4576
rect 14047 4573 14059 4607
rect 15286 4604 15292 4616
rect 15247 4576 15292 4604
rect 14001 4567 14059 4573
rect 15286 4564 15292 4576
rect 15344 4564 15350 4616
rect 17589 4607 17647 4613
rect 17589 4573 17601 4607
rect 17635 4604 17647 4607
rect 17954 4604 17960 4616
rect 17635 4576 17960 4604
rect 17635 4573 17647 4576
rect 17589 4567 17647 4573
rect 17954 4564 17960 4576
rect 18012 4564 18018 4616
rect 21361 4607 21419 4613
rect 21361 4573 21373 4607
rect 21407 4573 21419 4607
rect 21361 4567 21419 4573
rect 3326 4496 3332 4548
rect 3384 4536 3390 4548
rect 8570 4536 8576 4548
rect 3384 4508 8576 4536
rect 3384 4496 3390 4508
rect 8570 4496 8576 4508
rect 8628 4496 8634 4548
rect 9858 4496 9864 4548
rect 9916 4536 9922 4548
rect 10134 4536 10140 4548
rect 9916 4508 10140 4536
rect 9916 4496 9922 4508
rect 10134 4496 10140 4508
rect 10192 4496 10198 4548
rect 10778 4536 10784 4548
rect 10739 4508 10784 4536
rect 10778 4496 10784 4508
rect 10836 4496 10842 4548
rect 11793 4539 11851 4545
rect 11793 4505 11805 4539
rect 11839 4536 11851 4539
rect 12250 4536 12256 4548
rect 11839 4508 12256 4536
rect 11839 4505 11851 4508
rect 11793 4499 11851 4505
rect 12250 4496 12256 4508
rect 12308 4496 12314 4548
rect 17862 4496 17868 4548
rect 17920 4536 17926 4548
rect 20990 4536 20996 4548
rect 17920 4508 18092 4536
rect 17920 4496 17926 4508
rect 198 4428 204 4480
rect 256 4468 262 4480
rect 8846 4468 8852 4480
rect 256 4440 8852 4468
rect 256 4428 262 4440
rect 8846 4428 8852 4440
rect 8904 4428 8910 4480
rect 11882 4468 11888 4480
rect 11843 4440 11888 4468
rect 11882 4428 11888 4440
rect 11940 4428 11946 4480
rect 13906 4428 13912 4480
rect 13964 4468 13970 4480
rect 14553 4471 14611 4477
rect 14553 4468 14565 4471
rect 13964 4440 14565 4468
rect 13964 4428 13970 4440
rect 14553 4437 14565 4440
rect 14599 4468 14611 4471
rect 14826 4468 14832 4480
rect 14599 4440 14832 4468
rect 14599 4437 14611 4440
rect 14553 4431 14611 4437
rect 14826 4428 14832 4440
rect 14884 4428 14890 4480
rect 16669 4471 16727 4477
rect 16669 4437 16681 4471
rect 16715 4468 16727 4471
rect 16850 4468 16856 4480
rect 16715 4440 16856 4468
rect 16715 4437 16727 4440
rect 16669 4431 16727 4437
rect 16850 4428 16856 4440
rect 16908 4428 16914 4480
rect 17954 4468 17960 4480
rect 17915 4440 17960 4468
rect 17954 4428 17960 4440
rect 18012 4428 18018 4480
rect 18064 4468 18092 4508
rect 18984 4508 20996 4536
rect 18984 4468 19012 4508
rect 20990 4496 20996 4508
rect 21048 4496 21054 4548
rect 21376 4536 21404 4567
rect 21450 4564 21456 4616
rect 21508 4604 21514 4616
rect 22922 4604 22928 4616
rect 21508 4576 21601 4604
rect 22883 4576 22928 4604
rect 21508 4564 21514 4576
rect 22922 4564 22928 4576
rect 22980 4564 22986 4616
rect 23109 4607 23167 4613
rect 23109 4573 23121 4607
rect 23155 4573 23167 4607
rect 23109 4567 23167 4573
rect 21634 4536 21640 4548
rect 21376 4508 21640 4536
rect 21634 4496 21640 4508
rect 21692 4496 21698 4548
rect 21726 4496 21732 4548
rect 21784 4536 21790 4548
rect 21913 4539 21971 4545
rect 21913 4536 21925 4539
rect 21784 4508 21925 4536
rect 21784 4496 21790 4508
rect 21913 4505 21925 4508
rect 21959 4536 21971 4539
rect 23124 4536 23152 4567
rect 24118 4564 24124 4616
rect 24176 4604 24182 4616
rect 24581 4607 24639 4613
rect 24581 4604 24593 4607
rect 24176 4576 24593 4604
rect 24176 4564 24182 4576
rect 24581 4573 24593 4576
rect 24627 4573 24639 4607
rect 24581 4567 24639 4573
rect 21959 4508 23152 4536
rect 21959 4505 21971 4508
rect 21913 4499 21971 4505
rect 23566 4496 23572 4548
rect 23624 4536 23630 4548
rect 24029 4539 24087 4545
rect 24029 4536 24041 4539
rect 23624 4508 24041 4536
rect 23624 4496 23630 4508
rect 24029 4505 24041 4508
rect 24075 4505 24087 4539
rect 24029 4499 24087 4505
rect 19978 4468 19984 4480
rect 18064 4440 19012 4468
rect 19939 4440 19984 4468
rect 19978 4428 19984 4440
rect 20036 4428 20042 4480
rect 22094 4428 22100 4480
rect 22152 4468 22158 4480
rect 22373 4471 22431 4477
rect 22373 4468 22385 4471
rect 22152 4440 22385 4468
rect 22152 4428 22158 4440
rect 22373 4437 22385 4440
rect 22419 4468 22431 4471
rect 22465 4471 22523 4477
rect 22465 4468 22477 4471
rect 22419 4440 22477 4468
rect 22419 4437 22431 4440
rect 22373 4431 22431 4437
rect 22465 4437 22477 4440
rect 22511 4437 22523 4471
rect 22465 4431 22523 4437
rect 24670 4428 24676 4480
rect 24728 4468 24734 4480
rect 25038 4468 25044 4480
rect 24728 4440 25044 4468
rect 24728 4428 24734 4440
rect 25038 4428 25044 4440
rect 25096 4428 25102 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 2406 4224 2412 4276
rect 2464 4264 2470 4276
rect 2501 4267 2559 4273
rect 2501 4264 2513 4267
rect 2464 4236 2513 4264
rect 2464 4224 2470 4236
rect 2501 4233 2513 4236
rect 2547 4264 2559 4267
rect 2590 4264 2596 4276
rect 2547 4236 2596 4264
rect 2547 4233 2559 4236
rect 2501 4227 2559 4233
rect 2590 4224 2596 4236
rect 2648 4224 2654 4276
rect 5905 4267 5963 4273
rect 5905 4264 5917 4267
rect 3988 4236 5917 4264
rect 1210 4156 1216 4208
rect 1268 4196 1274 4208
rect 3988 4196 4016 4236
rect 5905 4233 5917 4236
rect 5951 4264 5963 4267
rect 5994 4264 6000 4276
rect 5951 4236 6000 4264
rect 5951 4233 5963 4236
rect 5905 4227 5963 4233
rect 5994 4224 6000 4236
rect 6052 4224 6058 4276
rect 9674 4264 9680 4276
rect 9635 4236 9680 4264
rect 9674 4224 9680 4236
rect 9732 4224 9738 4276
rect 11885 4267 11943 4273
rect 11885 4233 11897 4267
rect 11931 4264 11943 4267
rect 12158 4264 12164 4276
rect 11931 4236 12164 4264
rect 11931 4233 11943 4236
rect 11885 4227 11943 4233
rect 12158 4224 12164 4236
rect 12216 4224 12222 4276
rect 13909 4267 13967 4273
rect 12268 4236 13124 4264
rect 1268 4168 4016 4196
rect 1268 4156 1274 4168
rect 9214 4156 9220 4208
rect 9272 4196 9278 4208
rect 10781 4199 10839 4205
rect 9272 4168 10272 4196
rect 9272 4156 9278 4168
rect 2041 4131 2099 4137
rect 2041 4097 2053 4131
rect 2087 4128 2099 4131
rect 2130 4128 2136 4140
rect 2087 4100 2136 4128
rect 2087 4097 2099 4100
rect 2041 4091 2099 4097
rect 2130 4088 2136 4100
rect 2188 4088 2194 4140
rect 3970 4128 3976 4140
rect 3931 4100 3976 4128
rect 3970 4088 3976 4100
rect 4028 4088 4034 4140
rect 6270 4088 6276 4140
rect 6328 4128 6334 4140
rect 10244 4137 10272 4168
rect 10781 4165 10793 4199
rect 10827 4196 10839 4199
rect 10962 4196 10968 4208
rect 10827 4168 10968 4196
rect 10827 4165 10839 4168
rect 10781 4159 10839 4165
rect 10962 4156 10968 4168
rect 11020 4156 11026 4208
rect 12268 4196 12296 4236
rect 11072 4168 12296 4196
rect 7009 4131 7067 4137
rect 7009 4128 7021 4131
rect 6328 4100 7021 4128
rect 6328 4088 6334 4100
rect 7009 4097 7021 4100
rect 7055 4128 7067 4131
rect 10229 4131 10287 4137
rect 7055 4100 7328 4128
rect 7055 4097 7067 4100
rect 7009 4091 7067 4097
rect 3881 4063 3939 4069
rect 3881 4029 3893 4063
rect 3927 4060 3939 4063
rect 4706 4060 4712 4072
rect 3927 4032 4712 4060
rect 3927 4029 3939 4032
rect 3881 4023 3939 4029
rect 4706 4020 4712 4032
rect 4764 4020 4770 4072
rect 7193 4063 7251 4069
rect 7193 4029 7205 4063
rect 7239 4029 7251 4063
rect 7300 4060 7328 4100
rect 10229 4097 10241 4131
rect 10275 4097 10287 4131
rect 10229 4091 10287 4097
rect 7466 4069 7472 4072
rect 7449 4063 7472 4069
rect 7449 4060 7461 4063
rect 7300 4032 7461 4060
rect 7193 4023 7251 4029
rect 7449 4029 7461 4032
rect 7524 4060 7530 4072
rect 7524 4032 7597 4060
rect 7449 4023 7472 4029
rect 1854 3992 1860 4004
rect 1767 3964 1860 3992
rect 1854 3952 1860 3964
rect 1912 3992 1918 4004
rect 2866 3992 2872 4004
rect 1912 3964 2872 3992
rect 1912 3952 1918 3964
rect 2866 3952 2872 3964
rect 2924 3952 2930 4004
rect 3513 3995 3571 4001
rect 3513 3961 3525 3995
rect 3559 3992 3571 3995
rect 4218 3995 4276 4001
rect 4218 3992 4230 3995
rect 3559 3964 4230 3992
rect 3559 3961 3571 3964
rect 3513 3955 3571 3961
rect 4218 3961 4230 3964
rect 4264 3992 4276 3995
rect 6086 3992 6092 4004
rect 4264 3964 6092 3992
rect 4264 3961 4276 3964
rect 4218 3955 4276 3961
rect 6086 3952 6092 3964
rect 6144 3952 6150 4004
rect 7006 3952 7012 4004
rect 7064 3992 7070 4004
rect 7208 3992 7236 4023
rect 7466 4020 7472 4023
rect 7524 4020 7530 4032
rect 9950 4020 9956 4072
rect 10008 4060 10014 4072
rect 10045 4063 10103 4069
rect 10045 4060 10057 4063
rect 10008 4032 10057 4060
rect 10008 4020 10014 4032
rect 10045 4029 10057 4032
rect 10091 4060 10103 4063
rect 11072 4060 11100 4168
rect 12894 4156 12900 4208
rect 12952 4196 12958 4208
rect 13096 4196 13124 4236
rect 13909 4233 13921 4267
rect 13955 4264 13967 4267
rect 13998 4264 14004 4276
rect 13955 4236 14004 4264
rect 13955 4233 13967 4236
rect 13909 4227 13967 4233
rect 13998 4224 14004 4236
rect 14056 4224 14062 4276
rect 15565 4267 15623 4273
rect 15565 4233 15577 4267
rect 15611 4233 15623 4267
rect 15565 4227 15623 4233
rect 14458 4196 14464 4208
rect 12952 4168 13032 4196
rect 13096 4168 14464 4196
rect 12952 4156 12958 4168
rect 11149 4131 11207 4137
rect 11149 4097 11161 4131
rect 11195 4128 11207 4131
rect 11422 4128 11428 4140
rect 11195 4100 11428 4128
rect 11195 4097 11207 4100
rect 11149 4091 11207 4097
rect 11422 4088 11428 4100
rect 11480 4088 11486 4140
rect 12618 4128 12624 4140
rect 11532 4100 12624 4128
rect 10091 4032 11100 4060
rect 11241 4063 11299 4069
rect 10091 4029 10103 4032
rect 10045 4023 10103 4029
rect 11241 4029 11253 4063
rect 11287 4060 11299 4063
rect 11330 4060 11336 4072
rect 11287 4032 11336 4060
rect 11287 4029 11299 4032
rect 11241 4023 11299 4029
rect 11330 4020 11336 4032
rect 11388 4020 11394 4072
rect 8110 3992 8116 4004
rect 7064 3964 8116 3992
rect 7064 3952 7070 3964
rect 8110 3952 8116 3964
rect 8168 3952 8174 4004
rect 8386 3952 8392 4004
rect 8444 3992 8450 4004
rect 9493 3995 9551 4001
rect 9493 3992 9505 3995
rect 8444 3964 9505 3992
rect 8444 3952 8450 3964
rect 9493 3961 9505 3964
rect 9539 3992 9551 3995
rect 10137 3995 10195 4001
rect 10137 3992 10149 3995
rect 9539 3964 10149 3992
rect 9539 3961 9551 3964
rect 9493 3955 9551 3961
rect 10137 3961 10149 3964
rect 10183 3992 10195 3995
rect 11532 3992 11560 4100
rect 12618 4088 12624 4100
rect 12676 4088 12682 4140
rect 13004 4137 13032 4168
rect 14458 4156 14464 4168
rect 14516 4156 14522 4208
rect 14642 4156 14648 4208
rect 14700 4156 14706 4208
rect 15580 4196 15608 4227
rect 15746 4224 15752 4276
rect 15804 4264 15810 4276
rect 16022 4264 16028 4276
rect 15804 4236 16028 4264
rect 15804 4224 15810 4236
rect 16022 4224 16028 4236
rect 16080 4224 16086 4276
rect 16206 4224 16212 4276
rect 16264 4264 16270 4276
rect 18414 4264 18420 4276
rect 16264 4236 17448 4264
rect 18375 4236 18420 4264
rect 16264 4224 16270 4236
rect 15838 4196 15844 4208
rect 15580 4168 15844 4196
rect 15838 4156 15844 4168
rect 15896 4156 15902 4208
rect 16482 4156 16488 4208
rect 16540 4156 16546 4208
rect 12989 4131 13047 4137
rect 12989 4097 13001 4131
rect 13035 4097 13047 4131
rect 14550 4128 14556 4140
rect 14511 4100 14556 4128
rect 12989 4091 13047 4097
rect 14550 4088 14556 4100
rect 14608 4088 14614 4140
rect 14660 4128 14688 4156
rect 14918 4128 14924 4140
rect 14660 4100 14924 4128
rect 14918 4088 14924 4100
rect 14976 4088 14982 4140
rect 15105 4131 15163 4137
rect 15105 4097 15117 4131
rect 15151 4128 15163 4131
rect 15562 4128 15568 4140
rect 15151 4100 15568 4128
rect 15151 4097 15163 4100
rect 15105 4091 15163 4097
rect 15562 4088 15568 4100
rect 15620 4088 15626 4140
rect 16209 4131 16267 4137
rect 16209 4097 16221 4131
rect 16255 4128 16267 4131
rect 16298 4128 16304 4140
rect 16255 4100 16304 4128
rect 16255 4097 16267 4100
rect 16209 4091 16267 4097
rect 16298 4088 16304 4100
rect 16356 4088 16362 4140
rect 16500 4128 16528 4156
rect 17420 4128 17448 4236
rect 18414 4224 18420 4236
rect 18472 4224 18478 4276
rect 19426 4264 19432 4276
rect 19387 4236 19432 4264
rect 19426 4224 19432 4236
rect 19484 4224 19490 4276
rect 20806 4224 20812 4276
rect 20864 4264 20870 4276
rect 21085 4267 21143 4273
rect 21085 4264 21097 4267
rect 20864 4236 21097 4264
rect 20864 4224 20870 4236
rect 21085 4233 21097 4236
rect 21131 4264 21143 4267
rect 21634 4264 21640 4276
rect 21131 4236 21640 4264
rect 21131 4233 21143 4236
rect 21085 4227 21143 4233
rect 21634 4224 21640 4236
rect 21692 4224 21698 4276
rect 22649 4267 22707 4273
rect 22649 4233 22661 4267
rect 22695 4264 22707 4267
rect 22922 4264 22928 4276
rect 22695 4236 22928 4264
rect 22695 4233 22707 4236
rect 22649 4227 22707 4233
rect 22922 4224 22928 4236
rect 22980 4264 22986 4276
rect 22980 4236 24900 4264
rect 22980 4224 22986 4236
rect 17865 4199 17923 4205
rect 17865 4165 17877 4199
rect 17911 4196 17923 4199
rect 18322 4196 18328 4208
rect 17911 4168 18328 4196
rect 17911 4165 17923 4168
rect 17865 4159 17923 4165
rect 18322 4156 18328 4168
rect 18380 4156 18386 4208
rect 19444 4196 19472 4224
rect 19076 4168 19472 4196
rect 19889 4199 19947 4205
rect 18141 4131 18199 4137
rect 18141 4128 18153 4131
rect 16500 4100 16712 4128
rect 17420 4100 18153 4128
rect 12526 4020 12532 4072
rect 12584 4060 12590 4072
rect 12897 4063 12955 4069
rect 12897 4060 12909 4063
rect 12584 4032 12909 4060
rect 12584 4020 12590 4032
rect 12897 4029 12909 4032
rect 12943 4060 12955 4063
rect 13538 4060 13544 4072
rect 12943 4032 13544 4060
rect 12943 4029 12955 4032
rect 12897 4023 12955 4029
rect 13538 4020 13544 4032
rect 13596 4020 13602 4072
rect 14366 4060 14372 4072
rect 14327 4032 14372 4060
rect 14366 4020 14372 4032
rect 14424 4060 14430 4072
rect 14642 4060 14648 4072
rect 14424 4032 14648 4060
rect 14424 4020 14430 4032
rect 14642 4020 14648 4032
rect 14700 4020 14706 4072
rect 15473 4063 15531 4069
rect 15473 4029 15485 4063
rect 15519 4060 15531 4063
rect 16025 4063 16083 4069
rect 16025 4060 16037 4063
rect 15519 4032 16037 4060
rect 15519 4029 15531 4032
rect 15473 4023 15531 4029
rect 16025 4029 16037 4032
rect 16071 4060 16083 4063
rect 16390 4060 16396 4072
rect 16071 4032 16396 4060
rect 16071 4029 16083 4032
rect 16025 4023 16083 4029
rect 16390 4020 16396 4032
rect 16448 4020 16454 4072
rect 16684 4069 16712 4100
rect 18141 4097 18153 4100
rect 18187 4128 18199 4131
rect 18233 4131 18291 4137
rect 18233 4128 18245 4131
rect 18187 4100 18245 4128
rect 18187 4097 18199 4100
rect 18141 4091 18199 4097
rect 18233 4097 18245 4100
rect 18279 4097 18291 4131
rect 18233 4091 18291 4097
rect 18782 4088 18788 4140
rect 18840 4128 18846 4140
rect 19076 4137 19104 4168
rect 19889 4165 19901 4199
rect 19935 4196 19947 4199
rect 20162 4196 20168 4208
rect 19935 4168 20168 4196
rect 19935 4165 19947 4168
rect 19889 4159 19947 4165
rect 20162 4156 20168 4168
rect 20220 4196 20226 4208
rect 20220 4168 20576 4196
rect 20220 4156 20226 4168
rect 18877 4131 18935 4137
rect 18877 4128 18889 4131
rect 18840 4100 18889 4128
rect 18840 4088 18846 4100
rect 18877 4097 18889 4100
rect 18923 4097 18935 4131
rect 18877 4091 18935 4097
rect 19061 4131 19119 4137
rect 19061 4097 19073 4131
rect 19107 4097 19119 4131
rect 20438 4128 20444 4140
rect 20399 4100 20444 4128
rect 19061 4091 19119 4097
rect 20438 4088 20444 4100
rect 20496 4088 20502 4140
rect 20548 4137 20576 4168
rect 21726 4156 21732 4208
rect 21784 4196 21790 4208
rect 22370 4196 22376 4208
rect 21784 4168 22376 4196
rect 21784 4156 21790 4168
rect 22204 4137 22232 4168
rect 22370 4156 22376 4168
rect 22428 4196 22434 4208
rect 23750 4196 23756 4208
rect 22428 4168 23756 4196
rect 22428 4156 22434 4168
rect 23750 4156 23756 4168
rect 23808 4156 23814 4208
rect 23934 4156 23940 4208
rect 23992 4196 23998 4208
rect 24872 4196 24900 4236
rect 25774 4224 25780 4276
rect 25832 4264 25838 4276
rect 26145 4267 26203 4273
rect 26145 4264 26157 4267
rect 25832 4236 26157 4264
rect 25832 4224 25838 4236
rect 26145 4233 26157 4236
rect 26191 4264 26203 4267
rect 26234 4264 26240 4276
rect 26191 4236 26240 4264
rect 26191 4233 26203 4236
rect 26145 4227 26203 4233
rect 26234 4224 26240 4236
rect 26292 4224 26298 4276
rect 25866 4196 25872 4208
rect 23992 4168 24808 4196
rect 24872 4168 25872 4196
rect 23992 4156 23998 4168
rect 20533 4131 20591 4137
rect 20533 4097 20545 4131
rect 20579 4097 20591 4131
rect 20533 4091 20591 4097
rect 22189 4131 22247 4137
rect 22189 4097 22201 4131
rect 22235 4097 22247 4131
rect 22189 4091 22247 4097
rect 22554 4088 22560 4140
rect 22612 4128 22618 4140
rect 22925 4131 22983 4137
rect 22925 4128 22937 4131
rect 22612 4100 22937 4128
rect 22612 4088 22618 4100
rect 22925 4097 22937 4100
rect 22971 4097 22983 4131
rect 22925 4091 22983 4097
rect 24121 4131 24179 4137
rect 24121 4097 24133 4131
rect 24167 4128 24179 4131
rect 24210 4128 24216 4140
rect 24167 4100 24216 4128
rect 24167 4097 24179 4100
rect 24121 4091 24179 4097
rect 24210 4088 24216 4100
rect 24268 4088 24274 4140
rect 24305 4131 24363 4137
rect 24305 4097 24317 4131
rect 24351 4128 24363 4131
rect 24670 4128 24676 4140
rect 24351 4100 24676 4128
rect 24351 4097 24363 4100
rect 24305 4091 24363 4097
rect 24670 4088 24676 4100
rect 24728 4088 24734 4140
rect 24780 4128 24808 4168
rect 25866 4156 25872 4168
rect 25924 4156 25930 4208
rect 25041 4131 25099 4137
rect 25041 4128 25053 4131
rect 24780 4100 25053 4128
rect 25041 4097 25053 4100
rect 25087 4097 25099 4131
rect 25041 4091 25099 4097
rect 16669 4063 16727 4069
rect 16669 4029 16681 4063
rect 16715 4060 16727 4063
rect 16942 4060 16948 4072
rect 16715 4032 16948 4060
rect 16715 4029 16727 4032
rect 16669 4023 16727 4029
rect 16942 4020 16948 4032
rect 17000 4060 17006 4072
rect 17000 4032 24164 4060
rect 17000 4020 17006 4032
rect 24136 4004 24164 4032
rect 24578 4020 24584 4072
rect 24636 4060 24642 4072
rect 24946 4060 24952 4072
rect 24636 4032 24952 4060
rect 24636 4020 24642 4032
rect 24946 4020 24952 4032
rect 25004 4020 25010 4072
rect 25222 4060 25228 4072
rect 25183 4032 25228 4060
rect 25222 4020 25228 4032
rect 25280 4060 25286 4072
rect 25777 4063 25835 4069
rect 25777 4060 25789 4063
rect 25280 4032 25789 4060
rect 25280 4020 25286 4032
rect 25777 4029 25789 4032
rect 25823 4029 25835 4063
rect 25777 4023 25835 4029
rect 10183 3964 11560 3992
rect 12253 3995 12311 4001
rect 10183 3961 10195 3964
rect 10137 3955 10195 3961
rect 12253 3961 12265 3995
rect 12299 3992 12311 3995
rect 12805 3995 12863 4001
rect 12805 3992 12817 3995
rect 12299 3964 12817 3992
rect 12299 3961 12311 3964
rect 12253 3955 12311 3961
rect 12805 3961 12817 3964
rect 12851 3992 12863 3995
rect 14090 3992 14096 4004
rect 12851 3964 14096 3992
rect 12851 3961 12863 3964
rect 12805 3955 12863 3961
rect 14090 3952 14096 3964
rect 14148 3952 14154 4004
rect 15562 3952 15568 4004
rect 15620 3992 15626 4004
rect 15933 3995 15991 4001
rect 15933 3992 15945 3995
rect 15620 3964 15945 3992
rect 15620 3952 15626 3964
rect 15933 3961 15945 3964
rect 15979 3961 15991 3995
rect 15933 3955 15991 3961
rect 17497 3995 17555 4001
rect 17497 3961 17509 3995
rect 17543 3992 17555 3995
rect 18690 3992 18696 4004
rect 17543 3964 18696 3992
rect 17543 3961 17555 3964
rect 17497 3955 17555 3961
rect 18690 3952 18696 3964
rect 18748 3952 18754 4004
rect 20622 3992 20628 4004
rect 19996 3964 20628 3992
rect 1397 3927 1455 3933
rect 1397 3893 1409 3927
rect 1443 3924 1455 3927
rect 1578 3924 1584 3936
rect 1443 3896 1584 3924
rect 1443 3893 1455 3896
rect 1397 3887 1455 3893
rect 1578 3884 1584 3896
rect 1636 3884 1642 3936
rect 1765 3927 1823 3933
rect 1765 3893 1777 3927
rect 1811 3924 1823 3927
rect 2314 3924 2320 3936
rect 1811 3896 2320 3924
rect 1811 3893 1823 3896
rect 1765 3887 1823 3893
rect 2314 3884 2320 3896
rect 2372 3884 2378 3936
rect 2958 3924 2964 3936
rect 2919 3896 2964 3924
rect 2958 3884 2964 3896
rect 3016 3884 3022 3936
rect 5350 3924 5356 3936
rect 5311 3896 5356 3924
rect 5350 3884 5356 3896
rect 5408 3884 5414 3936
rect 6362 3924 6368 3936
rect 6323 3896 6368 3924
rect 6362 3884 6368 3896
rect 6420 3884 6426 3936
rect 8294 3884 8300 3936
rect 8352 3924 8358 3936
rect 8573 3927 8631 3933
rect 8573 3924 8585 3927
rect 8352 3896 8585 3924
rect 8352 3884 8358 3896
rect 8573 3893 8585 3896
rect 8619 3893 8631 3927
rect 9122 3924 9128 3936
rect 9083 3896 9128 3924
rect 8573 3887 8631 3893
rect 9122 3884 9128 3896
rect 9180 3924 9186 3936
rect 9950 3924 9956 3936
rect 9180 3896 9956 3924
rect 9180 3884 9186 3896
rect 9950 3884 9956 3896
rect 10008 3884 10014 3936
rect 11422 3924 11428 3936
rect 11383 3896 11428 3924
rect 11422 3884 11428 3896
rect 11480 3884 11486 3936
rect 12437 3927 12495 3933
rect 12437 3893 12449 3927
rect 12483 3924 12495 3927
rect 12618 3924 12624 3936
rect 12483 3896 12624 3924
rect 12483 3893 12495 3896
rect 12437 3887 12495 3893
rect 12618 3884 12624 3896
rect 12676 3884 12682 3936
rect 13446 3924 13452 3936
rect 13407 3896 13452 3924
rect 13446 3884 13452 3896
rect 13504 3924 13510 3936
rect 13814 3924 13820 3936
rect 13504 3896 13820 3924
rect 13504 3884 13510 3896
rect 13814 3884 13820 3896
rect 13872 3884 13878 3936
rect 13998 3924 14004 3936
rect 13959 3896 14004 3924
rect 13998 3884 14004 3896
rect 14056 3884 14062 3936
rect 14461 3927 14519 3933
rect 14461 3893 14473 3927
rect 14507 3924 14519 3927
rect 14734 3924 14740 3936
rect 14507 3896 14740 3924
rect 14507 3893 14519 3896
rect 14461 3887 14519 3893
rect 14734 3884 14740 3896
rect 14792 3884 14798 3936
rect 16942 3924 16948 3936
rect 16903 3896 16948 3924
rect 16942 3884 16948 3896
rect 17000 3884 17006 3936
rect 18141 3927 18199 3933
rect 18141 3893 18153 3927
rect 18187 3924 18199 3927
rect 18782 3924 18788 3936
rect 18187 3896 18788 3924
rect 18187 3893 18199 3896
rect 18141 3887 18199 3893
rect 18782 3884 18788 3896
rect 18840 3884 18846 3936
rect 19996 3933 20024 3964
rect 20622 3952 20628 3964
rect 20680 3952 20686 4004
rect 21913 3995 21971 4001
rect 21913 3992 21925 3995
rect 21376 3964 21925 3992
rect 21376 3936 21404 3964
rect 21913 3961 21925 3964
rect 21959 3961 21971 3995
rect 21913 3955 21971 3961
rect 22005 3995 22063 4001
rect 22005 3961 22017 3995
rect 22051 3992 22063 3995
rect 22278 3992 22284 4004
rect 22051 3964 22284 3992
rect 22051 3961 22063 3964
rect 22005 3955 22063 3961
rect 22278 3952 22284 3964
rect 22336 3952 22342 4004
rect 23477 3995 23535 4001
rect 23477 3961 23489 3995
rect 23523 3992 23535 3995
rect 23523 3964 24072 3992
rect 23523 3961 23535 3964
rect 23477 3955 23535 3961
rect 19981 3927 20039 3933
rect 19981 3893 19993 3927
rect 20027 3893 20039 3927
rect 20346 3924 20352 3936
rect 20307 3896 20352 3924
rect 19981 3887 20039 3893
rect 20346 3884 20352 3896
rect 20404 3884 20410 3936
rect 21358 3924 21364 3936
rect 21319 3896 21364 3924
rect 21358 3884 21364 3896
rect 21416 3884 21422 3936
rect 21545 3927 21603 3933
rect 21545 3893 21557 3927
rect 21591 3924 21603 3927
rect 21818 3924 21824 3936
rect 21591 3896 21824 3924
rect 21591 3893 21603 3896
rect 21545 3887 21603 3893
rect 21818 3884 21824 3896
rect 21876 3884 21882 3936
rect 23658 3924 23664 3936
rect 23619 3896 23664 3924
rect 23658 3884 23664 3896
rect 23716 3884 23722 3936
rect 24044 3933 24072 3964
rect 24118 3952 24124 4004
rect 24176 3952 24182 4004
rect 24765 3995 24823 4001
rect 24765 3961 24777 3995
rect 24811 3992 24823 3995
rect 24854 3992 24860 4004
rect 24811 3964 24860 3992
rect 24811 3961 24823 3964
rect 24765 3955 24823 3961
rect 24854 3952 24860 3964
rect 24912 3952 24918 4004
rect 24029 3927 24087 3933
rect 24029 3893 24041 3927
rect 24075 3924 24087 3927
rect 24210 3924 24216 3936
rect 24075 3896 24216 3924
rect 24075 3893 24087 3896
rect 24029 3887 24087 3893
rect 24210 3884 24216 3896
rect 24268 3884 24274 3936
rect 25406 3924 25412 3936
rect 25367 3896 25412 3924
rect 25406 3884 25412 3896
rect 25464 3884 25470 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1397 3723 1455 3729
rect 1397 3689 1409 3723
rect 1443 3720 1455 3723
rect 1486 3720 1492 3732
rect 1443 3692 1492 3720
rect 1443 3689 1455 3692
rect 1397 3683 1455 3689
rect 1486 3680 1492 3692
rect 1544 3680 1550 3732
rect 1762 3720 1768 3732
rect 1723 3692 1768 3720
rect 1762 3680 1768 3692
rect 1820 3680 1826 3732
rect 1857 3723 1915 3729
rect 1857 3689 1869 3723
rect 1903 3720 1915 3723
rect 2222 3720 2228 3732
rect 1903 3692 2228 3720
rect 1903 3689 1915 3692
rect 1857 3683 1915 3689
rect 1578 3612 1584 3664
rect 1636 3652 1642 3664
rect 1872 3652 1900 3683
rect 2222 3680 2228 3692
rect 2280 3680 2286 3732
rect 2314 3680 2320 3732
rect 2372 3720 2378 3732
rect 2409 3723 2467 3729
rect 2409 3720 2421 3723
rect 2372 3692 2421 3720
rect 2372 3680 2378 3692
rect 2409 3689 2421 3692
rect 2455 3689 2467 3723
rect 5534 3720 5540 3732
rect 2409 3683 2467 3689
rect 3436 3692 5540 3720
rect 1636 3624 1900 3652
rect 1636 3612 1642 3624
rect 2130 3612 2136 3664
rect 2188 3652 2194 3664
rect 3436 3661 3464 3692
rect 5534 3680 5540 3692
rect 5592 3680 5598 3732
rect 6089 3723 6147 3729
rect 6089 3689 6101 3723
rect 6135 3720 6147 3723
rect 6270 3720 6276 3732
rect 6135 3692 6276 3720
rect 6135 3689 6147 3692
rect 6089 3683 6147 3689
rect 6270 3680 6276 3692
rect 6328 3680 6334 3732
rect 6457 3723 6515 3729
rect 6457 3689 6469 3723
rect 6503 3720 6515 3723
rect 6546 3720 6552 3732
rect 6503 3692 6552 3720
rect 6503 3689 6515 3692
rect 6457 3683 6515 3689
rect 6546 3680 6552 3692
rect 6604 3680 6610 3732
rect 7466 3680 7472 3732
rect 7524 3720 7530 3732
rect 7653 3723 7711 3729
rect 7653 3720 7665 3723
rect 7524 3692 7665 3720
rect 7524 3680 7530 3692
rect 7653 3689 7665 3692
rect 7699 3689 7711 3723
rect 7834 3720 7840 3732
rect 7795 3692 7840 3720
rect 7653 3683 7711 3689
rect 2777 3655 2835 3661
rect 2777 3652 2789 3655
rect 2188 3624 2789 3652
rect 2188 3612 2194 3624
rect 2777 3621 2789 3624
rect 2823 3652 2835 3655
rect 3421 3655 3479 3661
rect 3421 3652 3433 3655
rect 2823 3624 3433 3652
rect 2823 3621 2835 3624
rect 2777 3615 2835 3621
rect 3421 3621 3433 3624
rect 3467 3621 3479 3655
rect 3421 3615 3479 3621
rect 3881 3655 3939 3661
rect 3881 3621 3893 3655
rect 3927 3652 3939 3655
rect 4154 3652 4160 3664
rect 3927 3624 4160 3652
rect 3927 3621 3939 3624
rect 3881 3615 3939 3621
rect 4154 3612 4160 3624
rect 4212 3652 4218 3664
rect 4332 3655 4390 3661
rect 4332 3652 4344 3655
rect 4212 3624 4344 3652
rect 4212 3612 4218 3624
rect 4332 3621 4344 3624
rect 4378 3652 4390 3655
rect 5350 3652 5356 3664
rect 4378 3624 5356 3652
rect 4378 3621 4390 3624
rect 4332 3615 4390 3621
rect 5350 3612 5356 3624
rect 5408 3612 5414 3664
rect 3970 3544 3976 3596
rect 4028 3584 4034 3596
rect 4065 3587 4123 3593
rect 4065 3584 4077 3587
rect 4028 3556 4077 3584
rect 4028 3544 4034 3556
rect 4065 3553 4077 3556
rect 4111 3584 4123 3587
rect 4706 3584 4712 3596
rect 4111 3556 4712 3584
rect 4111 3553 4123 3556
rect 4065 3547 4123 3553
rect 4706 3544 4712 3556
rect 4764 3544 4770 3596
rect 6564 3593 6592 3680
rect 6638 3612 6644 3664
rect 6696 3652 6702 3664
rect 6825 3655 6883 3661
rect 6825 3652 6837 3655
rect 6696 3624 6837 3652
rect 6696 3612 6702 3624
rect 6825 3621 6837 3624
rect 6871 3621 6883 3655
rect 7668 3652 7696 3683
rect 7834 3680 7840 3692
rect 7892 3680 7898 3732
rect 8202 3720 8208 3732
rect 8115 3692 8208 3720
rect 8202 3680 8208 3692
rect 8260 3720 8266 3732
rect 9122 3720 9128 3732
rect 8260 3692 9128 3720
rect 8260 3680 8266 3692
rect 9122 3680 9128 3692
rect 9180 3680 9186 3732
rect 9674 3720 9680 3732
rect 9635 3692 9680 3720
rect 9674 3680 9680 3692
rect 9732 3680 9738 3732
rect 9950 3680 9956 3732
rect 10008 3720 10014 3732
rect 10045 3723 10103 3729
rect 10045 3720 10057 3723
rect 10008 3692 10057 3720
rect 10008 3680 10014 3692
rect 10045 3689 10057 3692
rect 10091 3689 10103 3723
rect 10045 3683 10103 3689
rect 10962 3680 10968 3732
rect 11020 3720 11026 3732
rect 11241 3723 11299 3729
rect 11241 3720 11253 3723
rect 11020 3692 11253 3720
rect 11020 3680 11026 3692
rect 11241 3689 11253 3692
rect 11287 3720 11299 3723
rect 12526 3720 12532 3732
rect 11287 3692 12020 3720
rect 12487 3692 12532 3720
rect 11287 3689 11299 3692
rect 11241 3683 11299 3689
rect 11606 3652 11612 3664
rect 7668 3624 8340 3652
rect 11567 3624 11612 3652
rect 6825 3615 6883 3621
rect 6549 3587 6607 3593
rect 6549 3553 6561 3587
rect 6595 3553 6607 3587
rect 8312 3584 8340 3624
rect 11606 3612 11612 3624
rect 11664 3612 11670 3664
rect 11992 3652 12020 3692
rect 12526 3680 12532 3692
rect 12584 3680 12590 3732
rect 12802 3720 12808 3732
rect 12763 3692 12808 3720
rect 12802 3680 12808 3692
rect 12860 3680 12866 3732
rect 13170 3680 13176 3732
rect 13228 3680 13234 3732
rect 13265 3723 13323 3729
rect 13265 3689 13277 3723
rect 13311 3720 13323 3723
rect 13722 3720 13728 3732
rect 13311 3692 13728 3720
rect 13311 3689 13323 3692
rect 13265 3683 13323 3689
rect 13722 3680 13728 3692
rect 13780 3680 13786 3732
rect 15289 3723 15347 3729
rect 15289 3689 15301 3723
rect 15335 3720 15347 3723
rect 15654 3720 15660 3732
rect 15335 3692 15660 3720
rect 15335 3689 15347 3692
rect 15289 3683 15347 3689
rect 15654 3680 15660 3692
rect 15712 3680 15718 3732
rect 15749 3723 15807 3729
rect 15749 3689 15761 3723
rect 15795 3720 15807 3723
rect 16853 3723 16911 3729
rect 16853 3720 16865 3723
rect 15795 3692 16865 3720
rect 15795 3689 15807 3692
rect 15749 3683 15807 3689
rect 16853 3689 16865 3692
rect 16899 3720 16911 3723
rect 16942 3720 16948 3732
rect 16899 3692 16948 3720
rect 16899 3689 16911 3692
rect 16853 3683 16911 3689
rect 16942 3680 16948 3692
rect 17000 3680 17006 3732
rect 17126 3680 17132 3732
rect 17184 3720 17190 3732
rect 17313 3723 17371 3729
rect 17313 3720 17325 3723
rect 17184 3692 17325 3720
rect 17184 3680 17190 3692
rect 17313 3689 17325 3692
rect 17359 3689 17371 3723
rect 17313 3683 17371 3689
rect 18046 3680 18052 3732
rect 18104 3720 18110 3732
rect 18874 3720 18880 3732
rect 18104 3692 18880 3720
rect 18104 3680 18110 3692
rect 18874 3680 18880 3692
rect 18932 3680 18938 3732
rect 19426 3680 19432 3732
rect 19484 3720 19490 3732
rect 19889 3723 19947 3729
rect 19889 3720 19901 3723
rect 19484 3692 19901 3720
rect 19484 3680 19490 3692
rect 19889 3689 19901 3692
rect 19935 3689 19947 3723
rect 19889 3683 19947 3689
rect 21361 3723 21419 3729
rect 21361 3689 21373 3723
rect 21407 3720 21419 3723
rect 22002 3720 22008 3732
rect 21407 3692 22008 3720
rect 21407 3689 21419 3692
rect 21361 3683 21419 3689
rect 22002 3680 22008 3692
rect 22060 3680 22066 3732
rect 22370 3720 22376 3732
rect 22331 3692 22376 3720
rect 22370 3680 22376 3692
rect 22428 3680 22434 3732
rect 22830 3720 22836 3732
rect 22791 3692 22836 3720
rect 22830 3680 22836 3692
rect 22888 3680 22894 3732
rect 22925 3723 22983 3729
rect 22925 3689 22937 3723
rect 22971 3720 22983 3723
rect 23106 3720 23112 3732
rect 22971 3692 23112 3720
rect 22971 3689 22983 3692
rect 22925 3683 22983 3689
rect 23106 3680 23112 3692
rect 23164 3680 23170 3732
rect 23474 3680 23480 3732
rect 23532 3720 23538 3732
rect 24029 3723 24087 3729
rect 24029 3720 24041 3723
rect 23532 3692 24041 3720
rect 23532 3680 23538 3692
rect 24029 3689 24041 3692
rect 24075 3689 24087 3723
rect 24394 3720 24400 3732
rect 24355 3692 24400 3720
rect 24029 3683 24087 3689
rect 24394 3680 24400 3692
rect 24452 3680 24458 3732
rect 24489 3723 24547 3729
rect 24489 3689 24501 3723
rect 24535 3720 24547 3723
rect 24535 3692 24808 3720
rect 24535 3689 24547 3692
rect 24489 3683 24547 3689
rect 13188 3652 13216 3680
rect 16298 3652 16304 3664
rect 11992 3624 13216 3652
rect 16259 3624 16304 3652
rect 16298 3612 16304 3624
rect 16356 3612 16362 3664
rect 16758 3652 16764 3664
rect 16719 3624 16764 3652
rect 16758 3612 16764 3624
rect 16816 3652 16822 3664
rect 17221 3655 17279 3661
rect 17221 3652 17233 3655
rect 16816 3624 17233 3652
rect 16816 3612 16822 3624
rect 17221 3621 17233 3624
rect 17267 3621 17279 3655
rect 18782 3652 18788 3664
rect 18743 3624 18788 3652
rect 17221 3615 17279 3621
rect 18782 3612 18788 3624
rect 18840 3612 18846 3664
rect 21269 3655 21327 3661
rect 21269 3621 21281 3655
rect 21315 3652 21327 3655
rect 21818 3652 21824 3664
rect 21315 3624 21824 3652
rect 21315 3621 21327 3624
rect 21269 3615 21327 3621
rect 21818 3612 21824 3624
rect 21876 3612 21882 3664
rect 21913 3655 21971 3661
rect 21913 3621 21925 3655
rect 21959 3652 21971 3655
rect 22278 3652 22284 3664
rect 21959 3624 22284 3652
rect 21959 3621 21971 3624
rect 21913 3615 21971 3621
rect 22278 3612 22284 3624
rect 22336 3612 22342 3664
rect 8312 3556 8432 3584
rect 6549 3547 6607 3553
rect 2041 3519 2099 3525
rect 2041 3485 2053 3519
rect 2087 3516 2099 3519
rect 2130 3516 2136 3528
rect 2087 3488 2136 3516
rect 2087 3485 2099 3488
rect 2041 3479 2099 3485
rect 2130 3476 2136 3488
rect 2188 3476 2194 3528
rect 2958 3516 2964 3528
rect 2919 3488 2964 3516
rect 2958 3476 2964 3488
rect 3016 3476 3022 3528
rect 7742 3476 7748 3528
rect 7800 3516 7806 3528
rect 8404 3525 8432 3556
rect 9858 3544 9864 3596
rect 9916 3584 9922 3596
rect 10689 3587 10747 3593
rect 10689 3584 10701 3587
rect 9916 3556 10701 3584
rect 9916 3544 9922 3556
rect 8297 3519 8355 3525
rect 8297 3516 8309 3519
rect 7800 3488 8309 3516
rect 7800 3476 7806 3488
rect 8297 3485 8309 3488
rect 8343 3485 8355 3519
rect 8297 3479 8355 3485
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3516 8447 3519
rect 8478 3516 8484 3528
rect 8435 3488 8484 3516
rect 8435 3485 8447 3488
rect 8389 3479 8447 3485
rect 8478 3476 8484 3488
rect 8536 3516 8542 3528
rect 9033 3519 9091 3525
rect 9033 3516 9045 3519
rect 8536 3488 9045 3516
rect 8536 3476 8542 3488
rect 9033 3485 9045 3488
rect 9079 3516 9091 3519
rect 9214 3516 9220 3528
rect 9079 3488 9220 3516
rect 9079 3485 9091 3488
rect 9033 3479 9091 3485
rect 9214 3476 9220 3488
rect 9272 3476 9278 3528
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10244 3525 10272 3556
rect 10689 3553 10701 3556
rect 10735 3584 10747 3587
rect 11057 3587 11115 3593
rect 11057 3584 11069 3587
rect 10735 3556 11069 3584
rect 10735 3553 10747 3556
rect 10689 3547 10747 3553
rect 11057 3553 11069 3556
rect 11103 3584 11115 3587
rect 11103 3556 11836 3584
rect 11103 3553 11115 3556
rect 11057 3547 11115 3553
rect 10137 3519 10195 3525
rect 10137 3516 10149 3519
rect 10008 3488 10149 3516
rect 10008 3476 10014 3488
rect 10137 3485 10149 3488
rect 10183 3485 10195 3519
rect 10137 3479 10195 3485
rect 10229 3519 10287 3525
rect 10229 3485 10241 3519
rect 10275 3485 10287 3519
rect 11698 3516 11704 3528
rect 11659 3488 11704 3516
rect 10229 3479 10287 3485
rect 11698 3476 11704 3488
rect 11756 3476 11762 3528
rect 11808 3525 11836 3556
rect 12250 3544 12256 3596
rect 12308 3584 12314 3596
rect 13173 3587 13231 3593
rect 13173 3584 13185 3587
rect 12308 3556 13185 3584
rect 12308 3544 12314 3556
rect 13173 3553 13185 3556
rect 13219 3584 13231 3587
rect 13262 3584 13268 3596
rect 13219 3556 13268 3584
rect 13219 3553 13231 3556
rect 13173 3547 13231 3553
rect 13262 3544 13268 3556
rect 13320 3544 13326 3596
rect 15105 3587 15163 3593
rect 15105 3553 15117 3587
rect 15151 3584 15163 3587
rect 15470 3584 15476 3596
rect 15151 3556 15476 3584
rect 15151 3553 15163 3556
rect 15105 3547 15163 3553
rect 15470 3544 15476 3556
rect 15528 3584 15534 3596
rect 15657 3587 15715 3593
rect 15657 3584 15669 3587
rect 15528 3556 15669 3584
rect 15528 3544 15534 3556
rect 15657 3553 15669 3556
rect 15703 3553 15715 3587
rect 15657 3547 15715 3553
rect 19150 3544 19156 3596
rect 19208 3584 19214 3596
rect 23753 3587 23811 3593
rect 19208 3556 23704 3584
rect 19208 3544 19214 3556
rect 11793 3519 11851 3525
rect 11793 3485 11805 3519
rect 11839 3485 11851 3519
rect 11793 3479 11851 3485
rect 13357 3519 13415 3525
rect 13357 3485 13369 3519
rect 13403 3516 13415 3519
rect 14001 3519 14059 3525
rect 14001 3516 14013 3519
rect 13403 3488 14013 3516
rect 13403 3485 13415 3488
rect 13357 3479 13415 3485
rect 14001 3485 14013 3488
rect 14047 3516 14059 3519
rect 14369 3519 14427 3525
rect 14369 3516 14381 3519
rect 14047 3488 14381 3516
rect 14047 3485 14059 3488
rect 14001 3479 14059 3485
rect 14369 3485 14381 3488
rect 14415 3516 14427 3519
rect 14550 3516 14556 3528
rect 14415 3488 14556 3516
rect 14415 3485 14427 3488
rect 14369 3479 14427 3485
rect 8202 3448 8208 3460
rect 5092 3420 8208 3448
rect 3878 3340 3884 3392
rect 3936 3380 3942 3392
rect 5092 3380 5120 3420
rect 8202 3408 8208 3420
rect 8260 3408 8266 3460
rect 12526 3408 12532 3460
rect 12584 3448 12590 3460
rect 13372 3448 13400 3479
rect 14550 3476 14556 3488
rect 14608 3476 14614 3528
rect 15838 3516 15844 3528
rect 15799 3488 15844 3516
rect 15838 3476 15844 3488
rect 15896 3476 15902 3528
rect 16850 3476 16856 3528
rect 16908 3516 16914 3528
rect 17405 3519 17463 3525
rect 17405 3516 17417 3519
rect 16908 3488 17417 3516
rect 16908 3476 16914 3488
rect 17405 3485 17417 3488
rect 17451 3485 17463 3519
rect 18969 3519 19027 3525
rect 18969 3516 18981 3519
rect 17405 3479 17463 3485
rect 18064 3488 18981 3516
rect 12584 3420 13400 3448
rect 12584 3408 12590 3420
rect 5442 3380 5448 3392
rect 3936 3352 5120 3380
rect 5403 3352 5448 3380
rect 3936 3340 3942 3352
rect 5442 3340 5448 3352
rect 5500 3340 5506 3392
rect 7377 3383 7435 3389
rect 7377 3349 7389 3383
rect 7423 3380 7435 3383
rect 7466 3380 7472 3392
rect 7423 3352 7472 3380
rect 7423 3349 7435 3352
rect 7377 3343 7435 3349
rect 7466 3340 7472 3352
rect 7524 3340 7530 3392
rect 9493 3383 9551 3389
rect 9493 3349 9505 3383
rect 9539 3380 9551 3383
rect 9858 3380 9864 3392
rect 9539 3352 9864 3380
rect 9539 3349 9551 3352
rect 9493 3343 9551 3349
rect 9858 3340 9864 3352
rect 9916 3340 9922 3392
rect 12802 3340 12808 3392
rect 12860 3380 12866 3392
rect 13630 3380 13636 3392
rect 12860 3352 13636 3380
rect 12860 3340 12866 3352
rect 13630 3340 13636 3352
rect 13688 3340 13694 3392
rect 14366 3340 14372 3392
rect 14424 3380 14430 3392
rect 17678 3380 17684 3392
rect 14424 3352 17684 3380
rect 14424 3340 14430 3352
rect 17678 3340 17684 3352
rect 17736 3340 17742 3392
rect 17770 3340 17776 3392
rect 17828 3380 17834 3392
rect 18064 3389 18092 3488
rect 18969 3485 18981 3488
rect 19015 3485 19027 3519
rect 21450 3516 21456 3528
rect 21411 3488 21456 3516
rect 18969 3479 19027 3485
rect 21450 3476 21456 3488
rect 21508 3476 21514 3528
rect 21726 3476 21732 3528
rect 21784 3516 21790 3528
rect 23106 3516 23112 3528
rect 21784 3488 22876 3516
rect 23067 3488 23112 3516
rect 21784 3476 21790 3488
rect 18414 3448 18420 3460
rect 18375 3420 18420 3448
rect 18414 3408 18420 3420
rect 18472 3408 18478 3460
rect 19613 3451 19671 3457
rect 19613 3417 19625 3451
rect 19659 3448 19671 3451
rect 20070 3448 20076 3460
rect 19659 3420 20076 3448
rect 19659 3417 19671 3420
rect 19613 3411 19671 3417
rect 20070 3408 20076 3420
rect 20128 3408 20134 3460
rect 20346 3408 20352 3460
rect 20404 3448 20410 3460
rect 20901 3451 20959 3457
rect 20901 3448 20913 3451
rect 20404 3420 20913 3448
rect 20404 3408 20410 3420
rect 20901 3417 20913 3420
rect 20947 3448 20959 3451
rect 22002 3448 22008 3460
rect 20947 3420 22008 3448
rect 20947 3417 20959 3420
rect 20901 3411 20959 3417
rect 22002 3408 22008 3420
rect 22060 3408 22066 3460
rect 22848 3448 22876 3488
rect 23106 3476 23112 3488
rect 23164 3476 23170 3528
rect 23676 3516 23704 3556
rect 23753 3553 23765 3587
rect 23799 3584 23811 3587
rect 24302 3584 24308 3596
rect 23799 3556 24308 3584
rect 23799 3553 23811 3556
rect 23753 3547 23811 3553
rect 24302 3544 24308 3556
rect 24360 3544 24366 3596
rect 24412 3584 24440 3680
rect 24780 3652 24808 3692
rect 25130 3680 25136 3732
rect 25188 3720 25194 3732
rect 25409 3723 25467 3729
rect 25409 3720 25421 3723
rect 25188 3692 25421 3720
rect 25188 3680 25194 3692
rect 25409 3689 25421 3692
rect 25455 3689 25467 3723
rect 26234 3720 26240 3732
rect 26195 3692 26240 3720
rect 25409 3683 25467 3689
rect 26234 3680 26240 3692
rect 26292 3680 26298 3732
rect 25148 3652 25176 3680
rect 24780 3624 25176 3652
rect 25777 3587 25835 3593
rect 25777 3584 25789 3587
rect 24412 3556 25789 3584
rect 25777 3553 25789 3556
rect 25823 3553 25835 3587
rect 25777 3547 25835 3553
rect 24581 3519 24639 3525
rect 24581 3516 24593 3519
rect 23676 3488 24593 3516
rect 24581 3485 24593 3488
rect 24627 3516 24639 3519
rect 24854 3516 24860 3528
rect 24627 3488 24860 3516
rect 24627 3485 24639 3488
rect 24581 3479 24639 3485
rect 24854 3476 24860 3488
rect 24912 3476 24918 3528
rect 23124 3448 23152 3476
rect 22848 3420 23152 3448
rect 24118 3408 24124 3460
rect 24176 3448 24182 3460
rect 25041 3451 25099 3457
rect 25041 3448 25053 3451
rect 24176 3420 25053 3448
rect 24176 3408 24182 3420
rect 25041 3417 25053 3420
rect 25087 3417 25099 3451
rect 25041 3411 25099 3417
rect 18049 3383 18107 3389
rect 18049 3380 18061 3383
rect 17828 3352 18061 3380
rect 17828 3340 17834 3352
rect 18049 3349 18061 3352
rect 18095 3349 18107 3383
rect 20254 3380 20260 3392
rect 20215 3352 20260 3380
rect 18049 3343 18107 3349
rect 20254 3340 20260 3352
rect 20312 3340 20318 3392
rect 20717 3383 20775 3389
rect 20717 3349 20729 3383
rect 20763 3380 20775 3383
rect 21266 3380 21272 3392
rect 20763 3352 21272 3380
rect 20763 3349 20775 3352
rect 20717 3343 20775 3349
rect 21266 3340 21272 3352
rect 21324 3380 21330 3392
rect 21634 3380 21640 3392
rect 21324 3352 21640 3380
rect 21324 3340 21330 3352
rect 21634 3340 21640 3352
rect 21692 3340 21698 3392
rect 22462 3380 22468 3392
rect 22423 3352 22468 3380
rect 22462 3340 22468 3352
rect 22520 3340 22526 3392
rect 24210 3340 24216 3392
rect 24268 3380 24274 3392
rect 25682 3380 25688 3392
rect 24268 3352 25688 3380
rect 24268 3340 24274 3352
rect 25682 3340 25688 3352
rect 25740 3340 25746 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1397 3179 1455 3185
rect 1397 3145 1409 3179
rect 1443 3176 1455 3179
rect 2038 3176 2044 3188
rect 1443 3148 2044 3176
rect 1443 3145 1455 3148
rect 1397 3139 1455 3145
rect 2038 3136 2044 3148
rect 2096 3136 2102 3188
rect 3605 3179 3663 3185
rect 3605 3145 3617 3179
rect 3651 3176 3663 3179
rect 4338 3176 4344 3188
rect 3651 3148 4344 3176
rect 3651 3145 3663 3148
rect 3605 3139 3663 3145
rect 4338 3136 4344 3148
rect 4396 3136 4402 3188
rect 5166 3176 5172 3188
rect 5127 3148 5172 3176
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 5534 3136 5540 3188
rect 5592 3176 5598 3188
rect 6549 3179 6607 3185
rect 6549 3176 6561 3179
rect 5592 3148 6561 3176
rect 5592 3136 5598 3148
rect 6549 3145 6561 3148
rect 6595 3145 6607 3179
rect 6549 3139 6607 3145
rect 7101 3179 7159 3185
rect 7101 3145 7113 3179
rect 7147 3176 7159 3179
rect 7834 3176 7840 3188
rect 7147 3148 7840 3176
rect 7147 3145 7159 3148
rect 7101 3139 7159 3145
rect 1762 3068 1768 3120
rect 1820 3108 1826 3120
rect 2777 3111 2835 3117
rect 2777 3108 2789 3111
rect 1820 3080 2789 3108
rect 1820 3068 1826 3080
rect 2777 3077 2789 3080
rect 2823 3077 2835 3111
rect 2777 3071 2835 3077
rect 3418 3068 3424 3120
rect 3476 3108 3482 3120
rect 7116 3108 7144 3139
rect 7834 3136 7840 3148
rect 7892 3136 7898 3188
rect 8478 3136 8484 3188
rect 8536 3176 8542 3188
rect 8573 3179 8631 3185
rect 8573 3176 8585 3179
rect 8536 3148 8585 3176
rect 8536 3136 8542 3148
rect 8573 3145 8585 3148
rect 8619 3145 8631 3179
rect 8573 3139 8631 3145
rect 8662 3136 8668 3188
rect 8720 3176 8726 3188
rect 9585 3179 9643 3185
rect 9585 3176 9597 3179
rect 8720 3148 9597 3176
rect 8720 3136 8726 3148
rect 9585 3145 9597 3148
rect 9631 3176 9643 3179
rect 9950 3176 9956 3188
rect 9631 3148 9956 3176
rect 9631 3145 9643 3148
rect 9585 3139 9643 3145
rect 9950 3136 9956 3148
rect 10008 3136 10014 3188
rect 11054 3176 11060 3188
rect 11015 3148 11060 3176
rect 11054 3136 11060 3148
rect 11112 3136 11118 3188
rect 11606 3136 11612 3188
rect 11664 3176 11670 3188
rect 11977 3179 12035 3185
rect 11977 3176 11989 3179
rect 11664 3148 11989 3176
rect 11664 3136 11670 3148
rect 11977 3145 11989 3148
rect 12023 3145 12035 3179
rect 14366 3176 14372 3188
rect 11977 3139 12035 3145
rect 12452 3148 14372 3176
rect 9214 3108 9220 3120
rect 3476 3080 7144 3108
rect 9175 3080 9220 3108
rect 3476 3068 3482 3080
rect 9214 3068 9220 3080
rect 9272 3068 9278 3120
rect 11698 3108 11704 3120
rect 11611 3080 11704 3108
rect 11698 3068 11704 3080
rect 11756 3108 11762 3120
rect 12452 3108 12480 3148
rect 14366 3136 14372 3148
rect 14424 3136 14430 3188
rect 16574 3136 16580 3188
rect 16632 3176 16638 3188
rect 16850 3176 16856 3188
rect 16632 3148 16856 3176
rect 16632 3136 16638 3148
rect 16850 3136 16856 3148
rect 16908 3176 16914 3188
rect 17037 3179 17095 3185
rect 17037 3176 17049 3179
rect 16908 3148 17049 3176
rect 16908 3136 16914 3148
rect 17037 3145 17049 3148
rect 17083 3145 17095 3179
rect 18046 3176 18052 3188
rect 18007 3148 18052 3176
rect 17037 3139 17095 3145
rect 18046 3136 18052 3148
rect 18104 3136 18110 3188
rect 18782 3136 18788 3188
rect 18840 3176 18846 3188
rect 19061 3179 19119 3185
rect 19061 3176 19073 3179
rect 18840 3148 19073 3176
rect 18840 3136 18846 3148
rect 19061 3145 19073 3148
rect 19107 3145 19119 3179
rect 19061 3139 19119 3145
rect 19334 3136 19340 3188
rect 19392 3176 19398 3188
rect 19613 3179 19671 3185
rect 19613 3176 19625 3179
rect 19392 3148 19625 3176
rect 19392 3136 19398 3148
rect 19613 3145 19625 3148
rect 19659 3145 19671 3179
rect 19613 3139 19671 3145
rect 20717 3179 20775 3185
rect 20717 3145 20729 3179
rect 20763 3176 20775 3179
rect 20898 3176 20904 3188
rect 20763 3148 20904 3176
rect 20763 3145 20775 3148
rect 20717 3139 20775 3145
rect 20898 3136 20904 3148
rect 20956 3136 20962 3188
rect 21174 3176 21180 3188
rect 21135 3148 21180 3176
rect 21174 3136 21180 3148
rect 21232 3136 21238 3188
rect 22557 3179 22615 3185
rect 22557 3145 22569 3179
rect 22603 3176 22615 3179
rect 22830 3176 22836 3188
rect 22603 3148 22836 3176
rect 22603 3145 22615 3148
rect 22557 3139 22615 3145
rect 22830 3136 22836 3148
rect 22888 3136 22894 3188
rect 22925 3179 22983 3185
rect 22925 3145 22937 3179
rect 22971 3176 22983 3179
rect 23014 3176 23020 3188
rect 22971 3148 23020 3176
rect 22971 3145 22983 3148
rect 22925 3139 22983 3145
rect 23014 3136 23020 3148
rect 23072 3136 23078 3188
rect 23477 3179 23535 3185
rect 23477 3145 23489 3179
rect 23523 3176 23535 3179
rect 23750 3176 23756 3188
rect 23523 3148 23756 3176
rect 23523 3145 23535 3148
rect 23477 3139 23535 3145
rect 23750 3136 23756 3148
rect 23808 3136 23814 3188
rect 24765 3179 24823 3185
rect 24765 3145 24777 3179
rect 24811 3176 24823 3179
rect 24854 3176 24860 3188
rect 24811 3148 24860 3176
rect 24811 3145 24823 3148
rect 24765 3139 24823 3145
rect 24854 3136 24860 3148
rect 24912 3136 24918 3188
rect 25038 3176 25044 3188
rect 24999 3148 25044 3176
rect 25038 3136 25044 3148
rect 25096 3136 25102 3188
rect 26050 3176 26056 3188
rect 26011 3148 26056 3176
rect 26050 3136 26056 3148
rect 26108 3136 26114 3188
rect 26326 3176 26332 3188
rect 26287 3148 26332 3176
rect 26326 3136 26332 3148
rect 26384 3136 26390 3188
rect 11756 3080 12480 3108
rect 13817 3111 13875 3117
rect 11756 3068 11762 3080
rect 13817 3077 13829 3111
rect 13863 3108 13875 3111
rect 13906 3108 13912 3120
rect 13863 3080 13912 3108
rect 13863 3077 13875 3080
rect 13817 3071 13875 3077
rect 13906 3068 13912 3080
rect 13964 3068 13970 3120
rect 19444 3080 20208 3108
rect 2041 3043 2099 3049
rect 2041 3009 2053 3043
rect 2087 3040 2099 3043
rect 2130 3040 2136 3052
rect 2087 3012 2136 3040
rect 2087 3009 2099 3012
rect 2041 3003 2099 3009
rect 2130 3000 2136 3012
rect 2188 3000 2194 3052
rect 3510 3040 3516 3052
rect 3423 3012 3516 3040
rect 3510 3000 3516 3012
rect 3568 3040 3574 3052
rect 4154 3040 4160 3052
rect 3568 3012 4160 3040
rect 3568 3000 3574 3012
rect 4154 3000 4160 3012
rect 4212 3000 4218 3052
rect 5813 3043 5871 3049
rect 5813 3009 5825 3043
rect 5859 3040 5871 3043
rect 5859 3012 6316 3040
rect 5859 3009 5871 3012
rect 5813 3003 5871 3009
rect 2225 2975 2283 2981
rect 2225 2941 2237 2975
rect 2271 2972 2283 2975
rect 4246 2972 4252 2984
rect 2271 2944 4252 2972
rect 2271 2941 2283 2944
rect 2225 2935 2283 2941
rect 4246 2932 4252 2944
rect 4304 2932 4310 2984
rect 4709 2975 4767 2981
rect 4709 2941 4721 2975
rect 4755 2972 4767 2975
rect 5629 2975 5687 2981
rect 5629 2972 5641 2975
rect 4755 2944 5641 2972
rect 4755 2941 4767 2944
rect 4709 2935 4767 2941
rect 5629 2941 5641 2944
rect 5675 2972 5687 2975
rect 6086 2972 6092 2984
rect 5675 2944 6092 2972
rect 5675 2941 5687 2944
rect 5629 2935 5687 2941
rect 6086 2932 6092 2944
rect 6144 2932 6150 2984
rect 6288 2981 6316 3012
rect 7006 3000 7012 3052
rect 7064 3040 7070 3052
rect 7193 3043 7251 3049
rect 7193 3040 7205 3043
rect 7064 3012 7205 3040
rect 7064 3000 7070 3012
rect 7193 3009 7205 3012
rect 7239 3009 7251 3043
rect 7193 3003 7251 3009
rect 17126 3000 17132 3052
rect 17184 3040 17190 3052
rect 17405 3043 17463 3049
rect 17405 3040 17417 3043
rect 17184 3012 17417 3040
rect 17184 3000 17190 3012
rect 17405 3009 17417 3012
rect 17451 3009 17463 3043
rect 18601 3043 18659 3049
rect 18601 3040 18613 3043
rect 17405 3003 17463 3009
rect 17788 3012 18613 3040
rect 17788 2984 17816 3012
rect 18601 3009 18613 3012
rect 18647 3040 18659 3043
rect 18874 3040 18880 3052
rect 18647 3012 18880 3040
rect 18647 3009 18659 3012
rect 18601 3003 18659 3009
rect 18874 3000 18880 3012
rect 18932 3040 18938 3052
rect 19444 3049 19472 3080
rect 19429 3043 19487 3049
rect 19429 3040 19441 3043
rect 18932 3012 19441 3040
rect 18932 3000 18938 3012
rect 19429 3009 19441 3012
rect 19475 3009 19487 3043
rect 20070 3040 20076 3052
rect 20031 3012 20076 3040
rect 19429 3003 19487 3009
rect 20070 3000 20076 3012
rect 20128 3000 20134 3052
rect 20180 3049 20208 3080
rect 20254 3068 20260 3120
rect 20312 3108 20318 3120
rect 21726 3108 21732 3120
rect 20312 3080 21732 3108
rect 20312 3068 20318 3080
rect 21726 3068 21732 3080
rect 21784 3108 21790 3120
rect 23658 3108 23664 3120
rect 21784 3080 21864 3108
rect 23619 3080 23664 3108
rect 21784 3068 21790 3080
rect 21836 3049 21864 3080
rect 23658 3068 23664 3080
rect 23716 3068 23722 3120
rect 20165 3043 20223 3049
rect 20165 3009 20177 3043
rect 20211 3009 20223 3043
rect 20165 3003 20223 3009
rect 21821 3043 21879 3049
rect 21821 3009 21833 3043
rect 21867 3009 21879 3043
rect 21821 3003 21879 3009
rect 23106 3000 23112 3052
rect 23164 3040 23170 3052
rect 24305 3043 24363 3049
rect 24305 3040 24317 3043
rect 23164 3012 24317 3040
rect 23164 3000 23170 3012
rect 24305 3009 24317 3012
rect 24351 3040 24363 3043
rect 25056 3040 25084 3136
rect 24351 3012 25084 3040
rect 24351 3009 24363 3012
rect 24305 3003 24363 3009
rect 6273 2975 6331 2981
rect 6273 2941 6285 2975
rect 6319 2972 6331 2975
rect 9677 2975 9735 2981
rect 6319 2944 7503 2972
rect 6319 2941 6331 2944
rect 6273 2935 6331 2941
rect 7475 2916 7503 2944
rect 9677 2941 9689 2975
rect 9723 2972 9735 2975
rect 11974 2972 11980 2984
rect 9723 2944 11980 2972
rect 9723 2941 9735 2944
rect 9677 2935 9735 2941
rect 1762 2904 1768 2916
rect 1675 2876 1768 2904
rect 1762 2864 1768 2876
rect 1820 2904 1826 2916
rect 2501 2907 2559 2913
rect 2501 2904 2513 2907
rect 1820 2876 2513 2904
rect 1820 2864 1826 2876
rect 2501 2873 2513 2876
rect 2547 2904 2559 2907
rect 2774 2904 2780 2916
rect 2547 2876 2780 2904
rect 2547 2873 2559 2876
rect 2501 2867 2559 2873
rect 2774 2864 2780 2876
rect 2832 2864 2838 2916
rect 3970 2904 3976 2916
rect 3931 2876 3976 2904
rect 3970 2864 3976 2876
rect 4028 2864 4034 2916
rect 7466 2913 7472 2916
rect 5077 2907 5135 2913
rect 5077 2873 5089 2907
rect 5123 2904 5135 2907
rect 5537 2907 5595 2913
rect 5537 2904 5549 2907
rect 5123 2876 5549 2904
rect 5123 2873 5135 2876
rect 5077 2867 5135 2873
rect 5537 2873 5549 2876
rect 5583 2904 5595 2907
rect 5583 2876 6224 2904
rect 5583 2873 5595 2876
rect 5537 2867 5595 2873
rect 1670 2796 1676 2848
rect 1728 2836 1734 2848
rect 1857 2839 1915 2845
rect 1857 2836 1869 2839
rect 1728 2808 1869 2836
rect 1728 2796 1734 2808
rect 1857 2805 1869 2808
rect 1903 2836 1915 2839
rect 2225 2839 2283 2845
rect 2225 2836 2237 2839
rect 1903 2808 2237 2836
rect 1903 2805 1915 2808
rect 1857 2799 1915 2805
rect 2225 2805 2237 2808
rect 2271 2805 2283 2839
rect 2225 2799 2283 2805
rect 4065 2839 4123 2845
rect 4065 2805 4077 2839
rect 4111 2836 4123 2839
rect 4246 2836 4252 2848
rect 4111 2808 4252 2836
rect 4111 2805 4123 2808
rect 4065 2799 4123 2805
rect 4246 2796 4252 2808
rect 4304 2796 4310 2848
rect 6196 2836 6224 2876
rect 7460 2867 7472 2913
rect 7524 2904 7530 2916
rect 7926 2904 7932 2916
rect 7524 2876 7932 2904
rect 7466 2864 7472 2867
rect 7524 2864 7530 2876
rect 7926 2864 7932 2876
rect 7984 2864 7990 2916
rect 9692 2848 9720 2935
rect 11974 2932 11980 2944
rect 12032 2972 12038 2984
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 12032 2944 12449 2972
rect 12032 2932 12038 2944
rect 12437 2941 12449 2944
rect 12483 2941 12495 2975
rect 15102 2972 15108 2984
rect 15063 2944 15108 2972
rect 12437 2935 12495 2941
rect 15102 2932 15108 2944
rect 15160 2932 15166 2984
rect 17770 2972 17776 2984
rect 17731 2944 17776 2972
rect 17770 2932 17776 2944
rect 17828 2932 17834 2984
rect 17954 2932 17960 2984
rect 18012 2972 18018 2984
rect 18414 2972 18420 2984
rect 18012 2944 18420 2972
rect 18012 2932 18018 2944
rect 18414 2932 18420 2944
rect 18472 2932 18478 2984
rect 18509 2975 18567 2981
rect 18509 2941 18521 2975
rect 18555 2972 18567 2975
rect 18690 2972 18696 2984
rect 18555 2944 18696 2972
rect 18555 2941 18567 2944
rect 18509 2935 18567 2941
rect 18690 2932 18696 2944
rect 18748 2932 18754 2984
rect 20898 2932 20904 2984
rect 20956 2972 20962 2984
rect 21545 2975 21603 2981
rect 21545 2972 21557 2975
rect 20956 2944 21557 2972
rect 20956 2932 20962 2944
rect 21545 2941 21557 2944
rect 21591 2941 21603 2975
rect 21545 2935 21603 2941
rect 23842 2932 23848 2984
rect 23900 2972 23906 2984
rect 24118 2972 24124 2984
rect 23900 2944 23980 2972
rect 24079 2944 24124 2972
rect 23900 2932 23906 2944
rect 9858 2864 9864 2916
rect 9916 2913 9922 2916
rect 9916 2907 9980 2913
rect 9916 2873 9934 2907
rect 9968 2904 9980 2907
rect 11054 2904 11060 2916
rect 9968 2876 11060 2904
rect 9968 2873 9980 2876
rect 9916 2867 9980 2873
rect 9916 2864 9922 2867
rect 11054 2864 11060 2876
rect 11112 2864 11118 2916
rect 12710 2913 12716 2916
rect 12704 2867 12716 2913
rect 12768 2904 12774 2916
rect 15378 2913 15384 2916
rect 14645 2907 14703 2913
rect 12768 2876 12804 2904
rect 12710 2864 12716 2867
rect 12768 2864 12774 2876
rect 14645 2873 14657 2907
rect 14691 2904 14703 2907
rect 15350 2907 15384 2913
rect 15350 2904 15362 2907
rect 14691 2876 15362 2904
rect 14691 2873 14703 2876
rect 14645 2867 14703 2873
rect 15350 2873 15362 2876
rect 15436 2904 15442 2916
rect 15436 2876 15498 2904
rect 15350 2867 15384 2873
rect 15378 2864 15384 2867
rect 15436 2864 15442 2876
rect 15838 2864 15844 2916
rect 15896 2864 15902 2916
rect 19981 2907 20039 2913
rect 19981 2873 19993 2907
rect 20027 2904 20039 2907
rect 20714 2904 20720 2916
rect 20027 2876 20720 2904
rect 20027 2873 20039 2876
rect 19981 2867 20039 2873
rect 20714 2864 20720 2876
rect 20772 2864 20778 2916
rect 20990 2864 20996 2916
rect 21048 2904 21054 2916
rect 21085 2907 21143 2913
rect 21085 2904 21097 2907
rect 21048 2876 21097 2904
rect 21048 2864 21054 2876
rect 21085 2873 21097 2876
rect 21131 2904 21143 2907
rect 21637 2907 21695 2913
rect 21637 2904 21649 2907
rect 21131 2876 21649 2904
rect 21131 2873 21143 2876
rect 21085 2867 21143 2873
rect 21637 2873 21649 2876
rect 21683 2873 21695 2907
rect 21637 2867 21695 2873
rect 23474 2864 23480 2916
rect 23532 2904 23538 2916
rect 23952 2904 23980 2944
rect 24118 2932 24124 2944
rect 24176 2932 24182 2984
rect 25225 2975 25283 2981
rect 25225 2941 25237 2975
rect 25271 2972 25283 2975
rect 26050 2972 26056 2984
rect 25271 2944 26056 2972
rect 25271 2941 25283 2944
rect 25225 2935 25283 2941
rect 26050 2932 26056 2944
rect 26108 2932 26114 2984
rect 24029 2907 24087 2913
rect 24029 2904 24041 2907
rect 23532 2876 23888 2904
rect 23952 2876 24041 2904
rect 23532 2864 23538 2876
rect 6454 2836 6460 2848
rect 6196 2808 6460 2836
rect 6454 2796 6460 2808
rect 6512 2796 6518 2848
rect 9674 2796 9680 2848
rect 9732 2796 9738 2848
rect 13906 2796 13912 2848
rect 13964 2836 13970 2848
rect 14274 2836 14280 2848
rect 13964 2808 14280 2836
rect 13964 2796 13970 2808
rect 14274 2796 14280 2808
rect 14332 2796 14338 2848
rect 14918 2836 14924 2848
rect 14879 2808 14924 2836
rect 14918 2796 14924 2808
rect 14976 2836 14982 2848
rect 15856 2836 15884 2864
rect 23860 2848 23888 2876
rect 24029 2873 24041 2876
rect 24075 2873 24087 2907
rect 25498 2904 25504 2916
rect 25459 2876 25504 2904
rect 24029 2867 24087 2873
rect 25498 2864 25504 2876
rect 25556 2864 25562 2916
rect 16485 2839 16543 2845
rect 16485 2836 16497 2839
rect 14976 2808 16497 2836
rect 14976 2796 14982 2808
rect 16485 2805 16497 2808
rect 16531 2805 16543 2839
rect 16485 2799 16543 2805
rect 23842 2796 23848 2848
rect 23900 2796 23906 2848
rect 24854 2796 24860 2848
rect 24912 2836 24918 2848
rect 25038 2836 25044 2848
rect 24912 2808 25044 2836
rect 24912 2796 24918 2808
rect 25038 2796 25044 2808
rect 25096 2796 25102 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1578 2592 1584 2644
rect 1636 2632 1642 2644
rect 1949 2635 2007 2641
rect 1949 2632 1961 2635
rect 1636 2604 1961 2632
rect 1636 2592 1642 2604
rect 1949 2601 1961 2604
rect 1995 2601 2007 2635
rect 1949 2595 2007 2601
rect 2777 2635 2835 2641
rect 2777 2601 2789 2635
rect 2823 2632 2835 2635
rect 3326 2632 3332 2644
rect 2823 2604 3332 2632
rect 2823 2601 2835 2604
rect 2777 2595 2835 2601
rect 3326 2592 3332 2604
rect 3384 2592 3390 2644
rect 3510 2632 3516 2644
rect 3471 2604 3516 2632
rect 3510 2592 3516 2604
rect 3568 2592 3574 2644
rect 5258 2592 5264 2644
rect 5316 2632 5322 2644
rect 6273 2635 6331 2641
rect 6273 2632 6285 2635
rect 5316 2604 6285 2632
rect 5316 2592 5322 2604
rect 6273 2601 6285 2604
rect 6319 2601 6331 2635
rect 6273 2595 6331 2601
rect 7926 2592 7932 2644
rect 7984 2632 7990 2644
rect 8573 2635 8631 2641
rect 8573 2632 8585 2635
rect 7984 2604 8585 2632
rect 7984 2592 7990 2604
rect 8573 2601 8585 2604
rect 8619 2601 8631 2635
rect 9582 2632 9588 2644
rect 9543 2604 9588 2632
rect 8573 2595 8631 2601
rect 9582 2592 9588 2604
rect 9640 2592 9646 2644
rect 11054 2592 11060 2644
rect 11112 2632 11118 2644
rect 11425 2635 11483 2641
rect 11425 2632 11437 2635
rect 11112 2604 11437 2632
rect 11112 2592 11118 2604
rect 11425 2601 11437 2604
rect 11471 2632 11483 2635
rect 12342 2632 12348 2644
rect 11471 2604 12348 2632
rect 11471 2601 11483 2604
rect 11425 2595 11483 2601
rect 12342 2592 12348 2604
rect 12400 2592 12406 2644
rect 14829 2635 14887 2641
rect 14829 2601 14841 2635
rect 14875 2632 14887 2635
rect 15470 2632 15476 2644
rect 14875 2604 15148 2632
rect 15431 2604 15476 2632
rect 14875 2601 14887 2604
rect 14829 2595 14887 2601
rect 1670 2564 1676 2576
rect 1631 2536 1676 2564
rect 1670 2524 1676 2536
rect 1728 2524 1734 2576
rect 4706 2564 4712 2576
rect 4356 2536 4712 2564
rect 4356 2505 4384 2536
rect 4706 2524 4712 2536
rect 4764 2564 4770 2576
rect 7466 2573 7472 2576
rect 6733 2567 6791 2573
rect 4764 2536 5212 2564
rect 4764 2524 4770 2536
rect 4341 2499 4399 2505
rect 4341 2465 4353 2499
rect 4387 2465 4399 2499
rect 4608 2499 4666 2505
rect 4608 2496 4620 2499
rect 4341 2459 4399 2465
rect 4448 2468 4620 2496
rect 2866 2428 2872 2440
rect 2827 2400 2872 2428
rect 2866 2388 2872 2400
rect 2924 2388 2930 2440
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2428 3111 2431
rect 3510 2428 3516 2440
rect 3099 2400 3516 2428
rect 3099 2397 3111 2400
rect 3053 2391 3111 2397
rect 3510 2388 3516 2400
rect 3568 2388 3574 2440
rect 3881 2431 3939 2437
rect 3881 2397 3893 2431
rect 3927 2428 3939 2431
rect 4448 2428 4476 2468
rect 4608 2465 4620 2468
rect 4654 2496 4666 2499
rect 5074 2496 5080 2508
rect 4654 2468 5080 2496
rect 4654 2465 4666 2468
rect 4608 2459 4666 2465
rect 5074 2456 5080 2468
rect 5132 2456 5138 2508
rect 5184 2496 5212 2536
rect 6733 2533 6745 2567
rect 6779 2564 6791 2567
rect 7460 2564 7472 2573
rect 6779 2536 7472 2564
rect 6779 2533 6791 2536
rect 6733 2527 6791 2533
rect 7460 2527 7472 2536
rect 7466 2524 7472 2527
rect 7524 2524 7530 2576
rect 9217 2567 9275 2573
rect 9217 2533 9229 2567
rect 9263 2564 9275 2567
rect 10312 2567 10370 2573
rect 10312 2564 10324 2567
rect 9263 2536 10324 2564
rect 9263 2533 9275 2536
rect 9217 2527 9275 2533
rect 10312 2533 10324 2536
rect 10358 2564 10370 2567
rect 10778 2564 10784 2576
rect 10358 2536 10784 2564
rect 10358 2533 10370 2536
rect 10312 2527 10370 2533
rect 10778 2524 10784 2536
rect 10836 2524 10842 2576
rect 10870 2524 10876 2576
rect 10928 2564 10934 2576
rect 11698 2564 11704 2576
rect 10928 2536 11704 2564
rect 10928 2524 10934 2536
rect 11698 2524 11704 2536
rect 11756 2524 11762 2576
rect 12437 2567 12495 2573
rect 12437 2533 12449 2567
rect 12483 2564 12495 2567
rect 13142 2567 13200 2573
rect 13142 2564 13154 2567
rect 12483 2536 13154 2564
rect 12483 2533 12495 2536
rect 12437 2527 12495 2533
rect 13142 2533 13154 2536
rect 13188 2564 13200 2567
rect 14918 2564 14924 2576
rect 13188 2536 14924 2564
rect 13188 2533 13200 2536
rect 13142 2527 13200 2533
rect 14918 2524 14924 2536
rect 14976 2524 14982 2576
rect 15120 2564 15148 2604
rect 15470 2592 15476 2604
rect 15528 2592 15534 2644
rect 15933 2635 15991 2641
rect 15933 2601 15945 2635
rect 15979 2632 15991 2635
rect 17034 2632 17040 2644
rect 15979 2604 17040 2632
rect 15979 2601 15991 2604
rect 15933 2595 15991 2601
rect 15948 2564 15976 2595
rect 17034 2592 17040 2604
rect 17092 2592 17098 2644
rect 18322 2632 18328 2644
rect 18283 2604 18328 2632
rect 18322 2592 18328 2604
rect 18380 2592 18386 2644
rect 18785 2635 18843 2641
rect 18785 2601 18797 2635
rect 18831 2632 18843 2635
rect 20806 2632 20812 2644
rect 18831 2604 20812 2632
rect 18831 2601 18843 2604
rect 18785 2595 18843 2601
rect 15120 2536 15976 2564
rect 18141 2567 18199 2573
rect 18141 2533 18153 2567
rect 18187 2564 18199 2567
rect 18800 2564 18828 2595
rect 20806 2592 20812 2604
rect 20864 2592 20870 2644
rect 21174 2632 21180 2644
rect 21135 2604 21180 2632
rect 21174 2592 21180 2604
rect 21232 2592 21238 2644
rect 23014 2632 23020 2644
rect 22975 2604 23020 2632
rect 23014 2592 23020 2604
rect 23072 2592 23078 2644
rect 24029 2635 24087 2641
rect 24029 2601 24041 2635
rect 24075 2632 24087 2635
rect 24762 2632 24768 2644
rect 24075 2604 24768 2632
rect 24075 2601 24087 2604
rect 24029 2595 24087 2601
rect 24762 2592 24768 2604
rect 24820 2592 24826 2644
rect 25038 2632 25044 2644
rect 24999 2604 25044 2632
rect 25038 2592 25044 2604
rect 25096 2592 25102 2644
rect 26326 2592 26332 2644
rect 26384 2632 26390 2644
rect 26421 2635 26479 2641
rect 26421 2632 26433 2635
rect 26384 2604 26433 2632
rect 26384 2592 26390 2604
rect 26421 2601 26433 2604
rect 26467 2601 26479 2635
rect 26421 2595 26479 2601
rect 18187 2536 18828 2564
rect 18187 2533 18199 2536
rect 18141 2527 18199 2533
rect 19426 2524 19432 2576
rect 19484 2564 19490 2576
rect 19886 2564 19892 2576
rect 19484 2536 19892 2564
rect 19484 2524 19490 2536
rect 19886 2524 19892 2536
rect 19944 2524 19950 2576
rect 20898 2524 20904 2576
rect 20956 2564 20962 2576
rect 21637 2567 21695 2573
rect 21637 2564 21649 2567
rect 20956 2536 21649 2564
rect 20956 2524 20962 2536
rect 21637 2533 21649 2536
rect 21683 2533 21695 2567
rect 21637 2527 21695 2533
rect 23845 2567 23903 2573
rect 23845 2533 23857 2567
rect 23891 2564 23903 2567
rect 24118 2564 24124 2576
rect 23891 2536 24124 2564
rect 23891 2533 23903 2536
rect 23845 2527 23903 2533
rect 24118 2524 24124 2536
rect 24176 2524 24182 2576
rect 24486 2564 24492 2576
rect 24447 2536 24492 2564
rect 24486 2524 24492 2536
rect 24544 2564 24550 2576
rect 25409 2567 25467 2573
rect 25409 2564 25421 2567
rect 24544 2536 25421 2564
rect 24544 2524 24550 2536
rect 25409 2533 25421 2536
rect 25455 2533 25467 2567
rect 25590 2564 25596 2576
rect 25551 2536 25596 2564
rect 25409 2527 25467 2533
rect 25590 2524 25596 2536
rect 25648 2524 25654 2576
rect 7006 2496 7012 2508
rect 5184 2468 7012 2496
rect 7006 2456 7012 2468
rect 7064 2496 7070 2508
rect 7193 2499 7251 2505
rect 7193 2496 7205 2499
rect 7064 2468 7205 2496
rect 7064 2456 7070 2468
rect 7193 2465 7205 2468
rect 7239 2465 7251 2499
rect 7193 2459 7251 2465
rect 9030 2456 9036 2508
rect 9088 2496 9094 2508
rect 9490 2496 9496 2508
rect 9088 2468 9496 2496
rect 9088 2456 9094 2468
rect 9490 2456 9496 2468
rect 9548 2456 9554 2508
rect 9674 2456 9680 2508
rect 9732 2496 9738 2508
rect 10045 2499 10103 2505
rect 10045 2496 10057 2499
rect 9732 2468 10057 2496
rect 9732 2456 9738 2468
rect 10045 2465 10057 2468
rect 10091 2465 10103 2499
rect 10045 2459 10103 2465
rect 12897 2499 12955 2505
rect 12897 2465 12909 2499
rect 12943 2496 12955 2499
rect 15102 2496 15108 2508
rect 12943 2468 15108 2496
rect 12943 2465 12955 2468
rect 12897 2459 12955 2465
rect 15102 2456 15108 2468
rect 15160 2456 15166 2508
rect 15841 2499 15899 2505
rect 15841 2465 15853 2499
rect 15887 2496 15899 2499
rect 15887 2468 16620 2496
rect 15887 2465 15899 2468
rect 15841 2459 15899 2465
rect 12066 2428 12072 2440
rect 3927 2400 4476 2428
rect 12027 2400 12072 2428
rect 3927 2397 3939 2400
rect 3881 2391 3939 2397
rect 12066 2388 12072 2400
rect 12124 2388 12130 2440
rect 16117 2431 16175 2437
rect 16117 2397 16129 2431
rect 16163 2428 16175 2431
rect 16482 2428 16488 2440
rect 16163 2400 16488 2428
rect 16163 2397 16175 2400
rect 16117 2391 16175 2397
rect 2406 2360 2412 2372
rect 2367 2332 2412 2360
rect 2406 2320 2412 2332
rect 2464 2320 2470 2372
rect 14274 2360 14280 2372
rect 14235 2332 14280 2360
rect 14274 2320 14280 2332
rect 14332 2320 14338 2372
rect 15289 2363 15347 2369
rect 15289 2329 15301 2363
rect 15335 2360 15347 2363
rect 15378 2360 15384 2372
rect 15335 2332 15384 2360
rect 15335 2329 15347 2332
rect 15289 2323 15347 2329
rect 15378 2320 15384 2332
rect 15436 2360 15442 2372
rect 16132 2360 16160 2391
rect 16482 2388 16488 2400
rect 16540 2388 16546 2440
rect 15436 2332 16160 2360
rect 15436 2320 15442 2332
rect 5721 2295 5779 2301
rect 5721 2261 5733 2295
rect 5767 2292 5779 2295
rect 6546 2292 6552 2304
rect 5767 2264 6552 2292
rect 5767 2261 5779 2264
rect 5721 2255 5779 2261
rect 6546 2252 6552 2264
rect 6604 2252 6610 2304
rect 15470 2252 15476 2304
rect 15528 2292 15534 2304
rect 16114 2292 16120 2304
rect 15528 2264 16120 2292
rect 15528 2252 15534 2264
rect 16114 2252 16120 2264
rect 16172 2252 16178 2304
rect 16592 2301 16620 2468
rect 16942 2456 16948 2508
rect 17000 2496 17006 2508
rect 17037 2499 17095 2505
rect 17037 2496 17049 2499
rect 17000 2468 17049 2496
rect 17000 2456 17006 2468
rect 17037 2465 17049 2468
rect 17083 2465 17095 2499
rect 18693 2499 18751 2505
rect 18693 2496 18705 2499
rect 17037 2459 17095 2465
rect 17696 2468 18705 2496
rect 16577 2295 16635 2301
rect 16577 2261 16589 2295
rect 16623 2292 16635 2295
rect 16666 2292 16672 2304
rect 16623 2264 16672 2292
rect 16623 2261 16635 2264
rect 16577 2255 16635 2261
rect 16666 2252 16672 2264
rect 16724 2252 16730 2304
rect 16942 2292 16948 2304
rect 16903 2264 16948 2292
rect 16942 2252 16948 2264
rect 17000 2252 17006 2304
rect 17126 2252 17132 2304
rect 17184 2292 17190 2304
rect 17221 2295 17279 2301
rect 17221 2292 17233 2295
rect 17184 2264 17233 2292
rect 17184 2252 17190 2264
rect 17221 2261 17233 2264
rect 17267 2261 17279 2295
rect 17221 2255 17279 2261
rect 17586 2252 17592 2304
rect 17644 2292 17650 2304
rect 17696 2301 17724 2468
rect 18693 2465 18705 2468
rect 18739 2465 18751 2499
rect 18693 2459 18751 2465
rect 19794 2456 19800 2508
rect 19852 2496 19858 2508
rect 19981 2499 20039 2505
rect 19981 2496 19993 2499
rect 19852 2468 19993 2496
rect 19852 2456 19858 2468
rect 19981 2465 19993 2468
rect 20027 2465 20039 2499
rect 19981 2459 20039 2465
rect 21545 2499 21603 2505
rect 21545 2465 21557 2499
rect 21591 2465 21603 2499
rect 21545 2459 21603 2465
rect 22833 2499 22891 2505
rect 22833 2465 22845 2499
rect 22879 2496 22891 2499
rect 22922 2496 22928 2508
rect 22879 2468 22928 2496
rect 22879 2465 22891 2468
rect 22833 2459 22891 2465
rect 18874 2388 18880 2440
rect 18932 2428 18938 2440
rect 19337 2431 19395 2437
rect 19337 2428 19349 2431
rect 18932 2400 19349 2428
rect 18932 2388 18938 2400
rect 19337 2397 19349 2400
rect 19383 2397 19395 2431
rect 20530 2428 20536 2440
rect 20491 2400 20536 2428
rect 19337 2391 19395 2397
rect 20530 2388 20536 2400
rect 20588 2428 20594 2440
rect 21560 2428 21588 2459
rect 22922 2456 22928 2468
rect 22980 2496 22986 2508
rect 23385 2499 23443 2505
rect 23385 2496 23397 2499
rect 22980 2468 23397 2496
rect 22980 2456 22986 2468
rect 23385 2465 23397 2468
rect 23431 2465 23443 2499
rect 23385 2459 23443 2465
rect 24210 2456 24216 2508
rect 24268 2496 24274 2508
rect 24397 2499 24455 2505
rect 24397 2496 24409 2499
rect 24268 2468 24409 2496
rect 24268 2456 24274 2468
rect 24397 2465 24409 2468
rect 24443 2496 24455 2499
rect 26053 2499 26111 2505
rect 26053 2496 26065 2499
rect 24443 2468 26065 2496
rect 24443 2465 24455 2468
rect 24397 2459 24455 2465
rect 26053 2465 26065 2468
rect 26099 2465 26111 2499
rect 26053 2459 26111 2465
rect 21726 2428 21732 2440
rect 20588 2400 21588 2428
rect 21687 2400 21732 2428
rect 20588 2388 20594 2400
rect 21726 2388 21732 2400
rect 21784 2428 21790 2440
rect 22189 2431 22247 2437
rect 22189 2428 22201 2431
rect 21784 2400 22201 2428
rect 21784 2388 21790 2400
rect 22189 2397 22201 2400
rect 22235 2428 22247 2431
rect 22557 2431 22615 2437
rect 22557 2428 22569 2431
rect 22235 2400 22569 2428
rect 22235 2397 22247 2400
rect 22189 2391 22247 2397
rect 22557 2397 22569 2400
rect 22603 2397 22615 2431
rect 22557 2391 22615 2397
rect 24673 2431 24731 2437
rect 24673 2397 24685 2431
rect 24719 2428 24731 2431
rect 25038 2428 25044 2440
rect 24719 2400 25044 2428
rect 24719 2397 24731 2400
rect 24673 2391 24731 2397
rect 25038 2388 25044 2400
rect 25096 2388 25102 2440
rect 17681 2295 17739 2301
rect 17681 2292 17693 2295
rect 17644 2264 17693 2292
rect 17644 2252 17650 2264
rect 17681 2261 17693 2264
rect 17727 2261 17739 2295
rect 19794 2292 19800 2304
rect 19755 2264 19800 2292
rect 17681 2255 17739 2261
rect 19794 2252 19800 2264
rect 19852 2252 19858 2304
rect 20162 2292 20168 2304
rect 20123 2264 20168 2292
rect 20162 2252 20168 2264
rect 20220 2252 20226 2304
rect 20898 2292 20904 2304
rect 20859 2264 20904 2292
rect 20898 2252 20904 2264
rect 20956 2252 20962 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 7742 552 7748 604
rect 7800 592 7806 604
rect 7834 592 7840 604
rect 7800 564 7840 592
rect 7800 552 7806 564
rect 7834 552 7840 564
rect 7892 552 7898 604
rect 11882 552 11888 604
rect 11940 592 11946 604
rect 12250 592 12256 604
rect 11940 564 12256 592
rect 11940 552 11946 564
rect 12250 552 12256 564
rect 12308 552 12314 604
<< via1 >>
rect 2872 27412 2924 27464
rect 3792 27412 3844 27464
rect 21088 26800 21140 26852
rect 24676 26800 24728 26852
rect 20076 26392 20128 26444
rect 24768 26392 24820 26444
rect 11888 26324 11940 26376
rect 17960 26324 18012 26376
rect 8300 26188 8352 26240
rect 18236 26188 18288 26240
rect 7748 26120 7800 26172
rect 17132 26120 17184 26172
rect 8760 26052 8812 26104
rect 18328 26052 18380 26104
rect 7840 25984 7892 26036
rect 13084 25984 13136 26036
rect 13176 25984 13228 26036
rect 24676 25984 24728 26036
rect 8944 25916 8996 25968
rect 16580 25916 16632 25968
rect 17224 25916 17276 25968
rect 22376 25916 22428 25968
rect 6368 25848 6420 25900
rect 17776 25848 17828 25900
rect 8852 25780 8904 25832
rect 19524 25780 19576 25832
rect 22468 25780 22520 25832
rect 26516 25780 26568 25832
rect 7472 25712 7524 25764
rect 18880 25712 18932 25764
rect 18972 25712 19024 25764
rect 25872 25712 25924 25764
rect 9128 25644 9180 25696
rect 21272 25644 21324 25696
rect 22192 25644 22244 25696
rect 24768 25644 24820 25696
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 8944 25440 8996 25492
rect 17224 25440 17276 25492
rect 19984 25440 20036 25492
rect 14648 25372 14700 25424
rect 15660 25372 15712 25424
rect 15936 25372 15988 25424
rect 24768 25440 24820 25492
rect 24584 25372 24636 25424
rect 1400 25347 1452 25356
rect 1400 25313 1409 25347
rect 1409 25313 1443 25347
rect 1443 25313 1452 25347
rect 1400 25304 1452 25313
rect 8668 25304 8720 25356
rect 9312 25304 9364 25356
rect 9588 25304 9640 25356
rect 10968 25347 11020 25356
rect 10968 25313 10977 25347
rect 10977 25313 11011 25347
rect 11011 25313 11020 25347
rect 10968 25304 11020 25313
rect 11612 25304 11664 25356
rect 11796 25304 11848 25356
rect 12992 25347 13044 25356
rect 12992 25313 13001 25347
rect 13001 25313 13035 25347
rect 13035 25313 13044 25347
rect 12992 25304 13044 25313
rect 13912 25304 13964 25356
rect 15752 25304 15804 25356
rect 17132 25347 17184 25356
rect 13820 25236 13872 25288
rect 15936 25279 15988 25288
rect 15936 25245 15945 25279
rect 15945 25245 15979 25279
rect 15979 25245 15988 25279
rect 16120 25279 16172 25288
rect 15936 25236 15988 25245
rect 16120 25245 16129 25279
rect 16129 25245 16163 25279
rect 16163 25245 16172 25279
rect 16120 25236 16172 25245
rect 16488 25236 16540 25288
rect 17132 25313 17141 25347
rect 17141 25313 17175 25347
rect 17175 25313 17184 25347
rect 17132 25304 17184 25313
rect 18880 25347 18932 25356
rect 18880 25313 18889 25347
rect 18889 25313 18923 25347
rect 18923 25313 18932 25347
rect 18880 25304 18932 25313
rect 20628 25304 20680 25356
rect 21180 25304 21232 25356
rect 22744 25347 22796 25356
rect 22744 25313 22753 25347
rect 22753 25313 22787 25347
rect 22787 25313 22796 25347
rect 22744 25304 22796 25313
rect 22928 25304 22980 25356
rect 24032 25304 24084 25356
rect 7104 25168 7156 25220
rect 9772 25168 9824 25220
rect 11796 25168 11848 25220
rect 2780 25100 2832 25152
rect 7380 25100 7432 25152
rect 13176 25143 13228 25152
rect 13176 25109 13185 25143
rect 13185 25109 13219 25143
rect 13219 25109 13228 25143
rect 13544 25143 13596 25152
rect 13176 25100 13228 25109
rect 13544 25109 13553 25143
rect 13553 25109 13587 25143
rect 13587 25109 13596 25143
rect 13544 25100 13596 25109
rect 13912 25143 13964 25152
rect 13912 25109 13921 25143
rect 13921 25109 13955 25143
rect 13955 25109 13964 25143
rect 13912 25100 13964 25109
rect 14740 25100 14792 25152
rect 15292 25143 15344 25152
rect 15292 25109 15301 25143
rect 15301 25109 15335 25143
rect 15335 25109 15344 25143
rect 15292 25100 15344 25109
rect 15476 25143 15528 25152
rect 15476 25109 15485 25143
rect 15485 25109 15519 25143
rect 15519 25109 15528 25143
rect 15476 25100 15528 25109
rect 17224 25168 17276 25220
rect 22468 25236 22520 25288
rect 23020 25279 23072 25288
rect 23020 25245 23029 25279
rect 23029 25245 23063 25279
rect 23063 25245 23072 25279
rect 23020 25236 23072 25245
rect 23572 25236 23624 25288
rect 16764 25100 16816 25152
rect 16856 25100 16908 25152
rect 18972 25168 19024 25220
rect 21824 25168 21876 25220
rect 25044 25211 25096 25220
rect 25044 25177 25053 25211
rect 25053 25177 25087 25211
rect 25087 25177 25096 25211
rect 25044 25168 25096 25177
rect 18052 25143 18104 25152
rect 18052 25109 18061 25143
rect 18061 25109 18095 25143
rect 18095 25109 18104 25143
rect 18052 25100 18104 25109
rect 20996 25143 21048 25152
rect 20996 25109 21005 25143
rect 21005 25109 21039 25143
rect 21039 25109 21048 25143
rect 20996 25100 21048 25109
rect 23480 25100 23532 25152
rect 24124 25100 24176 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 1584 24939 1636 24948
rect 1584 24905 1593 24939
rect 1593 24905 1627 24939
rect 1627 24905 1636 24939
rect 1584 24896 1636 24905
rect 7104 24939 7156 24948
rect 7104 24905 7113 24939
rect 7113 24905 7147 24939
rect 7147 24905 7156 24939
rect 7104 24896 7156 24905
rect 7656 24939 7708 24948
rect 7656 24905 7665 24939
rect 7665 24905 7699 24939
rect 7699 24905 7708 24939
rect 7656 24896 7708 24905
rect 8760 24939 8812 24948
rect 8760 24905 8769 24939
rect 8769 24905 8803 24939
rect 8803 24905 8812 24939
rect 8760 24896 8812 24905
rect 9312 24896 9364 24948
rect 13912 24896 13964 24948
rect 14648 24896 14700 24948
rect 8668 24828 8720 24880
rect 9956 24828 10008 24880
rect 10692 24828 10744 24880
rect 14924 24828 14976 24880
rect 16856 24896 16908 24948
rect 17224 24896 17276 24948
rect 22652 24896 22704 24948
rect 22928 24896 22980 24948
rect 9496 24760 9548 24812
rect 11428 24803 11480 24812
rect 7564 24692 7616 24744
rect 8760 24692 8812 24744
rect 11152 24735 11204 24744
rect 11152 24701 11161 24735
rect 11161 24701 11195 24735
rect 11195 24701 11204 24735
rect 11152 24692 11204 24701
rect 11428 24769 11437 24803
rect 11437 24769 11471 24803
rect 11471 24769 11480 24803
rect 11428 24760 11480 24769
rect 11612 24760 11664 24812
rect 11980 24760 12032 24812
rect 13636 24803 13688 24812
rect 13636 24769 13645 24803
rect 13645 24769 13679 24803
rect 13679 24769 13688 24803
rect 13636 24760 13688 24769
rect 15476 24828 15528 24880
rect 16304 24828 16356 24880
rect 18052 24828 18104 24880
rect 19984 24828 20036 24880
rect 22192 24828 22244 24880
rect 16856 24803 16908 24812
rect 16856 24769 16865 24803
rect 16865 24769 16899 24803
rect 16899 24769 16908 24803
rect 16856 24760 16908 24769
rect 17132 24760 17184 24812
rect 12256 24692 12308 24744
rect 13084 24692 13136 24744
rect 13544 24692 13596 24744
rect 15108 24735 15160 24744
rect 15108 24701 15117 24735
rect 15117 24701 15151 24735
rect 15151 24701 15160 24735
rect 15108 24692 15160 24701
rect 15752 24692 15804 24744
rect 15936 24692 15988 24744
rect 18236 24803 18288 24812
rect 18236 24769 18245 24803
rect 18245 24769 18279 24803
rect 18279 24769 18288 24803
rect 18236 24760 18288 24769
rect 21180 24760 21232 24812
rect 22468 24803 22520 24812
rect 22468 24769 22477 24803
rect 22477 24769 22511 24803
rect 22511 24769 22520 24803
rect 22468 24760 22520 24769
rect 22652 24803 22704 24812
rect 22652 24769 22661 24803
rect 22661 24769 22695 24803
rect 22695 24769 22704 24803
rect 22652 24760 22704 24769
rect 23020 24760 23072 24812
rect 25044 24803 25096 24812
rect 25044 24769 25053 24803
rect 25053 24769 25087 24803
rect 25087 24769 25096 24803
rect 25044 24760 25096 24769
rect 13268 24624 13320 24676
rect 16028 24624 16080 24676
rect 1400 24556 1452 24608
rect 2044 24599 2096 24608
rect 2044 24565 2053 24599
rect 2053 24565 2087 24599
rect 2087 24565 2096 24599
rect 2044 24556 2096 24565
rect 2412 24599 2464 24608
rect 2412 24565 2421 24599
rect 2421 24565 2455 24599
rect 2455 24565 2464 24599
rect 2412 24556 2464 24565
rect 2504 24556 2556 24608
rect 3056 24599 3108 24608
rect 3056 24565 3065 24599
rect 3065 24565 3099 24599
rect 3099 24565 3108 24599
rect 3056 24556 3108 24565
rect 10968 24556 11020 24608
rect 11244 24599 11296 24608
rect 11244 24565 11253 24599
rect 11253 24565 11287 24599
rect 11287 24565 11296 24599
rect 11244 24556 11296 24565
rect 12164 24599 12216 24608
rect 12164 24565 12173 24599
rect 12173 24565 12207 24599
rect 12207 24565 12216 24599
rect 12164 24556 12216 24565
rect 12992 24599 13044 24608
rect 12992 24565 13001 24599
rect 13001 24565 13035 24599
rect 13035 24565 13044 24599
rect 12992 24556 13044 24565
rect 14740 24599 14792 24608
rect 14740 24565 14749 24599
rect 14749 24565 14783 24599
rect 14783 24565 14792 24599
rect 14740 24556 14792 24565
rect 15844 24599 15896 24608
rect 15844 24565 15853 24599
rect 15853 24565 15887 24599
rect 15887 24565 15896 24599
rect 15844 24556 15896 24565
rect 15936 24556 15988 24608
rect 19800 24735 19852 24744
rect 17132 24624 17184 24676
rect 19800 24701 19809 24735
rect 19809 24701 19843 24735
rect 19843 24701 19852 24735
rect 19800 24692 19852 24701
rect 19248 24624 19300 24676
rect 16672 24599 16724 24608
rect 16672 24565 16681 24599
rect 16681 24565 16715 24599
rect 16715 24565 16724 24599
rect 16672 24556 16724 24565
rect 16764 24599 16816 24608
rect 16764 24565 16773 24599
rect 16773 24565 16807 24599
rect 16807 24565 16816 24599
rect 17776 24599 17828 24608
rect 16764 24556 16816 24565
rect 17776 24565 17785 24599
rect 17785 24565 17819 24599
rect 17819 24565 17828 24599
rect 17776 24556 17828 24565
rect 18880 24599 18932 24608
rect 18880 24565 18889 24599
rect 18889 24565 18923 24599
rect 18923 24565 18932 24599
rect 18880 24556 18932 24565
rect 19340 24599 19392 24608
rect 19340 24565 19349 24599
rect 19349 24565 19383 24599
rect 19383 24565 19392 24599
rect 19340 24556 19392 24565
rect 20076 24556 20128 24608
rect 20996 24692 21048 24744
rect 21456 24692 21508 24744
rect 22928 24692 22980 24744
rect 21824 24667 21876 24676
rect 21824 24633 21833 24667
rect 21833 24633 21867 24667
rect 21867 24633 21876 24667
rect 21824 24624 21876 24633
rect 20536 24556 20588 24608
rect 20720 24599 20772 24608
rect 20720 24565 20729 24599
rect 20729 24565 20763 24599
rect 20763 24565 20772 24599
rect 20720 24556 20772 24565
rect 21088 24599 21140 24608
rect 21088 24565 21097 24599
rect 21097 24565 21131 24599
rect 21131 24565 21140 24599
rect 21088 24556 21140 24565
rect 21916 24556 21968 24608
rect 22560 24556 22612 24608
rect 24032 24624 24084 24676
rect 24584 24624 24636 24676
rect 23572 24556 23624 24608
rect 24676 24556 24728 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 1492 24352 1544 24404
rect 2688 24395 2740 24404
rect 2688 24361 2697 24395
rect 2697 24361 2731 24395
rect 2731 24361 2740 24395
rect 2688 24352 2740 24361
rect 6368 24395 6420 24404
rect 6368 24361 6377 24395
rect 6377 24361 6411 24395
rect 6411 24361 6420 24395
rect 6368 24352 6420 24361
rect 7748 24352 7800 24404
rect 8300 24395 8352 24404
rect 8300 24361 8309 24395
rect 8309 24361 8343 24395
rect 8343 24361 8352 24395
rect 8300 24352 8352 24361
rect 8852 24352 8904 24404
rect 11060 24352 11112 24404
rect 11612 24352 11664 24404
rect 12164 24352 12216 24404
rect 12440 24352 12492 24404
rect 18236 24352 18288 24404
rect 19984 24352 20036 24404
rect 21364 24352 21416 24404
rect 22468 24352 22520 24404
rect 7104 24284 7156 24336
rect 13544 24284 13596 24336
rect 16856 24284 16908 24336
rect 17408 24284 17460 24336
rect 23940 24284 23992 24336
rect 2136 24216 2188 24268
rect 2596 24216 2648 24268
rect 6184 24259 6236 24268
rect 6184 24225 6193 24259
rect 6193 24225 6227 24259
rect 6227 24225 6236 24259
rect 6184 24216 6236 24225
rect 7380 24259 7432 24268
rect 7380 24225 7389 24259
rect 7389 24225 7423 24259
rect 7423 24225 7432 24259
rect 7380 24216 7432 24225
rect 8484 24259 8536 24268
rect 8484 24225 8493 24259
rect 8493 24225 8527 24259
rect 8527 24225 8536 24259
rect 8484 24216 8536 24225
rect 10508 24259 10560 24268
rect 10508 24225 10517 24259
rect 10517 24225 10551 24259
rect 10551 24225 10560 24259
rect 10508 24216 10560 24225
rect 10876 24216 10928 24268
rect 12348 24216 12400 24268
rect 13452 24216 13504 24268
rect 15476 24216 15528 24268
rect 16028 24216 16080 24268
rect 10784 24191 10836 24200
rect 10784 24157 10793 24191
rect 10793 24157 10827 24191
rect 10827 24157 10836 24191
rect 10784 24148 10836 24157
rect 12072 24148 12124 24200
rect 13360 24148 13412 24200
rect 3516 24080 3568 24132
rect 9680 24080 9732 24132
rect 11428 24080 11480 24132
rect 13544 24080 13596 24132
rect 15568 24148 15620 24200
rect 16212 24148 16264 24200
rect 16672 24080 16724 24132
rect 17040 24080 17092 24132
rect 17500 24216 17552 24268
rect 17960 24216 18012 24268
rect 20352 24216 20404 24268
rect 21272 24216 21324 24268
rect 22744 24216 22796 24268
rect 23756 24259 23808 24268
rect 23756 24225 23765 24259
rect 23765 24225 23799 24259
rect 23799 24225 23808 24259
rect 23756 24216 23808 24225
rect 23848 24259 23900 24268
rect 23848 24225 23857 24259
rect 23857 24225 23891 24259
rect 23891 24225 23900 24259
rect 24492 24259 24544 24268
rect 23848 24216 23900 24225
rect 24492 24225 24501 24259
rect 24501 24225 24535 24259
rect 24535 24225 24544 24259
rect 24492 24216 24544 24225
rect 24952 24259 25004 24268
rect 24952 24225 24961 24259
rect 24961 24225 24995 24259
rect 24995 24225 25004 24259
rect 24952 24216 25004 24225
rect 17316 24191 17368 24200
rect 17316 24157 17325 24191
rect 17325 24157 17359 24191
rect 17359 24157 17368 24191
rect 17316 24148 17368 24157
rect 18696 24191 18748 24200
rect 18696 24157 18705 24191
rect 18705 24157 18739 24191
rect 18739 24157 18748 24191
rect 18696 24148 18748 24157
rect 20720 24148 20772 24200
rect 18604 24080 18656 24132
rect 23296 24148 23348 24200
rect 22652 24080 22704 24132
rect 22836 24080 22888 24132
rect 25136 24123 25188 24132
rect 25136 24089 25145 24123
rect 25145 24089 25179 24123
rect 25179 24089 25188 24123
rect 25136 24080 25188 24089
rect 5264 24055 5316 24064
rect 5264 24021 5273 24055
rect 5273 24021 5307 24055
rect 5307 24021 5316 24055
rect 5264 24012 5316 24021
rect 6276 24012 6328 24064
rect 7196 24055 7248 24064
rect 7196 24021 7205 24055
rect 7205 24021 7239 24055
rect 7239 24021 7248 24055
rect 7196 24012 7248 24021
rect 9404 24055 9456 24064
rect 9404 24021 9413 24055
rect 9413 24021 9447 24055
rect 9447 24021 9456 24055
rect 9404 24012 9456 24021
rect 9772 24012 9824 24064
rect 11704 24055 11756 24064
rect 11704 24021 11713 24055
rect 11713 24021 11747 24055
rect 11747 24021 11756 24055
rect 11704 24012 11756 24021
rect 12808 24055 12860 24064
rect 12808 24021 12817 24055
rect 12817 24021 12851 24055
rect 12851 24021 12860 24055
rect 12808 24012 12860 24021
rect 13176 24012 13228 24064
rect 15292 24055 15344 24064
rect 15292 24021 15301 24055
rect 15301 24021 15335 24055
rect 15335 24021 15344 24055
rect 15292 24012 15344 24021
rect 16856 24055 16908 24064
rect 16856 24021 16865 24055
rect 16865 24021 16899 24055
rect 16899 24021 16908 24055
rect 16856 24012 16908 24021
rect 18144 24055 18196 24064
rect 18144 24021 18153 24055
rect 18153 24021 18187 24055
rect 18187 24021 18196 24055
rect 18144 24012 18196 24021
rect 20352 24055 20404 24064
rect 20352 24021 20361 24055
rect 20361 24021 20395 24055
rect 20395 24021 20404 24055
rect 20352 24012 20404 24021
rect 20904 24012 20956 24064
rect 21824 24012 21876 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 1676 23808 1728 23860
rect 2320 23808 2372 23860
rect 3516 23851 3568 23860
rect 3516 23817 3525 23851
rect 3525 23817 3559 23851
rect 3559 23817 3568 23851
rect 3516 23808 3568 23817
rect 7380 23808 7432 23860
rect 9128 23808 9180 23860
rect 9312 23851 9364 23860
rect 9312 23817 9321 23851
rect 9321 23817 9355 23851
rect 9355 23817 9364 23851
rect 9312 23808 9364 23817
rect 9864 23808 9916 23860
rect 11244 23808 11296 23860
rect 11520 23808 11572 23860
rect 4068 23740 4120 23792
rect 7472 23740 7524 23792
rect 8668 23740 8720 23792
rect 15476 23808 15528 23860
rect 16028 23851 16080 23860
rect 12716 23740 12768 23792
rect 13452 23783 13504 23792
rect 13452 23749 13461 23783
rect 13461 23749 13495 23783
rect 13495 23749 13504 23783
rect 13452 23740 13504 23749
rect 13636 23740 13688 23792
rect 14280 23740 14332 23792
rect 16028 23817 16037 23851
rect 16037 23817 16071 23851
rect 16071 23817 16080 23851
rect 16028 23808 16080 23817
rect 16764 23808 16816 23860
rect 21364 23808 21416 23860
rect 24952 23851 25004 23860
rect 24952 23817 24961 23851
rect 24961 23817 24995 23851
rect 24995 23817 25004 23851
rect 24952 23808 25004 23817
rect 26056 23808 26108 23860
rect 17316 23740 17368 23792
rect 20168 23783 20220 23792
rect 20168 23749 20177 23783
rect 20177 23749 20211 23783
rect 20211 23749 20220 23783
rect 20168 23740 20220 23749
rect 1952 23672 2004 23724
rect 2596 23672 2648 23724
rect 6092 23672 6144 23724
rect 8484 23672 8536 23724
rect 8944 23672 8996 23724
rect 9404 23672 9456 23724
rect 9956 23715 10008 23724
rect 9956 23681 9965 23715
rect 9965 23681 9999 23715
rect 9999 23681 10008 23715
rect 9956 23672 10008 23681
rect 12900 23715 12952 23724
rect 12900 23681 12909 23715
rect 12909 23681 12943 23715
rect 12943 23681 12952 23715
rect 12900 23672 12952 23681
rect 13360 23672 13412 23724
rect 1676 23604 1728 23656
rect 2136 23468 2188 23520
rect 2228 23468 2280 23520
rect 2688 23604 2740 23656
rect 5540 23604 5592 23656
rect 6184 23647 6236 23656
rect 6184 23613 6193 23647
rect 6193 23613 6227 23647
rect 6227 23613 6236 23647
rect 6184 23604 6236 23613
rect 7196 23604 7248 23656
rect 8300 23604 8352 23656
rect 10508 23604 10560 23656
rect 11060 23604 11112 23656
rect 11244 23647 11296 23656
rect 11244 23613 11253 23647
rect 11253 23613 11287 23647
rect 11287 23613 11296 23647
rect 11244 23604 11296 23613
rect 12440 23604 12492 23656
rect 5264 23536 5316 23588
rect 3516 23468 3568 23520
rect 4620 23468 4672 23520
rect 5448 23468 5500 23520
rect 10784 23536 10836 23588
rect 11520 23536 11572 23588
rect 14556 23604 14608 23656
rect 16120 23672 16172 23724
rect 16488 23672 16540 23724
rect 18604 23715 18656 23724
rect 16212 23604 16264 23656
rect 18604 23681 18613 23715
rect 18613 23681 18647 23715
rect 18647 23681 18656 23715
rect 18604 23672 18656 23681
rect 18972 23672 19024 23724
rect 22284 23715 22336 23724
rect 22284 23681 22293 23715
rect 22293 23681 22327 23715
rect 22327 23681 22336 23715
rect 22284 23672 22336 23681
rect 20904 23604 20956 23656
rect 24308 23715 24360 23724
rect 24308 23681 24317 23715
rect 24317 23681 24351 23715
rect 24351 23681 24360 23715
rect 24308 23672 24360 23681
rect 6368 23468 6420 23520
rect 8300 23468 8352 23520
rect 9680 23511 9732 23520
rect 9680 23477 9689 23511
rect 9689 23477 9723 23511
rect 9723 23477 9732 23511
rect 9680 23468 9732 23477
rect 11060 23511 11112 23520
rect 11060 23477 11069 23511
rect 11069 23477 11103 23511
rect 11103 23477 11112 23511
rect 11060 23468 11112 23477
rect 12808 23511 12860 23520
rect 12808 23477 12817 23511
rect 12817 23477 12851 23511
rect 12851 23477 12860 23511
rect 12808 23468 12860 23477
rect 13912 23468 13964 23520
rect 17776 23536 17828 23588
rect 18144 23536 18196 23588
rect 19156 23536 19208 23588
rect 20076 23536 20128 23588
rect 15108 23468 15160 23520
rect 16396 23468 16448 23520
rect 17500 23511 17552 23520
rect 17500 23477 17509 23511
rect 17509 23477 17543 23511
rect 17543 23477 17552 23511
rect 17500 23468 17552 23477
rect 18052 23468 18104 23520
rect 18788 23468 18840 23520
rect 19432 23468 19484 23520
rect 21272 23536 21324 23588
rect 24860 23604 24912 23656
rect 25228 23647 25280 23656
rect 25228 23613 25237 23647
rect 25237 23613 25271 23647
rect 25271 23613 25280 23647
rect 25228 23604 25280 23613
rect 23480 23536 23532 23588
rect 20260 23468 20312 23520
rect 22100 23511 22152 23520
rect 22100 23477 22109 23511
rect 22109 23477 22143 23511
rect 22143 23477 22152 23511
rect 22744 23511 22796 23520
rect 22100 23468 22152 23477
rect 22744 23477 22753 23511
rect 22753 23477 22787 23511
rect 22787 23477 22796 23511
rect 22744 23468 22796 23477
rect 23664 23511 23716 23520
rect 23664 23477 23673 23511
rect 23673 23477 23707 23511
rect 23707 23477 23716 23511
rect 23664 23468 23716 23477
rect 25412 23511 25464 23520
rect 25412 23477 25421 23511
rect 25421 23477 25455 23511
rect 25455 23477 25464 23511
rect 25412 23468 25464 23477
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 4068 23264 4120 23316
rect 5908 23264 5960 23316
rect 6552 23307 6604 23316
rect 6552 23273 6561 23307
rect 6561 23273 6595 23307
rect 6595 23273 6604 23307
rect 6552 23264 6604 23273
rect 11060 23307 11112 23316
rect 11060 23273 11069 23307
rect 11069 23273 11103 23307
rect 11103 23273 11112 23307
rect 11060 23264 11112 23273
rect 12164 23264 12216 23316
rect 13636 23307 13688 23316
rect 13636 23273 13645 23307
rect 13645 23273 13679 23307
rect 13679 23273 13688 23307
rect 13636 23264 13688 23273
rect 16764 23264 16816 23316
rect 16948 23264 17000 23316
rect 17224 23307 17276 23316
rect 17224 23273 17233 23307
rect 17233 23273 17267 23307
rect 17267 23273 17276 23307
rect 17224 23264 17276 23273
rect 18052 23307 18104 23316
rect 18052 23273 18061 23307
rect 18061 23273 18095 23307
rect 18095 23273 18104 23307
rect 18052 23264 18104 23273
rect 18420 23307 18472 23316
rect 18420 23273 18429 23307
rect 18429 23273 18463 23307
rect 18463 23273 18472 23307
rect 18420 23264 18472 23273
rect 20720 23264 20772 23316
rect 22008 23264 22060 23316
rect 23296 23307 23348 23316
rect 23296 23273 23305 23307
rect 23305 23273 23339 23307
rect 23339 23273 23348 23307
rect 23296 23264 23348 23273
rect 23480 23307 23532 23316
rect 23480 23273 23489 23307
rect 23489 23273 23523 23307
rect 23523 23273 23532 23307
rect 23480 23264 23532 23273
rect 24860 23307 24912 23316
rect 24860 23273 24869 23307
rect 24869 23273 24903 23307
rect 24903 23273 24912 23307
rect 24860 23264 24912 23273
rect 1676 23239 1728 23248
rect 1676 23205 1685 23239
rect 1685 23205 1719 23239
rect 1719 23205 1728 23239
rect 1676 23196 1728 23205
rect 2412 23196 2464 23248
rect 5540 23196 5592 23248
rect 6184 23196 6236 23248
rect 11796 23196 11848 23248
rect 12072 23196 12124 23248
rect 13544 23196 13596 23248
rect 14096 23239 14148 23248
rect 14096 23205 14105 23239
rect 14105 23205 14139 23239
rect 14139 23205 14148 23239
rect 14096 23196 14148 23205
rect 4896 23171 4948 23180
rect 4896 23137 4905 23171
rect 4905 23137 4939 23171
rect 4939 23137 4948 23171
rect 4896 23128 4948 23137
rect 7104 23128 7156 23180
rect 8116 23171 8168 23180
rect 8116 23137 8125 23171
rect 8125 23137 8159 23171
rect 8159 23137 8168 23171
rect 8116 23128 8168 23137
rect 2412 23060 2464 23112
rect 7012 23060 7064 23112
rect 8024 23060 8076 23112
rect 8300 23103 8352 23112
rect 8300 23069 8309 23103
rect 8309 23069 8343 23103
rect 8343 23069 8352 23103
rect 11152 23103 11204 23112
rect 8300 23060 8352 23069
rect 11152 23069 11161 23103
rect 11161 23069 11195 23103
rect 11195 23069 11204 23103
rect 11152 23060 11204 23069
rect 12440 23128 12492 23180
rect 14188 23128 14240 23180
rect 12072 23060 12124 23112
rect 12716 23103 12768 23112
rect 12716 23069 12725 23103
rect 12725 23069 12759 23103
rect 12759 23069 12768 23103
rect 12716 23060 12768 23069
rect 13360 23060 13412 23112
rect 13636 23060 13688 23112
rect 15936 23196 15988 23248
rect 19064 23196 19116 23248
rect 15568 23128 15620 23180
rect 17776 23128 17828 23180
rect 21364 23128 21416 23180
rect 24032 23196 24084 23248
rect 25320 23239 25372 23248
rect 25320 23205 25329 23239
rect 25329 23205 25363 23239
rect 25363 23205 25372 23239
rect 25320 23196 25372 23205
rect 25044 23171 25096 23180
rect 15476 23060 15528 23112
rect 15936 23103 15988 23112
rect 15936 23069 15945 23103
rect 15945 23069 15979 23103
rect 15979 23069 15988 23103
rect 15936 23060 15988 23069
rect 16580 23060 16632 23112
rect 5540 22992 5592 23044
rect 6736 22992 6788 23044
rect 2044 22967 2096 22976
rect 2044 22933 2053 22967
rect 2053 22933 2087 22967
rect 2087 22933 2096 22967
rect 2044 22924 2096 22933
rect 2596 22924 2648 22976
rect 4344 22967 4396 22976
rect 4344 22933 4353 22967
rect 4353 22933 4387 22967
rect 4387 22933 4396 22967
rect 4344 22924 4396 22933
rect 4804 22967 4856 22976
rect 4804 22933 4813 22967
rect 4813 22933 4847 22967
rect 4847 22933 4856 22967
rect 4804 22924 4856 22933
rect 6276 22924 6328 22976
rect 7472 22967 7524 22976
rect 7472 22933 7481 22967
rect 7481 22933 7515 22967
rect 7515 22933 7524 22967
rect 7472 22924 7524 22933
rect 8300 22924 8352 22976
rect 9680 22992 9732 23044
rect 10876 22992 10928 23044
rect 14740 22992 14792 23044
rect 16948 22992 17000 23044
rect 18972 23103 19024 23112
rect 18972 23069 18981 23103
rect 18981 23069 19015 23103
rect 19015 23069 19024 23103
rect 18972 23060 19024 23069
rect 19800 23103 19852 23112
rect 19800 23069 19809 23103
rect 19809 23069 19843 23103
rect 19843 23069 19852 23103
rect 19800 23060 19852 23069
rect 17684 22992 17736 23044
rect 22100 23060 22152 23112
rect 22284 23060 22336 23112
rect 23940 23103 23992 23112
rect 23940 23069 23949 23103
rect 23949 23069 23983 23103
rect 23983 23069 23992 23103
rect 23940 23060 23992 23069
rect 25044 23137 25053 23171
rect 25053 23137 25087 23171
rect 25087 23137 25096 23171
rect 25044 23128 25096 23137
rect 22468 23035 22520 23044
rect 22468 23001 22477 23035
rect 22477 23001 22511 23035
rect 22511 23001 22520 23035
rect 22468 22992 22520 23001
rect 23204 22992 23256 23044
rect 25320 23060 25372 23112
rect 9128 22924 9180 22976
rect 10692 22967 10744 22976
rect 10692 22933 10701 22967
rect 10701 22933 10735 22967
rect 10735 22933 10744 22967
rect 10692 22924 10744 22933
rect 11796 22967 11848 22976
rect 11796 22933 11805 22967
rect 11805 22933 11839 22967
rect 11839 22933 11848 22967
rect 11796 22924 11848 22933
rect 12164 22967 12216 22976
rect 12164 22933 12173 22967
rect 12173 22933 12207 22967
rect 12207 22933 12216 22967
rect 12164 22924 12216 22933
rect 14556 22967 14608 22976
rect 14556 22933 14565 22967
rect 14565 22933 14599 22967
rect 14599 22933 14608 22967
rect 14556 22924 14608 22933
rect 16212 22924 16264 22976
rect 16764 22967 16816 22976
rect 16764 22933 16773 22967
rect 16773 22933 16807 22967
rect 16807 22933 16816 22967
rect 16764 22924 16816 22933
rect 20168 22967 20220 22976
rect 20168 22933 20177 22967
rect 20177 22933 20211 22967
rect 20211 22933 20220 22967
rect 20168 22924 20220 22933
rect 20720 22967 20772 22976
rect 20720 22933 20729 22967
rect 20729 22933 20763 22967
rect 20763 22933 20772 22967
rect 20720 22924 20772 22933
rect 23020 22967 23072 22976
rect 23020 22933 23029 22967
rect 23029 22933 23063 22967
rect 23063 22933 23072 22967
rect 23020 22924 23072 22933
rect 24860 22924 24912 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 1584 22720 1636 22772
rect 3240 22720 3292 22772
rect 4988 22763 5040 22772
rect 4988 22729 4997 22763
rect 4997 22729 5031 22763
rect 5031 22729 5040 22763
rect 4988 22720 5040 22729
rect 6552 22763 6604 22772
rect 6552 22729 6561 22763
rect 6561 22729 6595 22763
rect 6595 22729 6604 22763
rect 6552 22720 6604 22729
rect 8116 22720 8168 22772
rect 5540 22584 5592 22636
rect 6092 22652 6144 22704
rect 6184 22627 6236 22636
rect 3148 22559 3200 22568
rect 3148 22525 3157 22559
rect 3157 22525 3191 22559
rect 3191 22525 3200 22559
rect 3148 22516 3200 22525
rect 2320 22448 2372 22500
rect 1584 22423 1636 22432
rect 1584 22389 1593 22423
rect 1593 22389 1627 22423
rect 1627 22389 1636 22423
rect 1584 22380 1636 22389
rect 2412 22423 2464 22432
rect 2412 22389 2421 22423
rect 2421 22389 2455 22423
rect 2455 22389 2464 22423
rect 2412 22380 2464 22389
rect 3332 22380 3384 22432
rect 6184 22593 6193 22627
rect 6193 22593 6227 22627
rect 6227 22593 6236 22627
rect 6184 22584 6236 22593
rect 6552 22516 6604 22568
rect 4988 22448 5040 22500
rect 7104 22448 7156 22500
rect 7288 22584 7340 22636
rect 7932 22627 7984 22636
rect 7932 22593 7941 22627
rect 7941 22593 7975 22627
rect 7975 22593 7984 22627
rect 7932 22584 7984 22593
rect 7472 22516 7524 22568
rect 8024 22448 8076 22500
rect 9404 22720 9456 22772
rect 11060 22720 11112 22772
rect 11428 22720 11480 22772
rect 9220 22584 9272 22636
rect 11244 22584 11296 22636
rect 12440 22720 12492 22772
rect 13636 22720 13688 22772
rect 14832 22720 14884 22772
rect 15568 22720 15620 22772
rect 16028 22720 16080 22772
rect 12348 22652 12400 22704
rect 12256 22584 12308 22636
rect 13544 22584 13596 22636
rect 9128 22516 9180 22568
rect 10692 22516 10744 22568
rect 13268 22516 13320 22568
rect 14464 22516 14516 22568
rect 9312 22448 9364 22500
rect 10508 22448 10560 22500
rect 12900 22448 12952 22500
rect 13360 22448 13412 22500
rect 16580 22720 16632 22772
rect 17224 22720 17276 22772
rect 19064 22763 19116 22772
rect 19064 22729 19073 22763
rect 19073 22729 19107 22763
rect 19107 22729 19116 22763
rect 19064 22720 19116 22729
rect 19616 22763 19668 22772
rect 19616 22729 19625 22763
rect 19625 22729 19659 22763
rect 19659 22729 19668 22763
rect 19616 22720 19668 22729
rect 20904 22720 20956 22772
rect 23848 22763 23900 22772
rect 23848 22729 23857 22763
rect 23857 22729 23891 22763
rect 23891 22729 23900 22763
rect 23848 22720 23900 22729
rect 14648 22584 14700 22636
rect 14924 22584 14976 22636
rect 15384 22584 15436 22636
rect 16488 22584 16540 22636
rect 15568 22559 15620 22568
rect 15568 22525 15577 22559
rect 15577 22525 15611 22559
rect 15611 22525 15620 22559
rect 15568 22516 15620 22525
rect 18696 22652 18748 22704
rect 16764 22584 16816 22636
rect 23572 22652 23624 22704
rect 23756 22652 23808 22704
rect 17316 22516 17368 22568
rect 19800 22584 19852 22636
rect 22100 22627 22152 22636
rect 22100 22593 22109 22627
rect 22109 22593 22143 22627
rect 22143 22593 22152 22627
rect 25044 22695 25096 22704
rect 25044 22661 25053 22695
rect 25053 22661 25087 22695
rect 25087 22661 25096 22695
rect 25044 22652 25096 22661
rect 22100 22584 22152 22593
rect 20352 22516 20404 22568
rect 20720 22516 20772 22568
rect 21732 22516 21784 22568
rect 23388 22516 23440 22568
rect 23572 22516 23624 22568
rect 23848 22516 23900 22568
rect 24860 22584 24912 22636
rect 18328 22448 18380 22500
rect 19524 22448 19576 22500
rect 4528 22380 4580 22432
rect 5080 22380 5132 22432
rect 6184 22380 6236 22432
rect 6644 22380 6696 22432
rect 7380 22423 7432 22432
rect 7380 22389 7389 22423
rect 7389 22389 7423 22423
rect 7423 22389 7432 22423
rect 7380 22380 7432 22389
rect 8852 22380 8904 22432
rect 11060 22380 11112 22432
rect 12440 22423 12492 22432
rect 12440 22389 12449 22423
rect 12449 22389 12483 22423
rect 12483 22389 12492 22423
rect 12440 22380 12492 22389
rect 13544 22423 13596 22432
rect 13544 22389 13553 22423
rect 13553 22389 13587 22423
rect 13587 22389 13596 22423
rect 13544 22380 13596 22389
rect 16304 22380 16356 22432
rect 17040 22423 17092 22432
rect 17040 22389 17049 22423
rect 17049 22389 17083 22423
rect 17083 22389 17092 22423
rect 17040 22380 17092 22389
rect 17776 22423 17828 22432
rect 17776 22389 17785 22423
rect 17785 22389 17819 22423
rect 17819 22389 17828 22423
rect 17776 22380 17828 22389
rect 18144 22380 18196 22432
rect 19248 22380 19300 22432
rect 21364 22380 21416 22432
rect 21548 22380 21600 22432
rect 23204 22380 23256 22432
rect 23388 22380 23440 22432
rect 24032 22423 24084 22432
rect 24032 22389 24041 22423
rect 24041 22389 24075 22423
rect 24075 22389 24084 22423
rect 24032 22380 24084 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 2872 22176 2924 22228
rect 1584 22040 1636 22092
rect 2688 22040 2740 22092
rect 5080 22176 5132 22228
rect 7288 22176 7340 22228
rect 7932 22176 7984 22228
rect 8668 22176 8720 22228
rect 9128 22176 9180 22228
rect 9496 22176 9548 22228
rect 12900 22219 12952 22228
rect 12900 22185 12909 22219
rect 12909 22185 12943 22219
rect 12943 22185 12952 22219
rect 12900 22176 12952 22185
rect 13268 22176 13320 22228
rect 13452 22176 13504 22228
rect 15568 22176 15620 22228
rect 7196 22108 7248 22160
rect 7656 22108 7708 22160
rect 4988 22040 5040 22092
rect 7288 22083 7340 22092
rect 7288 22049 7322 22083
rect 7322 22049 7340 22083
rect 7288 22040 7340 22049
rect 8668 22040 8720 22092
rect 10140 22040 10192 22092
rect 11152 22108 11204 22160
rect 12348 22108 12400 22160
rect 12440 22108 12492 22160
rect 11244 22083 11296 22092
rect 11244 22049 11278 22083
rect 11278 22049 11296 22083
rect 11244 22040 11296 22049
rect 11980 22040 12032 22092
rect 13728 22040 13780 22092
rect 14648 22040 14700 22092
rect 5172 22015 5224 22024
rect 5172 21981 5181 22015
rect 5181 21981 5215 22015
rect 5215 21981 5224 22015
rect 5172 21972 5224 21981
rect 5448 21972 5500 22024
rect 3608 21904 3660 21956
rect 4896 21904 4948 21956
rect 6644 21904 6696 21956
rect 8116 21972 8168 22024
rect 8392 21972 8444 22024
rect 9680 21972 9732 22024
rect 14096 21972 14148 22024
rect 21180 22176 21232 22228
rect 21548 22176 21600 22228
rect 21732 22176 21784 22228
rect 23940 22219 23992 22228
rect 23940 22185 23949 22219
rect 23949 22185 23983 22219
rect 23983 22185 23992 22219
rect 23940 22176 23992 22185
rect 24860 22176 24912 22228
rect 19064 22108 19116 22160
rect 20904 22151 20956 22160
rect 20904 22117 20913 22151
rect 20913 22117 20947 22151
rect 20947 22117 20956 22151
rect 20904 22108 20956 22117
rect 22100 22108 22152 22160
rect 17224 22083 17276 22092
rect 17224 22049 17233 22083
rect 17233 22049 17267 22083
rect 17267 22049 17276 22083
rect 17224 22040 17276 22049
rect 19524 22040 19576 22092
rect 22284 22083 22336 22092
rect 22284 22049 22293 22083
rect 22293 22049 22327 22083
rect 22327 22049 22336 22083
rect 22284 22040 22336 22049
rect 24032 22108 24084 22160
rect 24768 22040 24820 22092
rect 10692 21904 10744 21956
rect 15568 21972 15620 22024
rect 16304 21972 16356 22024
rect 15476 21904 15528 21956
rect 1400 21836 1452 21888
rect 3516 21879 3568 21888
rect 3516 21845 3525 21879
rect 3525 21845 3559 21879
rect 3559 21845 3568 21879
rect 3516 21836 3568 21845
rect 4160 21836 4212 21888
rect 6920 21836 6972 21888
rect 8392 21879 8444 21888
rect 8392 21845 8401 21879
rect 8401 21845 8435 21879
rect 8435 21845 8444 21879
rect 8392 21836 8444 21845
rect 9220 21879 9272 21888
rect 9220 21845 9229 21879
rect 9229 21845 9263 21879
rect 9263 21845 9272 21879
rect 9220 21836 9272 21845
rect 10968 21836 11020 21888
rect 11980 21836 12032 21888
rect 13636 21879 13688 21888
rect 13636 21845 13645 21879
rect 13645 21845 13679 21879
rect 13679 21845 13688 21879
rect 13636 21836 13688 21845
rect 15384 21836 15436 21888
rect 15844 21904 15896 21956
rect 16948 21972 17000 22024
rect 15936 21836 15988 21888
rect 16396 21836 16448 21888
rect 16856 21904 16908 21956
rect 17868 21972 17920 22024
rect 18328 21972 18380 22024
rect 18144 21879 18196 21888
rect 18144 21845 18153 21879
rect 18153 21845 18187 21879
rect 18187 21845 18196 21879
rect 18144 21836 18196 21845
rect 19248 21836 19300 21888
rect 22192 21972 22244 22024
rect 21824 21904 21876 21956
rect 23296 21972 23348 22024
rect 24952 21972 25004 22024
rect 23572 21904 23624 21956
rect 24032 21904 24084 21956
rect 20536 21836 20588 21888
rect 23940 21836 23992 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 3516 21632 3568 21684
rect 5172 21632 5224 21684
rect 6552 21632 6604 21684
rect 3056 21496 3108 21548
rect 4344 21496 4396 21548
rect 4712 21539 4764 21548
rect 4712 21505 4721 21539
rect 4721 21505 4755 21539
rect 4755 21505 4764 21539
rect 4712 21496 4764 21505
rect 1400 21471 1452 21480
rect 1400 21437 1409 21471
rect 1409 21437 1443 21471
rect 1443 21437 1452 21471
rect 1400 21428 1452 21437
rect 1584 21428 1636 21480
rect 5172 21496 5224 21548
rect 6092 21496 6144 21548
rect 6644 21496 6696 21548
rect 9680 21632 9732 21684
rect 9956 21632 10008 21684
rect 12256 21675 12308 21684
rect 12256 21641 12265 21675
rect 12265 21641 12299 21675
rect 12299 21641 12308 21675
rect 12256 21632 12308 21641
rect 12348 21632 12400 21684
rect 13728 21632 13780 21684
rect 14096 21632 14148 21684
rect 17224 21675 17276 21684
rect 17224 21641 17233 21675
rect 17233 21641 17267 21675
rect 17267 21641 17276 21675
rect 17224 21632 17276 21641
rect 21180 21675 21232 21684
rect 21180 21641 21189 21675
rect 21189 21641 21223 21675
rect 21223 21641 21232 21675
rect 21180 21632 21232 21641
rect 22192 21675 22244 21684
rect 22192 21641 22201 21675
rect 22201 21641 22235 21675
rect 22235 21641 22244 21675
rect 22192 21632 22244 21641
rect 23296 21632 23348 21684
rect 23756 21632 23808 21684
rect 24216 21632 24268 21684
rect 25412 21675 25464 21684
rect 25412 21641 25421 21675
rect 25421 21641 25455 21675
rect 25455 21641 25464 21675
rect 25412 21632 25464 21641
rect 17040 21564 17092 21616
rect 18328 21564 18380 21616
rect 19984 21564 20036 21616
rect 4988 21428 5040 21480
rect 6920 21428 6972 21480
rect 8392 21428 8444 21480
rect 9036 21428 9088 21480
rect 9220 21428 9272 21480
rect 13820 21496 13872 21548
rect 14924 21539 14976 21548
rect 14924 21505 14933 21539
rect 14933 21505 14967 21539
rect 14967 21505 14976 21539
rect 14924 21496 14976 21505
rect 16120 21496 16172 21548
rect 18604 21539 18656 21548
rect 18604 21505 18613 21539
rect 18613 21505 18647 21539
rect 18647 21505 18656 21539
rect 18604 21496 18656 21505
rect 19432 21496 19484 21548
rect 21456 21564 21508 21616
rect 20536 21496 20588 21548
rect 20720 21539 20772 21548
rect 20720 21505 20729 21539
rect 20729 21505 20763 21539
rect 20763 21505 20772 21539
rect 20720 21496 20772 21505
rect 21824 21539 21876 21548
rect 21824 21505 21833 21539
rect 21833 21505 21867 21539
rect 21867 21505 21876 21539
rect 21824 21496 21876 21505
rect 23940 21496 23992 21548
rect 1676 21403 1728 21412
rect 1676 21369 1685 21403
rect 1685 21369 1719 21403
rect 1719 21369 1728 21403
rect 1676 21360 1728 21369
rect 3240 21360 3292 21412
rect 7288 21360 7340 21412
rect 8668 21360 8720 21412
rect 10600 21360 10652 21412
rect 10968 21360 11020 21412
rect 2872 21292 2924 21344
rect 4160 21292 4212 21344
rect 5448 21292 5500 21344
rect 8852 21335 8904 21344
rect 8852 21301 8861 21335
rect 8861 21301 8895 21335
rect 8895 21301 8904 21335
rect 8852 21292 8904 21301
rect 11244 21292 11296 21344
rect 11428 21292 11480 21344
rect 14096 21360 14148 21412
rect 15384 21360 15436 21412
rect 23572 21428 23624 21480
rect 17960 21360 18012 21412
rect 23296 21360 23348 21412
rect 12440 21292 12492 21344
rect 13360 21292 13412 21344
rect 13820 21292 13872 21344
rect 14648 21292 14700 21344
rect 16120 21292 16172 21344
rect 16304 21335 16356 21344
rect 16304 21301 16313 21335
rect 16313 21301 16347 21335
rect 16347 21301 16356 21335
rect 16304 21292 16356 21301
rect 16948 21335 17000 21344
rect 16948 21301 16957 21335
rect 16957 21301 16991 21335
rect 16991 21301 17000 21335
rect 16948 21292 17000 21301
rect 18052 21335 18104 21344
rect 18052 21301 18061 21335
rect 18061 21301 18095 21335
rect 18095 21301 18104 21335
rect 18052 21292 18104 21301
rect 18328 21292 18380 21344
rect 19064 21335 19116 21344
rect 19064 21301 19073 21335
rect 19073 21301 19107 21335
rect 19107 21301 19116 21335
rect 19064 21292 19116 21301
rect 19524 21292 19576 21344
rect 20904 21292 20956 21344
rect 22284 21292 22336 21344
rect 23664 21335 23716 21344
rect 23664 21301 23673 21335
rect 23673 21301 23707 21335
rect 23707 21301 23716 21335
rect 23664 21292 23716 21301
rect 24768 21335 24820 21344
rect 24768 21301 24777 21335
rect 24777 21301 24811 21335
rect 24811 21301 24820 21335
rect 24768 21292 24820 21301
rect 25872 21292 25924 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 2412 21131 2464 21140
rect 2412 21097 2421 21131
rect 2421 21097 2455 21131
rect 2455 21097 2464 21131
rect 2412 21088 2464 21097
rect 6920 21131 6972 21140
rect 6920 21097 6929 21131
rect 6929 21097 6963 21131
rect 6963 21097 6972 21131
rect 6920 21088 6972 21097
rect 8208 21088 8260 21140
rect 1768 21020 1820 21072
rect 2688 21020 2740 21072
rect 4252 21020 4304 21072
rect 5172 21020 5224 21072
rect 8760 21020 8812 21072
rect 9220 21020 9272 21072
rect 2964 20952 3016 21004
rect 4896 20952 4948 21004
rect 8300 20952 8352 21004
rect 3056 20927 3108 20936
rect 3056 20893 3065 20927
rect 3065 20893 3099 20927
rect 3099 20893 3108 20927
rect 3056 20884 3108 20893
rect 9588 20952 9640 21004
rect 9680 20995 9732 21004
rect 9680 20961 9689 20995
rect 9689 20961 9723 20995
rect 9723 20961 9732 20995
rect 9956 20995 10008 21004
rect 9680 20952 9732 20961
rect 9956 20961 9990 20995
rect 9990 20961 10008 20995
rect 9956 20952 10008 20961
rect 13728 21088 13780 21140
rect 14096 21131 14148 21140
rect 14096 21097 14105 21131
rect 14105 21097 14139 21131
rect 14139 21097 14148 21131
rect 14096 21088 14148 21097
rect 14740 21131 14792 21140
rect 14740 21097 14749 21131
rect 14749 21097 14783 21131
rect 14783 21097 14792 21131
rect 14740 21088 14792 21097
rect 16580 21088 16632 21140
rect 18604 21088 18656 21140
rect 19432 21088 19484 21140
rect 20812 21088 20864 21140
rect 23296 21131 23348 21140
rect 23296 21097 23305 21131
rect 23305 21097 23339 21131
rect 23339 21097 23348 21131
rect 23296 21088 23348 21097
rect 23388 21088 23440 21140
rect 8760 20884 8812 20936
rect 9036 20884 9088 20936
rect 12164 20927 12216 20936
rect 12164 20893 12173 20927
rect 12173 20893 12207 20927
rect 12207 20893 12216 20927
rect 12164 20884 12216 20893
rect 14188 21020 14240 21072
rect 15384 21020 15436 21072
rect 16304 21020 16356 21072
rect 21180 21020 21232 21072
rect 24860 21088 24912 21140
rect 25412 21088 25464 21140
rect 24952 21020 25004 21072
rect 25320 21020 25372 21072
rect 13544 20952 13596 21004
rect 14096 20952 14148 21004
rect 16948 20952 17000 21004
rect 18604 20952 18656 21004
rect 20720 20952 20772 21004
rect 21824 20952 21876 21004
rect 23112 20952 23164 21004
rect 23664 20995 23716 21004
rect 23664 20961 23673 20995
rect 23673 20961 23707 20995
rect 23707 20961 23716 20995
rect 23664 20952 23716 20961
rect 14924 20884 14976 20936
rect 18972 20927 19024 20936
rect 18972 20893 18981 20927
rect 18981 20893 19015 20927
rect 19015 20893 19024 20927
rect 18972 20884 19024 20893
rect 20996 20884 21048 20936
rect 23480 20884 23532 20936
rect 24676 20884 24728 20936
rect 25044 20884 25096 20936
rect 11060 20859 11112 20868
rect 11060 20825 11069 20859
rect 11069 20825 11103 20859
rect 11103 20825 11112 20859
rect 11060 20816 11112 20825
rect 14188 20816 14240 20868
rect 1492 20748 1544 20800
rect 3700 20791 3752 20800
rect 3700 20757 3709 20791
rect 3709 20757 3743 20791
rect 3743 20757 3752 20791
rect 3700 20748 3752 20757
rect 4252 20791 4304 20800
rect 4252 20757 4261 20791
rect 4261 20757 4295 20791
rect 4295 20757 4304 20791
rect 4252 20748 4304 20757
rect 4344 20748 4396 20800
rect 5448 20748 5500 20800
rect 6828 20748 6880 20800
rect 12440 20748 12492 20800
rect 13360 20748 13412 20800
rect 15568 20748 15620 20800
rect 20904 20859 20956 20868
rect 20904 20825 20913 20859
rect 20913 20825 20947 20859
rect 20947 20825 20956 20859
rect 20904 20816 20956 20825
rect 18512 20748 18564 20800
rect 19616 20791 19668 20800
rect 19616 20757 19625 20791
rect 19625 20757 19659 20791
rect 19659 20757 19668 20791
rect 19616 20748 19668 20757
rect 19708 20748 19760 20800
rect 20352 20748 20404 20800
rect 20536 20748 20588 20800
rect 22100 20748 22152 20800
rect 22836 20791 22888 20800
rect 22836 20757 22845 20791
rect 22845 20757 22879 20791
rect 22879 20757 22888 20791
rect 22836 20748 22888 20757
rect 23296 20748 23348 20800
rect 23756 20748 23808 20800
rect 24860 20791 24912 20800
rect 24860 20757 24869 20791
rect 24869 20757 24903 20791
rect 24903 20757 24912 20791
rect 24860 20748 24912 20757
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 2688 20587 2740 20596
rect 2688 20553 2697 20587
rect 2697 20553 2731 20587
rect 2731 20553 2740 20587
rect 2688 20544 2740 20553
rect 2964 20587 3016 20596
rect 2964 20553 2973 20587
rect 2973 20553 3007 20587
rect 3007 20553 3016 20587
rect 2964 20544 3016 20553
rect 4160 20544 4212 20596
rect 4712 20587 4764 20596
rect 4712 20553 4721 20587
rect 4721 20553 4755 20587
rect 4755 20553 4764 20587
rect 4712 20544 4764 20553
rect 8300 20587 8352 20596
rect 8300 20553 8309 20587
rect 8309 20553 8343 20587
rect 8343 20553 8352 20587
rect 8300 20544 8352 20553
rect 9680 20544 9732 20596
rect 10692 20544 10744 20596
rect 10876 20544 10928 20596
rect 12440 20587 12492 20596
rect 12440 20553 12449 20587
rect 12449 20553 12483 20587
rect 12483 20553 12492 20587
rect 13544 20587 13596 20596
rect 12440 20544 12492 20553
rect 13544 20553 13553 20587
rect 13553 20553 13587 20587
rect 13587 20553 13596 20587
rect 13544 20544 13596 20553
rect 15292 20544 15344 20596
rect 15476 20544 15528 20596
rect 18052 20587 18104 20596
rect 18052 20553 18061 20587
rect 18061 20553 18095 20587
rect 18095 20553 18104 20587
rect 18052 20544 18104 20553
rect 18972 20544 19024 20596
rect 20720 20544 20772 20596
rect 20996 20587 21048 20596
rect 20996 20553 21005 20587
rect 21005 20553 21039 20587
rect 21039 20553 21048 20587
rect 20996 20544 21048 20553
rect 21180 20587 21232 20596
rect 21180 20553 21189 20587
rect 21189 20553 21223 20587
rect 21223 20553 21232 20587
rect 21180 20544 21232 20553
rect 22744 20544 22796 20596
rect 23572 20544 23624 20596
rect 25136 20544 25188 20596
rect 26240 20544 26292 20596
rect 2780 20476 2832 20528
rect 3056 20476 3108 20528
rect 6552 20476 6604 20528
rect 7012 20519 7064 20528
rect 7012 20485 7021 20519
rect 7021 20485 7055 20519
rect 7055 20485 7064 20519
rect 7012 20476 7064 20485
rect 11520 20476 11572 20528
rect 11704 20476 11756 20528
rect 17868 20476 17920 20528
rect 3516 20408 3568 20460
rect 4160 20408 4212 20460
rect 5080 20408 5132 20460
rect 9956 20408 10008 20460
rect 11980 20408 12032 20460
rect 14924 20408 14976 20460
rect 15384 20408 15436 20460
rect 16764 20451 16816 20460
rect 16764 20417 16773 20451
rect 16773 20417 16807 20451
rect 16807 20417 16816 20451
rect 16764 20408 16816 20417
rect 1768 20272 1820 20324
rect 1952 20315 2004 20324
rect 1952 20281 1961 20315
rect 1961 20281 1995 20315
rect 1995 20281 2004 20315
rect 1952 20272 2004 20281
rect 3332 20272 3384 20324
rect 1492 20204 1544 20256
rect 4160 20204 4212 20256
rect 7104 20340 7156 20392
rect 7564 20340 7616 20392
rect 10048 20340 10100 20392
rect 10784 20340 10836 20392
rect 12808 20383 12860 20392
rect 12808 20349 12817 20383
rect 12817 20349 12851 20383
rect 12851 20349 12860 20383
rect 12808 20340 12860 20349
rect 14740 20340 14792 20392
rect 17408 20340 17460 20392
rect 18512 20408 18564 20460
rect 19340 20408 19392 20460
rect 20168 20451 20220 20460
rect 20168 20417 20177 20451
rect 20177 20417 20211 20451
rect 20211 20417 20220 20451
rect 20168 20408 20220 20417
rect 23296 20408 23348 20460
rect 24676 20476 24728 20528
rect 24584 20408 24636 20460
rect 25320 20476 25372 20528
rect 25964 20519 26016 20528
rect 25964 20485 25973 20519
rect 25973 20485 26007 20519
rect 26007 20485 26016 20519
rect 25964 20476 26016 20485
rect 22008 20340 22060 20392
rect 24768 20340 24820 20392
rect 25228 20383 25280 20392
rect 25228 20349 25237 20383
rect 25237 20349 25271 20383
rect 25271 20349 25280 20383
rect 25228 20340 25280 20349
rect 4804 20272 4856 20324
rect 6552 20315 6604 20324
rect 6552 20281 6561 20315
rect 6561 20281 6595 20315
rect 6595 20281 6604 20315
rect 6552 20272 6604 20281
rect 8852 20272 8904 20324
rect 10692 20272 10744 20324
rect 11520 20272 11572 20324
rect 14188 20272 14240 20324
rect 15292 20272 15344 20324
rect 24952 20272 25004 20324
rect 5172 20204 5224 20256
rect 5448 20204 5500 20256
rect 6276 20204 6328 20256
rect 7564 20204 7616 20256
rect 9036 20204 9088 20256
rect 9956 20204 10008 20256
rect 13728 20204 13780 20256
rect 15200 20204 15252 20256
rect 15384 20204 15436 20256
rect 17776 20247 17828 20256
rect 17776 20213 17785 20247
rect 17785 20213 17819 20247
rect 17819 20213 17828 20247
rect 17776 20204 17828 20213
rect 19984 20247 20036 20256
rect 19984 20213 19993 20247
rect 19993 20213 20027 20247
rect 20027 20213 20036 20247
rect 19984 20204 20036 20213
rect 21640 20247 21692 20256
rect 21640 20213 21649 20247
rect 21649 20213 21683 20247
rect 21683 20213 21692 20247
rect 21640 20204 21692 20213
rect 23388 20247 23440 20256
rect 23388 20213 23397 20247
rect 23397 20213 23431 20247
rect 23431 20213 23440 20247
rect 23388 20204 23440 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 3332 20000 3384 20052
rect 6092 20043 6144 20052
rect 6092 20009 6101 20043
rect 6101 20009 6135 20043
rect 6135 20009 6144 20043
rect 6092 20000 6144 20009
rect 6736 20000 6788 20052
rect 7840 20000 7892 20052
rect 8024 20000 8076 20052
rect 8760 20043 8812 20052
rect 8760 20009 8769 20043
rect 8769 20009 8803 20043
rect 8803 20009 8812 20043
rect 8760 20000 8812 20009
rect 10784 20000 10836 20052
rect 11520 20043 11572 20052
rect 11520 20009 11529 20043
rect 11529 20009 11563 20043
rect 11563 20009 11572 20043
rect 11520 20000 11572 20009
rect 3148 19932 3200 19984
rect 3240 19864 3292 19916
rect 8944 19932 8996 19984
rect 10416 19932 10468 19984
rect 12348 20000 12400 20052
rect 13084 20043 13136 20052
rect 13084 20009 13093 20043
rect 13093 20009 13127 20043
rect 13127 20009 13136 20043
rect 13084 20000 13136 20009
rect 14188 20000 14240 20052
rect 14924 20000 14976 20052
rect 17868 20000 17920 20052
rect 18512 20000 18564 20052
rect 18972 20000 19024 20052
rect 21640 20000 21692 20052
rect 22468 20043 22520 20052
rect 22468 20009 22477 20043
rect 22477 20009 22511 20043
rect 22511 20009 22520 20043
rect 22468 20000 22520 20009
rect 23664 20000 23716 20052
rect 24492 20043 24544 20052
rect 24492 20009 24501 20043
rect 24501 20009 24535 20043
rect 24535 20009 24544 20043
rect 24492 20000 24544 20009
rect 24860 20000 24912 20052
rect 25412 20043 25464 20052
rect 25412 20009 25421 20043
rect 25421 20009 25455 20043
rect 25455 20009 25464 20043
rect 25412 20000 25464 20009
rect 11980 19932 12032 19984
rect 12992 19975 13044 19984
rect 12992 19941 13001 19975
rect 13001 19941 13035 19975
rect 13035 19941 13044 19975
rect 12992 19932 13044 19941
rect 16488 19932 16540 19984
rect 18052 19932 18104 19984
rect 20536 19932 20588 19984
rect 21272 19975 21324 19984
rect 4160 19864 4212 19916
rect 6920 19864 6972 19916
rect 2688 19796 2740 19848
rect 3056 19839 3108 19848
rect 3056 19805 3065 19839
rect 3065 19805 3099 19839
rect 3099 19805 3108 19839
rect 3056 19796 3108 19805
rect 3148 19796 3200 19848
rect 3792 19796 3844 19848
rect 4068 19839 4120 19848
rect 4068 19805 4077 19839
rect 4077 19805 4111 19839
rect 4111 19805 4120 19839
rect 4068 19796 4120 19805
rect 5080 19796 5132 19848
rect 6644 19796 6696 19848
rect 9772 19796 9824 19848
rect 11428 19796 11480 19848
rect 12440 19864 12492 19916
rect 13544 19907 13596 19916
rect 13544 19873 13553 19907
rect 13553 19873 13587 19907
rect 13587 19873 13596 19907
rect 13544 19864 13596 19873
rect 15200 19864 15252 19916
rect 15476 19864 15528 19916
rect 21272 19941 21281 19975
rect 21281 19941 21315 19975
rect 21315 19941 21324 19975
rect 21272 19932 21324 19941
rect 21824 19932 21876 19984
rect 22376 19932 22428 19984
rect 25228 19932 25280 19984
rect 11152 19728 11204 19780
rect 1676 19703 1728 19712
rect 1676 19669 1685 19703
rect 1685 19669 1719 19703
rect 1719 19669 1728 19703
rect 1676 19660 1728 19669
rect 2872 19660 2924 19712
rect 3792 19703 3844 19712
rect 3792 19669 3801 19703
rect 3801 19669 3835 19703
rect 3835 19669 3844 19703
rect 3792 19660 3844 19669
rect 5448 19703 5500 19712
rect 5448 19669 5457 19703
rect 5457 19669 5491 19703
rect 5491 19669 5500 19703
rect 5448 19660 5500 19669
rect 6368 19703 6420 19712
rect 6368 19669 6377 19703
rect 6377 19669 6411 19703
rect 6411 19669 6420 19703
rect 6368 19660 6420 19669
rect 11060 19703 11112 19712
rect 11060 19669 11069 19703
rect 11069 19669 11103 19703
rect 11103 19669 11112 19703
rect 11060 19660 11112 19669
rect 11888 19728 11940 19780
rect 12808 19796 12860 19848
rect 21364 19839 21416 19848
rect 21364 19805 21373 19839
rect 21373 19805 21407 19839
rect 21407 19805 21416 19839
rect 21364 19796 21416 19805
rect 22008 19864 22060 19916
rect 22284 19864 22336 19916
rect 22836 19907 22888 19916
rect 22836 19873 22845 19907
rect 22845 19873 22879 19907
rect 22879 19873 22888 19907
rect 22836 19864 22888 19873
rect 24032 19864 24084 19916
rect 21916 19796 21968 19848
rect 22744 19796 22796 19848
rect 22928 19839 22980 19848
rect 22928 19805 22937 19839
rect 22937 19805 22971 19839
rect 22971 19805 22980 19839
rect 22928 19796 22980 19805
rect 23112 19839 23164 19848
rect 23112 19805 23121 19839
rect 23121 19805 23155 19839
rect 23155 19805 23164 19839
rect 23112 19796 23164 19805
rect 23572 19796 23624 19848
rect 24584 19839 24636 19848
rect 24584 19805 24593 19839
rect 24593 19805 24627 19839
rect 24627 19805 24636 19839
rect 24584 19796 24636 19805
rect 12164 19728 12216 19780
rect 15292 19728 15344 19780
rect 21732 19728 21784 19780
rect 16580 19660 16632 19712
rect 17408 19703 17460 19712
rect 17408 19669 17417 19703
rect 17417 19669 17451 19703
rect 17451 19669 17460 19703
rect 17408 19660 17460 19669
rect 19248 19703 19300 19712
rect 19248 19669 19257 19703
rect 19257 19669 19291 19703
rect 19291 19669 19300 19703
rect 19248 19660 19300 19669
rect 20168 19660 20220 19712
rect 20536 19660 20588 19712
rect 21456 19660 21508 19712
rect 21916 19703 21968 19712
rect 21916 19669 21925 19703
rect 21925 19669 21959 19703
rect 21959 19669 21968 19703
rect 21916 19660 21968 19669
rect 22376 19703 22428 19712
rect 22376 19669 22385 19703
rect 22385 19669 22419 19703
rect 22419 19669 22428 19703
rect 22376 19660 22428 19669
rect 22468 19660 22520 19712
rect 23388 19660 23440 19712
rect 24032 19660 24084 19712
rect 24768 19660 24820 19712
rect 25044 19703 25096 19712
rect 25044 19669 25053 19703
rect 25053 19669 25087 19703
rect 25087 19669 25096 19703
rect 25044 19660 25096 19669
rect 26332 19660 26384 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 3240 19456 3292 19508
rect 8944 19456 8996 19508
rect 9772 19499 9824 19508
rect 9772 19465 9781 19499
rect 9781 19465 9815 19499
rect 9815 19465 9824 19499
rect 9772 19456 9824 19465
rect 12808 19499 12860 19508
rect 12808 19465 12817 19499
rect 12817 19465 12851 19499
rect 12851 19465 12860 19499
rect 12808 19456 12860 19465
rect 14648 19456 14700 19508
rect 16488 19499 16540 19508
rect 16488 19465 16497 19499
rect 16497 19465 16531 19499
rect 16531 19465 16540 19499
rect 16488 19456 16540 19465
rect 21364 19456 21416 19508
rect 22836 19456 22888 19508
rect 23572 19456 23624 19508
rect 23664 19456 23716 19508
rect 26148 19456 26200 19508
rect 1676 19388 1728 19440
rect 2688 19363 2740 19372
rect 2688 19329 2697 19363
rect 2697 19329 2731 19363
rect 2731 19329 2740 19363
rect 2688 19320 2740 19329
rect 3240 19320 3292 19372
rect 4160 19363 4212 19372
rect 4160 19329 4169 19363
rect 4169 19329 4203 19363
rect 4203 19329 4212 19363
rect 4160 19320 4212 19329
rect 5816 19363 5868 19372
rect 5816 19329 5825 19363
rect 5825 19329 5859 19363
rect 5859 19329 5868 19363
rect 5816 19320 5868 19329
rect 8116 19320 8168 19372
rect 8852 19363 8904 19372
rect 940 19116 992 19168
rect 4068 19295 4120 19304
rect 4068 19261 4077 19295
rect 4077 19261 4111 19295
rect 4111 19261 4120 19295
rect 4068 19252 4120 19261
rect 6644 19252 6696 19304
rect 7472 19252 7524 19304
rect 8852 19329 8861 19363
rect 8861 19329 8895 19363
rect 8895 19329 8904 19363
rect 8852 19320 8904 19329
rect 20812 19388 20864 19440
rect 22008 19388 22060 19440
rect 8668 19295 8720 19304
rect 2136 19184 2188 19236
rect 2780 19184 2832 19236
rect 2044 19159 2096 19168
rect 2044 19125 2053 19159
rect 2053 19125 2087 19159
rect 2087 19125 2096 19159
rect 2044 19116 2096 19125
rect 2872 19116 2924 19168
rect 3608 19159 3660 19168
rect 3608 19125 3617 19159
rect 3617 19125 3651 19159
rect 3651 19125 3660 19159
rect 3608 19116 3660 19125
rect 3976 19159 4028 19168
rect 3976 19125 3985 19159
rect 3985 19125 4019 19159
rect 4019 19125 4028 19159
rect 3976 19116 4028 19125
rect 4896 19116 4948 19168
rect 5356 19184 5408 19236
rect 6368 19184 6420 19236
rect 5172 19159 5224 19168
rect 5172 19125 5181 19159
rect 5181 19125 5215 19159
rect 5215 19125 5224 19159
rect 5172 19116 5224 19125
rect 5816 19116 5868 19168
rect 6552 19116 6604 19168
rect 7196 19116 7248 19168
rect 7380 19184 7432 19236
rect 8024 19184 8076 19236
rect 8668 19261 8677 19295
rect 8677 19261 8711 19295
rect 8711 19261 8720 19295
rect 8668 19252 8720 19261
rect 9588 19184 9640 19236
rect 8852 19116 8904 19168
rect 9956 19116 10008 19168
rect 10048 19116 10100 19168
rect 10232 19184 10284 19236
rect 12992 19252 13044 19304
rect 16764 19363 16816 19372
rect 16764 19329 16773 19363
rect 16773 19329 16807 19363
rect 16807 19329 16816 19363
rect 16764 19320 16816 19329
rect 16948 19295 17000 19304
rect 13636 19184 13688 19236
rect 11152 19116 11204 19168
rect 11428 19116 11480 19168
rect 11888 19159 11940 19168
rect 11888 19125 11897 19159
rect 11897 19125 11931 19159
rect 11931 19125 11940 19159
rect 11888 19116 11940 19125
rect 11980 19116 12032 19168
rect 13820 19116 13872 19168
rect 16948 19261 16957 19295
rect 16957 19261 16991 19295
rect 16991 19261 17000 19295
rect 16948 19252 17000 19261
rect 17500 19295 17552 19304
rect 17500 19261 17509 19295
rect 17509 19261 17543 19295
rect 17543 19261 17552 19295
rect 17500 19252 17552 19261
rect 19432 19252 19484 19304
rect 15660 19184 15712 19236
rect 19248 19184 19300 19236
rect 15752 19159 15804 19168
rect 15752 19125 15761 19159
rect 15761 19125 15795 19159
rect 15795 19125 15804 19159
rect 15752 19116 15804 19125
rect 18052 19116 18104 19168
rect 18328 19159 18380 19168
rect 18328 19125 18337 19159
rect 18337 19125 18371 19159
rect 18371 19125 18380 19159
rect 18328 19116 18380 19125
rect 19984 19116 20036 19168
rect 20996 19320 21048 19372
rect 21732 19363 21784 19372
rect 21732 19329 21741 19363
rect 21741 19329 21775 19363
rect 21775 19329 21784 19363
rect 21732 19320 21784 19329
rect 22560 19320 22612 19372
rect 25044 19388 25096 19440
rect 24584 19320 24636 19372
rect 25872 19320 25924 19372
rect 22744 19252 22796 19304
rect 24032 19295 24084 19304
rect 24032 19261 24041 19295
rect 24041 19261 24075 19295
rect 24075 19261 24084 19295
rect 24032 19252 24084 19261
rect 24124 19295 24176 19304
rect 24124 19261 24133 19295
rect 24133 19261 24167 19295
rect 24167 19261 24176 19295
rect 24124 19252 24176 19261
rect 25964 19252 26016 19304
rect 26240 19295 26292 19304
rect 26240 19261 26249 19295
rect 26249 19261 26283 19295
rect 26283 19261 26292 19295
rect 26240 19252 26292 19261
rect 20996 19184 21048 19236
rect 21916 19184 21968 19236
rect 21180 19159 21232 19168
rect 21180 19125 21189 19159
rect 21189 19125 21223 19159
rect 21223 19125 21232 19159
rect 21180 19116 21232 19125
rect 21456 19116 21508 19168
rect 23480 19116 23532 19168
rect 25136 19116 25188 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 2412 18955 2464 18964
rect 2412 18921 2421 18955
rect 2421 18921 2455 18955
rect 2455 18921 2464 18955
rect 2412 18912 2464 18921
rect 3608 18912 3660 18964
rect 3884 18912 3936 18964
rect 6828 18912 6880 18964
rect 8392 18912 8444 18964
rect 10048 18912 10100 18964
rect 12808 18912 12860 18964
rect 12992 18912 13044 18964
rect 15108 18955 15160 18964
rect 15108 18921 15117 18955
rect 15117 18921 15151 18955
rect 15151 18921 15160 18955
rect 15108 18912 15160 18921
rect 16212 18912 16264 18964
rect 2780 18887 2832 18896
rect 2780 18853 2789 18887
rect 2789 18853 2823 18887
rect 2823 18853 2832 18887
rect 2780 18844 2832 18853
rect 4344 18844 4396 18896
rect 5540 18844 5592 18896
rect 6920 18844 6972 18896
rect 7656 18844 7708 18896
rect 8944 18844 8996 18896
rect 10232 18844 10284 18896
rect 11520 18844 11572 18896
rect 18236 18912 18288 18964
rect 18420 18955 18472 18964
rect 18420 18921 18429 18955
rect 18429 18921 18463 18955
rect 18463 18921 18472 18955
rect 18420 18912 18472 18921
rect 18512 18912 18564 18964
rect 19248 18912 19300 18964
rect 19340 18912 19392 18964
rect 21272 18912 21324 18964
rect 21732 18912 21784 18964
rect 22376 18912 22428 18964
rect 24032 18912 24084 18964
rect 18052 18844 18104 18896
rect 21180 18844 21232 18896
rect 22560 18844 22612 18896
rect 24216 18844 24268 18896
rect 24860 18844 24912 18896
rect 4712 18776 4764 18828
rect 4804 18776 4856 18828
rect 6276 18776 6328 18828
rect 7104 18776 7156 18828
rect 7748 18776 7800 18828
rect 8484 18776 8536 18828
rect 9128 18776 9180 18828
rect 11060 18776 11112 18828
rect 11796 18776 11848 18828
rect 12256 18776 12308 18828
rect 12440 18819 12492 18828
rect 12440 18785 12474 18819
rect 12474 18785 12492 18819
rect 12440 18776 12492 18785
rect 15844 18776 15896 18828
rect 16028 18776 16080 18828
rect 16212 18776 16264 18828
rect 16948 18776 17000 18828
rect 17500 18776 17552 18828
rect 21088 18776 21140 18828
rect 21640 18776 21692 18828
rect 22192 18776 22244 18828
rect 24124 18776 24176 18828
rect 3424 18708 3476 18760
rect 5356 18708 5408 18760
rect 5816 18751 5868 18760
rect 5816 18717 5825 18751
rect 5825 18717 5859 18751
rect 5859 18717 5868 18751
rect 5816 18708 5868 18717
rect 7380 18751 7432 18760
rect 7380 18717 7389 18751
rect 7389 18717 7423 18751
rect 7423 18717 7432 18751
rect 7380 18708 7432 18717
rect 9588 18708 9640 18760
rect 2688 18640 2740 18692
rect 3148 18640 3200 18692
rect 4160 18640 4212 18692
rect 5448 18640 5500 18692
rect 2136 18615 2188 18624
rect 2136 18581 2145 18615
rect 2145 18581 2179 18615
rect 2179 18581 2188 18615
rect 2136 18572 2188 18581
rect 5264 18615 5316 18624
rect 5264 18581 5273 18615
rect 5273 18581 5307 18615
rect 5307 18581 5316 18615
rect 5264 18572 5316 18581
rect 5540 18572 5592 18624
rect 6828 18615 6880 18624
rect 6828 18581 6837 18615
rect 6837 18581 6871 18615
rect 6871 18581 6880 18615
rect 6828 18572 6880 18581
rect 8024 18572 8076 18624
rect 8300 18615 8352 18624
rect 8300 18581 8309 18615
rect 8309 18581 8343 18615
rect 8343 18581 8352 18615
rect 8300 18572 8352 18581
rect 9128 18615 9180 18624
rect 9128 18581 9137 18615
rect 9137 18581 9171 18615
rect 9171 18581 9180 18615
rect 9128 18572 9180 18581
rect 11796 18640 11848 18692
rect 14188 18708 14240 18760
rect 14648 18708 14700 18760
rect 13728 18640 13780 18692
rect 14740 18640 14792 18692
rect 16488 18708 16540 18760
rect 16764 18640 16816 18692
rect 11428 18572 11480 18624
rect 12440 18572 12492 18624
rect 15292 18615 15344 18624
rect 15292 18581 15301 18615
rect 15301 18581 15335 18615
rect 15335 18581 15344 18615
rect 15292 18572 15344 18581
rect 16672 18615 16724 18624
rect 16672 18581 16681 18615
rect 16681 18581 16715 18615
rect 16715 18581 16724 18615
rect 18604 18708 18656 18760
rect 19616 18708 19668 18760
rect 21364 18751 21416 18760
rect 21364 18717 21373 18751
rect 21373 18717 21407 18751
rect 21407 18717 21416 18751
rect 21364 18708 21416 18717
rect 21548 18751 21600 18760
rect 21548 18717 21557 18751
rect 21557 18717 21591 18751
rect 21591 18717 21600 18751
rect 21548 18708 21600 18717
rect 23020 18751 23072 18760
rect 23020 18717 23029 18751
rect 23029 18717 23063 18751
rect 23063 18717 23072 18751
rect 23020 18708 23072 18717
rect 23480 18708 23532 18760
rect 16672 18572 16724 18581
rect 18604 18572 18656 18624
rect 19432 18572 19484 18624
rect 21456 18640 21508 18692
rect 23940 18640 23992 18692
rect 24952 18640 25004 18692
rect 20904 18615 20956 18624
rect 20904 18581 20913 18615
rect 20913 18581 20947 18615
rect 20947 18581 20956 18615
rect 20904 18572 20956 18581
rect 23112 18572 23164 18624
rect 23388 18572 23440 18624
rect 23664 18572 23716 18624
rect 25136 18572 25188 18624
rect 26148 18615 26200 18624
rect 26148 18581 26157 18615
rect 26157 18581 26191 18615
rect 26191 18581 26200 18615
rect 26148 18572 26200 18581
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 2780 18368 2832 18420
rect 3148 18411 3200 18420
rect 3148 18377 3157 18411
rect 3157 18377 3191 18411
rect 3191 18377 3200 18411
rect 3148 18368 3200 18377
rect 3516 18368 3568 18420
rect 6736 18368 6788 18420
rect 7380 18368 7432 18420
rect 10692 18368 10744 18420
rect 11520 18411 11572 18420
rect 11520 18377 11529 18411
rect 11529 18377 11563 18411
rect 11563 18377 11572 18411
rect 11520 18368 11572 18377
rect 12808 18368 12860 18420
rect 13360 18411 13412 18420
rect 13360 18377 13369 18411
rect 13369 18377 13403 18411
rect 13403 18377 13412 18411
rect 13360 18368 13412 18377
rect 19064 18368 19116 18420
rect 21548 18368 21600 18420
rect 22100 18411 22152 18420
rect 22100 18377 22109 18411
rect 22109 18377 22143 18411
rect 22143 18377 22152 18411
rect 22100 18368 22152 18377
rect 2044 18232 2096 18284
rect 3700 18232 3752 18284
rect 12256 18343 12308 18352
rect 12256 18309 12265 18343
rect 12265 18309 12299 18343
rect 12299 18309 12308 18343
rect 12256 18300 12308 18309
rect 12900 18300 12952 18352
rect 2596 18164 2648 18216
rect 3976 18164 4028 18216
rect 4528 18232 4580 18284
rect 4988 18232 5040 18284
rect 5356 18232 5408 18284
rect 5816 18275 5868 18284
rect 5816 18241 5825 18275
rect 5825 18241 5859 18275
rect 5859 18241 5868 18275
rect 5816 18232 5868 18241
rect 10692 18232 10744 18284
rect 11428 18232 11480 18284
rect 16856 18343 16908 18352
rect 16856 18309 16865 18343
rect 16865 18309 16899 18343
rect 16899 18309 16908 18343
rect 16856 18300 16908 18309
rect 16948 18300 17000 18352
rect 22928 18343 22980 18352
rect 22928 18309 22937 18343
rect 22937 18309 22971 18343
rect 22971 18309 22980 18343
rect 22928 18300 22980 18309
rect 14740 18232 14792 18284
rect 15476 18275 15528 18284
rect 15476 18241 15485 18275
rect 15485 18241 15519 18275
rect 15519 18241 15528 18275
rect 15476 18232 15528 18241
rect 18604 18275 18656 18284
rect 18604 18241 18613 18275
rect 18613 18241 18647 18275
rect 18647 18241 18656 18275
rect 18604 18232 18656 18241
rect 4712 18207 4764 18216
rect 4712 18173 4721 18207
rect 4721 18173 4755 18207
rect 4755 18173 4764 18207
rect 4712 18164 4764 18173
rect 6368 18164 6420 18216
rect 7656 18164 7708 18216
rect 9588 18164 9640 18216
rect 6092 18096 6144 18148
rect 8024 18139 8076 18148
rect 8024 18105 8058 18139
rect 8058 18105 8076 18139
rect 8024 18096 8076 18105
rect 13544 18164 13596 18216
rect 16488 18164 16540 18216
rect 18236 18164 18288 18216
rect 23664 18232 23716 18284
rect 24952 18368 25004 18420
rect 25504 18368 25556 18420
rect 19984 18207 20036 18216
rect 19984 18173 20018 18207
rect 20018 18173 20036 18207
rect 16304 18096 16356 18148
rect 17500 18139 17552 18148
rect 17500 18105 17509 18139
rect 17509 18105 17543 18139
rect 17543 18105 17552 18139
rect 17500 18096 17552 18105
rect 18604 18096 18656 18148
rect 19340 18096 19392 18148
rect 19984 18164 20036 18173
rect 22376 18164 22428 18216
rect 23480 18164 23532 18216
rect 20904 18096 20956 18148
rect 21824 18096 21876 18148
rect 24216 18096 24268 18148
rect 26424 18096 26476 18148
rect 1676 18071 1728 18080
rect 1676 18037 1685 18071
rect 1685 18037 1719 18071
rect 1719 18037 1728 18071
rect 1676 18028 1728 18037
rect 4160 18028 4212 18080
rect 4804 18028 4856 18080
rect 5172 18028 5224 18080
rect 7104 18071 7156 18080
rect 7104 18037 7113 18071
rect 7113 18037 7147 18071
rect 7147 18037 7156 18071
rect 7104 18028 7156 18037
rect 8484 18028 8536 18080
rect 9128 18071 9180 18080
rect 9128 18037 9137 18071
rect 9137 18037 9171 18071
rect 9171 18037 9180 18071
rect 9128 18028 9180 18037
rect 10968 18071 11020 18080
rect 10968 18037 10977 18071
rect 10977 18037 11011 18071
rect 11011 18037 11020 18071
rect 10968 18028 11020 18037
rect 12992 18071 13044 18080
rect 12992 18037 13001 18071
rect 13001 18037 13035 18071
rect 13035 18037 13044 18071
rect 12992 18028 13044 18037
rect 13544 18071 13596 18080
rect 13544 18037 13553 18071
rect 13553 18037 13587 18071
rect 13587 18037 13596 18071
rect 13544 18028 13596 18037
rect 14648 18028 14700 18080
rect 15844 18028 15896 18080
rect 16396 18028 16448 18080
rect 17868 18071 17920 18080
rect 17868 18037 17877 18071
rect 17877 18037 17911 18071
rect 17911 18037 17920 18071
rect 17868 18028 17920 18037
rect 20720 18028 20772 18080
rect 21272 18028 21324 18080
rect 21456 18028 21508 18080
rect 23480 18071 23532 18080
rect 23480 18037 23489 18071
rect 23489 18037 23523 18071
rect 23523 18037 23532 18071
rect 23480 18028 23532 18037
rect 23756 18028 23808 18080
rect 24124 18028 24176 18080
rect 26240 18071 26292 18080
rect 26240 18037 26249 18071
rect 26249 18037 26283 18071
rect 26283 18037 26292 18071
rect 26240 18028 26292 18037
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 2596 17824 2648 17876
rect 3424 17867 3476 17876
rect 3424 17833 3433 17867
rect 3433 17833 3467 17867
rect 3467 17833 3476 17867
rect 3424 17824 3476 17833
rect 5448 17824 5500 17876
rect 6828 17824 6880 17876
rect 10692 17867 10744 17876
rect 10692 17833 10701 17867
rect 10701 17833 10735 17867
rect 10735 17833 10744 17867
rect 10692 17824 10744 17833
rect 12348 17824 12400 17876
rect 13544 17824 13596 17876
rect 14740 17824 14792 17876
rect 15292 17867 15344 17876
rect 15292 17833 15301 17867
rect 15301 17833 15335 17867
rect 15335 17833 15344 17867
rect 15292 17824 15344 17833
rect 5816 17756 5868 17808
rect 8024 17756 8076 17808
rect 10876 17756 10928 17808
rect 11520 17756 11572 17808
rect 11704 17799 11756 17808
rect 11704 17765 11713 17799
rect 11713 17765 11747 17799
rect 11747 17765 11756 17799
rect 11704 17756 11756 17765
rect 12440 17756 12492 17808
rect 13728 17756 13780 17808
rect 14004 17799 14056 17808
rect 14004 17765 14013 17799
rect 14013 17765 14047 17799
rect 14047 17765 14056 17799
rect 14004 17756 14056 17765
rect 15108 17756 15160 17808
rect 15936 17824 15988 17876
rect 17408 17824 17460 17876
rect 18420 17824 18472 17876
rect 19340 17824 19392 17876
rect 22192 17824 22244 17876
rect 22560 17824 22612 17876
rect 16856 17756 16908 17808
rect 19248 17756 19300 17808
rect 21456 17756 21508 17808
rect 22008 17756 22060 17808
rect 24032 17824 24084 17876
rect 26332 17867 26384 17876
rect 26332 17833 26341 17867
rect 26341 17833 26375 17867
rect 26375 17833 26384 17867
rect 26332 17824 26384 17833
rect 2780 17731 2832 17740
rect 2780 17697 2789 17731
rect 2789 17697 2823 17731
rect 2823 17697 2832 17731
rect 4436 17731 4488 17740
rect 2780 17688 2832 17697
rect 2228 17620 2280 17672
rect 2504 17620 2556 17672
rect 4436 17697 4470 17731
rect 4470 17697 4488 17731
rect 4436 17688 4488 17697
rect 6644 17688 6696 17740
rect 6828 17688 6880 17740
rect 7012 17731 7064 17740
rect 7012 17697 7021 17731
rect 7021 17697 7055 17731
rect 7055 17697 7064 17731
rect 7012 17688 7064 17697
rect 8116 17688 8168 17740
rect 9128 17688 9180 17740
rect 10416 17688 10468 17740
rect 13636 17688 13688 17740
rect 15292 17688 15344 17740
rect 15476 17688 15528 17740
rect 16488 17688 16540 17740
rect 17500 17688 17552 17740
rect 19524 17731 19576 17740
rect 19524 17697 19533 17731
rect 19533 17697 19567 17731
rect 19567 17697 19576 17731
rect 19524 17688 19576 17697
rect 21548 17688 21600 17740
rect 22468 17688 22520 17740
rect 23112 17756 23164 17808
rect 23664 17799 23716 17808
rect 23664 17765 23673 17799
rect 23673 17765 23707 17799
rect 23707 17765 23716 17799
rect 23664 17756 23716 17765
rect 24676 17756 24728 17808
rect 25228 17756 25280 17808
rect 22928 17731 22980 17740
rect 22928 17697 22937 17731
rect 22937 17697 22971 17731
rect 22971 17697 22980 17731
rect 22928 17688 22980 17697
rect 24768 17688 24820 17740
rect 2688 17552 2740 17604
rect 1952 17527 2004 17536
rect 1952 17493 1961 17527
rect 1961 17493 1995 17527
rect 1995 17493 2004 17527
rect 1952 17484 2004 17493
rect 2596 17484 2648 17536
rect 3608 17484 3660 17536
rect 6092 17620 6144 17672
rect 7472 17620 7524 17672
rect 10232 17663 10284 17672
rect 10232 17629 10241 17663
rect 10241 17629 10275 17663
rect 10275 17629 10284 17663
rect 10232 17620 10284 17629
rect 11060 17620 11112 17672
rect 12716 17620 12768 17672
rect 12992 17620 13044 17672
rect 7380 17552 7432 17604
rect 8852 17552 8904 17604
rect 9312 17595 9364 17604
rect 9312 17561 9321 17595
rect 9321 17561 9355 17595
rect 9355 17561 9364 17595
rect 9312 17552 9364 17561
rect 13636 17595 13688 17604
rect 13636 17561 13645 17595
rect 13645 17561 13679 17595
rect 13679 17561 13688 17595
rect 13636 17552 13688 17561
rect 14464 17620 14516 17672
rect 15752 17663 15804 17672
rect 15752 17629 15761 17663
rect 15761 17629 15795 17663
rect 15795 17629 15804 17663
rect 15752 17620 15804 17629
rect 16028 17620 16080 17672
rect 19708 17663 19760 17672
rect 19708 17629 19717 17663
rect 19717 17629 19751 17663
rect 19751 17629 19760 17663
rect 19708 17620 19760 17629
rect 21456 17663 21508 17672
rect 21456 17629 21465 17663
rect 21465 17629 21499 17663
rect 21499 17629 21508 17663
rect 21456 17620 21508 17629
rect 22008 17620 22060 17672
rect 23020 17663 23072 17672
rect 23020 17629 23029 17663
rect 23029 17629 23063 17663
rect 23063 17629 23072 17663
rect 23020 17620 23072 17629
rect 23112 17663 23164 17672
rect 23112 17629 23121 17663
rect 23121 17629 23155 17663
rect 23155 17629 23164 17663
rect 24676 17663 24728 17672
rect 23112 17620 23164 17629
rect 24676 17629 24685 17663
rect 24685 17629 24719 17663
rect 24719 17629 24728 17663
rect 24676 17620 24728 17629
rect 16672 17552 16724 17604
rect 19616 17552 19668 17604
rect 21180 17552 21232 17604
rect 24952 17552 25004 17604
rect 5080 17484 5132 17536
rect 6644 17527 6696 17536
rect 6644 17493 6653 17527
rect 6653 17493 6687 17527
rect 6687 17493 6696 17527
rect 6644 17484 6696 17493
rect 8208 17484 8260 17536
rect 8944 17527 8996 17536
rect 8944 17493 8953 17527
rect 8953 17493 8987 17527
rect 8987 17493 8996 17527
rect 8944 17484 8996 17493
rect 9680 17527 9732 17536
rect 9680 17493 9689 17527
rect 9689 17493 9723 17527
rect 9723 17493 9732 17527
rect 9680 17484 9732 17493
rect 12716 17484 12768 17536
rect 13084 17484 13136 17536
rect 13360 17484 13412 17536
rect 13820 17484 13872 17536
rect 16304 17527 16356 17536
rect 16304 17493 16313 17527
rect 16313 17493 16347 17527
rect 16347 17493 16356 17527
rect 16304 17484 16356 17493
rect 16764 17527 16816 17536
rect 16764 17493 16773 17527
rect 16773 17493 16807 17527
rect 16807 17493 16816 17527
rect 16764 17484 16816 17493
rect 18972 17527 19024 17536
rect 18972 17493 18981 17527
rect 18981 17493 19015 17527
rect 19015 17493 19024 17527
rect 18972 17484 19024 17493
rect 20996 17527 21048 17536
rect 20996 17493 21005 17527
rect 21005 17493 21039 17527
rect 21039 17493 21048 17527
rect 20996 17484 21048 17493
rect 24216 17484 24268 17536
rect 26148 17484 26200 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 2780 17323 2832 17332
rect 2780 17289 2789 17323
rect 2789 17289 2823 17323
rect 2823 17289 2832 17323
rect 2780 17280 2832 17289
rect 4436 17280 4488 17332
rect 7012 17280 7064 17332
rect 8024 17280 8076 17332
rect 9220 17280 9272 17332
rect 4620 17255 4672 17264
rect 4620 17221 4629 17255
rect 4629 17221 4663 17255
rect 4663 17221 4672 17255
rect 4620 17212 4672 17221
rect 1676 17144 1728 17196
rect 2964 17144 3016 17196
rect 3516 17144 3568 17196
rect 5080 17144 5132 17196
rect 9772 17212 9824 17264
rect 9956 17212 10008 17264
rect 10416 17255 10468 17264
rect 10416 17221 10425 17255
rect 10425 17221 10459 17255
rect 10459 17221 10468 17255
rect 10416 17212 10468 17221
rect 5264 17187 5316 17196
rect 5264 17153 5273 17187
rect 5273 17153 5307 17187
rect 5307 17153 5316 17187
rect 5264 17144 5316 17153
rect 6092 17144 6144 17196
rect 6276 17144 6328 17196
rect 9588 17144 9640 17196
rect 10232 17144 10284 17196
rect 11060 17280 11112 17332
rect 14188 17280 14240 17332
rect 15476 17280 15528 17332
rect 16304 17280 16356 17332
rect 16856 17280 16908 17332
rect 17960 17280 18012 17332
rect 19708 17323 19760 17332
rect 19708 17289 19717 17323
rect 19717 17289 19751 17323
rect 19751 17289 19760 17323
rect 19708 17280 19760 17289
rect 20076 17280 20128 17332
rect 23572 17280 23624 17332
rect 23756 17280 23808 17332
rect 24032 17280 24084 17332
rect 24768 17280 24820 17332
rect 12532 17212 12584 17264
rect 12808 17212 12860 17264
rect 13084 17212 13136 17264
rect 13268 17212 13320 17264
rect 11060 17144 11112 17196
rect 12256 17187 12308 17196
rect 12256 17153 12265 17187
rect 12265 17153 12299 17187
rect 12299 17153 12308 17187
rect 12256 17144 12308 17153
rect 13820 17144 13872 17196
rect 2596 17076 2648 17128
rect 3240 17076 3292 17128
rect 3424 17076 3476 17128
rect 7380 17076 7432 17128
rect 9312 17076 9364 17128
rect 10876 17119 10928 17128
rect 10876 17085 10885 17119
rect 10885 17085 10919 17119
rect 10919 17085 10928 17119
rect 10876 17076 10928 17085
rect 12716 17076 12768 17128
rect 17500 17212 17552 17264
rect 18972 17144 19024 17196
rect 17408 17119 17460 17128
rect 17408 17085 17417 17119
rect 17417 17085 17451 17119
rect 17451 17085 17460 17119
rect 17408 17076 17460 17085
rect 1124 17008 1176 17060
rect 2504 17051 2556 17060
rect 2504 17017 2513 17051
rect 2513 17017 2547 17051
rect 2547 17017 2556 17051
rect 2504 17008 2556 17017
rect 8392 17008 8444 17060
rect 12348 17008 12400 17060
rect 14464 17008 14516 17060
rect 15108 17008 15160 17060
rect 19248 17076 19300 17128
rect 21916 17212 21968 17264
rect 20904 17119 20956 17128
rect 20904 17085 20913 17119
rect 20913 17085 20947 17119
rect 20947 17085 20956 17119
rect 20904 17076 20956 17085
rect 22560 17076 22612 17128
rect 24216 17187 24268 17196
rect 24216 17153 24225 17187
rect 24225 17153 24259 17187
rect 24259 17153 24268 17187
rect 24216 17144 24268 17153
rect 24124 17119 24176 17128
rect 1676 16940 1728 16992
rect 1952 16940 2004 16992
rect 3056 16940 3108 16992
rect 3240 16940 3292 16992
rect 3608 16983 3660 16992
rect 3608 16949 3617 16983
rect 3617 16949 3651 16983
rect 3651 16949 3660 16983
rect 3608 16940 3660 16949
rect 4344 16940 4396 16992
rect 4712 16983 4764 16992
rect 4712 16949 4721 16983
rect 4721 16949 4755 16983
rect 4755 16949 4764 16983
rect 4712 16940 4764 16949
rect 8668 16940 8720 16992
rect 9128 16983 9180 16992
rect 9128 16949 9137 16983
rect 9137 16949 9171 16983
rect 9171 16949 9180 16983
rect 9128 16940 9180 16949
rect 9220 16940 9272 16992
rect 10784 16940 10836 16992
rect 12440 16983 12492 16992
rect 12440 16949 12449 16983
rect 12449 16949 12483 16983
rect 12483 16949 12492 16983
rect 12440 16940 12492 16949
rect 18512 16983 18564 16992
rect 18512 16949 18521 16983
rect 18521 16949 18555 16983
rect 18555 16949 18564 16983
rect 18512 16940 18564 16949
rect 18972 16940 19024 16992
rect 20444 16983 20496 16992
rect 20444 16949 20453 16983
rect 20453 16949 20487 16983
rect 20487 16949 20496 16983
rect 20444 16940 20496 16949
rect 22376 17008 22428 17060
rect 23112 17008 23164 17060
rect 24124 17085 24133 17119
rect 24133 17085 24167 17119
rect 24167 17085 24176 17119
rect 24124 17076 24176 17085
rect 24400 17008 24452 17060
rect 21364 16940 21416 16992
rect 22008 16940 22060 16992
rect 22560 16940 22612 16992
rect 22836 16940 22888 16992
rect 22928 16983 22980 16992
rect 22928 16949 22937 16983
rect 22937 16949 22971 16983
rect 22971 16949 22980 16983
rect 22928 16940 22980 16949
rect 24308 16940 24360 16992
rect 25228 16940 25280 16992
rect 25412 16983 25464 16992
rect 25412 16949 25421 16983
rect 25421 16949 25455 16983
rect 25455 16949 25464 16983
rect 25412 16940 25464 16949
rect 25504 16940 25556 16992
rect 26148 16983 26200 16992
rect 26148 16949 26157 16983
rect 26157 16949 26191 16983
rect 26191 16949 26200 16983
rect 26148 16940 26200 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 2688 16736 2740 16788
rect 2780 16736 2832 16788
rect 3516 16779 3568 16788
rect 3516 16745 3525 16779
rect 3525 16745 3559 16779
rect 3559 16745 3568 16779
rect 3516 16736 3568 16745
rect 6092 16736 6144 16788
rect 8024 16736 8076 16788
rect 9864 16736 9916 16788
rect 10692 16736 10744 16788
rect 11704 16736 11756 16788
rect 12900 16736 12952 16788
rect 13544 16736 13596 16788
rect 14004 16779 14056 16788
rect 14004 16745 14013 16779
rect 14013 16745 14047 16779
rect 14047 16745 14056 16779
rect 14004 16736 14056 16745
rect 14188 16779 14240 16788
rect 14188 16745 14197 16779
rect 14197 16745 14231 16779
rect 14231 16745 14240 16779
rect 14188 16736 14240 16745
rect 15752 16736 15804 16788
rect 16672 16736 16724 16788
rect 17224 16779 17276 16788
rect 17224 16745 17233 16779
rect 17233 16745 17267 16779
rect 17267 16745 17276 16779
rect 17224 16736 17276 16745
rect 18052 16779 18104 16788
rect 18052 16745 18061 16779
rect 18061 16745 18095 16779
rect 18095 16745 18104 16779
rect 18052 16736 18104 16745
rect 19524 16736 19576 16788
rect 20720 16736 20772 16788
rect 21916 16736 21968 16788
rect 23020 16736 23072 16788
rect 23112 16736 23164 16788
rect 1768 16711 1820 16720
rect 1768 16677 1777 16711
rect 1777 16677 1811 16711
rect 1811 16677 1820 16711
rect 1768 16668 1820 16677
rect 5448 16668 5500 16720
rect 6644 16668 6696 16720
rect 9312 16711 9364 16720
rect 9312 16677 9321 16711
rect 9321 16677 9355 16711
rect 9355 16677 9364 16711
rect 9312 16668 9364 16677
rect 11612 16668 11664 16720
rect 15108 16711 15160 16720
rect 2136 16600 2188 16652
rect 2412 16600 2464 16652
rect 3240 16600 3292 16652
rect 4712 16600 4764 16652
rect 5356 16600 5408 16652
rect 2044 16575 2096 16584
rect 2044 16541 2053 16575
rect 2053 16541 2087 16575
rect 2087 16541 2096 16575
rect 2044 16532 2096 16541
rect 4620 16575 4672 16584
rect 4620 16541 4629 16575
rect 4629 16541 4663 16575
rect 4663 16541 4672 16575
rect 4620 16532 4672 16541
rect 3424 16464 3476 16516
rect 5264 16464 5316 16516
rect 2504 16396 2556 16448
rect 4068 16439 4120 16448
rect 4068 16405 4077 16439
rect 4077 16405 4111 16439
rect 4111 16405 4120 16439
rect 4068 16396 4120 16405
rect 7104 16600 7156 16652
rect 8208 16600 8260 16652
rect 8300 16643 8352 16652
rect 8300 16609 8309 16643
rect 8309 16609 8343 16643
rect 8343 16609 8352 16643
rect 8300 16600 8352 16609
rect 10232 16600 10284 16652
rect 11428 16600 11480 16652
rect 6276 16575 6328 16584
rect 6276 16541 6285 16575
rect 6285 16541 6319 16575
rect 6319 16541 6328 16575
rect 6276 16532 6328 16541
rect 6644 16532 6696 16584
rect 6920 16532 6972 16584
rect 6276 16396 6328 16448
rect 6920 16396 6972 16448
rect 10324 16575 10376 16584
rect 10324 16541 10333 16575
rect 10333 16541 10367 16575
rect 10367 16541 10376 16575
rect 10324 16532 10376 16541
rect 11796 16600 11848 16652
rect 11980 16643 12032 16652
rect 11980 16609 12014 16643
rect 12014 16609 12032 16643
rect 15108 16677 15117 16711
rect 15117 16677 15151 16711
rect 15151 16677 15160 16711
rect 15108 16668 15160 16677
rect 16028 16668 16080 16720
rect 18144 16668 18196 16720
rect 18604 16668 18656 16720
rect 20444 16668 20496 16720
rect 22008 16668 22060 16720
rect 15844 16643 15896 16652
rect 11980 16600 12032 16609
rect 15844 16609 15853 16643
rect 15853 16609 15887 16643
rect 15887 16609 15896 16643
rect 15844 16600 15896 16609
rect 17040 16643 17092 16652
rect 17040 16609 17049 16643
rect 17049 16609 17083 16643
rect 17083 16609 17092 16643
rect 17040 16600 17092 16609
rect 10600 16464 10652 16516
rect 7196 16439 7248 16448
rect 7196 16405 7205 16439
rect 7205 16405 7239 16439
rect 7239 16405 7248 16439
rect 7196 16396 7248 16405
rect 9128 16396 9180 16448
rect 10692 16439 10744 16448
rect 10692 16405 10701 16439
rect 10701 16405 10735 16439
rect 10735 16405 10744 16439
rect 10692 16396 10744 16405
rect 13728 16532 13780 16584
rect 15936 16575 15988 16584
rect 15936 16541 15945 16575
rect 15945 16541 15979 16575
rect 15979 16541 15988 16575
rect 15936 16532 15988 16541
rect 14740 16464 14792 16516
rect 17500 16532 17552 16584
rect 19248 16600 19300 16652
rect 21456 16600 21508 16652
rect 21548 16600 21600 16652
rect 18144 16575 18196 16584
rect 18144 16541 18153 16575
rect 18153 16541 18187 16575
rect 18187 16541 18196 16575
rect 18144 16532 18196 16541
rect 20904 16575 20956 16584
rect 20904 16541 20913 16575
rect 20913 16541 20947 16575
rect 20947 16541 20956 16575
rect 20904 16532 20956 16541
rect 16396 16464 16448 16516
rect 17408 16464 17460 16516
rect 23112 16464 23164 16516
rect 23756 16736 23808 16788
rect 24400 16779 24452 16788
rect 24400 16745 24409 16779
rect 24409 16745 24443 16779
rect 24443 16745 24452 16779
rect 24400 16736 24452 16745
rect 25228 16711 25280 16720
rect 25228 16677 25237 16711
rect 25237 16677 25271 16711
rect 25271 16677 25280 16711
rect 25228 16668 25280 16677
rect 23756 16643 23808 16652
rect 23756 16609 23765 16643
rect 23765 16609 23799 16643
rect 23799 16609 23808 16643
rect 23756 16600 23808 16609
rect 25688 16643 25740 16652
rect 25688 16609 25697 16643
rect 25697 16609 25731 16643
rect 25731 16609 25740 16643
rect 25688 16600 25740 16609
rect 24032 16575 24084 16584
rect 24032 16541 24041 16575
rect 24041 16541 24075 16575
rect 24075 16541 24084 16575
rect 24032 16532 24084 16541
rect 24860 16532 24912 16584
rect 24124 16464 24176 16516
rect 24308 16464 24360 16516
rect 16672 16396 16724 16448
rect 17684 16439 17736 16448
rect 17684 16405 17693 16439
rect 17693 16405 17727 16439
rect 17727 16405 17736 16439
rect 17684 16396 17736 16405
rect 19524 16439 19576 16448
rect 19524 16405 19533 16439
rect 19533 16405 19567 16439
rect 19567 16405 19576 16439
rect 19524 16396 19576 16405
rect 23296 16396 23348 16448
rect 23756 16396 23808 16448
rect 24676 16396 24728 16448
rect 25688 16396 25740 16448
rect 26148 16396 26200 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 5264 16192 5316 16244
rect 8208 16192 8260 16244
rect 8852 16192 8904 16244
rect 9864 16192 9916 16244
rect 9956 16192 10008 16244
rect 10324 16192 10376 16244
rect 12348 16192 12400 16244
rect 13728 16192 13780 16244
rect 14740 16192 14792 16244
rect 16028 16192 16080 16244
rect 16396 16192 16448 16244
rect 17040 16235 17092 16244
rect 17040 16201 17049 16235
rect 17049 16201 17083 16235
rect 17083 16201 17092 16235
rect 17040 16192 17092 16201
rect 17500 16235 17552 16244
rect 17500 16201 17509 16235
rect 17509 16201 17543 16235
rect 17543 16201 17552 16235
rect 17500 16192 17552 16201
rect 20720 16235 20772 16244
rect 20720 16201 20729 16235
rect 20729 16201 20763 16235
rect 20763 16201 20772 16235
rect 20720 16192 20772 16201
rect 23112 16235 23164 16244
rect 23112 16201 23121 16235
rect 23121 16201 23155 16235
rect 23155 16201 23164 16235
rect 23112 16192 23164 16201
rect 23756 16192 23808 16244
rect 24860 16192 24912 16244
rect 25228 16192 25280 16244
rect 2872 16124 2924 16176
rect 3884 16124 3936 16176
rect 4712 16167 4764 16176
rect 4712 16133 4721 16167
rect 4721 16133 4755 16167
rect 4755 16133 4764 16167
rect 4712 16124 4764 16133
rect 5724 16124 5776 16176
rect 6276 16124 6328 16176
rect 8392 16124 8444 16176
rect 8760 16124 8812 16176
rect 2044 16099 2096 16108
rect 2044 16065 2053 16099
rect 2053 16065 2087 16099
rect 2087 16065 2096 16099
rect 2044 16056 2096 16065
rect 3424 16056 3476 16108
rect 6920 16056 6972 16108
rect 4620 15988 4672 16040
rect 5080 15988 5132 16040
rect 5448 15988 5500 16040
rect 6828 15988 6880 16040
rect 7104 15988 7156 16040
rect 8760 15988 8812 16040
rect 9128 16099 9180 16108
rect 9128 16065 9137 16099
rect 9137 16065 9171 16099
rect 9171 16065 9180 16099
rect 9128 16056 9180 16065
rect 9220 16056 9272 16108
rect 11060 16124 11112 16176
rect 10784 16099 10836 16108
rect 10784 16065 10793 16099
rect 10793 16065 10827 16099
rect 10827 16065 10836 16099
rect 10784 16056 10836 16065
rect 9036 15988 9088 16040
rect 10600 16031 10652 16040
rect 1308 15920 1360 15972
rect 1032 15852 1084 15904
rect 1676 15920 1728 15972
rect 2320 15920 2372 15972
rect 2596 15852 2648 15904
rect 3148 15895 3200 15904
rect 3148 15861 3157 15895
rect 3157 15861 3191 15895
rect 3191 15861 3200 15895
rect 3148 15852 3200 15861
rect 3516 15895 3568 15904
rect 3516 15861 3525 15895
rect 3525 15861 3559 15895
rect 3559 15861 3568 15895
rect 3516 15852 3568 15861
rect 3884 15852 3936 15904
rect 5080 15895 5132 15904
rect 5080 15861 5089 15895
rect 5089 15861 5123 15895
rect 5123 15861 5132 15895
rect 5080 15852 5132 15861
rect 8852 15920 8904 15972
rect 10048 15963 10100 15972
rect 10048 15929 10057 15963
rect 10057 15929 10091 15963
rect 10091 15929 10100 15963
rect 10048 15920 10100 15929
rect 10232 15920 10284 15972
rect 5264 15852 5316 15904
rect 6828 15852 6880 15904
rect 7104 15895 7156 15904
rect 7104 15861 7113 15895
rect 7113 15861 7147 15895
rect 7147 15861 7156 15895
rect 7104 15852 7156 15861
rect 7564 15895 7616 15904
rect 7564 15861 7573 15895
rect 7573 15861 7607 15895
rect 7607 15861 7616 15895
rect 7564 15852 7616 15861
rect 8484 15852 8536 15904
rect 9036 15895 9088 15904
rect 9036 15861 9045 15895
rect 9045 15861 9079 15895
rect 9079 15861 9088 15895
rect 9036 15852 9088 15861
rect 9496 15852 9548 15904
rect 10600 15997 10609 16031
rect 10609 15997 10643 16031
rect 10643 15997 10652 16031
rect 10600 15988 10652 15997
rect 13820 16124 13872 16176
rect 14096 16124 14148 16176
rect 12900 16056 12952 16108
rect 26240 16124 26292 16176
rect 19248 16056 19300 16108
rect 21916 16056 21968 16108
rect 22192 16056 22244 16108
rect 13820 16031 13872 16040
rect 10692 15895 10744 15904
rect 10692 15861 10701 15895
rect 10701 15861 10735 15895
rect 10735 15861 10744 15895
rect 10692 15852 10744 15861
rect 11428 15852 11480 15904
rect 13820 15997 13829 16031
rect 13829 15997 13863 16031
rect 13863 15997 13872 16031
rect 13820 15988 13872 15997
rect 16948 15988 17000 16040
rect 17684 15988 17736 16040
rect 18144 15988 18196 16040
rect 20996 15988 21048 16040
rect 22008 15988 22060 16040
rect 14740 15920 14792 15972
rect 18604 15920 18656 15972
rect 22192 15920 22244 15972
rect 17224 15852 17276 15904
rect 17408 15852 17460 15904
rect 17684 15852 17736 15904
rect 19340 15852 19392 15904
rect 20628 15852 20680 15904
rect 22928 15988 22980 16040
rect 23848 16056 23900 16108
rect 25044 16056 25096 16108
rect 24676 15988 24728 16040
rect 25596 15988 25648 16040
rect 24860 15920 24912 15972
rect 22560 15852 22612 15904
rect 23572 15852 23624 15904
rect 23848 15852 23900 15904
rect 26240 15852 26292 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 2688 15691 2740 15700
rect 2688 15657 2697 15691
rect 2697 15657 2731 15691
rect 2731 15657 2740 15691
rect 2688 15648 2740 15657
rect 3148 15648 3200 15700
rect 5080 15648 5132 15700
rect 5448 15648 5500 15700
rect 5724 15691 5776 15700
rect 5724 15657 5733 15691
rect 5733 15657 5767 15691
rect 5767 15657 5776 15691
rect 5724 15648 5776 15657
rect 6092 15691 6144 15700
rect 6092 15657 6101 15691
rect 6101 15657 6135 15691
rect 6135 15657 6144 15691
rect 6092 15648 6144 15657
rect 4068 15580 4120 15632
rect 4896 15580 4948 15632
rect 5264 15580 5316 15632
rect 8944 15648 8996 15700
rect 9220 15691 9272 15700
rect 9220 15657 9229 15691
rect 9229 15657 9263 15691
rect 9263 15657 9272 15691
rect 9220 15648 9272 15657
rect 9680 15691 9732 15700
rect 9680 15657 9689 15691
rect 9689 15657 9723 15691
rect 9723 15657 9732 15691
rect 9680 15648 9732 15657
rect 9864 15648 9916 15700
rect 10784 15648 10836 15700
rect 11980 15648 12032 15700
rect 12716 15648 12768 15700
rect 14372 15648 14424 15700
rect 16488 15648 16540 15700
rect 19432 15648 19484 15700
rect 20996 15648 21048 15700
rect 21640 15648 21692 15700
rect 22192 15648 22244 15700
rect 25044 15691 25096 15700
rect 5172 15512 5224 15564
rect 2320 15444 2372 15496
rect 2964 15444 3016 15496
rect 3424 15444 3476 15496
rect 5264 15487 5316 15496
rect 5264 15453 5273 15487
rect 5273 15453 5307 15487
rect 5307 15453 5316 15487
rect 5264 15444 5316 15453
rect 1860 15376 1912 15428
rect 2504 15376 2556 15428
rect 3148 15376 3200 15428
rect 4712 15419 4764 15428
rect 4712 15385 4721 15419
rect 4721 15385 4755 15419
rect 4755 15385 4764 15419
rect 4712 15376 4764 15385
rect 2044 15351 2096 15360
rect 2044 15317 2053 15351
rect 2053 15317 2087 15351
rect 2087 15317 2096 15351
rect 2044 15308 2096 15317
rect 2596 15308 2648 15360
rect 6276 15580 6328 15632
rect 8300 15623 8352 15632
rect 8300 15589 8309 15623
rect 8309 15589 8343 15623
rect 8343 15589 8352 15623
rect 8300 15580 8352 15589
rect 11152 15580 11204 15632
rect 13728 15580 13780 15632
rect 15844 15623 15896 15632
rect 15844 15589 15853 15623
rect 15853 15589 15887 15623
rect 15887 15589 15896 15623
rect 15844 15580 15896 15589
rect 20720 15580 20772 15632
rect 25044 15657 25053 15691
rect 25053 15657 25087 15691
rect 25087 15657 25096 15691
rect 25044 15648 25096 15657
rect 26332 15648 26384 15700
rect 23756 15580 23808 15632
rect 24676 15580 24728 15632
rect 6092 15512 6144 15564
rect 6368 15512 6420 15564
rect 9128 15512 9180 15564
rect 9772 15376 9824 15428
rect 11796 15512 11848 15564
rect 16488 15555 16540 15564
rect 16488 15521 16497 15555
rect 16497 15521 16531 15555
rect 16531 15521 16540 15555
rect 16488 15512 16540 15521
rect 13636 15487 13688 15496
rect 13636 15453 13645 15487
rect 13645 15453 13679 15487
rect 13679 15453 13688 15487
rect 13636 15444 13688 15453
rect 16672 15487 16724 15496
rect 7288 15308 7340 15360
rect 7656 15351 7708 15360
rect 7656 15317 7665 15351
rect 7665 15317 7699 15351
rect 7699 15317 7708 15351
rect 7656 15308 7708 15317
rect 8300 15308 8352 15360
rect 9496 15308 9548 15360
rect 12808 15308 12860 15360
rect 16672 15453 16681 15487
rect 16681 15453 16715 15487
rect 16715 15453 16724 15487
rect 16672 15444 16724 15453
rect 21548 15512 21600 15564
rect 22928 15555 22980 15564
rect 22928 15521 22937 15555
rect 22937 15521 22971 15555
rect 22971 15521 22980 15555
rect 22928 15512 22980 15521
rect 17960 15444 18012 15496
rect 18420 15444 18472 15496
rect 19708 15487 19760 15496
rect 19708 15453 19717 15487
rect 19717 15453 19751 15487
rect 19751 15453 19760 15487
rect 19708 15444 19760 15453
rect 17500 15376 17552 15428
rect 21180 15376 21232 15428
rect 22008 15444 22060 15496
rect 23020 15487 23072 15496
rect 23020 15453 23029 15487
rect 23029 15453 23063 15487
rect 23063 15453 23072 15487
rect 23020 15444 23072 15453
rect 23848 15444 23900 15496
rect 24032 15444 24084 15496
rect 25228 15444 25280 15496
rect 14648 15351 14700 15360
rect 14648 15317 14657 15351
rect 14657 15317 14691 15351
rect 14691 15317 14700 15351
rect 14648 15308 14700 15317
rect 15292 15308 15344 15360
rect 15936 15308 15988 15360
rect 17868 15308 17920 15360
rect 18604 15308 18656 15360
rect 19524 15308 19576 15360
rect 20904 15351 20956 15360
rect 20904 15317 20913 15351
rect 20913 15317 20947 15351
rect 20947 15317 20956 15351
rect 20904 15308 20956 15317
rect 23112 15308 23164 15360
rect 23388 15308 23440 15360
rect 25688 15308 25740 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 3056 15104 3108 15156
rect 5264 15104 5316 15156
rect 8760 15104 8812 15156
rect 11060 15104 11112 15156
rect 11152 15104 11204 15156
rect 12348 15104 12400 15156
rect 16396 15104 16448 15156
rect 2320 15079 2372 15088
rect 2320 15045 2329 15079
rect 2329 15045 2363 15079
rect 2363 15045 2372 15079
rect 2320 15036 2372 15045
rect 9128 15079 9180 15088
rect 9128 15045 9137 15079
rect 9137 15045 9171 15079
rect 9171 15045 9180 15079
rect 9128 15036 9180 15045
rect 12532 15036 12584 15088
rect 13820 15036 13872 15088
rect 1584 14900 1636 14952
rect 3792 14900 3844 14952
rect 1768 14875 1820 14884
rect 1768 14841 1777 14875
rect 1777 14841 1811 14875
rect 1811 14841 1820 14875
rect 1768 14832 1820 14841
rect 2504 14832 2556 14884
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 6920 14900 6972 14952
rect 4712 14764 4764 14816
rect 5080 14807 5132 14816
rect 5080 14773 5089 14807
rect 5089 14773 5123 14807
rect 5123 14773 5132 14807
rect 5080 14764 5132 14773
rect 6276 14807 6328 14816
rect 6276 14773 6285 14807
rect 6285 14773 6319 14807
rect 6319 14773 6328 14807
rect 6276 14764 6328 14773
rect 6368 14764 6420 14816
rect 6920 14764 6972 14816
rect 7564 14832 7616 14884
rect 10048 14900 10100 14952
rect 10784 14900 10836 14952
rect 11060 14900 11112 14952
rect 17040 14968 17092 15020
rect 17408 14968 17460 15020
rect 18236 15104 18288 15156
rect 18420 15104 18472 15156
rect 20444 15147 20496 15156
rect 20444 15113 20453 15147
rect 20453 15113 20487 15147
rect 20487 15113 20496 15147
rect 20444 15104 20496 15113
rect 20720 15104 20772 15156
rect 22376 15147 22428 15156
rect 22376 15113 22385 15147
rect 22385 15113 22419 15147
rect 22419 15113 22428 15147
rect 22376 15104 22428 15113
rect 23020 15147 23072 15156
rect 23020 15113 23029 15147
rect 23029 15113 23063 15147
rect 23063 15113 23072 15147
rect 23020 15104 23072 15113
rect 24676 15147 24728 15156
rect 24676 15113 24685 15147
rect 24685 15113 24719 15147
rect 24719 15113 24728 15147
rect 24676 15104 24728 15113
rect 26332 15147 26384 15156
rect 26332 15113 26341 15147
rect 26341 15113 26375 15147
rect 26375 15113 26384 15147
rect 26332 15104 26384 15113
rect 23572 15036 23624 15088
rect 19248 14968 19300 15020
rect 19432 14968 19484 15020
rect 24124 15011 24176 15020
rect 24124 14977 24133 15011
rect 24133 14977 24167 15011
rect 24167 14977 24176 15011
rect 24124 14968 24176 14977
rect 13912 14900 13964 14952
rect 14096 14900 14148 14952
rect 15568 14900 15620 14952
rect 15936 14900 15988 14952
rect 16396 14900 16448 14952
rect 17684 14900 17736 14952
rect 18604 14900 18656 14952
rect 20628 14900 20680 14952
rect 9772 14832 9824 14884
rect 14372 14832 14424 14884
rect 19340 14832 19392 14884
rect 19708 14832 19760 14884
rect 8116 14764 8168 14816
rect 8208 14807 8260 14816
rect 8208 14773 8217 14807
rect 8217 14773 8251 14807
rect 8251 14773 8260 14807
rect 10692 14807 10744 14816
rect 8208 14764 8260 14773
rect 10692 14773 10701 14807
rect 10701 14773 10735 14807
rect 10735 14773 10744 14807
rect 10692 14764 10744 14773
rect 11796 14807 11848 14816
rect 11796 14773 11805 14807
rect 11805 14773 11839 14807
rect 11839 14773 11848 14807
rect 11796 14764 11848 14773
rect 12440 14764 12492 14816
rect 13636 14764 13688 14816
rect 13728 14764 13780 14816
rect 14096 14764 14148 14816
rect 15568 14764 15620 14816
rect 16488 14807 16540 14816
rect 16488 14773 16497 14807
rect 16497 14773 16531 14807
rect 16531 14773 16540 14807
rect 16488 14764 16540 14773
rect 17040 14807 17092 14816
rect 17040 14773 17049 14807
rect 17049 14773 17083 14807
rect 17083 14773 17092 14807
rect 17040 14764 17092 14773
rect 18236 14764 18288 14816
rect 22008 14900 22060 14952
rect 25412 14900 25464 14952
rect 21180 14832 21232 14884
rect 23020 14832 23072 14884
rect 22928 14764 22980 14816
rect 24032 14807 24084 14816
rect 24032 14773 24041 14807
rect 24041 14773 24075 14807
rect 24075 14773 24084 14807
rect 24032 14764 24084 14773
rect 24952 14832 25004 14884
rect 25688 14764 25740 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1400 14603 1452 14612
rect 1400 14569 1409 14603
rect 1409 14569 1443 14603
rect 1443 14569 1452 14603
rect 1400 14560 1452 14569
rect 2504 14603 2556 14612
rect 2504 14569 2513 14603
rect 2513 14569 2547 14603
rect 2547 14569 2556 14603
rect 2504 14560 2556 14569
rect 3056 14560 3108 14612
rect 5356 14560 5408 14612
rect 7104 14560 7156 14612
rect 9220 14603 9272 14612
rect 9220 14569 9229 14603
rect 9229 14569 9263 14603
rect 9263 14569 9272 14603
rect 9220 14560 9272 14569
rect 9588 14560 9640 14612
rect 13268 14560 13320 14612
rect 13544 14560 13596 14612
rect 16488 14560 16540 14612
rect 17500 14560 17552 14612
rect 17960 14603 18012 14612
rect 17960 14569 17969 14603
rect 17969 14569 18003 14603
rect 18003 14569 18012 14603
rect 17960 14560 18012 14569
rect 19340 14603 19392 14612
rect 19340 14569 19349 14603
rect 19349 14569 19383 14603
rect 19383 14569 19392 14603
rect 19340 14560 19392 14569
rect 19984 14560 20036 14612
rect 20628 14560 20680 14612
rect 21180 14560 21232 14612
rect 21916 14560 21968 14612
rect 22928 14560 22980 14612
rect 1676 14492 1728 14544
rect 2412 14492 2464 14544
rect 3792 14492 3844 14544
rect 4896 14492 4948 14544
rect 5448 14492 5500 14544
rect 7196 14492 7248 14544
rect 7380 14492 7432 14544
rect 8024 14535 8076 14544
rect 8024 14501 8033 14535
rect 8033 14501 8067 14535
rect 8067 14501 8076 14535
rect 8024 14492 8076 14501
rect 10692 14535 10744 14544
rect 10692 14501 10726 14535
rect 10726 14501 10744 14535
rect 10692 14492 10744 14501
rect 15476 14492 15528 14544
rect 15752 14492 15804 14544
rect 17224 14492 17276 14544
rect 18144 14492 18196 14544
rect 18420 14492 18472 14544
rect 21364 14492 21416 14544
rect 4712 14424 4764 14476
rect 8116 14467 8168 14476
rect 8116 14433 8125 14467
rect 8125 14433 8159 14467
rect 8159 14433 8168 14467
rect 8116 14424 8168 14433
rect 9312 14424 9364 14476
rect 11704 14424 11756 14476
rect 12532 14424 12584 14476
rect 16396 14424 16448 14476
rect 16856 14424 16908 14476
rect 17960 14424 18012 14476
rect 18972 14424 19024 14476
rect 20076 14424 20128 14476
rect 21640 14467 21692 14476
rect 21640 14433 21649 14467
rect 21649 14433 21683 14467
rect 21683 14433 21692 14467
rect 21640 14424 21692 14433
rect 23296 14492 23348 14544
rect 1860 14399 1912 14408
rect 1860 14365 1869 14399
rect 1869 14365 1903 14399
rect 1903 14365 1912 14399
rect 1860 14356 1912 14365
rect 2504 14356 2556 14408
rect 3976 14356 4028 14408
rect 6276 14356 6328 14408
rect 8208 14356 8260 14408
rect 8760 14356 8812 14408
rect 9772 14356 9824 14408
rect 12440 14399 12492 14408
rect 12440 14365 12449 14399
rect 12449 14365 12483 14399
rect 12483 14365 12492 14399
rect 12440 14356 12492 14365
rect 1032 14288 1084 14340
rect 5540 14288 5592 14340
rect 7012 14288 7064 14340
rect 7932 14288 7984 14340
rect 8024 14288 8076 14340
rect 12808 14331 12860 14340
rect 12808 14297 12817 14331
rect 12817 14297 12851 14331
rect 12851 14297 12860 14331
rect 15844 14356 15896 14408
rect 12808 14288 12860 14297
rect 13544 14288 13596 14340
rect 15476 14288 15528 14340
rect 16672 14288 16724 14340
rect 17224 14356 17276 14408
rect 18604 14399 18656 14408
rect 18604 14365 18613 14399
rect 18613 14365 18647 14399
rect 18647 14365 18656 14399
rect 18604 14356 18656 14365
rect 22284 14356 22336 14408
rect 24032 14560 24084 14612
rect 24584 14560 24636 14612
rect 26148 14560 26200 14612
rect 23572 14492 23624 14544
rect 24124 14535 24176 14544
rect 24124 14501 24158 14535
rect 24158 14501 24176 14535
rect 24124 14492 24176 14501
rect 24860 14492 24912 14544
rect 26332 14560 26384 14612
rect 23848 14399 23900 14408
rect 23848 14365 23857 14399
rect 23857 14365 23891 14399
rect 23891 14365 23900 14399
rect 23848 14356 23900 14365
rect 2964 14220 3016 14272
rect 5356 14220 5408 14272
rect 6368 14220 6420 14272
rect 7840 14220 7892 14272
rect 8760 14263 8812 14272
rect 8760 14229 8769 14263
rect 8769 14229 8803 14263
rect 8803 14229 8812 14263
rect 8760 14220 8812 14229
rect 9772 14220 9824 14272
rect 9956 14220 10008 14272
rect 12900 14263 12952 14272
rect 12900 14229 12909 14263
rect 12909 14229 12943 14263
rect 12943 14229 12952 14263
rect 12900 14220 12952 14229
rect 14004 14263 14056 14272
rect 14004 14229 14013 14263
rect 14013 14229 14047 14263
rect 14047 14229 14056 14263
rect 14004 14220 14056 14229
rect 14096 14220 14148 14272
rect 14648 14263 14700 14272
rect 14648 14229 14657 14263
rect 14657 14229 14691 14263
rect 14691 14229 14700 14263
rect 14648 14220 14700 14229
rect 15292 14220 15344 14272
rect 21548 14220 21600 14272
rect 25228 14263 25280 14272
rect 25228 14229 25237 14263
rect 25237 14229 25271 14263
rect 25271 14229 25280 14263
rect 25228 14220 25280 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 2504 14016 2556 14068
rect 3148 14016 3200 14068
rect 4252 14059 4304 14068
rect 4252 14025 4261 14059
rect 4261 14025 4295 14059
rect 4295 14025 4304 14059
rect 4252 14016 4304 14025
rect 5172 14059 5224 14068
rect 5172 14025 5181 14059
rect 5181 14025 5215 14059
rect 5215 14025 5224 14059
rect 5172 14016 5224 14025
rect 8484 14059 8536 14068
rect 8484 14025 8493 14059
rect 8493 14025 8527 14059
rect 8527 14025 8536 14059
rect 8484 14016 8536 14025
rect 10048 14059 10100 14068
rect 10048 14025 10057 14059
rect 10057 14025 10091 14059
rect 10091 14025 10100 14059
rect 10048 14016 10100 14025
rect 10692 14016 10744 14068
rect 11796 14016 11848 14068
rect 13268 14016 13320 14068
rect 13728 14016 13780 14068
rect 14372 14016 14424 14068
rect 16856 14016 16908 14068
rect 17224 14016 17276 14068
rect 18052 14016 18104 14068
rect 18236 14016 18288 14068
rect 20812 14059 20864 14068
rect 20812 14025 20821 14059
rect 20821 14025 20855 14059
rect 20855 14025 20864 14059
rect 20812 14016 20864 14025
rect 23112 14016 23164 14068
rect 24860 14016 24912 14068
rect 25688 14059 25740 14068
rect 25688 14025 25697 14059
rect 25697 14025 25731 14059
rect 25731 14025 25740 14059
rect 25688 14016 25740 14025
rect 26332 14059 26384 14068
rect 26332 14025 26341 14059
rect 26341 14025 26375 14059
rect 26375 14025 26384 14059
rect 26332 14016 26384 14025
rect 2688 13948 2740 14000
rect 4712 13991 4764 14000
rect 4712 13957 4721 13991
rect 4721 13957 4755 13991
rect 4755 13957 4764 13991
rect 4712 13948 4764 13957
rect 6828 13991 6880 14000
rect 1584 13923 1636 13932
rect 1584 13889 1593 13923
rect 1593 13889 1627 13923
rect 1627 13889 1636 13923
rect 1584 13880 1636 13889
rect 2780 13880 2832 13932
rect 6828 13957 6837 13991
rect 6837 13957 6871 13991
rect 6871 13957 6880 13991
rect 6828 13948 6880 13957
rect 6920 13948 6972 14000
rect 8300 13948 8352 14000
rect 2320 13812 2372 13864
rect 2964 13812 3016 13864
rect 2504 13744 2556 13796
rect 4712 13812 4764 13864
rect 6276 13880 6328 13932
rect 7288 13923 7340 13932
rect 7288 13889 7297 13923
rect 7297 13889 7331 13923
rect 7331 13889 7340 13923
rect 7288 13880 7340 13889
rect 8944 13923 8996 13932
rect 5908 13812 5960 13864
rect 2780 13676 2832 13728
rect 3240 13676 3292 13728
rect 5540 13719 5592 13728
rect 5540 13685 5549 13719
rect 5549 13685 5583 13719
rect 5583 13685 5592 13719
rect 5540 13676 5592 13685
rect 6368 13812 6420 13864
rect 8944 13889 8953 13923
rect 8953 13889 8987 13923
rect 8987 13889 8996 13923
rect 8944 13880 8996 13889
rect 9588 13948 9640 14000
rect 9956 13948 10008 14000
rect 15384 13948 15436 14000
rect 15844 13948 15896 14000
rect 11704 13880 11756 13932
rect 12256 13880 12308 13932
rect 10968 13812 11020 13864
rect 11428 13855 11480 13864
rect 11428 13821 11437 13855
rect 11437 13821 11471 13855
rect 11471 13821 11480 13855
rect 11428 13812 11480 13821
rect 6092 13744 6144 13796
rect 6276 13744 6328 13796
rect 9404 13744 9456 13796
rect 12532 13744 12584 13796
rect 13912 13744 13964 13796
rect 14004 13744 14056 13796
rect 8760 13676 8812 13728
rect 9680 13676 9732 13728
rect 10692 13676 10744 13728
rect 14188 13676 14240 13728
rect 16672 13880 16724 13932
rect 16856 13855 16908 13864
rect 16856 13821 16865 13855
rect 16865 13821 16899 13855
rect 16899 13821 16908 13855
rect 16856 13812 16908 13821
rect 17224 13812 17276 13864
rect 17960 13948 18012 14000
rect 22284 13991 22336 14000
rect 17684 13880 17736 13932
rect 20720 13923 20772 13932
rect 20720 13889 20729 13923
rect 20729 13889 20763 13923
rect 20763 13889 20772 13923
rect 21364 13923 21416 13932
rect 20720 13880 20772 13889
rect 18052 13855 18104 13864
rect 18052 13821 18061 13855
rect 18061 13821 18095 13855
rect 18095 13821 18104 13855
rect 18052 13812 18104 13821
rect 18144 13812 18196 13864
rect 21364 13889 21373 13923
rect 21373 13889 21407 13923
rect 21407 13889 21416 13923
rect 21364 13880 21416 13889
rect 22284 13957 22293 13991
rect 22293 13957 22327 13991
rect 22327 13957 22336 13991
rect 22284 13948 22336 13957
rect 26240 13880 26292 13932
rect 21732 13812 21784 13864
rect 21916 13855 21968 13864
rect 21916 13821 21925 13855
rect 21925 13821 21959 13855
rect 21959 13821 21968 13855
rect 21916 13812 21968 13821
rect 22100 13812 22152 13864
rect 15844 13676 15896 13728
rect 16396 13719 16448 13728
rect 16396 13685 16405 13719
rect 16405 13685 16439 13719
rect 16439 13685 16448 13719
rect 16396 13676 16448 13685
rect 18420 13676 18472 13728
rect 23940 13855 23992 13864
rect 23940 13821 23974 13855
rect 23974 13821 23992 13855
rect 23572 13744 23624 13796
rect 23940 13812 23992 13821
rect 23848 13744 23900 13796
rect 23756 13676 23808 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 5540 13472 5592 13524
rect 5724 13515 5776 13524
rect 5724 13481 5733 13515
rect 5733 13481 5767 13515
rect 5767 13481 5776 13515
rect 5724 13472 5776 13481
rect 7196 13472 7248 13524
rect 7472 13472 7524 13524
rect 8944 13472 8996 13524
rect 9220 13515 9272 13524
rect 9220 13481 9229 13515
rect 9229 13481 9263 13515
rect 9263 13481 9272 13515
rect 9220 13472 9272 13481
rect 10968 13472 11020 13524
rect 12532 13472 12584 13524
rect 13268 13472 13320 13524
rect 16028 13472 16080 13524
rect 17500 13472 17552 13524
rect 17592 13472 17644 13524
rect 17960 13472 18012 13524
rect 20352 13472 20404 13524
rect 21088 13472 21140 13524
rect 21640 13515 21692 13524
rect 21640 13481 21649 13515
rect 21649 13481 21683 13515
rect 21683 13481 21692 13515
rect 21640 13472 21692 13481
rect 23940 13472 23992 13524
rect 25044 13472 25096 13524
rect 26332 13472 26384 13524
rect 2044 13404 2096 13456
rect 3976 13404 4028 13456
rect 6736 13404 6788 13456
rect 8300 13404 8352 13456
rect 9956 13447 10008 13456
rect 9956 13413 9990 13447
rect 9990 13413 10008 13447
rect 9956 13404 10008 13413
rect 10600 13404 10652 13456
rect 10784 13404 10836 13456
rect 11796 13404 11848 13456
rect 13544 13404 13596 13456
rect 13820 13404 13872 13456
rect 14464 13404 14516 13456
rect 15384 13404 15436 13456
rect 17684 13447 17736 13456
rect 17684 13413 17693 13447
rect 17693 13413 17727 13447
rect 17727 13413 17736 13447
rect 17684 13404 17736 13413
rect 18604 13404 18656 13456
rect 20076 13404 20128 13456
rect 21364 13404 21416 13456
rect 22284 13404 22336 13456
rect 22560 13404 22612 13456
rect 1492 13336 1544 13388
rect 1676 13379 1728 13388
rect 1676 13345 1710 13379
rect 1710 13345 1728 13379
rect 1676 13336 1728 13345
rect 4712 13268 4764 13320
rect 5356 13336 5408 13388
rect 5448 13336 5500 13388
rect 8392 13336 8444 13388
rect 8760 13336 8812 13388
rect 9220 13336 9272 13388
rect 9588 13336 9640 13388
rect 12164 13336 12216 13388
rect 7932 13268 7984 13320
rect 13912 13336 13964 13388
rect 15200 13336 15252 13388
rect 15568 13379 15620 13388
rect 15568 13345 15602 13379
rect 15602 13345 15620 13379
rect 15568 13336 15620 13345
rect 18236 13379 18288 13388
rect 18236 13345 18245 13379
rect 18245 13345 18279 13379
rect 18279 13345 18288 13379
rect 18236 13336 18288 13345
rect 12808 13311 12860 13320
rect 3148 13200 3200 13252
rect 2964 13132 3016 13184
rect 3332 13175 3384 13184
rect 3332 13141 3341 13175
rect 3341 13141 3375 13175
rect 3375 13141 3384 13175
rect 3332 13132 3384 13141
rect 3700 13175 3752 13184
rect 3700 13141 3709 13175
rect 3709 13141 3743 13175
rect 3743 13141 3752 13175
rect 3700 13132 3752 13141
rect 8392 13200 8444 13252
rect 9588 13200 9640 13252
rect 10784 13200 10836 13252
rect 12808 13277 12817 13311
rect 12817 13277 12851 13311
rect 12851 13277 12860 13311
rect 12808 13268 12860 13277
rect 14188 13311 14240 13320
rect 14188 13277 14197 13311
rect 14197 13277 14231 13311
rect 14231 13277 14240 13311
rect 14188 13268 14240 13277
rect 18420 13311 18472 13320
rect 18420 13277 18429 13311
rect 18429 13277 18463 13311
rect 18463 13277 18472 13311
rect 18420 13268 18472 13277
rect 20812 13336 20864 13388
rect 22008 13336 22060 13388
rect 23572 13336 23624 13388
rect 21824 13268 21876 13320
rect 25044 13311 25096 13320
rect 25044 13277 25053 13311
rect 25053 13277 25087 13311
rect 25087 13277 25096 13311
rect 25044 13268 25096 13277
rect 11796 13200 11848 13252
rect 24768 13200 24820 13252
rect 8300 13132 8352 13184
rect 11060 13175 11112 13184
rect 11060 13141 11069 13175
rect 11069 13141 11103 13175
rect 11103 13141 11112 13175
rect 11060 13132 11112 13141
rect 11152 13132 11204 13184
rect 16672 13175 16724 13184
rect 16672 13141 16681 13175
rect 16681 13141 16715 13175
rect 16715 13141 16724 13175
rect 16672 13132 16724 13141
rect 24124 13132 24176 13184
rect 25596 13175 25648 13184
rect 25596 13141 25605 13175
rect 25605 13141 25639 13175
rect 25639 13141 25648 13175
rect 25596 13132 25648 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 1860 12928 1912 12980
rect 3976 12971 4028 12980
rect 1584 12835 1636 12844
rect 1584 12801 1593 12835
rect 1593 12801 1627 12835
rect 1627 12801 1636 12835
rect 1584 12792 1636 12801
rect 3976 12937 3985 12971
rect 3985 12937 4019 12971
rect 4019 12937 4028 12971
rect 3976 12928 4028 12937
rect 4896 12971 4948 12980
rect 4896 12937 4905 12971
rect 4905 12937 4939 12971
rect 4939 12937 4948 12971
rect 4896 12928 4948 12937
rect 6644 12971 6696 12980
rect 6644 12937 6653 12971
rect 6653 12937 6687 12971
rect 6687 12937 6696 12971
rect 6644 12928 6696 12937
rect 7564 12928 7616 12980
rect 9588 12928 9640 12980
rect 9864 12971 9916 12980
rect 9864 12937 9873 12971
rect 9873 12937 9907 12971
rect 9907 12937 9916 12971
rect 9864 12928 9916 12937
rect 9956 12928 10008 12980
rect 11704 12928 11756 12980
rect 12164 12928 12216 12980
rect 12532 12928 12584 12980
rect 3608 12724 3660 12776
rect 3884 12724 3936 12776
rect 1952 12656 2004 12708
rect 3056 12656 3108 12708
rect 5356 12792 5408 12844
rect 1216 12588 1268 12640
rect 1400 12588 1452 12640
rect 1676 12588 1728 12640
rect 2688 12588 2740 12640
rect 3516 12631 3568 12640
rect 3516 12597 3525 12631
rect 3525 12597 3559 12631
rect 3559 12597 3568 12631
rect 3516 12588 3568 12597
rect 3608 12588 3660 12640
rect 4436 12588 4488 12640
rect 4712 12631 4764 12640
rect 4712 12597 4721 12631
rect 4721 12597 4755 12631
rect 4755 12597 4764 12631
rect 4712 12588 4764 12597
rect 4988 12656 5040 12708
rect 6736 12860 6788 12912
rect 7656 12792 7708 12844
rect 9956 12792 10008 12844
rect 10692 12792 10744 12844
rect 7380 12724 7432 12776
rect 8300 12767 8352 12776
rect 8300 12733 8309 12767
rect 8309 12733 8343 12767
rect 8343 12733 8352 12767
rect 8300 12724 8352 12733
rect 9220 12724 9272 12776
rect 10048 12724 10100 12776
rect 10600 12724 10652 12776
rect 6644 12656 6696 12708
rect 10692 12656 10744 12708
rect 11336 12835 11388 12844
rect 11336 12801 11345 12835
rect 11345 12801 11379 12835
rect 11379 12801 11388 12835
rect 11336 12792 11388 12801
rect 12716 12792 12768 12844
rect 13268 12792 13320 12844
rect 14740 12928 14792 12980
rect 15292 12928 15344 12980
rect 16304 12928 16356 12980
rect 17500 12971 17552 12980
rect 17500 12937 17509 12971
rect 17509 12937 17543 12971
rect 17543 12937 17552 12971
rect 17500 12928 17552 12937
rect 18420 12971 18472 12980
rect 18420 12937 18429 12971
rect 18429 12937 18463 12971
rect 18463 12937 18472 12971
rect 18420 12928 18472 12937
rect 20996 12971 21048 12980
rect 20996 12937 21005 12971
rect 21005 12937 21039 12971
rect 21039 12937 21048 12971
rect 20996 12928 21048 12937
rect 23756 12928 23808 12980
rect 24768 12971 24820 12980
rect 24768 12937 24777 12971
rect 24777 12937 24811 12971
rect 24811 12937 24820 12971
rect 24768 12928 24820 12937
rect 25136 12928 25188 12980
rect 26240 12928 26292 12980
rect 15568 12860 15620 12912
rect 15660 12860 15712 12912
rect 15844 12860 15896 12912
rect 15384 12835 15436 12844
rect 15384 12801 15393 12835
rect 15393 12801 15427 12835
rect 15427 12801 15436 12835
rect 15384 12792 15436 12801
rect 16212 12835 16264 12844
rect 16212 12801 16221 12835
rect 16221 12801 16255 12835
rect 16255 12801 16264 12835
rect 16212 12792 16264 12801
rect 12440 12724 12492 12776
rect 10784 12631 10836 12640
rect 10784 12597 10793 12631
rect 10793 12597 10827 12631
rect 10827 12597 10836 12631
rect 10784 12588 10836 12597
rect 12624 12656 12676 12708
rect 13544 12724 13596 12776
rect 15108 12724 15160 12776
rect 15476 12724 15528 12776
rect 20076 12860 20128 12912
rect 24676 12860 24728 12912
rect 18236 12724 18288 12776
rect 21640 12835 21692 12844
rect 21640 12801 21649 12835
rect 21649 12801 21683 12835
rect 21683 12801 21692 12835
rect 21640 12792 21692 12801
rect 23204 12792 23256 12844
rect 25044 12835 25096 12844
rect 20260 12724 20312 12776
rect 20996 12724 21048 12776
rect 22284 12724 22336 12776
rect 23112 12724 23164 12776
rect 24124 12724 24176 12776
rect 13268 12631 13320 12640
rect 13268 12597 13277 12631
rect 13277 12597 13311 12631
rect 13311 12597 13320 12631
rect 13268 12588 13320 12597
rect 15200 12631 15252 12640
rect 15200 12597 15209 12631
rect 15209 12597 15243 12631
rect 15243 12597 15252 12631
rect 15200 12588 15252 12597
rect 16304 12656 16356 12708
rect 23572 12656 23624 12708
rect 25044 12801 25053 12835
rect 25053 12801 25087 12835
rect 25087 12801 25096 12835
rect 25044 12792 25096 12801
rect 25504 12835 25556 12844
rect 25504 12801 25513 12835
rect 25513 12801 25547 12835
rect 25547 12801 25556 12835
rect 25504 12792 25556 12801
rect 25136 12724 25188 12776
rect 25596 12724 25648 12776
rect 18052 12588 18104 12640
rect 20536 12588 20588 12640
rect 20812 12631 20864 12640
rect 20812 12597 20821 12631
rect 20821 12597 20855 12631
rect 20855 12597 20864 12631
rect 20812 12588 20864 12597
rect 21180 12588 21232 12640
rect 23388 12588 23440 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 1400 12427 1452 12436
rect 1400 12393 1409 12427
rect 1409 12393 1443 12427
rect 1443 12393 1452 12427
rect 1400 12384 1452 12393
rect 2136 12384 2188 12436
rect 3424 12427 3476 12436
rect 3424 12393 3433 12427
rect 3433 12393 3467 12427
rect 3467 12393 3476 12427
rect 3424 12384 3476 12393
rect 4160 12384 4212 12436
rect 6736 12384 6788 12436
rect 7463 12384 7515 12436
rect 8024 12384 8076 12436
rect 9128 12427 9180 12436
rect 1676 12112 1728 12164
rect 2044 12112 2096 12164
rect 1400 12044 1452 12096
rect 2688 12316 2740 12368
rect 5540 12316 5592 12368
rect 6276 12316 6328 12368
rect 9128 12393 9137 12427
rect 9137 12393 9171 12427
rect 9171 12393 9180 12427
rect 9128 12384 9180 12393
rect 9680 12384 9732 12436
rect 11244 12384 11296 12436
rect 12440 12384 12492 12436
rect 12716 12384 12768 12436
rect 15108 12427 15160 12436
rect 15108 12393 15117 12427
rect 15117 12393 15151 12427
rect 15151 12393 15160 12427
rect 15108 12384 15160 12393
rect 15200 12384 15252 12436
rect 16396 12384 16448 12436
rect 16672 12384 16724 12436
rect 17500 12384 17552 12436
rect 21364 12384 21416 12436
rect 9036 12316 9088 12368
rect 9864 12359 9916 12368
rect 9864 12325 9873 12359
rect 9873 12325 9907 12359
rect 9907 12325 9916 12359
rect 9864 12316 9916 12325
rect 9956 12316 10008 12368
rect 10232 12316 10284 12368
rect 3884 12248 3936 12300
rect 4252 12248 4304 12300
rect 5448 12291 5500 12300
rect 5448 12257 5457 12291
rect 5457 12257 5491 12291
rect 5491 12257 5500 12291
rect 5448 12248 5500 12257
rect 3056 12223 3108 12232
rect 3056 12189 3065 12223
rect 3065 12189 3099 12223
rect 3099 12189 3108 12223
rect 3056 12180 3108 12189
rect 3608 12180 3660 12232
rect 6920 12248 6972 12300
rect 7840 12248 7892 12300
rect 9128 12248 9180 12300
rect 10784 12316 10836 12368
rect 11428 12316 11480 12368
rect 11244 12291 11296 12300
rect 11244 12257 11253 12291
rect 11253 12257 11287 12291
rect 11287 12257 11296 12291
rect 11244 12248 11296 12257
rect 12164 12248 12216 12300
rect 14004 12248 14056 12300
rect 7104 12180 7156 12232
rect 7564 12180 7616 12232
rect 7748 12180 7800 12232
rect 8484 12223 8536 12232
rect 8484 12189 8493 12223
rect 8493 12189 8527 12223
rect 8527 12189 8536 12223
rect 8484 12180 8536 12189
rect 8668 12223 8720 12232
rect 8668 12189 8677 12223
rect 8677 12189 8711 12223
rect 8711 12189 8720 12223
rect 8668 12180 8720 12189
rect 9864 12180 9916 12232
rect 10140 12180 10192 12232
rect 4988 12087 5040 12096
rect 4988 12053 4997 12087
rect 4997 12053 5031 12087
rect 5031 12053 5040 12087
rect 4988 12044 5040 12053
rect 5356 12087 5408 12096
rect 5356 12053 5365 12087
rect 5365 12053 5399 12087
rect 5399 12053 5408 12087
rect 11152 12112 11204 12164
rect 11888 12180 11940 12232
rect 12256 12112 12308 12164
rect 13728 12112 13780 12164
rect 17868 12316 17920 12368
rect 18420 12316 18472 12368
rect 14740 12248 14792 12300
rect 15384 12248 15436 12300
rect 16856 12248 16908 12300
rect 19524 12291 19576 12300
rect 19524 12257 19533 12291
rect 19533 12257 19567 12291
rect 19567 12257 19576 12291
rect 19524 12248 19576 12257
rect 15936 12180 15988 12232
rect 20076 12180 20128 12232
rect 20904 12180 20956 12232
rect 21180 12180 21232 12232
rect 22284 12384 22336 12436
rect 22836 12427 22888 12436
rect 22836 12393 22845 12427
rect 22845 12393 22879 12427
rect 22879 12393 22888 12427
rect 22836 12384 22888 12393
rect 23296 12384 23348 12436
rect 24308 12384 24360 12436
rect 25044 12384 25096 12436
rect 26332 12384 26384 12436
rect 23204 12316 23256 12368
rect 24952 12316 25004 12368
rect 23848 12248 23900 12300
rect 24860 12248 24912 12300
rect 22376 12180 22428 12232
rect 21456 12112 21508 12164
rect 22744 12112 22796 12164
rect 5356 12044 5408 12053
rect 7104 12044 7156 12096
rect 8024 12087 8076 12096
rect 8024 12053 8033 12087
rect 8033 12053 8067 12087
rect 8067 12053 8076 12087
rect 8024 12044 8076 12053
rect 9772 12044 9824 12096
rect 12992 12044 13044 12096
rect 14096 12044 14148 12096
rect 14464 12044 14516 12096
rect 15936 12087 15988 12096
rect 15936 12053 15945 12087
rect 15945 12053 15979 12087
rect 15979 12053 15988 12087
rect 15936 12044 15988 12053
rect 16672 12044 16724 12096
rect 17408 12087 17460 12096
rect 17408 12053 17417 12087
rect 17417 12053 17451 12087
rect 17451 12053 17460 12087
rect 17408 12044 17460 12053
rect 18972 12087 19024 12096
rect 18972 12053 18981 12087
rect 18981 12053 19015 12087
rect 19015 12053 19024 12087
rect 18972 12044 19024 12053
rect 20444 12044 20496 12096
rect 22008 12044 22060 12096
rect 24768 12044 24820 12096
rect 25504 12044 25556 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 3240 11840 3292 11892
rect 5540 11883 5592 11892
rect 5540 11849 5549 11883
rect 5549 11849 5583 11883
rect 5583 11849 5592 11883
rect 5540 11840 5592 11849
rect 3424 11772 3476 11824
rect 9128 11840 9180 11892
rect 9772 11840 9824 11892
rect 10324 11883 10376 11892
rect 10324 11849 10333 11883
rect 10333 11849 10367 11883
rect 10367 11849 10376 11883
rect 10324 11840 10376 11849
rect 10876 11840 10928 11892
rect 11888 11883 11940 11892
rect 11888 11849 11897 11883
rect 11897 11849 11931 11883
rect 11931 11849 11940 11883
rect 11888 11840 11940 11849
rect 13636 11840 13688 11892
rect 16212 11840 16264 11892
rect 16396 11883 16448 11892
rect 16396 11849 16405 11883
rect 16405 11849 16439 11883
rect 16439 11849 16448 11883
rect 16396 11840 16448 11849
rect 17500 11883 17552 11892
rect 17500 11849 17509 11883
rect 17509 11849 17543 11883
rect 17543 11849 17552 11883
rect 17500 11840 17552 11849
rect 3608 11704 3660 11756
rect 2228 11636 2280 11688
rect 4160 11679 4212 11688
rect 4160 11645 4169 11679
rect 4169 11645 4203 11679
rect 4203 11645 4212 11679
rect 14096 11772 14148 11824
rect 16580 11772 16632 11824
rect 21272 11772 21324 11824
rect 23572 11840 23624 11892
rect 25320 11840 25372 11892
rect 21916 11772 21968 11824
rect 7288 11747 7340 11756
rect 7288 11713 7297 11747
rect 7297 11713 7331 11747
rect 7331 11713 7340 11747
rect 7288 11704 7340 11713
rect 4160 11636 4212 11645
rect 7104 11636 7156 11688
rect 9680 11704 9732 11756
rect 9496 11636 9548 11688
rect 9772 11636 9824 11688
rect 10876 11704 10928 11756
rect 15936 11704 15988 11756
rect 16856 11704 16908 11756
rect 18604 11747 18656 11756
rect 18604 11713 18613 11747
rect 18613 11713 18647 11747
rect 18647 11713 18656 11747
rect 18604 11704 18656 11713
rect 11612 11636 11664 11688
rect 11888 11636 11940 11688
rect 12072 11636 12124 11688
rect 12256 11636 12308 11688
rect 13912 11636 13964 11688
rect 14556 11636 14608 11688
rect 3884 11568 3936 11620
rect 5448 11568 5500 11620
rect 8116 11568 8168 11620
rect 2596 11543 2648 11552
rect 2596 11509 2605 11543
rect 2605 11509 2639 11543
rect 2639 11509 2648 11543
rect 2596 11500 2648 11509
rect 3424 11500 3476 11552
rect 4252 11500 4304 11552
rect 6184 11543 6236 11552
rect 6184 11509 6193 11543
rect 6193 11509 6227 11543
rect 6227 11509 6236 11543
rect 6184 11500 6236 11509
rect 6828 11543 6880 11552
rect 6828 11509 6837 11543
rect 6837 11509 6871 11543
rect 6871 11509 6880 11543
rect 6828 11500 6880 11509
rect 7012 11500 7064 11552
rect 7656 11500 7708 11552
rect 7840 11543 7892 11552
rect 7840 11509 7849 11543
rect 7849 11509 7883 11543
rect 7883 11509 7892 11543
rect 7840 11500 7892 11509
rect 8208 11543 8260 11552
rect 8208 11509 8217 11543
rect 8217 11509 8251 11543
rect 8251 11509 8260 11543
rect 8208 11500 8260 11509
rect 8300 11500 8352 11552
rect 8484 11500 8536 11552
rect 10876 11568 10928 11620
rect 11060 11568 11112 11620
rect 12164 11611 12216 11620
rect 10784 11543 10836 11552
rect 10784 11509 10793 11543
rect 10793 11509 10827 11543
rect 10827 11509 10836 11543
rect 10784 11500 10836 11509
rect 11152 11500 11204 11552
rect 12164 11577 12173 11611
rect 12173 11577 12207 11611
rect 12207 11577 12216 11611
rect 12164 11568 12216 11577
rect 13176 11568 13228 11620
rect 16764 11636 16816 11688
rect 20260 11704 20312 11756
rect 20444 11747 20496 11756
rect 20444 11713 20453 11747
rect 20453 11713 20487 11747
rect 20487 11713 20496 11747
rect 20444 11704 20496 11713
rect 21456 11747 21508 11756
rect 19984 11636 20036 11688
rect 21456 11713 21465 11747
rect 21465 11713 21499 11747
rect 21499 11713 21508 11747
rect 21456 11704 21508 11713
rect 22008 11747 22060 11756
rect 22008 11713 22017 11747
rect 22017 11713 22051 11747
rect 22051 11713 22060 11747
rect 22008 11704 22060 11713
rect 23756 11772 23808 11824
rect 20904 11636 20956 11688
rect 22468 11636 22520 11688
rect 24860 11636 24912 11688
rect 25228 11679 25280 11688
rect 25228 11645 25237 11679
rect 25237 11645 25271 11679
rect 25271 11645 25280 11679
rect 25228 11636 25280 11645
rect 15660 11568 15712 11620
rect 14740 11500 14792 11552
rect 15476 11543 15528 11552
rect 15476 11509 15485 11543
rect 15485 11509 15519 11543
rect 15519 11509 15528 11543
rect 15476 11500 15528 11509
rect 15568 11500 15620 11552
rect 16672 11568 16724 11620
rect 15844 11500 15896 11552
rect 17224 11568 17276 11620
rect 17316 11568 17368 11620
rect 17500 11568 17552 11620
rect 17960 11568 18012 11620
rect 20076 11568 20128 11620
rect 20628 11568 20680 11620
rect 18052 11543 18104 11552
rect 18052 11509 18061 11543
rect 18061 11509 18095 11543
rect 18095 11509 18104 11543
rect 18052 11500 18104 11509
rect 20812 11500 20864 11552
rect 21180 11500 21232 11552
rect 23756 11568 23808 11620
rect 23572 11500 23624 11552
rect 25504 11500 25556 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 2688 11296 2740 11348
rect 2780 11296 2832 11348
rect 3332 11296 3384 11348
rect 3884 11339 3936 11348
rect 3884 11305 3893 11339
rect 3893 11305 3927 11339
rect 3927 11305 3936 11339
rect 3884 11296 3936 11305
rect 5540 11296 5592 11348
rect 6368 11296 6420 11348
rect 7748 11339 7800 11348
rect 7748 11305 7757 11339
rect 7757 11305 7791 11339
rect 7791 11305 7800 11339
rect 7748 11296 7800 11305
rect 8576 11339 8628 11348
rect 8576 11305 8585 11339
rect 8585 11305 8619 11339
rect 8619 11305 8628 11339
rect 8576 11296 8628 11305
rect 9312 11296 9364 11348
rect 11060 11296 11112 11348
rect 11520 11296 11572 11348
rect 12440 11296 12492 11348
rect 12808 11296 12860 11348
rect 13176 11339 13228 11348
rect 13176 11305 13185 11339
rect 13185 11305 13219 11339
rect 13219 11305 13228 11339
rect 13176 11296 13228 11305
rect 16488 11296 16540 11348
rect 18236 11296 18288 11348
rect 20168 11296 20220 11348
rect 20628 11296 20680 11348
rect 21916 11339 21968 11348
rect 21916 11305 21925 11339
rect 21925 11305 21959 11339
rect 21959 11305 21968 11339
rect 21916 11296 21968 11305
rect 22008 11296 22060 11348
rect 22652 11339 22704 11348
rect 22652 11305 22661 11339
rect 22661 11305 22695 11339
rect 22695 11305 22704 11339
rect 22652 11296 22704 11305
rect 23204 11296 23256 11348
rect 3056 11228 3108 11280
rect 3608 11228 3660 11280
rect 5356 11228 5408 11280
rect 7012 11228 7064 11280
rect 8484 11271 8536 11280
rect 8484 11237 8493 11271
rect 8493 11237 8527 11271
rect 8527 11237 8536 11271
rect 8484 11228 8536 11237
rect 3148 11160 3200 11212
rect 3700 11160 3752 11212
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 2504 11092 2556 11144
rect 3884 11092 3936 11144
rect 2688 11024 2740 11076
rect 2872 11024 2924 11076
rect 3332 11024 3384 11076
rect 3700 11024 3752 11076
rect 4160 11160 4212 11212
rect 4712 11160 4764 11212
rect 6644 11092 6696 11144
rect 10600 11203 10652 11212
rect 10600 11169 10609 11203
rect 10609 11169 10643 11203
rect 10643 11169 10652 11203
rect 10600 11160 10652 11169
rect 11520 11160 11572 11212
rect 12256 11228 12308 11280
rect 14004 11271 14056 11280
rect 14004 11237 14013 11271
rect 14013 11237 14047 11271
rect 14047 11237 14056 11271
rect 14004 11228 14056 11237
rect 14556 11228 14608 11280
rect 18604 11271 18656 11280
rect 12072 11203 12124 11212
rect 12072 11169 12106 11203
rect 12106 11169 12124 11203
rect 12072 11160 12124 11169
rect 15568 11160 15620 11212
rect 17408 11160 17460 11212
rect 18604 11237 18638 11271
rect 18638 11237 18656 11271
rect 18604 11228 18656 11237
rect 20444 11228 20496 11280
rect 20720 11228 20772 11280
rect 18880 11160 18932 11212
rect 19892 11160 19944 11212
rect 21364 11203 21416 11212
rect 21364 11169 21373 11203
rect 21373 11169 21407 11203
rect 21407 11169 21416 11203
rect 21364 11160 21416 11169
rect 5448 11067 5500 11076
rect 5448 11033 5457 11067
rect 5457 11033 5491 11067
rect 5491 11033 5500 11067
rect 5448 11024 5500 11033
rect 6276 11024 6328 11076
rect 7840 11092 7892 11144
rect 8484 11092 8536 11144
rect 8668 11092 8720 11144
rect 10876 11135 10928 11144
rect 10876 11101 10885 11135
rect 10885 11101 10919 11135
rect 10919 11101 10928 11135
rect 10876 11092 10928 11101
rect 11336 11092 11388 11144
rect 12992 11092 13044 11144
rect 15292 11092 15344 11144
rect 15384 11092 15436 11144
rect 18236 11092 18288 11144
rect 9404 11024 9456 11076
rect 6368 10999 6420 11008
rect 6368 10965 6377 10999
rect 6377 10965 6411 10999
rect 6411 10965 6420 10999
rect 6368 10956 6420 10965
rect 8668 10956 8720 11008
rect 10232 11067 10284 11076
rect 10232 11033 10241 11067
rect 10241 11033 10275 11067
rect 10275 11033 10284 11067
rect 10232 11024 10284 11033
rect 11244 11067 11296 11076
rect 11244 11033 11253 11067
rect 11253 11033 11287 11067
rect 11287 11033 11296 11067
rect 11244 11024 11296 11033
rect 12164 10956 12216 11008
rect 13176 10956 13228 11008
rect 14188 10956 14240 11008
rect 17960 11024 18012 11076
rect 20076 11092 20128 11144
rect 21916 11092 21968 11144
rect 22376 11160 22428 11212
rect 23848 11296 23900 11348
rect 24032 11296 24084 11348
rect 24860 11296 24912 11348
rect 26332 11296 26384 11348
rect 23940 11271 23992 11280
rect 23940 11237 23974 11271
rect 23974 11237 23992 11271
rect 23940 11228 23992 11237
rect 25964 11160 26016 11212
rect 20352 11024 20404 11076
rect 21180 11024 21232 11076
rect 22468 11024 22520 11076
rect 20720 10999 20772 11008
rect 20720 10965 20729 10999
rect 20729 10965 20763 10999
rect 20763 10965 20772 10999
rect 20720 10956 20772 10965
rect 23112 10956 23164 11008
rect 23388 10999 23440 11008
rect 23388 10965 23397 10999
rect 23397 10965 23431 10999
rect 23431 10965 23440 10999
rect 23388 10956 23440 10965
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 1768 10752 1820 10804
rect 2504 10795 2556 10804
rect 2504 10761 2513 10795
rect 2513 10761 2547 10795
rect 2547 10761 2556 10795
rect 2504 10752 2556 10761
rect 5264 10752 5316 10804
rect 6276 10795 6328 10804
rect 1952 10616 2004 10668
rect 2964 10616 3016 10668
rect 1032 10548 1084 10600
rect 2412 10548 2464 10600
rect 3700 10548 3752 10600
rect 3608 10480 3660 10532
rect 2504 10412 2556 10464
rect 4436 10548 4488 10600
rect 6276 10761 6285 10795
rect 6285 10761 6319 10795
rect 6319 10761 6328 10795
rect 6276 10752 6328 10761
rect 8116 10752 8168 10804
rect 9680 10752 9732 10804
rect 10508 10752 10560 10804
rect 11060 10795 11112 10804
rect 11060 10761 11069 10795
rect 11069 10761 11103 10795
rect 11103 10761 11112 10795
rect 11060 10752 11112 10761
rect 11336 10795 11388 10804
rect 11336 10761 11345 10795
rect 11345 10761 11379 10795
rect 11379 10761 11388 10795
rect 11336 10752 11388 10761
rect 12164 10795 12216 10804
rect 12164 10761 12173 10795
rect 12173 10761 12207 10795
rect 12207 10761 12216 10795
rect 12164 10752 12216 10761
rect 13452 10795 13504 10804
rect 13452 10761 13461 10795
rect 13461 10761 13495 10795
rect 13495 10761 13504 10795
rect 13452 10752 13504 10761
rect 5724 10727 5776 10736
rect 5724 10693 5733 10727
rect 5733 10693 5767 10727
rect 5767 10693 5776 10727
rect 5724 10684 5776 10693
rect 6920 10616 6972 10668
rect 12072 10684 12124 10736
rect 12808 10684 12860 10736
rect 14556 10752 14608 10804
rect 15568 10795 15620 10804
rect 15568 10761 15577 10795
rect 15577 10761 15611 10795
rect 15611 10761 15620 10795
rect 15568 10752 15620 10761
rect 16396 10795 16448 10804
rect 16396 10761 16405 10795
rect 16405 10761 16439 10795
rect 16439 10761 16448 10795
rect 16396 10752 16448 10761
rect 18696 10752 18748 10804
rect 19064 10752 19116 10804
rect 19524 10795 19576 10804
rect 19524 10761 19533 10795
rect 19533 10761 19567 10795
rect 19567 10761 19576 10795
rect 19524 10752 19576 10761
rect 21364 10752 21416 10804
rect 22376 10752 22428 10804
rect 22836 10752 22888 10804
rect 6276 10548 6328 10600
rect 13176 10616 13228 10668
rect 3976 10412 4028 10464
rect 4712 10480 4764 10532
rect 8576 10480 8628 10532
rect 9588 10548 9640 10600
rect 15292 10684 15344 10736
rect 19800 10684 19852 10736
rect 19892 10684 19944 10736
rect 21088 10727 21140 10736
rect 21088 10693 21097 10727
rect 21097 10693 21131 10727
rect 21131 10693 21140 10727
rect 21088 10684 21140 10693
rect 14096 10616 14148 10668
rect 14556 10659 14608 10668
rect 14556 10625 14565 10659
rect 14565 10625 14599 10659
rect 14599 10625 14608 10659
rect 14556 10616 14608 10625
rect 16304 10616 16356 10668
rect 16856 10616 16908 10668
rect 20260 10616 20312 10668
rect 20812 10616 20864 10668
rect 21640 10616 21692 10668
rect 22100 10659 22152 10668
rect 22100 10625 22109 10659
rect 22109 10625 22143 10659
rect 22143 10625 22152 10659
rect 23940 10752 23992 10804
rect 22100 10616 22152 10625
rect 9128 10480 9180 10532
rect 11244 10480 11296 10532
rect 6828 10455 6880 10464
rect 6828 10421 6837 10455
rect 6837 10421 6871 10455
rect 6871 10421 6880 10455
rect 6828 10412 6880 10421
rect 12716 10412 12768 10464
rect 12900 10455 12952 10464
rect 12900 10421 12909 10455
rect 12909 10421 12943 10455
rect 12943 10421 12952 10455
rect 12900 10412 12952 10421
rect 13452 10480 13504 10532
rect 18512 10548 18564 10600
rect 19800 10548 19852 10600
rect 20720 10548 20772 10600
rect 22560 10480 22612 10532
rect 15936 10412 15988 10464
rect 16212 10455 16264 10464
rect 16212 10421 16221 10455
rect 16221 10421 16255 10455
rect 16255 10421 16264 10455
rect 16212 10412 16264 10421
rect 16856 10455 16908 10464
rect 16856 10421 16865 10455
rect 16865 10421 16899 10455
rect 16899 10421 16908 10455
rect 16856 10412 16908 10421
rect 18972 10412 19024 10464
rect 24860 10548 24912 10600
rect 24032 10412 24084 10464
rect 25504 10412 25556 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 1952 10251 2004 10260
rect 1952 10217 1961 10251
rect 1961 10217 1995 10251
rect 1995 10217 2004 10251
rect 1952 10208 2004 10217
rect 2780 10208 2832 10260
rect 3148 10208 3200 10260
rect 6368 10208 6420 10260
rect 8024 10208 8076 10260
rect 8576 10251 8628 10260
rect 8576 10217 8585 10251
rect 8585 10217 8619 10251
rect 8619 10217 8628 10251
rect 8576 10208 8628 10217
rect 10692 10251 10744 10260
rect 10692 10217 10701 10251
rect 10701 10217 10735 10251
rect 10735 10217 10744 10251
rect 10692 10208 10744 10217
rect 10876 10208 10928 10260
rect 3516 10140 3568 10192
rect 4436 10183 4488 10192
rect 4436 10149 4445 10183
rect 4445 10149 4479 10183
rect 4479 10149 4488 10183
rect 4436 10140 4488 10149
rect 8116 10140 8168 10192
rect 9220 10183 9272 10192
rect 9220 10149 9229 10183
rect 9229 10149 9263 10183
rect 9263 10149 9272 10183
rect 9220 10140 9272 10149
rect 10784 10140 10836 10192
rect 11060 10140 11112 10192
rect 11336 10140 11388 10192
rect 12900 10208 12952 10260
rect 14004 10208 14056 10260
rect 15384 10208 15436 10260
rect 16948 10208 17000 10260
rect 14648 10140 14700 10192
rect 16304 10140 16356 10192
rect 16488 10140 16540 10192
rect 1952 10072 2004 10124
rect 2780 10115 2832 10124
rect 2780 10081 2789 10115
rect 2789 10081 2823 10115
rect 2823 10081 2832 10115
rect 2780 10072 2832 10081
rect 4068 10072 4120 10124
rect 4804 10072 4856 10124
rect 9312 10072 9364 10124
rect 9772 10072 9824 10124
rect 10324 10072 10376 10124
rect 11520 10115 11572 10124
rect 11520 10081 11529 10115
rect 11529 10081 11563 10115
rect 11563 10081 11572 10115
rect 11520 10072 11572 10081
rect 12624 10072 12676 10124
rect 12900 10072 12952 10124
rect 13820 10072 13872 10124
rect 18052 10208 18104 10260
rect 19248 10251 19300 10260
rect 18144 10115 18196 10124
rect 18144 10081 18153 10115
rect 18153 10081 18187 10115
rect 18187 10081 18196 10115
rect 19248 10217 19257 10251
rect 19257 10217 19291 10251
rect 19291 10217 19300 10251
rect 19248 10208 19300 10217
rect 19432 10208 19484 10260
rect 20352 10208 20404 10260
rect 20536 10208 20588 10260
rect 21456 10208 21508 10260
rect 21640 10208 21692 10260
rect 23112 10208 23164 10260
rect 23756 10208 23808 10260
rect 23940 10208 23992 10260
rect 24676 10208 24728 10260
rect 24768 10251 24820 10260
rect 24768 10217 24777 10251
rect 24777 10217 24811 10251
rect 24811 10217 24820 10251
rect 24768 10208 24820 10217
rect 25320 10208 25372 10260
rect 25504 10251 25556 10260
rect 25504 10217 25513 10251
rect 25513 10217 25547 10251
rect 25547 10217 25556 10251
rect 25504 10208 25556 10217
rect 26424 10208 26476 10260
rect 20260 10183 20312 10192
rect 20260 10149 20269 10183
rect 20269 10149 20303 10183
rect 20303 10149 20312 10183
rect 20260 10140 20312 10149
rect 18144 10072 18196 10081
rect 19248 10072 19300 10124
rect 20628 10072 20680 10124
rect 21916 10140 21968 10192
rect 20996 10072 21048 10124
rect 1124 9936 1176 9988
rect 2964 10004 3016 10056
rect 3976 10004 4028 10056
rect 4712 10047 4764 10056
rect 4712 10013 4721 10047
rect 4721 10013 4755 10047
rect 4755 10013 4764 10047
rect 4712 10004 4764 10013
rect 6276 10047 6328 10056
rect 6276 10013 6285 10047
rect 6285 10013 6319 10047
rect 6319 10013 6328 10047
rect 6276 10004 6328 10013
rect 7656 10047 7708 10056
rect 7656 10013 7665 10047
rect 7665 10013 7699 10047
rect 7699 10013 7708 10047
rect 7656 10004 7708 10013
rect 2228 9911 2280 9920
rect 2228 9877 2237 9911
rect 2237 9877 2271 9911
rect 2271 9877 2280 9911
rect 2228 9868 2280 9877
rect 3884 9979 3936 9988
rect 3884 9945 3893 9979
rect 3893 9945 3927 9979
rect 3927 9945 3936 9979
rect 3884 9936 3936 9945
rect 6644 9936 6696 9988
rect 7196 9979 7248 9988
rect 7196 9945 7205 9979
rect 7205 9945 7239 9979
rect 7239 9945 7248 9979
rect 7196 9936 7248 9945
rect 9496 9936 9548 9988
rect 14188 10004 14240 10056
rect 15292 10047 15344 10056
rect 15292 10013 15301 10047
rect 15301 10013 15335 10047
rect 15335 10013 15344 10047
rect 15292 10004 15344 10013
rect 19156 10004 19208 10056
rect 19984 10004 20036 10056
rect 20168 10004 20220 10056
rect 20720 10004 20772 10056
rect 12808 9936 12860 9988
rect 23388 10072 23440 10124
rect 23756 10115 23808 10124
rect 23756 10081 23765 10115
rect 23765 10081 23799 10115
rect 23799 10081 23808 10115
rect 23756 10072 23808 10081
rect 24952 10115 25004 10124
rect 24952 10081 24961 10115
rect 24961 10081 24995 10115
rect 24995 10081 25004 10115
rect 24952 10072 25004 10081
rect 25596 10072 25648 10124
rect 22468 10004 22520 10056
rect 23848 10004 23900 10056
rect 23480 9936 23532 9988
rect 24676 10004 24728 10056
rect 2872 9868 2924 9920
rect 3516 9911 3568 9920
rect 3516 9877 3525 9911
rect 3525 9877 3559 9911
rect 3559 9877 3568 9911
rect 3516 9868 3568 9877
rect 4620 9868 4672 9920
rect 7288 9868 7340 9920
rect 8668 9868 8720 9920
rect 13452 9911 13504 9920
rect 13452 9877 13461 9911
rect 13461 9877 13495 9911
rect 13495 9877 13504 9911
rect 13452 9868 13504 9877
rect 14648 9911 14700 9920
rect 14648 9877 14657 9911
rect 14657 9877 14691 9911
rect 14691 9877 14700 9911
rect 14648 9868 14700 9877
rect 16764 9868 16816 9920
rect 17224 9911 17276 9920
rect 17224 9877 17233 9911
rect 17233 9877 17267 9911
rect 17267 9877 17276 9911
rect 17224 9868 17276 9877
rect 17316 9868 17368 9920
rect 18052 9868 18104 9920
rect 22008 9868 22060 9920
rect 24768 9868 24820 9920
rect 24952 9868 25004 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 2136 9664 2188 9716
rect 2504 9664 2556 9716
rect 4436 9707 4488 9716
rect 4436 9673 4445 9707
rect 4445 9673 4479 9707
rect 4479 9673 4488 9707
rect 4436 9664 4488 9673
rect 1952 9639 2004 9648
rect 1952 9605 1961 9639
rect 1961 9605 1995 9639
rect 1995 9605 2004 9639
rect 1952 9596 2004 9605
rect 6368 9664 6420 9716
rect 6276 9639 6328 9648
rect 6276 9605 6285 9639
rect 6285 9605 6319 9639
rect 6319 9605 6328 9639
rect 6276 9596 6328 9605
rect 1308 9460 1360 9512
rect 4620 9528 4672 9580
rect 7104 9664 7156 9716
rect 11336 9664 11388 9716
rect 8484 9528 8536 9580
rect 12808 9664 12860 9716
rect 13820 9707 13872 9716
rect 13820 9673 13829 9707
rect 13829 9673 13863 9707
rect 13863 9673 13872 9707
rect 13820 9664 13872 9673
rect 14004 9707 14056 9716
rect 14004 9673 14013 9707
rect 14013 9673 14047 9707
rect 14047 9673 14056 9707
rect 14004 9664 14056 9673
rect 14464 9664 14516 9716
rect 15660 9664 15712 9716
rect 15844 9664 15896 9716
rect 16488 9664 16540 9716
rect 16856 9664 16908 9716
rect 13728 9596 13780 9648
rect 13084 9571 13136 9580
rect 13084 9537 13093 9571
rect 13093 9537 13127 9571
rect 13127 9537 13136 9571
rect 13084 9528 13136 9537
rect 14924 9596 14976 9648
rect 15568 9639 15620 9648
rect 15568 9605 15577 9639
rect 15577 9605 15611 9639
rect 15611 9605 15620 9639
rect 15568 9596 15620 9605
rect 14556 9571 14608 9580
rect 14556 9537 14565 9571
rect 14565 9537 14599 9571
rect 14599 9537 14608 9571
rect 14556 9528 14608 9537
rect 16304 9596 16356 9648
rect 16672 9596 16724 9648
rect 18144 9664 18196 9716
rect 19156 9707 19208 9716
rect 19156 9673 19165 9707
rect 19165 9673 19199 9707
rect 19199 9673 19208 9707
rect 19156 9664 19208 9673
rect 19248 9664 19300 9716
rect 22100 9707 22152 9716
rect 22100 9673 22109 9707
rect 22109 9673 22143 9707
rect 22143 9673 22152 9707
rect 22100 9664 22152 9673
rect 18328 9596 18380 9648
rect 15936 9528 15988 9580
rect 2964 9460 3016 9512
rect 5632 9503 5684 9512
rect 5632 9469 5641 9503
rect 5641 9469 5675 9503
rect 5675 9469 5684 9503
rect 5632 9460 5684 9469
rect 7932 9460 7984 9512
rect 8944 9503 8996 9512
rect 8944 9469 8953 9503
rect 8953 9469 8987 9503
rect 8987 9469 8996 9503
rect 8944 9460 8996 9469
rect 9588 9460 9640 9512
rect 12440 9460 12492 9512
rect 13452 9460 13504 9512
rect 15844 9460 15896 9512
rect 17316 9503 17368 9512
rect 17316 9469 17333 9503
rect 17333 9469 17367 9503
rect 17367 9469 17368 9503
rect 17316 9460 17368 9469
rect 18236 9460 18288 9512
rect 20628 9639 20680 9648
rect 20628 9605 20637 9639
rect 20637 9605 20671 9639
rect 20671 9605 20680 9639
rect 20628 9596 20680 9605
rect 23388 9596 23440 9648
rect 24032 9664 24084 9716
rect 25596 9707 25648 9716
rect 25596 9673 25605 9707
rect 25605 9673 25639 9707
rect 25639 9673 25648 9707
rect 25596 9664 25648 9673
rect 24860 9596 24912 9648
rect 26424 9639 26476 9648
rect 26424 9605 26433 9639
rect 26433 9605 26467 9639
rect 26467 9605 26476 9639
rect 26424 9596 26476 9605
rect 20720 9503 20772 9512
rect 20720 9469 20729 9503
rect 20729 9469 20763 9503
rect 20763 9469 20772 9503
rect 20720 9460 20772 9469
rect 22652 9460 22704 9512
rect 23112 9460 23164 9512
rect 2320 9392 2372 9444
rect 6092 9392 6144 9444
rect 9220 9392 9272 9444
rect 15016 9392 15068 9444
rect 15292 9392 15344 9444
rect 3608 9324 3660 9376
rect 4804 9324 4856 9376
rect 5540 9367 5592 9376
rect 5540 9333 5549 9367
rect 5549 9333 5583 9367
rect 5583 9333 5592 9367
rect 5540 9324 5592 9333
rect 7472 9367 7524 9376
rect 7472 9333 7481 9367
rect 7481 9333 7515 9367
rect 7515 9333 7524 9367
rect 7472 9324 7524 9333
rect 7564 9324 7616 9376
rect 8484 9367 8536 9376
rect 8484 9333 8493 9367
rect 8493 9333 8527 9367
rect 8527 9333 8536 9367
rect 8484 9324 8536 9333
rect 8576 9324 8628 9376
rect 8944 9324 8996 9376
rect 9404 9324 9456 9376
rect 10692 9324 10744 9376
rect 11060 9367 11112 9376
rect 11060 9333 11069 9367
rect 11069 9333 11103 9367
rect 11103 9333 11112 9367
rect 11060 9324 11112 9333
rect 12072 9324 12124 9376
rect 12900 9367 12952 9376
rect 12900 9333 12909 9367
rect 12909 9333 12943 9367
rect 12943 9333 12952 9367
rect 12900 9324 12952 9333
rect 13820 9324 13872 9376
rect 14648 9324 14700 9376
rect 15200 9324 15252 9376
rect 17868 9392 17920 9444
rect 19432 9392 19484 9444
rect 19984 9392 20036 9444
rect 22008 9392 22060 9444
rect 22560 9392 22612 9444
rect 22928 9392 22980 9444
rect 17500 9324 17552 9376
rect 18144 9324 18196 9376
rect 20812 9324 20864 9376
rect 25596 9528 25648 9580
rect 25964 9528 26016 9580
rect 24768 9460 24820 9512
rect 25780 9392 25832 9444
rect 23940 9324 23992 9376
rect 25320 9324 25372 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 1860 9120 1912 9172
rect 2320 9120 2372 9172
rect 3884 9120 3936 9172
rect 4068 9163 4120 9172
rect 4068 9129 4077 9163
rect 4077 9129 4111 9163
rect 4111 9129 4120 9163
rect 4068 9120 4120 9129
rect 4160 9120 4212 9172
rect 4712 9120 4764 9172
rect 5632 9120 5684 9172
rect 9404 9120 9456 9172
rect 9588 9120 9640 9172
rect 9956 9120 10008 9172
rect 3332 9052 3384 9104
rect 6368 9095 6420 9104
rect 6368 9061 6402 9095
rect 6402 9061 6420 9095
rect 6368 9052 6420 9061
rect 9312 9052 9364 9104
rect 9496 9095 9548 9104
rect 9496 9061 9505 9095
rect 9505 9061 9539 9095
rect 9539 9061 9548 9095
rect 9496 9052 9548 9061
rect 11244 9120 11296 9172
rect 11796 9120 11848 9172
rect 13728 9120 13780 9172
rect 14924 9120 14976 9172
rect 15844 9120 15896 9172
rect 19984 9163 20036 9172
rect 14740 9052 14792 9104
rect 16304 9052 16356 9104
rect 17316 9095 17368 9104
rect 17316 9061 17325 9095
rect 17325 9061 17359 9095
rect 17359 9061 17368 9095
rect 17316 9052 17368 9061
rect 18972 9052 19024 9104
rect 19984 9129 19993 9163
rect 19993 9129 20027 9163
rect 20027 9129 20036 9163
rect 19984 9120 20036 9129
rect 21364 9163 21416 9172
rect 21364 9129 21373 9163
rect 21373 9129 21407 9163
rect 21407 9129 21416 9163
rect 21364 9120 21416 9129
rect 23020 9120 23072 9172
rect 23480 9163 23532 9172
rect 23480 9129 23489 9163
rect 23489 9129 23523 9163
rect 23523 9129 23532 9163
rect 23480 9120 23532 9129
rect 24124 9120 24176 9172
rect 25320 9120 25372 9172
rect 26148 9120 26200 9172
rect 26424 9120 26476 9172
rect 2780 9027 2832 9036
rect 2780 8993 2789 9027
rect 2789 8993 2823 9027
rect 2823 8993 2832 9027
rect 2780 8984 2832 8993
rect 3976 8984 4028 9036
rect 2964 8959 3016 8968
rect 2964 8925 2973 8959
rect 2973 8925 3007 8959
rect 3007 8925 3016 8959
rect 2964 8916 3016 8925
rect 4160 8916 4212 8968
rect 5080 8984 5132 9036
rect 6184 8984 6236 9036
rect 8484 8984 8536 9036
rect 11336 8984 11388 9036
rect 13912 8984 13964 9036
rect 15568 9027 15620 9036
rect 15568 8993 15602 9027
rect 15602 8993 15620 9027
rect 15568 8984 15620 8993
rect 17500 8984 17552 9036
rect 23296 9052 23348 9104
rect 22836 9027 22888 9036
rect 4620 8959 4672 8968
rect 4620 8925 4629 8959
rect 4629 8925 4663 8959
rect 4663 8925 4672 8959
rect 4620 8916 4672 8925
rect 1584 8848 1636 8900
rect 3608 8848 3660 8900
rect 5632 8891 5684 8900
rect 5632 8857 5641 8891
rect 5641 8857 5675 8891
rect 5675 8857 5684 8891
rect 5632 8848 5684 8857
rect 3148 8780 3200 8832
rect 4252 8780 4304 8832
rect 4620 8780 4672 8832
rect 8576 8959 8628 8968
rect 8576 8925 8585 8959
rect 8585 8925 8619 8959
rect 8619 8925 8628 8959
rect 8576 8916 8628 8925
rect 9772 8916 9824 8968
rect 10232 8959 10284 8968
rect 10232 8925 10241 8959
rect 10241 8925 10275 8959
rect 10275 8925 10284 8959
rect 11520 8959 11572 8968
rect 10232 8916 10284 8925
rect 11520 8925 11529 8959
rect 11529 8925 11563 8959
rect 11563 8925 11572 8959
rect 11520 8916 11572 8925
rect 12900 8916 12952 8968
rect 14188 8916 14240 8968
rect 14280 8916 14332 8968
rect 15200 8916 15252 8968
rect 9680 8891 9732 8900
rect 9680 8857 9689 8891
rect 9689 8857 9723 8891
rect 9723 8857 9732 8891
rect 9680 8848 9732 8857
rect 14464 8848 14516 8900
rect 14924 8848 14976 8900
rect 17316 8916 17368 8968
rect 17868 8959 17920 8968
rect 17868 8925 17877 8959
rect 17877 8925 17911 8959
rect 17911 8925 17920 8959
rect 17868 8916 17920 8925
rect 19524 8916 19576 8968
rect 22836 8993 22845 9027
rect 22845 8993 22879 9027
rect 22879 8993 22888 9027
rect 22836 8984 22888 8993
rect 24400 9027 24452 9036
rect 24400 8993 24409 9027
rect 24409 8993 24443 9027
rect 24443 8993 24452 9027
rect 24400 8984 24452 8993
rect 24860 8984 24912 9036
rect 21456 8959 21508 8968
rect 21456 8925 21465 8959
rect 21465 8925 21499 8959
rect 21499 8925 21508 8959
rect 21456 8916 21508 8925
rect 22928 8916 22980 8968
rect 20812 8848 20864 8900
rect 24952 8848 25004 8900
rect 7288 8780 7340 8832
rect 8208 8780 8260 8832
rect 13084 8780 13136 8832
rect 13728 8780 13780 8832
rect 14188 8780 14240 8832
rect 16304 8780 16356 8832
rect 17868 8780 17920 8832
rect 18236 8780 18288 8832
rect 20904 8823 20956 8832
rect 20904 8789 20913 8823
rect 20913 8789 20947 8823
rect 20947 8789 20956 8823
rect 20904 8780 20956 8789
rect 22468 8823 22520 8832
rect 22468 8789 22477 8823
rect 22477 8789 22511 8823
rect 22511 8789 22520 8823
rect 22468 8780 22520 8789
rect 23940 8780 23992 8832
rect 24124 8780 24176 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 2688 8619 2740 8628
rect 2688 8585 2697 8619
rect 2697 8585 2731 8619
rect 2731 8585 2740 8619
rect 2688 8576 2740 8585
rect 4896 8576 4948 8628
rect 6368 8576 6420 8628
rect 7288 8576 7340 8628
rect 10232 8576 10284 8628
rect 11796 8619 11848 8628
rect 11796 8585 11805 8619
rect 11805 8585 11839 8619
rect 11839 8585 11848 8619
rect 11796 8576 11848 8585
rect 12900 8576 12952 8628
rect 13912 8619 13964 8628
rect 13912 8585 13921 8619
rect 13921 8585 13955 8619
rect 13955 8585 13964 8619
rect 13912 8576 13964 8585
rect 15384 8619 15436 8628
rect 15384 8585 15393 8619
rect 15393 8585 15427 8619
rect 15427 8585 15436 8619
rect 15384 8576 15436 8585
rect 17316 8576 17368 8628
rect 17500 8576 17552 8628
rect 18972 8576 19024 8628
rect 19524 8576 19576 8628
rect 20444 8619 20496 8628
rect 20444 8585 20453 8619
rect 20453 8585 20487 8619
rect 20487 8585 20496 8619
rect 20444 8576 20496 8585
rect 21364 8576 21416 8628
rect 23020 8576 23072 8628
rect 23664 8619 23716 8628
rect 23664 8585 23673 8619
rect 23673 8585 23707 8619
rect 23707 8585 23716 8619
rect 23664 8576 23716 8585
rect 24860 8576 24912 8628
rect 24952 8576 25004 8628
rect 26148 8619 26200 8628
rect 26148 8585 26157 8619
rect 26157 8585 26191 8619
rect 26191 8585 26200 8619
rect 26148 8576 26200 8585
rect 2964 8508 3016 8560
rect 7196 8508 7248 8560
rect 12808 8508 12860 8560
rect 2412 8440 2464 8492
rect 2872 8440 2924 8492
rect 3976 8440 4028 8492
rect 8484 8483 8536 8492
rect 1584 8372 1636 8424
rect 2228 8372 2280 8424
rect 3516 8372 3568 8424
rect 4068 8372 4120 8424
rect 1952 8304 2004 8356
rect 2964 8304 3016 8356
rect 3240 8304 3292 8356
rect 4160 8347 4212 8356
rect 4160 8313 4169 8347
rect 4169 8313 4203 8347
rect 4203 8313 4212 8347
rect 4160 8304 4212 8313
rect 2228 8236 2280 8288
rect 2872 8236 2924 8288
rect 3148 8279 3200 8288
rect 3148 8245 3157 8279
rect 3157 8245 3191 8279
rect 3191 8245 3200 8279
rect 3148 8236 3200 8245
rect 3332 8236 3384 8288
rect 3700 8279 3752 8288
rect 3700 8245 3709 8279
rect 3709 8245 3743 8279
rect 3743 8245 3752 8279
rect 3700 8236 3752 8245
rect 4436 8304 4488 8356
rect 6644 8347 6696 8356
rect 6644 8313 6653 8347
rect 6653 8313 6687 8347
rect 6687 8313 6696 8347
rect 7104 8372 7156 8424
rect 8484 8449 8493 8483
rect 8493 8449 8527 8483
rect 8527 8449 8536 8483
rect 8484 8440 8536 8449
rect 11336 8483 11388 8492
rect 11336 8449 11345 8483
rect 11345 8449 11379 8483
rect 11379 8449 11388 8483
rect 11336 8440 11388 8449
rect 15200 8508 15252 8560
rect 16580 8508 16632 8560
rect 13084 8483 13136 8492
rect 8852 8372 8904 8424
rect 9588 8372 9640 8424
rect 11244 8415 11296 8424
rect 11244 8381 11253 8415
rect 11253 8381 11287 8415
rect 11287 8381 11296 8415
rect 11244 8372 11296 8381
rect 11796 8372 11848 8424
rect 13084 8449 13093 8483
rect 13093 8449 13127 8483
rect 13127 8449 13136 8483
rect 13084 8440 13136 8449
rect 15016 8440 15068 8492
rect 15568 8440 15620 8492
rect 16764 8440 16816 8492
rect 17316 8440 17368 8492
rect 19340 8508 19392 8560
rect 23296 8508 23348 8560
rect 13452 8372 13504 8424
rect 13636 8372 13688 8424
rect 13912 8372 13964 8424
rect 6644 8304 6696 8313
rect 9128 8304 9180 8356
rect 9772 8347 9824 8356
rect 9772 8313 9781 8347
rect 9781 8313 9815 8347
rect 9815 8313 9824 8347
rect 9772 8304 9824 8313
rect 10600 8347 10652 8356
rect 10600 8313 10609 8347
rect 10609 8313 10643 8347
rect 10643 8313 10652 8347
rect 10600 8304 10652 8313
rect 11888 8304 11940 8356
rect 12808 8347 12860 8356
rect 12808 8313 12817 8347
rect 12817 8313 12851 8347
rect 12851 8313 12860 8347
rect 12808 8304 12860 8313
rect 17684 8372 17736 8424
rect 21456 8440 21508 8492
rect 22376 8440 22428 8492
rect 22652 8440 22704 8492
rect 24124 8483 24176 8492
rect 24124 8449 24133 8483
rect 24133 8449 24167 8483
rect 24167 8449 24176 8483
rect 24124 8440 24176 8449
rect 24860 8440 24912 8492
rect 19616 8372 19668 8424
rect 20720 8372 20772 8424
rect 23664 8372 23716 8424
rect 25228 8415 25280 8424
rect 25228 8381 25237 8415
rect 25237 8381 25271 8415
rect 25271 8381 25280 8415
rect 25228 8372 25280 8381
rect 14464 8304 14516 8356
rect 15016 8304 15068 8356
rect 16764 8347 16816 8356
rect 16764 8313 16773 8347
rect 16773 8313 16807 8347
rect 16807 8313 16816 8347
rect 16764 8304 16816 8313
rect 18236 8304 18288 8356
rect 4620 8236 4672 8288
rect 8024 8236 8076 8288
rect 11060 8236 11112 8288
rect 12900 8236 12952 8288
rect 20444 8304 20496 8356
rect 19340 8236 19392 8288
rect 20536 8236 20588 8288
rect 22836 8304 22888 8356
rect 20720 8236 20772 8288
rect 22652 8279 22704 8288
rect 22652 8245 22661 8279
rect 22661 8245 22695 8279
rect 22695 8245 22704 8279
rect 22652 8236 22704 8245
rect 23388 8279 23440 8288
rect 23388 8245 23397 8279
rect 23397 8245 23431 8279
rect 23431 8245 23440 8279
rect 23388 8236 23440 8245
rect 25412 8279 25464 8288
rect 25412 8245 25421 8279
rect 25421 8245 25455 8279
rect 25455 8245 25464 8279
rect 25412 8236 25464 8245
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1400 8032 1452 8084
rect 1676 8032 1728 8084
rect 2320 8032 2372 8084
rect 3608 8032 3660 8084
rect 4436 8032 4488 8084
rect 5448 8032 5500 8084
rect 5540 8032 5592 8084
rect 5816 8075 5868 8084
rect 5816 8041 5825 8075
rect 5825 8041 5859 8075
rect 5859 8041 5868 8075
rect 5816 8032 5868 8041
rect 8392 8075 8444 8084
rect 8392 8041 8401 8075
rect 8401 8041 8435 8075
rect 8435 8041 8444 8075
rect 8392 8032 8444 8041
rect 9312 8032 9364 8084
rect 10692 8032 10744 8084
rect 11336 8075 11388 8084
rect 11336 8041 11345 8075
rect 11345 8041 11379 8075
rect 11379 8041 11388 8075
rect 11336 8032 11388 8041
rect 4712 7964 4764 8016
rect 12348 8032 12400 8084
rect 13084 8032 13136 8084
rect 13820 8032 13872 8084
rect 2872 7896 2924 7948
rect 4528 7896 4580 7948
rect 5264 7896 5316 7948
rect 7288 7896 7340 7948
rect 12256 7939 12308 7948
rect 12256 7905 12265 7939
rect 12265 7905 12299 7939
rect 12299 7905 12308 7939
rect 12256 7896 12308 7905
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 5356 7871 5408 7880
rect 5356 7837 5365 7871
rect 5365 7837 5399 7871
rect 5399 7837 5408 7871
rect 5356 7828 5408 7837
rect 6460 7828 6512 7880
rect 6828 7871 6880 7880
rect 6828 7837 6837 7871
rect 6837 7837 6871 7871
rect 6871 7837 6880 7871
rect 6828 7828 6880 7837
rect 7104 7828 7156 7880
rect 8484 7871 8536 7880
rect 8484 7837 8493 7871
rect 8493 7837 8527 7871
rect 8527 7837 8536 7871
rect 8484 7828 8536 7837
rect 5080 7760 5132 7812
rect 8116 7760 8168 7812
rect 9772 7760 9824 7812
rect 11060 7828 11112 7880
rect 12348 7871 12400 7880
rect 12348 7837 12357 7871
rect 12357 7837 12391 7871
rect 12391 7837 12400 7871
rect 12348 7828 12400 7837
rect 13176 7964 13228 8016
rect 14464 8032 14516 8084
rect 15292 8075 15344 8084
rect 15292 8041 15301 8075
rect 15301 8041 15335 8075
rect 15335 8041 15344 8075
rect 15292 8032 15344 8041
rect 16304 8032 16356 8084
rect 17776 8032 17828 8084
rect 18788 8075 18840 8084
rect 18788 8041 18797 8075
rect 18797 8041 18831 8075
rect 18831 8041 18840 8075
rect 18788 8032 18840 8041
rect 18972 8032 19024 8084
rect 21456 8032 21508 8084
rect 22928 8075 22980 8084
rect 22928 8041 22937 8075
rect 22937 8041 22971 8075
rect 22971 8041 22980 8075
rect 22928 8032 22980 8041
rect 23296 8075 23348 8084
rect 23296 8041 23305 8075
rect 23305 8041 23339 8075
rect 23339 8041 23348 8075
rect 23296 8032 23348 8041
rect 24032 8075 24084 8084
rect 24032 8041 24041 8075
rect 24041 8041 24075 8075
rect 24075 8041 24084 8075
rect 24032 8032 24084 8041
rect 24216 8032 24268 8084
rect 26148 8032 26200 8084
rect 26424 8032 26476 8084
rect 13636 7896 13688 7948
rect 14096 7964 14148 8016
rect 15016 7964 15068 8016
rect 16396 7964 16448 8016
rect 18328 8007 18380 8016
rect 18328 7973 18337 8007
rect 18337 7973 18371 8007
rect 18371 7973 18380 8007
rect 18328 7964 18380 7973
rect 20076 7964 20128 8016
rect 22008 7964 22060 8016
rect 13912 7939 13964 7948
rect 13912 7905 13921 7939
rect 13921 7905 13955 7939
rect 13955 7905 13964 7939
rect 13912 7896 13964 7905
rect 13728 7828 13780 7880
rect 14096 7871 14148 7880
rect 14096 7837 14105 7871
rect 14105 7837 14139 7871
rect 14139 7837 14148 7871
rect 14096 7828 14148 7837
rect 13084 7760 13136 7812
rect 13820 7760 13872 7812
rect 15568 7896 15620 7948
rect 14924 7828 14976 7880
rect 17684 7828 17736 7880
rect 18420 7828 18472 7880
rect 3332 7735 3384 7744
rect 3332 7701 3341 7735
rect 3341 7701 3375 7735
rect 3375 7701 3384 7735
rect 3332 7692 3384 7701
rect 4436 7692 4488 7744
rect 6092 7735 6144 7744
rect 6092 7701 6101 7735
rect 6101 7701 6135 7735
rect 6135 7701 6144 7735
rect 6092 7692 6144 7701
rect 6920 7692 6972 7744
rect 7932 7735 7984 7744
rect 7932 7701 7941 7735
rect 7941 7701 7975 7735
rect 7975 7701 7984 7735
rect 7932 7692 7984 7701
rect 9956 7735 10008 7744
rect 9956 7701 9965 7735
rect 9965 7701 9999 7735
rect 9999 7701 10008 7735
rect 9956 7692 10008 7701
rect 10048 7692 10100 7744
rect 11888 7692 11940 7744
rect 15660 7760 15712 7812
rect 18880 7896 18932 7948
rect 23388 7939 23440 7948
rect 23388 7905 23397 7939
rect 23397 7905 23431 7939
rect 23431 7905 23440 7939
rect 23388 7896 23440 7905
rect 23572 7896 23624 7948
rect 23756 7896 23808 7948
rect 25228 7896 25280 7948
rect 19248 7871 19300 7880
rect 19248 7837 19257 7871
rect 19257 7837 19291 7871
rect 19291 7837 19300 7871
rect 19248 7828 19300 7837
rect 19340 7871 19392 7880
rect 19340 7837 19349 7871
rect 19349 7837 19383 7871
rect 19383 7837 19392 7871
rect 19340 7828 19392 7837
rect 20812 7828 20864 7880
rect 24952 7871 25004 7880
rect 24952 7837 24961 7871
rect 24961 7837 24995 7871
rect 24995 7837 25004 7871
rect 24952 7828 25004 7837
rect 24860 7760 24912 7812
rect 14464 7735 14516 7744
rect 14464 7701 14473 7735
rect 14473 7701 14507 7735
rect 14507 7701 14516 7735
rect 14464 7692 14516 7701
rect 18604 7735 18656 7744
rect 18604 7701 18613 7735
rect 18613 7701 18647 7735
rect 18647 7701 18656 7735
rect 18604 7692 18656 7701
rect 20536 7735 20588 7744
rect 20536 7701 20545 7735
rect 20545 7701 20579 7735
rect 20579 7701 20588 7735
rect 20536 7692 20588 7701
rect 23296 7692 23348 7744
rect 25320 7692 25372 7744
rect 25504 7735 25556 7744
rect 25504 7701 25513 7735
rect 25513 7701 25547 7735
rect 25547 7701 25556 7735
rect 25504 7692 25556 7701
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 1584 7488 1636 7540
rect 2320 7488 2372 7540
rect 3148 7488 3200 7540
rect 5448 7531 5500 7540
rect 5448 7497 5457 7531
rect 5457 7497 5491 7531
rect 5491 7497 5500 7531
rect 5448 7488 5500 7497
rect 8392 7488 8444 7540
rect 9772 7531 9824 7540
rect 9772 7497 9781 7531
rect 9781 7497 9815 7531
rect 9815 7497 9824 7531
rect 9772 7488 9824 7497
rect 11336 7488 11388 7540
rect 12348 7488 12400 7540
rect 12624 7488 12676 7540
rect 13636 7488 13688 7540
rect 13912 7488 13964 7540
rect 15568 7531 15620 7540
rect 15568 7497 15577 7531
rect 15577 7497 15611 7531
rect 15611 7497 15620 7531
rect 15568 7488 15620 7497
rect 15844 7531 15896 7540
rect 15844 7497 15853 7531
rect 15853 7497 15887 7531
rect 15887 7497 15896 7531
rect 15844 7488 15896 7497
rect 17500 7531 17552 7540
rect 17500 7497 17509 7531
rect 17509 7497 17543 7531
rect 17543 7497 17552 7531
rect 17500 7488 17552 7497
rect 17776 7488 17828 7540
rect 18972 7488 19024 7540
rect 19340 7531 19392 7540
rect 19340 7497 19349 7531
rect 19349 7497 19383 7531
rect 19383 7497 19392 7531
rect 20076 7531 20128 7540
rect 19340 7488 19392 7497
rect 20076 7497 20085 7531
rect 20085 7497 20119 7531
rect 20119 7497 20128 7531
rect 20076 7488 20128 7497
rect 23388 7531 23440 7540
rect 23388 7497 23397 7531
rect 23397 7497 23431 7531
rect 23431 7497 23440 7531
rect 23388 7488 23440 7497
rect 23940 7531 23992 7540
rect 23940 7497 23949 7531
rect 23949 7497 23983 7531
rect 23983 7497 23992 7531
rect 23940 7488 23992 7497
rect 26424 7531 26476 7540
rect 26424 7497 26433 7531
rect 26433 7497 26467 7531
rect 26467 7497 26476 7531
rect 26424 7488 26476 7497
rect 7012 7420 7064 7472
rect 12164 7463 12216 7472
rect 12164 7429 12173 7463
rect 12173 7429 12207 7463
rect 12207 7429 12216 7463
rect 12164 7420 12216 7429
rect 12900 7420 12952 7472
rect 13820 7420 13872 7472
rect 4436 7395 4488 7404
rect 4436 7361 4445 7395
rect 4445 7361 4479 7395
rect 4479 7361 4488 7395
rect 4436 7352 4488 7361
rect 8024 7395 8076 7404
rect 3332 7284 3384 7336
rect 3608 7284 3660 7336
rect 8024 7361 8033 7395
rect 8033 7361 8067 7395
rect 8067 7361 8076 7395
rect 8024 7352 8076 7361
rect 8116 7395 8168 7404
rect 8116 7361 8125 7395
rect 8125 7361 8159 7395
rect 8159 7361 8168 7395
rect 8116 7352 8168 7361
rect 12716 7352 12768 7404
rect 13176 7352 13228 7404
rect 13912 7352 13964 7404
rect 14280 7352 14332 7404
rect 14464 7395 14516 7404
rect 14464 7361 14473 7395
rect 14473 7361 14507 7395
rect 14507 7361 14516 7395
rect 14464 7352 14516 7361
rect 19248 7420 19300 7472
rect 20260 7352 20312 7404
rect 21456 7352 21508 7404
rect 21916 7352 21968 7404
rect 22928 7420 22980 7472
rect 5540 7284 5592 7336
rect 7932 7327 7984 7336
rect 7932 7293 7941 7327
rect 7941 7293 7975 7327
rect 7975 7293 7984 7327
rect 7932 7284 7984 7293
rect 8668 7284 8720 7336
rect 9588 7284 9640 7336
rect 9956 7284 10008 7336
rect 12440 7284 12492 7336
rect 2688 7216 2740 7268
rect 5080 7216 5132 7268
rect 7104 7259 7156 7268
rect 7104 7225 7113 7259
rect 7113 7225 7147 7259
rect 7147 7225 7156 7259
rect 7104 7216 7156 7225
rect 8392 7216 8444 7268
rect 8852 7216 8904 7268
rect 11060 7216 11112 7268
rect 11152 7216 11204 7268
rect 15844 7284 15896 7336
rect 17408 7284 17460 7336
rect 18236 7284 18288 7336
rect 18788 7284 18840 7336
rect 22008 7284 22060 7336
rect 23756 7284 23808 7336
rect 23940 7284 23992 7336
rect 24860 7352 24912 7404
rect 24952 7284 25004 7336
rect 25504 7327 25556 7336
rect 25504 7293 25513 7327
rect 25513 7293 25547 7327
rect 25547 7293 25556 7327
rect 25504 7284 25556 7293
rect 1860 7191 1912 7200
rect 1860 7157 1869 7191
rect 1869 7157 1903 7191
rect 1903 7157 1912 7191
rect 1860 7148 1912 7157
rect 2872 7148 2924 7200
rect 3148 7148 3200 7200
rect 4252 7148 4304 7200
rect 5264 7148 5316 7200
rect 6276 7148 6328 7200
rect 6460 7191 6512 7200
rect 6460 7157 6469 7191
rect 6469 7157 6503 7191
rect 6503 7157 6512 7191
rect 6460 7148 6512 7157
rect 7288 7148 7340 7200
rect 9220 7148 9272 7200
rect 9588 7148 9640 7200
rect 12532 7148 12584 7200
rect 12900 7191 12952 7200
rect 12900 7157 12909 7191
rect 12909 7157 12943 7191
rect 12943 7157 12952 7191
rect 12900 7148 12952 7157
rect 14280 7148 14332 7200
rect 17592 7216 17644 7268
rect 18604 7259 18656 7268
rect 18604 7225 18613 7259
rect 18613 7225 18647 7259
rect 18647 7225 18656 7259
rect 18604 7216 18656 7225
rect 14464 7148 14516 7200
rect 16396 7191 16448 7200
rect 16396 7157 16405 7191
rect 16405 7157 16439 7191
rect 16439 7157 16448 7191
rect 16396 7148 16448 7157
rect 18328 7148 18380 7200
rect 19340 7148 19392 7200
rect 20444 7148 20496 7200
rect 20628 7148 20680 7200
rect 24124 7216 24176 7268
rect 22008 7148 22060 7200
rect 22192 7148 22244 7200
rect 22284 7148 22336 7200
rect 23756 7148 23808 7200
rect 25964 7148 26016 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 4436 6944 4488 6996
rect 7472 6944 7524 6996
rect 10692 6944 10744 6996
rect 12256 6944 12308 6996
rect 12440 6987 12492 6996
rect 12440 6953 12449 6987
rect 12449 6953 12483 6987
rect 12483 6953 12492 6987
rect 13084 6987 13136 6996
rect 12440 6944 12492 6953
rect 13084 6953 13093 6987
rect 13093 6953 13127 6987
rect 13127 6953 13136 6987
rect 13084 6944 13136 6953
rect 13268 6944 13320 6996
rect 14096 6944 14148 6996
rect 17592 6944 17644 6996
rect 18880 6944 18932 6996
rect 19248 6944 19300 6996
rect 20260 6987 20312 6996
rect 20260 6953 20269 6987
rect 20269 6953 20303 6987
rect 20303 6953 20312 6987
rect 20260 6944 20312 6953
rect 21916 6987 21968 6996
rect 21916 6953 21925 6987
rect 21925 6953 21959 6987
rect 21959 6953 21968 6987
rect 21916 6944 21968 6953
rect 26148 6944 26200 6996
rect 8024 6876 8076 6928
rect 1400 6808 1452 6860
rect 1584 6808 1636 6860
rect 3608 6808 3660 6860
rect 4896 6808 4948 6860
rect 5540 6808 5592 6860
rect 6828 6808 6880 6860
rect 6920 6808 6972 6860
rect 13728 6876 13780 6928
rect 13820 6876 13872 6928
rect 9772 6808 9824 6860
rect 11336 6808 11388 6860
rect 14648 6876 14700 6928
rect 14832 6876 14884 6928
rect 16396 6876 16448 6928
rect 15844 6808 15896 6860
rect 16212 6808 16264 6860
rect 19156 6876 19208 6928
rect 23112 6876 23164 6928
rect 24860 6876 24912 6928
rect 25044 6876 25096 6928
rect 19432 6851 19484 6860
rect 4620 6740 4672 6792
rect 3148 6604 3200 6656
rect 3424 6647 3476 6656
rect 3424 6613 3433 6647
rect 3433 6613 3467 6647
rect 3467 6613 3476 6647
rect 3424 6604 3476 6613
rect 3884 6647 3936 6656
rect 3884 6613 3893 6647
rect 3893 6613 3927 6647
rect 3927 6613 3936 6647
rect 3884 6604 3936 6613
rect 4252 6604 4304 6656
rect 7472 6740 7524 6792
rect 8116 6740 8168 6792
rect 9588 6740 9640 6792
rect 7932 6672 7984 6724
rect 5540 6604 5592 6656
rect 6092 6604 6144 6656
rect 8392 6647 8444 6656
rect 8392 6613 8401 6647
rect 8401 6613 8435 6647
rect 8435 6613 8444 6647
rect 8392 6604 8444 6613
rect 9220 6604 9272 6656
rect 9312 6604 9364 6656
rect 13176 6783 13228 6792
rect 13176 6749 13185 6783
rect 13185 6749 13219 6783
rect 13219 6749 13228 6783
rect 13176 6740 13228 6749
rect 14096 6740 14148 6792
rect 15476 6783 15528 6792
rect 15476 6749 15485 6783
rect 15485 6749 15519 6783
rect 15519 6749 15528 6783
rect 15476 6740 15528 6749
rect 16672 6783 16724 6792
rect 16120 6672 16172 6724
rect 16672 6749 16681 6783
rect 16681 6749 16715 6783
rect 16715 6749 16724 6783
rect 16672 6740 16724 6749
rect 19432 6817 19441 6851
rect 19441 6817 19475 6851
rect 19475 6817 19484 6851
rect 19432 6808 19484 6817
rect 21272 6851 21324 6860
rect 21272 6817 21281 6851
rect 21281 6817 21315 6851
rect 21315 6817 21324 6851
rect 21272 6808 21324 6817
rect 18604 6740 18656 6792
rect 18788 6740 18840 6792
rect 19616 6783 19668 6792
rect 19616 6749 19625 6783
rect 19625 6749 19659 6783
rect 19659 6749 19668 6783
rect 19616 6740 19668 6749
rect 20720 6740 20772 6792
rect 21824 6740 21876 6792
rect 23296 6783 23348 6792
rect 23296 6749 23305 6783
rect 23305 6749 23339 6783
rect 23339 6749 23348 6783
rect 23296 6740 23348 6749
rect 16856 6672 16908 6724
rect 20444 6672 20496 6724
rect 20996 6672 21048 6724
rect 21732 6672 21784 6724
rect 24768 6672 24820 6724
rect 25228 6672 25280 6724
rect 25872 6672 25924 6724
rect 10416 6604 10468 6656
rect 11060 6604 11112 6656
rect 12900 6604 12952 6656
rect 14832 6604 14884 6656
rect 16396 6604 16448 6656
rect 20628 6647 20680 6656
rect 20628 6613 20637 6647
rect 20637 6613 20671 6647
rect 20671 6613 20680 6647
rect 20628 6604 20680 6613
rect 21364 6604 21416 6656
rect 24860 6604 24912 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 3608 6400 3660 6452
rect 1584 6264 1636 6316
rect 4068 6400 4120 6452
rect 9772 6443 9824 6452
rect 9772 6409 9781 6443
rect 9781 6409 9815 6443
rect 9815 6409 9824 6443
rect 9772 6400 9824 6409
rect 13820 6400 13872 6452
rect 16948 6400 17000 6452
rect 17776 6443 17828 6452
rect 4436 6332 4488 6384
rect 6460 6332 6512 6384
rect 17776 6409 17785 6443
rect 17785 6409 17819 6443
rect 17819 6409 17828 6443
rect 17776 6400 17828 6409
rect 18328 6332 18380 6384
rect 1768 6196 1820 6248
rect 2136 6196 2188 6248
rect 2688 6171 2740 6180
rect 2688 6137 2700 6171
rect 2700 6137 2740 6171
rect 2688 6128 2740 6137
rect 4896 6196 4948 6248
rect 5264 6239 5316 6248
rect 5264 6205 5273 6239
rect 5273 6205 5307 6239
rect 5307 6205 5316 6239
rect 5264 6196 5316 6205
rect 5540 6196 5592 6248
rect 8116 6196 8168 6248
rect 10416 6196 10468 6248
rect 11520 6196 11572 6248
rect 11980 6196 12032 6248
rect 7104 6128 7156 6180
rect 1768 6060 1820 6112
rect 5356 6103 5408 6112
rect 5356 6069 5365 6103
rect 5365 6069 5399 6103
rect 5399 6069 5408 6103
rect 5356 6060 5408 6069
rect 7472 6060 7524 6112
rect 8024 6060 8076 6112
rect 13176 6196 13228 6248
rect 16304 6264 16356 6316
rect 18604 6400 18656 6452
rect 21824 6443 21876 6452
rect 21824 6409 21833 6443
rect 21833 6409 21867 6443
rect 21867 6409 21876 6443
rect 21824 6400 21876 6409
rect 23112 6443 23164 6452
rect 23112 6409 23121 6443
rect 23121 6409 23155 6443
rect 23155 6409 23164 6443
rect 23112 6400 23164 6409
rect 23388 6443 23440 6452
rect 23388 6409 23397 6443
rect 23397 6409 23431 6443
rect 23431 6409 23440 6443
rect 23388 6400 23440 6409
rect 25044 6443 25096 6452
rect 25044 6409 25053 6443
rect 25053 6409 25087 6443
rect 25087 6409 25096 6443
rect 25044 6400 25096 6409
rect 26148 6400 26200 6452
rect 15200 6128 15252 6180
rect 18420 6196 18472 6248
rect 19432 6264 19484 6316
rect 20536 6196 20588 6248
rect 23296 6196 23348 6248
rect 24860 6196 24912 6248
rect 9956 6060 10008 6112
rect 12164 6103 12216 6112
rect 12164 6069 12173 6103
rect 12173 6069 12207 6103
rect 12207 6069 12216 6103
rect 12164 6060 12216 6069
rect 13452 6060 13504 6112
rect 14372 6103 14424 6112
rect 14372 6069 14381 6103
rect 14381 6069 14415 6103
rect 14415 6069 14424 6103
rect 14372 6060 14424 6069
rect 15660 6060 15712 6112
rect 16212 6060 16264 6112
rect 16948 6060 17000 6112
rect 17500 6060 17552 6112
rect 19340 6128 19392 6180
rect 20168 6128 20220 6180
rect 23388 6128 23440 6180
rect 25044 6128 25096 6180
rect 18328 6060 18380 6112
rect 20076 6060 20128 6112
rect 22192 6060 22244 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 1860 5856 1912 5908
rect 3148 5856 3200 5908
rect 4252 5899 4304 5908
rect 4252 5865 4261 5899
rect 4261 5865 4295 5899
rect 4295 5865 4304 5899
rect 4252 5856 4304 5865
rect 4712 5899 4764 5908
rect 4712 5865 4721 5899
rect 4721 5865 4755 5899
rect 4755 5865 4764 5899
rect 4712 5856 4764 5865
rect 5080 5856 5132 5908
rect 6920 5856 6972 5908
rect 7932 5856 7984 5908
rect 9680 5899 9732 5908
rect 9680 5865 9689 5899
rect 9689 5865 9723 5899
rect 9723 5865 9732 5899
rect 9680 5856 9732 5865
rect 11520 5899 11572 5908
rect 11520 5865 11529 5899
rect 11529 5865 11563 5899
rect 11563 5865 11572 5899
rect 11520 5856 11572 5865
rect 13084 5856 13136 5908
rect 13268 5856 13320 5908
rect 13728 5856 13780 5908
rect 15292 5856 15344 5908
rect 15660 5899 15712 5908
rect 15660 5865 15669 5899
rect 15669 5865 15703 5899
rect 15703 5865 15712 5899
rect 15660 5856 15712 5865
rect 15936 5856 15988 5908
rect 16672 5899 16724 5908
rect 16672 5865 16681 5899
rect 16681 5865 16715 5899
rect 16715 5865 16724 5899
rect 16672 5856 16724 5865
rect 16856 5899 16908 5908
rect 16856 5865 16865 5899
rect 16865 5865 16899 5899
rect 16899 5865 16908 5899
rect 16856 5856 16908 5865
rect 17684 5899 17736 5908
rect 17684 5865 17693 5899
rect 17693 5865 17727 5899
rect 17727 5865 17736 5899
rect 17684 5856 17736 5865
rect 18236 5899 18288 5908
rect 18236 5865 18245 5899
rect 18245 5865 18279 5899
rect 18279 5865 18288 5899
rect 18236 5856 18288 5865
rect 21272 5856 21324 5908
rect 22008 5856 22060 5908
rect 22376 5856 22428 5908
rect 23388 5856 23440 5908
rect 23480 5856 23532 5908
rect 23756 5856 23808 5908
rect 25044 5899 25096 5908
rect 2872 5831 2924 5840
rect 2872 5797 2881 5831
rect 2881 5797 2915 5831
rect 2915 5797 2924 5831
rect 2872 5788 2924 5797
rect 3608 5788 3660 5840
rect 5540 5788 5592 5840
rect 7012 5788 7064 5840
rect 11152 5788 11204 5840
rect 12348 5788 12400 5840
rect 16580 5788 16632 5840
rect 19248 5788 19300 5840
rect 20904 5788 20956 5840
rect 21824 5831 21876 5840
rect 21824 5797 21858 5831
rect 21858 5797 21876 5831
rect 21824 5788 21876 5797
rect 23572 5788 23624 5840
rect 25044 5865 25053 5899
rect 25053 5865 25087 5899
rect 25087 5865 25096 5899
rect 25044 5856 25096 5865
rect 26148 5899 26200 5908
rect 26148 5865 26157 5899
rect 26157 5865 26191 5899
rect 26191 5865 26200 5899
rect 26148 5856 26200 5865
rect 1400 5720 1452 5772
rect 1952 5720 2004 5772
rect 4344 5720 4396 5772
rect 3976 5652 4028 5704
rect 4068 5652 4120 5704
rect 5080 5652 5132 5704
rect 6828 5720 6880 5772
rect 7288 5720 7340 5772
rect 10048 5763 10100 5772
rect 10048 5729 10057 5763
rect 10057 5729 10091 5763
rect 10091 5729 10100 5763
rect 10048 5720 10100 5729
rect 11888 5720 11940 5772
rect 12716 5720 12768 5772
rect 13176 5720 13228 5772
rect 14832 5720 14884 5772
rect 18236 5720 18288 5772
rect 19984 5720 20036 5772
rect 20536 5720 20588 5772
rect 20812 5720 20864 5772
rect 23296 5720 23348 5772
rect 23480 5720 23532 5772
rect 24768 5720 24820 5772
rect 6460 5695 6512 5704
rect 6460 5661 6469 5695
rect 6469 5661 6503 5695
rect 6503 5661 6512 5695
rect 6460 5652 6512 5661
rect 8024 5695 8076 5704
rect 8024 5661 8033 5695
rect 8033 5661 8067 5695
rect 8067 5661 8076 5695
rect 8024 5652 8076 5661
rect 11980 5695 12032 5704
rect 3148 5584 3200 5636
rect 5356 5584 5408 5636
rect 5816 5627 5868 5636
rect 5816 5593 5825 5627
rect 5825 5593 5859 5627
rect 5859 5593 5868 5627
rect 5816 5584 5868 5593
rect 9956 5584 10008 5636
rect 11980 5661 11989 5695
rect 11989 5661 12023 5695
rect 12023 5661 12032 5695
rect 11980 5652 12032 5661
rect 15844 5695 15896 5704
rect 15844 5661 15853 5695
rect 15853 5661 15887 5695
rect 15887 5661 15896 5695
rect 15844 5652 15896 5661
rect 17500 5652 17552 5704
rect 18420 5695 18472 5704
rect 18420 5661 18429 5695
rect 18429 5661 18463 5695
rect 18463 5661 18472 5695
rect 18420 5652 18472 5661
rect 19524 5652 19576 5704
rect 24584 5695 24636 5704
rect 24584 5661 24593 5695
rect 24593 5661 24627 5695
rect 24627 5661 24636 5695
rect 24584 5652 24636 5661
rect 16028 5584 16080 5636
rect 18788 5584 18840 5636
rect 19432 5584 19484 5636
rect 2504 5559 2556 5568
rect 2504 5525 2513 5559
rect 2513 5525 2547 5559
rect 2547 5525 2556 5559
rect 2504 5516 2556 5525
rect 2872 5516 2924 5568
rect 7012 5516 7064 5568
rect 8484 5559 8536 5568
rect 8484 5525 8493 5559
rect 8493 5525 8527 5559
rect 8527 5525 8536 5559
rect 8484 5516 8536 5525
rect 9220 5559 9272 5568
rect 9220 5525 9229 5559
rect 9229 5525 9263 5559
rect 9263 5525 9272 5559
rect 9220 5516 9272 5525
rect 10048 5516 10100 5568
rect 10600 5516 10652 5568
rect 11152 5559 11204 5568
rect 11152 5525 11161 5559
rect 11161 5525 11195 5559
rect 11195 5525 11204 5559
rect 11152 5516 11204 5525
rect 12164 5516 12216 5568
rect 14740 5516 14792 5568
rect 15384 5516 15436 5568
rect 15936 5516 15988 5568
rect 16488 5516 16540 5568
rect 19248 5516 19300 5568
rect 20168 5516 20220 5568
rect 24860 5516 24912 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 1952 5312 2004 5364
rect 3424 5312 3476 5364
rect 4344 5355 4396 5364
rect 4344 5321 4353 5355
rect 4353 5321 4387 5355
rect 4387 5321 4396 5355
rect 4344 5312 4396 5321
rect 4712 5355 4764 5364
rect 4712 5321 4721 5355
rect 4721 5321 4755 5355
rect 4755 5321 4764 5355
rect 4712 5312 4764 5321
rect 5080 5312 5132 5364
rect 5356 5312 5408 5364
rect 6920 5312 6972 5364
rect 8208 5312 8260 5364
rect 9956 5312 10008 5364
rect 11888 5355 11940 5364
rect 11888 5321 11897 5355
rect 11897 5321 11931 5355
rect 11931 5321 11940 5355
rect 11888 5312 11940 5321
rect 12992 5312 13044 5364
rect 13820 5355 13872 5364
rect 2504 5176 2556 5228
rect 2780 5176 2832 5228
rect 4068 5176 4120 5228
rect 5172 5176 5224 5228
rect 6460 5244 6512 5296
rect 8024 5244 8076 5296
rect 8576 5244 8628 5296
rect 10784 5244 10836 5296
rect 10968 5244 11020 5296
rect 12900 5244 12952 5296
rect 13820 5321 13829 5355
rect 13829 5321 13863 5355
rect 13863 5321 13872 5355
rect 13820 5312 13872 5321
rect 14280 5312 14332 5364
rect 15660 5312 15712 5364
rect 16580 5355 16632 5364
rect 16580 5321 16589 5355
rect 16589 5321 16623 5355
rect 16623 5321 16632 5355
rect 16580 5312 16632 5321
rect 18236 5355 18288 5364
rect 18236 5321 18245 5355
rect 18245 5321 18279 5355
rect 18279 5321 18288 5355
rect 18236 5312 18288 5321
rect 18328 5312 18380 5364
rect 21272 5355 21324 5364
rect 21272 5321 21281 5355
rect 21281 5321 21315 5355
rect 21315 5321 21324 5355
rect 21272 5312 21324 5321
rect 22100 5312 22152 5364
rect 23388 5312 23440 5364
rect 23664 5355 23716 5364
rect 23664 5321 23673 5355
rect 23673 5321 23707 5355
rect 23707 5321 23716 5355
rect 23664 5312 23716 5321
rect 24676 5355 24728 5364
rect 24676 5321 24685 5355
rect 24685 5321 24719 5355
rect 24719 5321 24728 5355
rect 24676 5312 24728 5321
rect 26240 5312 26292 5364
rect 15568 5287 15620 5296
rect 7472 5219 7524 5228
rect 7472 5185 7481 5219
rect 7481 5185 7515 5219
rect 7515 5185 7524 5219
rect 8208 5219 8260 5228
rect 7472 5176 7524 5185
rect 8208 5185 8217 5219
rect 8217 5185 8251 5219
rect 8251 5185 8260 5219
rect 8208 5176 8260 5185
rect 9220 5176 9272 5228
rect 10600 5176 10652 5228
rect 11244 5219 11296 5228
rect 11244 5185 11253 5219
rect 11253 5185 11287 5219
rect 11287 5185 11296 5219
rect 11244 5176 11296 5185
rect 11336 5176 11388 5228
rect 12992 5219 13044 5228
rect 1768 5151 1820 5160
rect 1768 5117 1777 5151
rect 1777 5117 1811 5151
rect 1811 5117 1820 5151
rect 1768 5108 1820 5117
rect 3148 5108 3200 5160
rect 3792 5108 3844 5160
rect 5816 5108 5868 5160
rect 7104 5108 7156 5160
rect 7840 5108 7892 5160
rect 3332 5083 3384 5092
rect 3332 5049 3341 5083
rect 3341 5049 3375 5083
rect 3375 5049 3384 5083
rect 3332 5040 3384 5049
rect 7288 5040 7340 5092
rect 1400 5015 1452 5024
rect 1400 4981 1409 5015
rect 1409 4981 1443 5015
rect 1443 4981 1452 5015
rect 1400 4972 1452 4981
rect 1676 4972 1728 5024
rect 2412 5015 2464 5024
rect 2412 4981 2421 5015
rect 2421 4981 2455 5015
rect 2455 4981 2464 5015
rect 2412 4972 2464 4981
rect 6276 4972 6328 5024
rect 6828 4972 6880 5024
rect 8024 5015 8076 5024
rect 8024 4981 8033 5015
rect 8033 4981 8067 5015
rect 8067 4981 8076 5015
rect 8668 5015 8720 5024
rect 8024 4972 8076 4981
rect 8668 4981 8677 5015
rect 8677 4981 8711 5015
rect 8711 4981 8720 5015
rect 8668 4972 8720 4981
rect 8852 4972 8904 5024
rect 9128 5108 9180 5160
rect 10048 5108 10100 5160
rect 10876 5108 10928 5160
rect 12992 5185 13001 5219
rect 13001 5185 13035 5219
rect 13035 5185 13044 5219
rect 12992 5176 13044 5185
rect 13728 5176 13780 5228
rect 15568 5253 15577 5287
rect 15577 5253 15611 5287
rect 15611 5253 15620 5287
rect 15568 5244 15620 5253
rect 15844 5244 15896 5296
rect 16028 5219 16080 5228
rect 16028 5185 16037 5219
rect 16037 5185 16071 5219
rect 16071 5185 16080 5219
rect 16028 5176 16080 5185
rect 23572 5244 23624 5296
rect 23848 5244 23900 5296
rect 24124 5244 24176 5296
rect 9496 5083 9548 5092
rect 9496 5049 9505 5083
rect 9505 5049 9539 5083
rect 9539 5049 9548 5083
rect 9496 5040 9548 5049
rect 11612 5040 11664 5092
rect 11888 5040 11940 5092
rect 13820 5108 13872 5160
rect 15384 5108 15436 5160
rect 15844 5108 15896 5160
rect 18696 5108 18748 5160
rect 9128 5015 9180 5024
rect 9128 4981 9137 5015
rect 9137 4981 9171 5015
rect 9171 4981 9180 5015
rect 9128 4972 9180 4981
rect 10784 4972 10836 5024
rect 11060 5015 11112 5024
rect 11060 4981 11069 5015
rect 11069 4981 11103 5015
rect 11103 4981 11112 5015
rect 11060 4972 11112 4981
rect 11520 4972 11572 5024
rect 12348 4972 12400 5024
rect 12440 5015 12492 5024
rect 12440 4981 12449 5015
rect 12449 4981 12483 5015
rect 12483 4981 12492 5015
rect 12992 5040 13044 5092
rect 13452 5040 13504 5092
rect 14280 5040 14332 5092
rect 14648 5040 14700 5092
rect 18328 5040 18380 5092
rect 19248 5040 19300 5092
rect 19432 5040 19484 5092
rect 21732 5108 21784 5160
rect 23756 5176 23808 5228
rect 25504 5219 25556 5228
rect 25504 5185 25513 5219
rect 25513 5185 25547 5219
rect 25547 5185 25556 5219
rect 25504 5176 25556 5185
rect 23664 5108 23716 5160
rect 25228 5151 25280 5160
rect 25228 5117 25237 5151
rect 25237 5117 25271 5151
rect 25271 5117 25280 5151
rect 25228 5108 25280 5117
rect 21824 5040 21876 5092
rect 24032 5083 24084 5092
rect 24032 5049 24041 5083
rect 24041 5049 24075 5083
rect 24075 5049 24084 5083
rect 24032 5040 24084 5049
rect 12440 4972 12492 4981
rect 20168 5015 20220 5024
rect 20168 4981 20177 5015
rect 20177 4981 20211 5015
rect 20211 4981 20220 5015
rect 20168 4972 20220 4981
rect 20720 5015 20772 5024
rect 20720 4981 20729 5015
rect 20729 4981 20763 5015
rect 20763 4981 20772 5015
rect 20720 4972 20772 4981
rect 21456 4972 21508 5024
rect 24860 4972 24912 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 1768 4768 1820 4820
rect 1952 4811 2004 4820
rect 1952 4777 1961 4811
rect 1961 4777 1995 4811
rect 1995 4777 2004 4811
rect 1952 4768 2004 4777
rect 2504 4811 2556 4820
rect 2504 4777 2513 4811
rect 2513 4777 2547 4811
rect 2547 4777 2556 4811
rect 2504 4768 2556 4777
rect 3240 4768 3292 4820
rect 4436 4811 4488 4820
rect 4436 4777 4445 4811
rect 4445 4777 4479 4811
rect 4479 4777 4488 4811
rect 4436 4768 4488 4777
rect 5540 4811 5592 4820
rect 5540 4777 5549 4811
rect 5549 4777 5583 4811
rect 5583 4777 5592 4811
rect 5540 4768 5592 4777
rect 7012 4768 7064 4820
rect 7288 4811 7340 4820
rect 7288 4777 7297 4811
rect 7297 4777 7331 4811
rect 7331 4777 7340 4811
rect 7288 4768 7340 4777
rect 2596 4700 2648 4752
rect 2780 4700 2832 4752
rect 3332 4700 3384 4752
rect 5816 4700 5868 4752
rect 6000 4700 6052 4752
rect 9128 4768 9180 4820
rect 8392 4743 8444 4752
rect 8392 4709 8401 4743
rect 8401 4709 8435 4743
rect 8435 4709 8444 4743
rect 8392 4700 8444 4709
rect 8484 4700 8536 4752
rect 9496 4768 9548 4820
rect 9772 4768 9824 4820
rect 10692 4768 10744 4820
rect 12348 4811 12400 4820
rect 12348 4777 12357 4811
rect 12357 4777 12391 4811
rect 12391 4777 12400 4811
rect 12348 4768 12400 4777
rect 12716 4768 12768 4820
rect 10968 4700 11020 4752
rect 11244 4700 11296 4752
rect 12900 4743 12952 4752
rect 12900 4709 12909 4743
rect 12909 4709 12943 4743
rect 12943 4709 12952 4743
rect 12900 4700 12952 4709
rect 4068 4632 4120 4684
rect 6368 4632 6420 4684
rect 7012 4632 7064 4684
rect 11336 4675 11388 4684
rect 11336 4641 11345 4675
rect 11345 4641 11379 4675
rect 11379 4641 11388 4675
rect 11336 4632 11388 4641
rect 2504 4564 2556 4616
rect 4528 4607 4580 4616
rect 4528 4573 4537 4607
rect 4537 4573 4571 4607
rect 4571 4573 4580 4607
rect 4528 4564 4580 4573
rect 4712 4607 4764 4616
rect 4712 4573 4721 4607
rect 4721 4573 4755 4607
rect 4755 4573 4764 4607
rect 4712 4564 4764 4573
rect 5448 4564 5500 4616
rect 6276 4607 6328 4616
rect 6276 4573 6285 4607
rect 6285 4573 6319 4607
rect 6319 4573 6328 4607
rect 6276 4564 6328 4573
rect 8208 4564 8260 4616
rect 9404 4564 9456 4616
rect 11152 4564 11204 4616
rect 12164 4564 12216 4616
rect 13636 4768 13688 4820
rect 14004 4768 14056 4820
rect 16028 4768 16080 4820
rect 19432 4811 19484 4820
rect 19432 4777 19441 4811
rect 19441 4777 19475 4811
rect 19475 4777 19484 4811
rect 19432 4768 19484 4777
rect 20260 4768 20312 4820
rect 15292 4700 15344 4752
rect 13820 4675 13872 4684
rect 13820 4641 13829 4675
rect 13829 4641 13863 4675
rect 13863 4641 13872 4675
rect 13820 4632 13872 4641
rect 16488 4632 16540 4684
rect 18696 4700 18748 4752
rect 21732 4768 21784 4820
rect 22284 4768 22336 4820
rect 18328 4675 18380 4684
rect 18328 4641 18362 4675
rect 18362 4641 18380 4675
rect 18328 4632 18380 4641
rect 21272 4675 21324 4684
rect 21272 4641 21281 4675
rect 21281 4641 21315 4675
rect 21315 4641 21324 4675
rect 21272 4632 21324 4641
rect 22560 4700 22612 4752
rect 23388 4768 23440 4820
rect 24124 4768 24176 4820
rect 24860 4768 24912 4820
rect 25596 4768 25648 4820
rect 26240 4811 26292 4820
rect 26240 4777 26249 4811
rect 26249 4777 26283 4811
rect 26283 4777 26292 4811
rect 26240 4768 26292 4777
rect 26332 4700 26384 4752
rect 23940 4632 23992 4684
rect 25044 4632 25096 4684
rect 25780 4675 25832 4684
rect 25780 4641 25789 4675
rect 25789 4641 25823 4675
rect 25823 4641 25832 4675
rect 25780 4632 25832 4641
rect 15292 4607 15344 4616
rect 15292 4573 15301 4607
rect 15301 4573 15335 4607
rect 15335 4573 15344 4607
rect 15292 4564 15344 4573
rect 17960 4564 18012 4616
rect 3332 4496 3384 4548
rect 8576 4496 8628 4548
rect 9864 4496 9916 4548
rect 10140 4496 10192 4548
rect 10784 4539 10836 4548
rect 10784 4505 10793 4539
rect 10793 4505 10827 4539
rect 10827 4505 10836 4539
rect 10784 4496 10836 4505
rect 12256 4496 12308 4548
rect 17868 4496 17920 4548
rect 204 4428 256 4480
rect 8852 4428 8904 4480
rect 11888 4471 11940 4480
rect 11888 4437 11897 4471
rect 11897 4437 11931 4471
rect 11931 4437 11940 4471
rect 11888 4428 11940 4437
rect 13912 4428 13964 4480
rect 14832 4428 14884 4480
rect 16856 4428 16908 4480
rect 17960 4471 18012 4480
rect 17960 4437 17969 4471
rect 17969 4437 18003 4471
rect 18003 4437 18012 4471
rect 17960 4428 18012 4437
rect 20996 4496 21048 4548
rect 21456 4607 21508 4616
rect 21456 4573 21465 4607
rect 21465 4573 21499 4607
rect 21499 4573 21508 4607
rect 22928 4607 22980 4616
rect 21456 4564 21508 4573
rect 22928 4573 22937 4607
rect 22937 4573 22971 4607
rect 22971 4573 22980 4607
rect 22928 4564 22980 4573
rect 21640 4496 21692 4548
rect 21732 4496 21784 4548
rect 24124 4564 24176 4616
rect 23572 4496 23624 4548
rect 19984 4471 20036 4480
rect 19984 4437 19993 4471
rect 19993 4437 20027 4471
rect 20027 4437 20036 4471
rect 19984 4428 20036 4437
rect 22100 4428 22152 4480
rect 24676 4428 24728 4480
rect 25044 4471 25096 4480
rect 25044 4437 25053 4471
rect 25053 4437 25087 4471
rect 25087 4437 25096 4471
rect 25044 4428 25096 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 2412 4224 2464 4276
rect 2596 4224 2648 4276
rect 1216 4156 1268 4208
rect 6000 4224 6052 4276
rect 9680 4267 9732 4276
rect 9680 4233 9689 4267
rect 9689 4233 9723 4267
rect 9723 4233 9732 4267
rect 9680 4224 9732 4233
rect 12164 4224 12216 4276
rect 9220 4156 9272 4208
rect 2136 4088 2188 4140
rect 3976 4131 4028 4140
rect 3976 4097 3985 4131
rect 3985 4097 4019 4131
rect 4019 4097 4028 4131
rect 3976 4088 4028 4097
rect 6276 4088 6328 4140
rect 10968 4156 11020 4208
rect 4712 4020 4764 4072
rect 7472 4063 7524 4072
rect 7472 4029 7495 4063
rect 7495 4029 7524 4063
rect 1860 3995 1912 4004
rect 1860 3961 1869 3995
rect 1869 3961 1903 3995
rect 1903 3961 1912 3995
rect 2872 3995 2924 4004
rect 1860 3952 1912 3961
rect 2872 3961 2881 3995
rect 2881 3961 2915 3995
rect 2915 3961 2924 3995
rect 2872 3952 2924 3961
rect 6092 3952 6144 4004
rect 7012 3952 7064 4004
rect 7472 4020 7524 4029
rect 9956 4020 10008 4072
rect 12900 4156 12952 4208
rect 14004 4224 14056 4276
rect 11428 4088 11480 4140
rect 11336 4020 11388 4072
rect 8116 3952 8168 4004
rect 8392 3952 8444 4004
rect 12624 4088 12676 4140
rect 14464 4156 14516 4208
rect 14648 4156 14700 4208
rect 15752 4224 15804 4276
rect 16028 4224 16080 4276
rect 16212 4224 16264 4276
rect 18420 4267 18472 4276
rect 15844 4156 15896 4208
rect 16488 4156 16540 4208
rect 14556 4131 14608 4140
rect 14556 4097 14565 4131
rect 14565 4097 14599 4131
rect 14599 4097 14608 4131
rect 14556 4088 14608 4097
rect 14924 4088 14976 4140
rect 15568 4088 15620 4140
rect 16304 4088 16356 4140
rect 18420 4233 18429 4267
rect 18429 4233 18463 4267
rect 18463 4233 18472 4267
rect 18420 4224 18472 4233
rect 19432 4267 19484 4276
rect 19432 4233 19441 4267
rect 19441 4233 19475 4267
rect 19475 4233 19484 4267
rect 19432 4224 19484 4233
rect 20812 4224 20864 4276
rect 21640 4224 21692 4276
rect 22928 4224 22980 4276
rect 18328 4156 18380 4208
rect 12532 4020 12584 4072
rect 13544 4020 13596 4072
rect 14372 4063 14424 4072
rect 14372 4029 14381 4063
rect 14381 4029 14415 4063
rect 14415 4029 14424 4063
rect 14372 4020 14424 4029
rect 14648 4020 14700 4072
rect 16396 4020 16448 4072
rect 18788 4088 18840 4140
rect 20168 4156 20220 4208
rect 20444 4131 20496 4140
rect 20444 4097 20453 4131
rect 20453 4097 20487 4131
rect 20487 4097 20496 4131
rect 20444 4088 20496 4097
rect 21732 4156 21784 4208
rect 22376 4156 22428 4208
rect 23756 4156 23808 4208
rect 23940 4156 23992 4208
rect 25780 4224 25832 4276
rect 26240 4224 26292 4276
rect 22560 4088 22612 4140
rect 24216 4088 24268 4140
rect 24676 4088 24728 4140
rect 25872 4156 25924 4208
rect 16948 4020 17000 4072
rect 24584 4020 24636 4072
rect 24952 4020 25004 4072
rect 25228 4063 25280 4072
rect 25228 4029 25237 4063
rect 25237 4029 25271 4063
rect 25271 4029 25280 4063
rect 25228 4020 25280 4029
rect 14096 3952 14148 4004
rect 15568 3952 15620 4004
rect 18696 3952 18748 4004
rect 1584 3884 1636 3936
rect 2320 3884 2372 3936
rect 2964 3927 3016 3936
rect 2964 3893 2973 3927
rect 2973 3893 3007 3927
rect 3007 3893 3016 3927
rect 2964 3884 3016 3893
rect 5356 3927 5408 3936
rect 5356 3893 5365 3927
rect 5365 3893 5399 3927
rect 5399 3893 5408 3927
rect 5356 3884 5408 3893
rect 6368 3927 6420 3936
rect 6368 3893 6377 3927
rect 6377 3893 6411 3927
rect 6411 3893 6420 3927
rect 6368 3884 6420 3893
rect 8300 3884 8352 3936
rect 9128 3927 9180 3936
rect 9128 3893 9137 3927
rect 9137 3893 9171 3927
rect 9171 3893 9180 3927
rect 9128 3884 9180 3893
rect 9956 3884 10008 3936
rect 11428 3927 11480 3936
rect 11428 3893 11437 3927
rect 11437 3893 11471 3927
rect 11471 3893 11480 3927
rect 11428 3884 11480 3893
rect 12624 3884 12676 3936
rect 13452 3927 13504 3936
rect 13452 3893 13461 3927
rect 13461 3893 13495 3927
rect 13495 3893 13504 3927
rect 13452 3884 13504 3893
rect 13820 3884 13872 3936
rect 14004 3927 14056 3936
rect 14004 3893 14013 3927
rect 14013 3893 14047 3927
rect 14047 3893 14056 3927
rect 14004 3884 14056 3893
rect 14740 3884 14792 3936
rect 16948 3927 17000 3936
rect 16948 3893 16957 3927
rect 16957 3893 16991 3927
rect 16991 3893 17000 3927
rect 16948 3884 17000 3893
rect 18788 3927 18840 3936
rect 18788 3893 18797 3927
rect 18797 3893 18831 3927
rect 18831 3893 18840 3927
rect 18788 3884 18840 3893
rect 20628 3952 20680 4004
rect 22284 3952 22336 4004
rect 20352 3927 20404 3936
rect 20352 3893 20361 3927
rect 20361 3893 20395 3927
rect 20395 3893 20404 3927
rect 20352 3884 20404 3893
rect 21364 3927 21416 3936
rect 21364 3893 21373 3927
rect 21373 3893 21407 3927
rect 21407 3893 21416 3927
rect 21364 3884 21416 3893
rect 21824 3884 21876 3936
rect 23664 3927 23716 3936
rect 23664 3893 23673 3927
rect 23673 3893 23707 3927
rect 23707 3893 23716 3927
rect 23664 3884 23716 3893
rect 24124 3952 24176 4004
rect 24860 3952 24912 4004
rect 24216 3884 24268 3936
rect 25412 3927 25464 3936
rect 25412 3893 25421 3927
rect 25421 3893 25455 3927
rect 25455 3893 25464 3927
rect 25412 3884 25464 3893
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 1492 3680 1544 3732
rect 1768 3723 1820 3732
rect 1768 3689 1777 3723
rect 1777 3689 1811 3723
rect 1811 3689 1820 3723
rect 1768 3680 1820 3689
rect 1584 3612 1636 3664
rect 2228 3680 2280 3732
rect 2320 3680 2372 3732
rect 2136 3612 2188 3664
rect 5540 3680 5592 3732
rect 6276 3680 6328 3732
rect 6552 3680 6604 3732
rect 7472 3680 7524 3732
rect 7840 3723 7892 3732
rect 4160 3612 4212 3664
rect 5356 3612 5408 3664
rect 3976 3544 4028 3596
rect 4712 3544 4764 3596
rect 6644 3612 6696 3664
rect 7840 3689 7849 3723
rect 7849 3689 7883 3723
rect 7883 3689 7892 3723
rect 7840 3680 7892 3689
rect 8208 3723 8260 3732
rect 8208 3689 8217 3723
rect 8217 3689 8251 3723
rect 8251 3689 8260 3723
rect 8208 3680 8260 3689
rect 9128 3680 9180 3732
rect 9680 3723 9732 3732
rect 9680 3689 9689 3723
rect 9689 3689 9723 3723
rect 9723 3689 9732 3723
rect 9680 3680 9732 3689
rect 9956 3680 10008 3732
rect 10968 3680 11020 3732
rect 12532 3723 12584 3732
rect 11612 3655 11664 3664
rect 11612 3621 11621 3655
rect 11621 3621 11655 3655
rect 11655 3621 11664 3655
rect 11612 3612 11664 3621
rect 12532 3689 12541 3723
rect 12541 3689 12575 3723
rect 12575 3689 12584 3723
rect 12532 3680 12584 3689
rect 12808 3723 12860 3732
rect 12808 3689 12817 3723
rect 12817 3689 12851 3723
rect 12851 3689 12860 3723
rect 12808 3680 12860 3689
rect 13176 3680 13228 3732
rect 13728 3680 13780 3732
rect 15660 3680 15712 3732
rect 16948 3680 17000 3732
rect 17132 3680 17184 3732
rect 18052 3680 18104 3732
rect 18880 3723 18932 3732
rect 18880 3689 18889 3723
rect 18889 3689 18923 3723
rect 18923 3689 18932 3723
rect 18880 3680 18932 3689
rect 19432 3680 19484 3732
rect 22008 3680 22060 3732
rect 22376 3723 22428 3732
rect 22376 3689 22385 3723
rect 22385 3689 22419 3723
rect 22419 3689 22428 3723
rect 22376 3680 22428 3689
rect 22836 3723 22888 3732
rect 22836 3689 22845 3723
rect 22845 3689 22879 3723
rect 22879 3689 22888 3723
rect 22836 3680 22888 3689
rect 23112 3680 23164 3732
rect 23480 3680 23532 3732
rect 24400 3723 24452 3732
rect 24400 3689 24409 3723
rect 24409 3689 24443 3723
rect 24443 3689 24452 3723
rect 24400 3680 24452 3689
rect 16304 3655 16356 3664
rect 16304 3621 16313 3655
rect 16313 3621 16347 3655
rect 16347 3621 16356 3655
rect 16304 3612 16356 3621
rect 16764 3655 16816 3664
rect 16764 3621 16773 3655
rect 16773 3621 16807 3655
rect 16807 3621 16816 3655
rect 16764 3612 16816 3621
rect 18788 3655 18840 3664
rect 18788 3621 18797 3655
rect 18797 3621 18831 3655
rect 18831 3621 18840 3655
rect 18788 3612 18840 3621
rect 21824 3612 21876 3664
rect 22284 3612 22336 3664
rect 2136 3476 2188 3528
rect 2964 3519 3016 3528
rect 2964 3485 2973 3519
rect 2973 3485 3007 3519
rect 3007 3485 3016 3519
rect 2964 3476 3016 3485
rect 7748 3476 7800 3528
rect 9864 3544 9916 3596
rect 8484 3476 8536 3528
rect 9220 3476 9272 3528
rect 9956 3476 10008 3528
rect 11704 3519 11756 3528
rect 11704 3485 11713 3519
rect 11713 3485 11747 3519
rect 11747 3485 11756 3519
rect 11704 3476 11756 3485
rect 12256 3544 12308 3596
rect 13268 3544 13320 3596
rect 15476 3544 15528 3596
rect 19156 3544 19208 3596
rect 3884 3340 3936 3392
rect 8208 3408 8260 3460
rect 12532 3408 12584 3460
rect 14556 3476 14608 3528
rect 15844 3519 15896 3528
rect 15844 3485 15853 3519
rect 15853 3485 15887 3519
rect 15887 3485 15896 3519
rect 15844 3476 15896 3485
rect 16856 3476 16908 3528
rect 5448 3383 5500 3392
rect 5448 3349 5457 3383
rect 5457 3349 5491 3383
rect 5491 3349 5500 3383
rect 5448 3340 5500 3349
rect 7472 3340 7524 3392
rect 9864 3340 9916 3392
rect 12808 3340 12860 3392
rect 13636 3340 13688 3392
rect 14372 3340 14424 3392
rect 17684 3340 17736 3392
rect 17776 3340 17828 3392
rect 21456 3519 21508 3528
rect 21456 3485 21465 3519
rect 21465 3485 21499 3519
rect 21499 3485 21508 3519
rect 21456 3476 21508 3485
rect 21732 3476 21784 3528
rect 23112 3519 23164 3528
rect 18420 3451 18472 3460
rect 18420 3417 18429 3451
rect 18429 3417 18463 3451
rect 18463 3417 18472 3451
rect 18420 3408 18472 3417
rect 20076 3408 20128 3460
rect 20352 3408 20404 3460
rect 22008 3408 22060 3460
rect 23112 3485 23121 3519
rect 23121 3485 23155 3519
rect 23155 3485 23164 3519
rect 23112 3476 23164 3485
rect 24308 3544 24360 3596
rect 25136 3680 25188 3732
rect 26240 3723 26292 3732
rect 26240 3689 26249 3723
rect 26249 3689 26283 3723
rect 26283 3689 26292 3723
rect 26240 3680 26292 3689
rect 24860 3476 24912 3528
rect 24124 3408 24176 3460
rect 20260 3383 20312 3392
rect 20260 3349 20269 3383
rect 20269 3349 20303 3383
rect 20303 3349 20312 3383
rect 20260 3340 20312 3349
rect 21272 3340 21324 3392
rect 21640 3340 21692 3392
rect 22468 3383 22520 3392
rect 22468 3349 22477 3383
rect 22477 3349 22511 3383
rect 22511 3349 22520 3383
rect 22468 3340 22520 3349
rect 24216 3340 24268 3392
rect 25688 3340 25740 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 2044 3136 2096 3188
rect 4344 3136 4396 3188
rect 5172 3179 5224 3188
rect 5172 3145 5181 3179
rect 5181 3145 5215 3179
rect 5215 3145 5224 3179
rect 5172 3136 5224 3145
rect 5540 3136 5592 3188
rect 1768 3068 1820 3120
rect 3424 3068 3476 3120
rect 7840 3136 7892 3188
rect 8484 3136 8536 3188
rect 8668 3136 8720 3188
rect 9956 3136 10008 3188
rect 11060 3179 11112 3188
rect 11060 3145 11069 3179
rect 11069 3145 11103 3179
rect 11103 3145 11112 3179
rect 11060 3136 11112 3145
rect 11612 3136 11664 3188
rect 9220 3111 9272 3120
rect 9220 3077 9229 3111
rect 9229 3077 9263 3111
rect 9263 3077 9272 3111
rect 9220 3068 9272 3077
rect 11704 3111 11756 3120
rect 11704 3077 11713 3111
rect 11713 3077 11747 3111
rect 11747 3077 11756 3111
rect 14372 3136 14424 3188
rect 16580 3136 16632 3188
rect 16856 3136 16908 3188
rect 18052 3179 18104 3188
rect 18052 3145 18061 3179
rect 18061 3145 18095 3179
rect 18095 3145 18104 3179
rect 18052 3136 18104 3145
rect 18788 3136 18840 3188
rect 19340 3136 19392 3188
rect 20904 3136 20956 3188
rect 21180 3179 21232 3188
rect 21180 3145 21189 3179
rect 21189 3145 21223 3179
rect 21223 3145 21232 3179
rect 21180 3136 21232 3145
rect 22836 3136 22888 3188
rect 23020 3136 23072 3188
rect 23756 3136 23808 3188
rect 24860 3136 24912 3188
rect 25044 3179 25096 3188
rect 25044 3145 25053 3179
rect 25053 3145 25087 3179
rect 25087 3145 25096 3179
rect 25044 3136 25096 3145
rect 26056 3179 26108 3188
rect 26056 3145 26065 3179
rect 26065 3145 26099 3179
rect 26099 3145 26108 3179
rect 26056 3136 26108 3145
rect 26332 3179 26384 3188
rect 26332 3145 26341 3179
rect 26341 3145 26375 3179
rect 26375 3145 26384 3179
rect 26332 3136 26384 3145
rect 11704 3068 11756 3077
rect 13912 3068 13964 3120
rect 2136 3000 2188 3052
rect 3516 3043 3568 3052
rect 3516 3009 3525 3043
rect 3525 3009 3559 3043
rect 3559 3009 3568 3043
rect 4160 3043 4212 3052
rect 3516 3000 3568 3009
rect 4160 3009 4169 3043
rect 4169 3009 4203 3043
rect 4203 3009 4212 3043
rect 4160 3000 4212 3009
rect 4252 2932 4304 2984
rect 6092 2932 6144 2984
rect 7012 3000 7064 3052
rect 17132 3000 17184 3052
rect 18880 3000 18932 3052
rect 20076 3043 20128 3052
rect 20076 3009 20085 3043
rect 20085 3009 20119 3043
rect 20119 3009 20128 3043
rect 20076 3000 20128 3009
rect 20260 3068 20312 3120
rect 21732 3068 21784 3120
rect 23664 3111 23716 3120
rect 23664 3077 23673 3111
rect 23673 3077 23707 3111
rect 23707 3077 23716 3111
rect 23664 3068 23716 3077
rect 23112 3000 23164 3052
rect 1768 2907 1820 2916
rect 1768 2873 1777 2907
rect 1777 2873 1811 2907
rect 1811 2873 1820 2907
rect 1768 2864 1820 2873
rect 2780 2864 2832 2916
rect 3976 2907 4028 2916
rect 3976 2873 3985 2907
rect 3985 2873 4019 2907
rect 4019 2873 4028 2907
rect 3976 2864 4028 2873
rect 1676 2796 1728 2848
rect 4252 2796 4304 2848
rect 7472 2907 7524 2916
rect 7472 2873 7506 2907
rect 7506 2873 7524 2907
rect 7472 2864 7524 2873
rect 7932 2864 7984 2916
rect 11980 2932 12032 2984
rect 15108 2975 15160 2984
rect 15108 2941 15117 2975
rect 15117 2941 15151 2975
rect 15151 2941 15160 2975
rect 15108 2932 15160 2941
rect 17776 2975 17828 2984
rect 17776 2941 17785 2975
rect 17785 2941 17819 2975
rect 17819 2941 17828 2975
rect 17776 2932 17828 2941
rect 17960 2932 18012 2984
rect 18420 2975 18472 2984
rect 18420 2941 18429 2975
rect 18429 2941 18463 2975
rect 18463 2941 18472 2975
rect 18420 2932 18472 2941
rect 18696 2932 18748 2984
rect 20904 2932 20956 2984
rect 23848 2932 23900 2984
rect 24124 2975 24176 2984
rect 9864 2864 9916 2916
rect 11060 2864 11112 2916
rect 12716 2907 12768 2916
rect 12716 2873 12750 2907
rect 12750 2873 12768 2907
rect 12716 2864 12768 2873
rect 15384 2907 15436 2916
rect 15384 2873 15396 2907
rect 15396 2873 15436 2907
rect 15384 2864 15436 2873
rect 15844 2864 15896 2916
rect 20720 2864 20772 2916
rect 20996 2864 21048 2916
rect 23480 2864 23532 2916
rect 24124 2941 24133 2975
rect 24133 2941 24167 2975
rect 24167 2941 24176 2975
rect 24124 2932 24176 2941
rect 26056 2932 26108 2984
rect 6460 2796 6512 2848
rect 9680 2796 9732 2848
rect 13912 2796 13964 2848
rect 14280 2796 14332 2848
rect 14924 2839 14976 2848
rect 14924 2805 14933 2839
rect 14933 2805 14967 2839
rect 14967 2805 14976 2839
rect 25504 2907 25556 2916
rect 25504 2873 25513 2907
rect 25513 2873 25547 2907
rect 25547 2873 25556 2907
rect 25504 2864 25556 2873
rect 14924 2796 14976 2805
rect 23848 2796 23900 2848
rect 24860 2796 24912 2848
rect 25044 2796 25096 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 1584 2592 1636 2644
rect 3332 2592 3384 2644
rect 3516 2635 3568 2644
rect 3516 2601 3525 2635
rect 3525 2601 3559 2635
rect 3559 2601 3568 2635
rect 3516 2592 3568 2601
rect 5264 2592 5316 2644
rect 7932 2592 7984 2644
rect 9588 2635 9640 2644
rect 9588 2601 9597 2635
rect 9597 2601 9631 2635
rect 9631 2601 9640 2635
rect 9588 2592 9640 2601
rect 11060 2592 11112 2644
rect 12348 2592 12400 2644
rect 15476 2635 15528 2644
rect 1676 2567 1728 2576
rect 1676 2533 1685 2567
rect 1685 2533 1719 2567
rect 1719 2533 1728 2567
rect 1676 2524 1728 2533
rect 4712 2524 4764 2576
rect 2872 2431 2924 2440
rect 2872 2397 2881 2431
rect 2881 2397 2915 2431
rect 2915 2397 2924 2431
rect 2872 2388 2924 2397
rect 3516 2388 3568 2440
rect 5080 2456 5132 2508
rect 7472 2567 7524 2576
rect 7472 2533 7506 2567
rect 7506 2533 7524 2567
rect 7472 2524 7524 2533
rect 10784 2524 10836 2576
rect 10876 2524 10928 2576
rect 11704 2524 11756 2576
rect 14924 2524 14976 2576
rect 15476 2601 15485 2635
rect 15485 2601 15519 2635
rect 15519 2601 15528 2635
rect 15476 2592 15528 2601
rect 17040 2592 17092 2644
rect 18328 2635 18380 2644
rect 18328 2601 18337 2635
rect 18337 2601 18371 2635
rect 18371 2601 18380 2635
rect 18328 2592 18380 2601
rect 20812 2592 20864 2644
rect 21180 2635 21232 2644
rect 21180 2601 21189 2635
rect 21189 2601 21223 2635
rect 21223 2601 21232 2635
rect 21180 2592 21232 2601
rect 23020 2635 23072 2644
rect 23020 2601 23029 2635
rect 23029 2601 23063 2635
rect 23063 2601 23072 2635
rect 23020 2592 23072 2601
rect 24768 2592 24820 2644
rect 25044 2635 25096 2644
rect 25044 2601 25053 2635
rect 25053 2601 25087 2635
rect 25087 2601 25096 2635
rect 25044 2592 25096 2601
rect 26332 2592 26384 2644
rect 19432 2524 19484 2576
rect 19892 2524 19944 2576
rect 20904 2524 20956 2576
rect 24124 2524 24176 2576
rect 24492 2567 24544 2576
rect 24492 2533 24501 2567
rect 24501 2533 24535 2567
rect 24535 2533 24544 2567
rect 24492 2524 24544 2533
rect 25596 2567 25648 2576
rect 25596 2533 25605 2567
rect 25605 2533 25639 2567
rect 25639 2533 25648 2567
rect 25596 2524 25648 2533
rect 7012 2456 7064 2508
rect 9036 2456 9088 2508
rect 9496 2456 9548 2508
rect 9680 2456 9732 2508
rect 15108 2456 15160 2508
rect 12072 2431 12124 2440
rect 12072 2397 12081 2431
rect 12081 2397 12115 2431
rect 12115 2397 12124 2431
rect 12072 2388 12124 2397
rect 2412 2363 2464 2372
rect 2412 2329 2421 2363
rect 2421 2329 2455 2363
rect 2455 2329 2464 2363
rect 2412 2320 2464 2329
rect 14280 2363 14332 2372
rect 14280 2329 14289 2363
rect 14289 2329 14323 2363
rect 14323 2329 14332 2363
rect 14280 2320 14332 2329
rect 15384 2320 15436 2372
rect 16488 2388 16540 2440
rect 6552 2252 6604 2304
rect 15476 2252 15528 2304
rect 16120 2252 16172 2304
rect 16948 2456 17000 2508
rect 16672 2252 16724 2304
rect 16948 2295 17000 2304
rect 16948 2261 16957 2295
rect 16957 2261 16991 2295
rect 16991 2261 17000 2295
rect 16948 2252 17000 2261
rect 17132 2252 17184 2304
rect 17592 2252 17644 2304
rect 19800 2456 19852 2508
rect 18880 2431 18932 2440
rect 18880 2397 18889 2431
rect 18889 2397 18923 2431
rect 18923 2397 18932 2431
rect 18880 2388 18932 2397
rect 20536 2431 20588 2440
rect 20536 2397 20545 2431
rect 20545 2397 20579 2431
rect 20579 2397 20588 2431
rect 22928 2456 22980 2508
rect 24216 2456 24268 2508
rect 21732 2431 21784 2440
rect 20536 2388 20588 2397
rect 21732 2397 21741 2431
rect 21741 2397 21775 2431
rect 21775 2397 21784 2431
rect 21732 2388 21784 2397
rect 25044 2388 25096 2440
rect 19800 2295 19852 2304
rect 19800 2261 19809 2295
rect 19809 2261 19843 2295
rect 19843 2261 19852 2295
rect 19800 2252 19852 2261
rect 20168 2295 20220 2304
rect 20168 2261 20177 2295
rect 20177 2261 20211 2295
rect 20211 2261 20220 2295
rect 20168 2252 20220 2261
rect 20904 2295 20956 2304
rect 20904 2261 20913 2295
rect 20913 2261 20947 2295
rect 20947 2261 20956 2295
rect 20904 2252 20956 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 7748 552 7800 604
rect 7840 552 7892 604
rect 11888 552 11940 604
rect 12256 552 12308 604
<< metal2 >>
rect 294 27520 350 28000
rect 846 27520 902 28000
rect 1398 27520 1454 28000
rect 1674 27704 1730 27713
rect 1674 27639 1730 27648
rect 308 22817 336 27520
rect 860 23361 888 27520
rect 1412 25514 1440 27520
rect 1490 27160 1546 27169
rect 1490 27095 1546 27104
rect 1320 25486 1440 25514
rect 1320 24426 1348 25486
rect 1400 25356 1452 25362
rect 1400 25298 1452 25304
rect 1412 24614 1440 25298
rect 1400 24608 1452 24614
rect 1400 24550 1452 24556
rect 1320 24398 1440 24426
rect 1504 24410 1532 27095
rect 1582 25936 1638 25945
rect 1582 25871 1638 25880
rect 1596 24954 1624 25871
rect 1584 24948 1636 24954
rect 1584 24890 1636 24896
rect 1582 24848 1638 24857
rect 1582 24783 1638 24792
rect 846 23352 902 23361
rect 846 23287 902 23296
rect 1412 22817 1440 24398
rect 1492 24404 1544 24410
rect 1492 24346 1544 24352
rect 294 22808 350 22817
rect 294 22743 350 22752
rect 1398 22808 1454 22817
rect 1596 22778 1624 24783
rect 1688 23866 1716 27639
rect 2042 27520 2098 28000
rect 2594 27520 2650 28000
rect 3146 27520 3202 28000
rect 3790 27520 3846 28000
rect 4342 27520 4398 28000
rect 4894 27520 4950 28000
rect 5538 27520 5594 28000
rect 6090 27520 6146 28000
rect 6642 27520 6698 28000
rect 7286 27520 7342 28000
rect 7838 27520 7894 28000
rect 8390 27520 8446 28000
rect 9034 27520 9090 28000
rect 9586 27520 9642 28000
rect 10138 27520 10194 28000
rect 10782 27520 10838 28000
rect 11334 27520 11390 28000
rect 11886 27520 11942 28000
rect 12530 27520 12586 28000
rect 13082 27520 13138 28000
rect 13634 27520 13690 28000
rect 14278 27520 14334 28000
rect 14830 27520 14886 28000
rect 15382 27520 15438 28000
rect 16026 27520 16082 28000
rect 16578 27520 16634 28000
rect 17130 27520 17186 28000
rect 17774 27520 17830 28000
rect 18326 27520 18382 28000
rect 18878 27520 18934 28000
rect 19522 27520 19578 28000
rect 20074 27520 20130 28000
rect 20626 27520 20682 28000
rect 21270 27520 21326 28000
rect 21822 27520 21878 28000
rect 22374 27520 22430 28000
rect 23018 27520 23074 28000
rect 23570 27520 23626 28000
rect 24122 27520 24178 28000
rect 24674 27704 24730 27713
rect 24674 27639 24730 27648
rect 2056 24800 2084 27520
rect 2608 26738 2636 27520
rect 2872 27464 2924 27470
rect 2872 27406 2924 27412
rect 1780 24772 2084 24800
rect 2148 26710 2636 26738
rect 1676 23860 1728 23866
rect 1676 23802 1728 23808
rect 1676 23656 1728 23662
rect 1676 23598 1728 23604
rect 1688 23254 1716 23598
rect 1676 23248 1728 23254
rect 1674 23216 1676 23225
rect 1728 23216 1730 23225
rect 1674 23151 1730 23160
rect 1398 22743 1454 22752
rect 1584 22772 1636 22778
rect 1584 22714 1636 22720
rect 1582 22536 1638 22545
rect 1582 22471 1638 22480
rect 1596 22438 1624 22471
rect 1584 22432 1636 22438
rect 1584 22374 1636 22380
rect 1584 22092 1636 22098
rect 1584 22034 1636 22040
rect 1400 21888 1452 21894
rect 1400 21830 1452 21836
rect 1412 21486 1440 21830
rect 1596 21486 1624 22034
rect 1400 21480 1452 21486
rect 1400 21422 1452 21428
rect 1584 21480 1636 21486
rect 1584 21422 1636 21428
rect 1412 20233 1440 21422
rect 1492 20800 1544 20806
rect 1492 20742 1544 20748
rect 1504 20262 1532 20742
rect 1492 20256 1544 20262
rect 1398 20224 1454 20233
rect 1492 20198 1544 20204
rect 1398 20159 1454 20168
rect 940 19168 992 19174
rect 940 19110 992 19116
rect 952 13161 980 19110
rect 1398 17640 1454 17649
rect 1398 17575 1454 17584
rect 1124 17060 1176 17066
rect 1124 17002 1176 17008
rect 1032 15904 1084 15910
rect 1032 15846 1084 15852
rect 1044 14346 1072 15846
rect 1032 14340 1084 14346
rect 1032 14282 1084 14288
rect 938 13152 994 13161
rect 938 13087 994 13096
rect 1044 10606 1072 14282
rect 1136 13705 1164 17002
rect 1412 16130 1440 17575
rect 1504 16153 1532 20198
rect 1228 16102 1440 16130
rect 1490 16144 1546 16153
rect 1122 13696 1178 13705
rect 1122 13631 1178 13640
rect 1032 10600 1084 10606
rect 1032 10542 1084 10548
rect 1136 9994 1164 13631
rect 1228 12646 1256 16102
rect 1490 16079 1546 16088
rect 1308 15972 1360 15978
rect 1308 15914 1360 15920
rect 1216 12640 1268 12646
rect 1216 12582 1268 12588
rect 1320 12322 1348 15914
rect 1596 15042 1624 21422
rect 1676 21412 1728 21418
rect 1676 21354 1728 21360
rect 1688 20369 1716 21354
rect 1780 21078 1808 24772
rect 2148 24698 2176 26710
rect 2318 26616 2374 26625
rect 2318 26551 2374 26560
rect 1872 24670 2176 24698
rect 1872 21457 1900 24670
rect 2044 24608 2096 24614
rect 2044 24550 2096 24556
rect 2056 24313 2084 24550
rect 2042 24304 2098 24313
rect 2042 24239 2098 24248
rect 2136 24268 2188 24274
rect 2136 24210 2188 24216
rect 1952 23724 2004 23730
rect 1952 23666 2004 23672
rect 1858 21448 1914 21457
rect 1858 21383 1914 21392
rect 1768 21072 1820 21078
rect 1768 21014 1820 21020
rect 1674 20360 1730 20369
rect 1964 20330 1992 23666
rect 2148 23526 2176 24210
rect 2332 23866 2360 26551
rect 2686 25392 2742 25401
rect 2686 25327 2742 25336
rect 2412 24608 2464 24614
rect 2412 24550 2464 24556
rect 2504 24608 2556 24614
rect 2504 24550 2556 24556
rect 2320 23860 2372 23866
rect 2320 23802 2372 23808
rect 2136 23520 2188 23526
rect 2136 23462 2188 23468
rect 2228 23520 2280 23526
rect 2228 23462 2280 23468
rect 2044 22976 2096 22982
rect 2044 22918 2096 22924
rect 1674 20295 1730 20304
rect 1768 20324 1820 20330
rect 1768 20266 1820 20272
rect 1952 20324 2004 20330
rect 1952 20266 2004 20272
rect 1676 19712 1728 19718
rect 1780 19700 1808 20266
rect 1728 19672 1808 19700
rect 1676 19654 1728 19660
rect 1688 19446 1716 19654
rect 1676 19440 1728 19446
rect 1676 19382 1728 19388
rect 2056 19174 2084 22918
rect 2148 22137 2176 23462
rect 2240 22409 2268 23462
rect 2424 23254 2452 24550
rect 2412 23248 2464 23254
rect 2412 23190 2464 23196
rect 2412 23112 2464 23118
rect 2412 23054 2464 23060
rect 2320 22500 2372 22506
rect 2320 22442 2372 22448
rect 2226 22400 2282 22409
rect 2226 22335 2282 22344
rect 2134 22128 2190 22137
rect 2134 22063 2190 22072
rect 2332 19825 2360 22442
rect 2424 22438 2452 23054
rect 2412 22432 2464 22438
rect 2412 22374 2464 22380
rect 2424 22273 2452 22374
rect 2410 22264 2466 22273
rect 2410 22199 2466 22208
rect 2410 21176 2466 21185
rect 2410 21111 2412 21120
rect 2464 21111 2466 21120
rect 2412 21082 2464 21088
rect 2410 21040 2466 21049
rect 2410 20975 2466 20984
rect 2318 19816 2374 19825
rect 2318 19751 2374 19760
rect 2318 19408 2374 19417
rect 2318 19343 2374 19352
rect 2136 19236 2188 19242
rect 2136 19178 2188 19184
rect 2044 19168 2096 19174
rect 2044 19110 2096 19116
rect 2056 18290 2084 19110
rect 2148 18630 2176 19178
rect 2136 18624 2188 18630
rect 2134 18592 2136 18601
rect 2188 18592 2190 18601
rect 2134 18527 2190 18536
rect 2044 18284 2096 18290
rect 2044 18226 2096 18232
rect 1676 18080 1728 18086
rect 1676 18022 1728 18028
rect 1688 17202 1716 18022
rect 2228 17672 2280 17678
rect 2228 17614 2280 17620
rect 1952 17536 2004 17542
rect 1952 17478 2004 17484
rect 1676 17196 1728 17202
rect 1676 17138 1728 17144
rect 1964 16998 1992 17478
rect 1676 16992 1728 16998
rect 1952 16992 2004 16998
rect 1728 16940 1808 16946
rect 1676 16934 1808 16940
rect 1952 16934 2004 16940
rect 1688 16918 1808 16934
rect 1780 16726 1808 16918
rect 1768 16720 1820 16726
rect 1766 16688 1768 16697
rect 1820 16688 1822 16697
rect 1766 16623 1822 16632
rect 1676 15972 1728 15978
rect 1676 15914 1728 15920
rect 1504 15014 1624 15042
rect 1398 14784 1454 14793
rect 1398 14719 1454 14728
rect 1412 14618 1440 14719
rect 1400 14612 1452 14618
rect 1400 14554 1452 14560
rect 1504 13512 1532 15014
rect 1584 14952 1636 14958
rect 1584 14894 1636 14900
rect 1596 13938 1624 14894
rect 1688 14657 1716 15914
rect 1860 15428 1912 15434
rect 1860 15370 1912 15376
rect 1768 14884 1820 14890
rect 1768 14826 1820 14832
rect 1674 14648 1730 14657
rect 1674 14583 1730 14592
rect 1676 14544 1728 14550
rect 1676 14486 1728 14492
rect 1688 13954 1716 14486
rect 1780 14113 1808 14826
rect 1872 14414 1900 15370
rect 1964 15337 1992 16934
rect 2136 16652 2188 16658
rect 2136 16594 2188 16600
rect 2044 16584 2096 16590
rect 2044 16526 2096 16532
rect 2056 16114 2084 16526
rect 2044 16108 2096 16114
rect 2044 16050 2096 16056
rect 2056 15366 2084 16050
rect 2044 15360 2096 15366
rect 1950 15328 2006 15337
rect 2044 15302 2096 15308
rect 1950 15263 2006 15272
rect 1860 14408 1912 14414
rect 1860 14350 1912 14356
rect 1766 14104 1822 14113
rect 1766 14039 1822 14048
rect 1584 13932 1636 13938
rect 1688 13926 1808 13954
rect 1584 13874 1636 13880
rect 1412 13484 1532 13512
rect 1412 12730 1440 13484
rect 1492 13388 1544 13394
rect 1596 13376 1624 13874
rect 1544 13348 1624 13376
rect 1492 13330 1544 13336
rect 1596 12850 1624 13348
rect 1676 13388 1728 13394
rect 1676 13330 1728 13336
rect 1584 12844 1636 12850
rect 1584 12786 1636 12792
rect 1412 12702 1532 12730
rect 1400 12640 1452 12646
rect 1400 12582 1452 12588
rect 1412 12442 1440 12582
rect 1400 12436 1452 12442
rect 1504 12424 1532 12702
rect 1688 12646 1716 13330
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 1504 12396 1624 12424
rect 1400 12378 1452 12384
rect 1320 12294 1532 12322
rect 1400 12096 1452 12102
rect 1400 12038 1452 12044
rect 1412 11234 1440 12038
rect 1320 11206 1440 11234
rect 1320 10962 1348 11206
rect 1400 11144 1452 11150
rect 1398 11112 1400 11121
rect 1452 11112 1454 11121
rect 1398 11047 1454 11056
rect 1320 10934 1440 10962
rect 1124 9988 1176 9994
rect 1124 9930 1176 9936
rect 1308 9512 1360 9518
rect 1308 9454 1360 9460
rect 1320 7868 1348 9454
rect 1412 8090 1440 10934
rect 1400 8084 1452 8090
rect 1400 8026 1452 8032
rect 1400 7880 1452 7886
rect 1320 7840 1400 7868
rect 1400 7822 1452 7828
rect 1412 6866 1440 7822
rect 1400 6860 1452 6866
rect 1400 6802 1452 6808
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 1412 5030 1440 5714
rect 1400 5024 1452 5030
rect 1400 4966 1452 4972
rect 662 4584 718 4593
rect 662 4519 718 4528
rect 204 4480 256 4486
rect 204 4422 256 4428
rect 216 480 244 4422
rect 676 480 704 4519
rect 1412 4321 1440 4966
rect 1398 4312 1454 4321
rect 1398 4247 1454 4256
rect 1216 4208 1268 4214
rect 1216 4150 1268 4156
rect 1228 480 1256 4150
rect 1504 3738 1532 12294
rect 1596 8906 1624 12396
rect 1676 12164 1728 12170
rect 1676 12106 1728 12112
rect 1688 10690 1716 12106
rect 1780 10810 1808 13926
rect 1872 13705 1900 14350
rect 1858 13696 1914 13705
rect 1858 13631 1914 13640
rect 2056 13462 2084 15302
rect 2148 15201 2176 16594
rect 2134 15192 2190 15201
rect 2134 15127 2190 15136
rect 2044 13456 2096 13462
rect 2044 13398 2096 13404
rect 2042 13288 2098 13297
rect 2042 13223 2098 13232
rect 1860 12980 1912 12986
rect 1860 12922 1912 12928
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 1688 10662 1808 10690
rect 1584 8900 1636 8906
rect 1584 8842 1636 8848
rect 1584 8424 1636 8430
rect 1584 8366 1636 8372
rect 1596 7546 1624 8366
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 1596 6322 1624 6802
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 1688 5114 1716 8026
rect 1780 6254 1808 10662
rect 1872 9178 1900 12922
rect 1952 12708 2004 12714
rect 1952 12650 2004 12656
rect 1964 12458 1992 12650
rect 2056 12594 2084 13223
rect 2148 12753 2176 15127
rect 2240 13682 2268 17614
rect 2332 15978 2360 19343
rect 2424 18970 2452 20975
rect 2516 20097 2544 24550
rect 2700 24410 2728 25327
rect 2780 25152 2832 25158
rect 2780 25094 2832 25100
rect 2688 24404 2740 24410
rect 2688 24346 2740 24352
rect 2596 24268 2648 24274
rect 2596 24210 2648 24216
rect 2608 23730 2636 24210
rect 2596 23724 2648 23730
rect 2596 23666 2648 23672
rect 2688 23656 2740 23662
rect 2688 23598 2740 23604
rect 2596 22976 2648 22982
rect 2596 22918 2648 22924
rect 2502 20088 2558 20097
rect 2502 20023 2558 20032
rect 2412 18964 2464 18970
rect 2412 18906 2464 18912
rect 2608 18222 2636 22918
rect 2700 22098 2728 23598
rect 2792 23089 2820 25094
rect 2778 23080 2834 23089
rect 2778 23015 2834 23024
rect 2884 22234 2912 27406
rect 3056 24608 3108 24614
rect 3056 24550 3108 24556
rect 2872 22228 2924 22234
rect 2872 22170 2924 22176
rect 2688 22092 2740 22098
rect 2688 22034 2740 22040
rect 2884 21350 2912 22170
rect 3068 21672 3096 24550
rect 3160 22658 3188 27520
rect 3804 27470 3832 27520
rect 3792 27464 3844 27470
rect 3792 27406 3844 27412
rect 4356 24834 4384 27520
rect 4908 24834 4936 27520
rect 4264 24806 4384 24834
rect 4448 24806 4936 24834
rect 3238 24168 3294 24177
rect 3238 24103 3294 24112
rect 3516 24132 3568 24138
rect 3252 22778 3280 24103
rect 3516 24074 3568 24080
rect 3528 23866 3556 24074
rect 3516 23860 3568 23866
rect 3516 23802 3568 23808
rect 4068 23792 4120 23798
rect 4068 23734 4120 23740
rect 3514 23624 3570 23633
rect 3514 23559 3570 23568
rect 3528 23526 3556 23559
rect 3516 23520 3568 23526
rect 3516 23462 3568 23468
rect 4080 23322 4108 23734
rect 4068 23316 4120 23322
rect 4068 23258 4120 23264
rect 3240 22772 3292 22778
rect 3240 22714 3292 22720
rect 4080 22658 4108 23258
rect 3160 22630 3280 22658
rect 3148 22568 3200 22574
rect 3146 22536 3148 22545
rect 3200 22536 3202 22545
rect 3146 22471 3202 22480
rect 3252 22273 3280 22630
rect 3988 22630 4108 22658
rect 3332 22432 3384 22438
rect 3332 22374 3384 22380
rect 3238 22264 3294 22273
rect 3238 22199 3294 22208
rect 3068 21644 3188 21672
rect 3056 21548 3108 21554
rect 3056 21490 3108 21496
rect 2962 21448 3018 21457
rect 2962 21383 3018 21392
rect 2872 21344 2924 21350
rect 2792 21304 2872 21332
rect 2688 21072 2740 21078
rect 2688 21014 2740 21020
rect 2700 20602 2728 21014
rect 2792 20618 2820 21304
rect 2872 21286 2924 21292
rect 2976 21010 3004 21383
rect 2964 21004 3016 21010
rect 2964 20946 3016 20952
rect 2688 20596 2740 20602
rect 2792 20590 2912 20618
rect 2976 20602 3004 20946
rect 3068 20942 3096 21490
rect 3056 20936 3108 20942
rect 3056 20878 3108 20884
rect 2688 20538 2740 20544
rect 2780 20528 2832 20534
rect 2780 20470 2832 20476
rect 2884 20482 2912 20590
rect 2964 20596 3016 20602
rect 2964 20538 3016 20544
rect 3068 20534 3096 20878
rect 3056 20528 3108 20534
rect 2688 19848 2740 19854
rect 2688 19790 2740 19796
rect 2700 19378 2728 19790
rect 2688 19372 2740 19378
rect 2688 19314 2740 19320
rect 2700 18698 2728 19314
rect 2792 19242 2820 20470
rect 2884 20454 3004 20482
rect 3056 20470 3108 20476
rect 2872 19712 2924 19718
rect 2872 19654 2924 19660
rect 2780 19236 2832 19242
rect 2780 19178 2832 19184
rect 2884 19174 2912 19654
rect 2976 19281 3004 20454
rect 3068 19854 3096 20470
rect 3160 19990 3188 21644
rect 3252 21418 3280 22199
rect 3240 21412 3292 21418
rect 3240 21354 3292 21360
rect 3344 20330 3372 22374
rect 3608 21956 3660 21962
rect 3608 21898 3660 21904
rect 3516 21888 3568 21894
rect 3516 21830 3568 21836
rect 3528 21690 3556 21830
rect 3516 21684 3568 21690
rect 3516 21626 3568 21632
rect 3422 21584 3478 21593
rect 3422 21519 3478 21528
rect 3332 20324 3384 20330
rect 3332 20266 3384 20272
rect 3344 20058 3372 20266
rect 3332 20052 3384 20058
rect 3332 19994 3384 20000
rect 3148 19984 3200 19990
rect 3148 19926 3200 19932
rect 3240 19916 3292 19922
rect 3240 19858 3292 19864
rect 3056 19848 3108 19854
rect 3056 19790 3108 19796
rect 3148 19848 3200 19854
rect 3148 19790 3200 19796
rect 3252 19802 3280 19858
rect 3436 19802 3464 21519
rect 3528 20466 3556 21626
rect 3516 20460 3568 20466
rect 3516 20402 3568 20408
rect 3514 19952 3570 19961
rect 3514 19887 3570 19896
rect 3160 19700 3188 19790
rect 3068 19672 3188 19700
rect 3252 19774 3464 19802
rect 2962 19272 3018 19281
rect 2962 19207 3018 19216
rect 2872 19168 2924 19174
rect 2872 19110 2924 19116
rect 2780 18896 2832 18902
rect 2780 18838 2832 18844
rect 2688 18692 2740 18698
rect 2688 18634 2740 18640
rect 2596 18216 2648 18222
rect 2596 18158 2648 18164
rect 2608 17882 2636 18158
rect 2596 17876 2648 17882
rect 2596 17818 2648 17824
rect 2504 17672 2556 17678
rect 2504 17614 2556 17620
rect 2516 17066 2544 17614
rect 2700 17610 2728 18634
rect 2792 18426 2820 18838
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 2780 17740 2832 17746
rect 2780 17682 2832 17688
rect 2688 17604 2740 17610
rect 2688 17546 2740 17552
rect 2596 17536 2648 17542
rect 2596 17478 2648 17484
rect 2608 17134 2636 17478
rect 2596 17128 2648 17134
rect 2596 17070 2648 17076
rect 2504 17060 2556 17066
rect 2504 17002 2556 17008
rect 2608 16674 2636 17070
rect 2700 16794 2728 17546
rect 2792 17338 2820 17682
rect 2780 17332 2832 17338
rect 2780 17274 2832 17280
rect 2792 16794 2820 17274
rect 2688 16788 2740 16794
rect 2688 16730 2740 16736
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 2412 16652 2464 16658
rect 2608 16646 2820 16674
rect 2412 16594 2464 16600
rect 2320 15972 2372 15978
rect 2320 15914 2372 15920
rect 2320 15496 2372 15502
rect 2320 15438 2372 15444
rect 2332 15094 2360 15438
rect 2320 15088 2372 15094
rect 2320 15030 2372 15036
rect 2332 13870 2360 15030
rect 2424 14550 2452 16594
rect 2504 16448 2556 16454
rect 2504 16390 2556 16396
rect 2516 15434 2544 16390
rect 2596 15904 2648 15910
rect 2596 15846 2648 15852
rect 2686 15872 2742 15881
rect 2504 15428 2556 15434
rect 2504 15370 2556 15376
rect 2608 15366 2636 15846
rect 2686 15807 2742 15816
rect 2700 15706 2728 15807
rect 2688 15700 2740 15706
rect 2688 15642 2740 15648
rect 2596 15360 2648 15366
rect 2596 15302 2648 15308
rect 2504 14884 2556 14890
rect 2504 14826 2556 14832
rect 2516 14618 2544 14826
rect 2504 14612 2556 14618
rect 2504 14554 2556 14560
rect 2412 14544 2464 14550
rect 2412 14486 2464 14492
rect 2516 14414 2544 14554
rect 2504 14408 2556 14414
rect 2504 14350 2556 14356
rect 2516 14074 2544 14350
rect 2504 14068 2556 14074
rect 2504 14010 2556 14016
rect 2688 14000 2740 14006
rect 2688 13942 2740 13948
rect 2320 13864 2372 13870
rect 2320 13806 2372 13812
rect 2504 13796 2556 13802
rect 2504 13738 2556 13744
rect 2240 13654 2360 13682
rect 2134 12744 2190 12753
rect 2134 12679 2190 12688
rect 2056 12566 2176 12594
rect 1964 12430 2084 12458
rect 2148 12442 2176 12566
rect 1950 12336 2006 12345
rect 1950 12271 2006 12280
rect 1964 10826 1992 12271
rect 2056 12170 2084 12430
rect 2136 12436 2188 12442
rect 2136 12378 2188 12384
rect 2332 12322 2360 13654
rect 2148 12294 2360 12322
rect 2044 12164 2096 12170
rect 2044 12106 2096 12112
rect 1964 10798 2084 10826
rect 1952 10668 2004 10674
rect 1952 10610 2004 10616
rect 1964 10266 1992 10610
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 1952 10124 2004 10130
rect 1952 10066 2004 10072
rect 1964 9654 1992 10066
rect 1952 9648 2004 9654
rect 1952 9590 2004 9596
rect 1860 9172 1912 9178
rect 1860 9114 1912 9120
rect 1964 8362 1992 9590
rect 1952 8356 2004 8362
rect 1952 8298 2004 8304
rect 1860 7200 1912 7206
rect 1860 7142 1912 7148
rect 1768 6248 1820 6254
rect 1768 6190 1820 6196
rect 1768 6112 1820 6118
rect 1768 6054 1820 6060
rect 1780 5166 1808 6054
rect 1872 5914 1900 7142
rect 1950 6896 2006 6905
rect 1950 6831 2006 6840
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 1964 5778 1992 6831
rect 1952 5772 2004 5778
rect 1952 5714 2004 5720
rect 1964 5522 1992 5714
rect 1872 5494 1992 5522
rect 1596 5086 1716 5114
rect 1768 5160 1820 5166
rect 1768 5102 1820 5108
rect 1596 3942 1624 5086
rect 1676 5024 1728 5030
rect 1676 4966 1728 4972
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1688 3754 1716 4966
rect 1872 4842 1900 5494
rect 1952 5364 2004 5370
rect 1952 5306 2004 5312
rect 1780 4826 1900 4842
rect 1964 4826 1992 5306
rect 1768 4820 1900 4826
rect 1820 4814 1900 4820
rect 1952 4820 2004 4826
rect 1768 4762 1820 4768
rect 1952 4762 2004 4768
rect 1858 4448 1914 4457
rect 1858 4383 1914 4392
rect 1872 4010 1900 4383
rect 1860 4004 1912 4010
rect 1860 3946 1912 3952
rect 1766 3768 1822 3777
rect 1492 3732 1544 3738
rect 1688 3726 1766 3754
rect 1766 3703 1768 3712
rect 1492 3674 1544 3680
rect 1820 3703 1822 3712
rect 1768 3674 1820 3680
rect 1584 3664 1636 3670
rect 1584 3606 1636 3612
rect 1596 3233 1624 3606
rect 1582 3224 1638 3233
rect 1582 3159 1638 3168
rect 1596 2650 1624 3159
rect 1780 3126 1808 3674
rect 2056 3194 2084 10798
rect 2148 9722 2176 12294
rect 2516 12186 2544 13738
rect 2700 12730 2728 13942
rect 2792 13938 2820 16646
rect 2884 16182 2912 19110
rect 3068 18306 3096 19672
rect 3252 19514 3280 19774
rect 3422 19680 3478 19689
rect 3422 19615 3478 19624
rect 3330 19544 3386 19553
rect 3240 19508 3292 19514
rect 3330 19479 3386 19488
rect 3240 19450 3292 19456
rect 3240 19372 3292 19378
rect 3240 19314 3292 19320
rect 3148 18692 3200 18698
rect 3148 18634 3200 18640
rect 3160 18426 3188 18634
rect 3148 18420 3200 18426
rect 3148 18362 3200 18368
rect 3068 18278 3188 18306
rect 2964 17196 3016 17202
rect 2964 17138 3016 17144
rect 2872 16176 2924 16182
rect 2872 16118 2924 16124
rect 2976 15502 3004 17138
rect 3056 16992 3108 16998
rect 3056 16934 3108 16940
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 2870 15328 2926 15337
rect 2870 15263 2926 15272
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2780 13728 2832 13734
rect 2780 13670 2832 13676
rect 2332 12158 2544 12186
rect 2608 12702 2728 12730
rect 2228 11688 2280 11694
rect 2228 11630 2280 11636
rect 2240 11529 2268 11630
rect 2226 11520 2282 11529
rect 2226 11455 2282 11464
rect 2332 10452 2360 12158
rect 2608 11642 2636 12702
rect 2688 12640 2740 12646
rect 2688 12582 2740 12588
rect 2700 12374 2728 12582
rect 2688 12368 2740 12374
rect 2688 12310 2740 12316
rect 2424 11614 2636 11642
rect 2424 10606 2452 11614
rect 2596 11552 2648 11558
rect 2792 11506 2820 13670
rect 2596 11494 2648 11500
rect 2504 11144 2556 11150
rect 2504 11086 2556 11092
rect 2516 10810 2544 11086
rect 2504 10804 2556 10810
rect 2504 10746 2556 10752
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2504 10464 2556 10470
rect 2332 10424 2452 10452
rect 2228 9920 2280 9926
rect 2228 9862 2280 9868
rect 2136 9716 2188 9722
rect 2136 9658 2188 9664
rect 2240 8430 2268 9862
rect 2320 9444 2372 9450
rect 2320 9386 2372 9392
rect 2332 9178 2360 9386
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2228 8424 2280 8430
rect 2228 8366 2280 8372
rect 2228 8288 2280 8294
rect 2228 8230 2280 8236
rect 2136 6248 2188 6254
rect 2136 6190 2188 6196
rect 2148 4146 2176 6190
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 2148 3670 2176 4082
rect 2240 3738 2268 8230
rect 2332 8090 2360 9114
rect 2424 8498 2452 10424
rect 2504 10406 2556 10412
rect 2516 10180 2544 10406
rect 2608 10305 2636 11494
rect 2700 11478 2820 11506
rect 2700 11354 2728 11478
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2688 11076 2740 11082
rect 2688 11018 2740 11024
rect 2594 10296 2650 10305
rect 2594 10231 2650 10240
rect 2516 10152 2636 10180
rect 2504 9716 2556 9722
rect 2504 9658 2556 9664
rect 2412 8492 2464 8498
rect 2412 8434 2464 8440
rect 2320 8084 2372 8090
rect 2320 8026 2372 8032
rect 2332 7546 2360 8026
rect 2320 7540 2372 7546
rect 2320 7482 2372 7488
rect 2516 6610 2544 9658
rect 2332 6582 2544 6610
rect 2332 3942 2360 6582
rect 2504 5568 2556 5574
rect 2504 5510 2556 5516
rect 2410 5400 2466 5409
rect 2410 5335 2466 5344
rect 2424 5030 2452 5335
rect 2516 5234 2544 5510
rect 2504 5228 2556 5234
rect 2504 5170 2556 5176
rect 2412 5024 2464 5030
rect 2412 4966 2464 4972
rect 2516 4826 2544 5170
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2516 4622 2544 4762
rect 2608 4758 2636 10152
rect 2700 8634 2728 11018
rect 2792 10266 2820 11290
rect 2884 11082 2912 15263
rect 2976 14498 3004 15438
rect 3068 15162 3096 16934
rect 3160 16017 3188 18278
rect 3252 17134 3280 19314
rect 3240 17128 3292 17134
rect 3240 17070 3292 17076
rect 3240 16992 3292 16998
rect 3240 16934 3292 16940
rect 3252 16658 3280 16934
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 3146 16008 3202 16017
rect 3146 15943 3202 15952
rect 3148 15904 3200 15910
rect 3148 15846 3200 15852
rect 3160 15706 3188 15846
rect 3148 15700 3200 15706
rect 3148 15642 3200 15648
rect 3148 15428 3200 15434
rect 3148 15370 3200 15376
rect 3056 15156 3108 15162
rect 3056 15098 3108 15104
rect 3068 14618 3096 15098
rect 3056 14612 3108 14618
rect 3056 14554 3108 14560
rect 2976 14470 3096 14498
rect 2964 14272 3016 14278
rect 2964 14214 3016 14220
rect 2976 13870 3004 14214
rect 2964 13864 3016 13870
rect 2964 13806 3016 13812
rect 2976 13190 3004 13806
rect 2964 13184 3016 13190
rect 2964 13126 3016 13132
rect 2872 11076 2924 11082
rect 2872 11018 2924 11024
rect 2870 10976 2926 10985
rect 2870 10911 2926 10920
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2780 10124 2832 10130
rect 2884 10112 2912 10911
rect 2976 10674 3004 13126
rect 3068 12714 3096 14470
rect 3160 14074 3188 15370
rect 3148 14068 3200 14074
rect 3148 14010 3200 14016
rect 3252 13734 3280 16594
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 3344 13546 3372 19479
rect 3436 18766 3464 19615
rect 3424 18760 3476 18766
rect 3424 18702 3476 18708
rect 3436 17882 3464 18702
rect 3528 18426 3556 19887
rect 3620 19174 3648 21898
rect 3882 21856 3938 21865
rect 3882 21791 3938 21800
rect 3700 20800 3752 20806
rect 3700 20742 3752 20748
rect 3608 19168 3660 19174
rect 3608 19110 3660 19116
rect 3620 18970 3648 19110
rect 3608 18964 3660 18970
rect 3608 18906 3660 18912
rect 3516 18420 3568 18426
rect 3516 18362 3568 18368
rect 3712 18290 3740 20742
rect 3790 20088 3846 20097
rect 3790 20023 3846 20032
rect 3804 19854 3832 20023
rect 3792 19848 3844 19854
rect 3792 19790 3844 19796
rect 3792 19712 3844 19718
rect 3792 19654 3844 19660
rect 3804 19417 3832 19654
rect 3790 19408 3846 19417
rect 3790 19343 3846 19352
rect 3896 18970 3924 21791
rect 3988 19174 4016 22630
rect 4160 21888 4212 21894
rect 4160 21830 4212 21836
rect 4172 21350 4200 21830
rect 4264 21593 4292 24806
rect 4344 22976 4396 22982
rect 4344 22918 4396 22924
rect 4250 21584 4306 21593
rect 4356 21554 4384 22918
rect 4250 21519 4306 21528
rect 4344 21548 4396 21554
rect 4344 21490 4396 21496
rect 4160 21344 4212 21350
rect 4066 21312 4122 21321
rect 4160 21286 4212 21292
rect 4066 21247 4122 21256
rect 4080 20505 4108 21247
rect 4172 20602 4200 21286
rect 4252 21072 4304 21078
rect 4250 21040 4252 21049
rect 4304 21040 4306 21049
rect 4250 20975 4306 20984
rect 4252 20800 4304 20806
rect 4252 20742 4304 20748
rect 4344 20800 4396 20806
rect 4344 20742 4396 20748
rect 4160 20596 4212 20602
rect 4160 20538 4212 20544
rect 4066 20496 4122 20505
rect 4066 20431 4122 20440
rect 4160 20460 4212 20466
rect 4160 20402 4212 20408
rect 4172 20262 4200 20402
rect 4160 20256 4212 20262
rect 4160 20198 4212 20204
rect 4172 19922 4200 20198
rect 4160 19916 4212 19922
rect 4160 19858 4212 19864
rect 4068 19848 4120 19854
rect 4068 19790 4120 19796
rect 4080 19553 4108 19790
rect 4066 19544 4122 19553
rect 4066 19479 4122 19488
rect 4066 19408 4122 19417
rect 4172 19378 4200 19858
rect 4066 19343 4122 19352
rect 4160 19372 4212 19378
rect 4080 19310 4108 19343
rect 4160 19314 4212 19320
rect 4068 19304 4120 19310
rect 4068 19246 4120 19252
rect 3976 19168 4028 19174
rect 3976 19110 4028 19116
rect 3884 18964 3936 18970
rect 3884 18906 3936 18912
rect 4172 18698 4200 19314
rect 4160 18692 4212 18698
rect 4160 18634 4212 18640
rect 4264 18578 4292 20742
rect 4356 18902 4384 20742
rect 4344 18896 4396 18902
rect 4344 18838 4396 18844
rect 4172 18550 4292 18578
rect 4066 18456 4122 18465
rect 4066 18391 4122 18400
rect 3700 18284 3752 18290
rect 3700 18226 3752 18232
rect 3976 18216 4028 18222
rect 3976 18158 4028 18164
rect 3988 18057 4016 18158
rect 3974 18048 4030 18057
rect 3974 17983 4030 17992
rect 3424 17876 3476 17882
rect 3424 17818 3476 17824
rect 3608 17536 3660 17542
rect 3608 17478 3660 17484
rect 3516 17196 3568 17202
rect 3516 17138 3568 17144
rect 3424 17128 3476 17134
rect 3424 17070 3476 17076
rect 3436 16674 3464 17070
rect 3528 16969 3556 17138
rect 3620 16998 3648 17478
rect 3974 17232 4030 17241
rect 3974 17167 4030 17176
rect 3698 17096 3754 17105
rect 3698 17031 3754 17040
rect 3608 16992 3660 16998
rect 3514 16960 3570 16969
rect 3608 16934 3660 16940
rect 3514 16895 3570 16904
rect 3528 16794 3556 16895
rect 3516 16788 3568 16794
rect 3516 16730 3568 16736
rect 3436 16646 3556 16674
rect 3424 16516 3476 16522
rect 3424 16458 3476 16464
rect 3436 16114 3464 16458
rect 3424 16108 3476 16114
rect 3424 16050 3476 16056
rect 3436 15502 3464 16050
rect 3528 15910 3556 16646
rect 3516 15904 3568 15910
rect 3516 15846 3568 15852
rect 3424 15496 3476 15502
rect 3424 15438 3476 15444
rect 3422 14648 3478 14657
rect 3422 14583 3478 14592
rect 3252 13518 3372 13546
rect 3148 13252 3200 13258
rect 3148 13194 3200 13200
rect 3160 13161 3188 13194
rect 3146 13152 3202 13161
rect 3146 13087 3202 13096
rect 3056 12708 3108 12714
rect 3056 12650 3108 12656
rect 3056 12232 3108 12238
rect 3056 12174 3108 12180
rect 3068 11286 3096 12174
rect 3252 11898 3280 13518
rect 3332 13184 3384 13190
rect 3332 13126 3384 13132
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 3238 11656 3294 11665
rect 3238 11591 3294 11600
rect 3056 11280 3108 11286
rect 3056 11222 3108 11228
rect 3148 11212 3200 11218
rect 3148 11154 3200 11160
rect 3054 10840 3110 10849
rect 3054 10775 3110 10784
rect 2964 10668 3016 10674
rect 2964 10610 3016 10616
rect 2832 10084 2912 10112
rect 2780 10066 2832 10072
rect 2964 10056 3016 10062
rect 2964 9998 3016 10004
rect 2872 9920 2924 9926
rect 2872 9862 2924 9868
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 2792 8945 2820 8978
rect 2778 8936 2834 8945
rect 2778 8871 2834 8880
rect 2884 8786 2912 9862
rect 2976 9518 3004 9998
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2792 8758 2912 8786
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 2700 7274 2728 8570
rect 2688 7268 2740 7274
rect 2688 7210 2740 7216
rect 2792 7041 2820 8758
rect 2976 8566 3004 8910
rect 2964 8560 3016 8566
rect 2964 8502 3016 8508
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 2884 8294 2912 8434
rect 2964 8356 3016 8362
rect 2964 8298 3016 8304
rect 2872 8288 2924 8294
rect 2872 8230 2924 8236
rect 2884 7954 2912 8230
rect 2872 7948 2924 7954
rect 2872 7890 2924 7896
rect 2884 7206 2912 7890
rect 2976 7324 3004 8298
rect 3068 7449 3096 10775
rect 3160 10266 3188 11154
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 3160 8294 3188 8774
rect 3252 8362 3280 11591
rect 3344 11354 3372 13126
rect 3436 12442 3464 14583
rect 3528 13841 3556 15846
rect 3514 13832 3570 13841
rect 3514 13767 3570 13776
rect 3620 13569 3648 16934
rect 3606 13560 3662 13569
rect 3606 13495 3662 13504
rect 3712 13274 3740 17031
rect 3884 16176 3936 16182
rect 3884 16118 3936 16124
rect 3896 15910 3924 16118
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 3792 14952 3844 14958
rect 3792 14894 3844 14900
rect 3804 14550 3832 14894
rect 3792 14544 3844 14550
rect 3792 14486 3844 14492
rect 3620 13246 3740 13274
rect 3620 12782 3648 13246
rect 3700 13184 3752 13190
rect 3700 13126 3752 13132
rect 3608 12776 3660 12782
rect 3608 12718 3660 12724
rect 3516 12640 3568 12646
rect 3516 12582 3568 12588
rect 3608 12640 3660 12646
rect 3608 12582 3660 12588
rect 3424 12436 3476 12442
rect 3424 12378 3476 12384
rect 3424 11824 3476 11830
rect 3422 11792 3424 11801
rect 3476 11792 3478 11801
rect 3422 11727 3478 11736
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3332 11348 3384 11354
rect 3332 11290 3384 11296
rect 3332 11076 3384 11082
rect 3332 11018 3384 11024
rect 3344 9110 3372 11018
rect 3332 9104 3384 9110
rect 3332 9046 3384 9052
rect 3240 8356 3292 8362
rect 3240 8298 3292 8304
rect 3344 8294 3372 9046
rect 3148 8288 3200 8294
rect 3332 8288 3384 8294
rect 3148 8230 3200 8236
rect 3238 8256 3294 8265
rect 3160 7546 3188 8230
rect 3332 8230 3384 8236
rect 3238 8191 3294 8200
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 3054 7440 3110 7449
rect 3054 7375 3110 7384
rect 2976 7296 3096 7324
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 2778 7032 2834 7041
rect 2778 6967 2834 6976
rect 2688 6180 2740 6186
rect 2740 6140 2820 6168
rect 2688 6122 2740 6128
rect 2792 5234 2820 6140
rect 3068 6089 3096 7296
rect 3148 7200 3200 7206
rect 3148 7142 3200 7148
rect 3160 6662 3188 7142
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 3054 6080 3110 6089
rect 3054 6015 3110 6024
rect 3160 5914 3188 6598
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 2872 5840 2924 5846
rect 2872 5782 2924 5788
rect 2884 5574 2912 5782
rect 3160 5642 3188 5850
rect 3148 5636 3200 5642
rect 3148 5578 3200 5584
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2780 5228 2832 5234
rect 2780 5170 2832 5176
rect 3148 5160 3200 5166
rect 3148 5102 3200 5108
rect 2596 4752 2648 4758
rect 2596 4694 2648 4700
rect 2780 4752 2832 4758
rect 2780 4694 2832 4700
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 2608 4282 2636 4694
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 2596 4276 2648 4282
rect 2596 4218 2648 4224
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 2332 3738 2360 3878
rect 2228 3732 2280 3738
rect 2228 3674 2280 3680
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 2136 3664 2188 3670
rect 2136 3606 2188 3612
rect 2148 3534 2176 3606
rect 2136 3528 2188 3534
rect 2136 3470 2188 3476
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 1768 3120 1820 3126
rect 1768 3062 1820 3068
rect 1858 3088 1914 3097
rect 2148 3058 2176 3470
rect 1858 3023 1914 3032
rect 2136 3052 2188 3058
rect 1768 2916 1820 2922
rect 1768 2858 1820 2864
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 1688 2582 1716 2790
rect 1676 2576 1728 2582
rect 1676 2518 1728 2524
rect 1688 921 1716 2518
rect 1780 1465 1808 2858
rect 1766 1456 1822 1465
rect 1766 1391 1822 1400
rect 1872 1306 1900 3023
rect 2136 2994 2188 3000
rect 2424 2689 2452 4218
rect 2792 2922 2820 4694
rect 2872 4004 2924 4010
rect 2872 3946 2924 3952
rect 2884 3505 2912 3946
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 3054 3904 3110 3913
rect 2976 3777 3004 3878
rect 3054 3839 3110 3848
rect 2962 3768 3018 3777
rect 2962 3703 3018 3712
rect 2964 3528 3016 3534
rect 2870 3496 2926 3505
rect 2964 3470 3016 3476
rect 2870 3431 2926 3440
rect 2780 2916 2832 2922
rect 2780 2858 2832 2864
rect 2410 2680 2466 2689
rect 2410 2615 2466 2624
rect 2318 2544 2374 2553
rect 2318 2479 2374 2488
rect 1780 1278 1900 1306
rect 1674 912 1730 921
rect 1674 847 1730 856
rect 1780 480 1808 1278
rect 2332 480 2360 2479
rect 2872 2440 2924 2446
rect 2410 2408 2466 2417
rect 2872 2382 2924 2388
rect 2410 2343 2412 2352
rect 2464 2343 2466 2352
rect 2412 2314 2464 2320
rect 2884 1737 2912 2382
rect 2870 1728 2926 1737
rect 2870 1663 2926 1672
rect 2976 1578 3004 3470
rect 2792 1550 3004 1578
rect 2792 1329 2820 1550
rect 3068 1442 3096 3839
rect 2884 1414 3096 1442
rect 2778 1320 2834 1329
rect 2778 1255 2834 1264
rect 2884 480 2912 1414
rect 202 0 258 480
rect 662 0 718 480
rect 1214 0 1270 480
rect 1766 0 1822 480
rect 2318 0 2374 480
rect 2870 0 2926 480
rect 3160 377 3188 5102
rect 3252 4826 3280 8191
rect 3332 7744 3384 7750
rect 3332 7686 3384 7692
rect 3344 7342 3372 7686
rect 3332 7336 3384 7342
rect 3332 7278 3384 7284
rect 3436 7154 3464 11494
rect 3528 10198 3556 12582
rect 3620 12238 3648 12582
rect 3608 12232 3660 12238
rect 3608 12174 3660 12180
rect 3608 11756 3660 11762
rect 3608 11698 3660 11704
rect 3620 11286 3648 11698
rect 3608 11280 3660 11286
rect 3608 11222 3660 11228
rect 3712 11218 3740 13126
rect 3896 12866 3924 15846
rect 3988 15484 4016 17167
rect 4080 16538 4108 18391
rect 4172 18086 4200 18550
rect 4160 18080 4212 18086
rect 4160 18022 4212 18028
rect 4172 17241 4200 18022
rect 4448 17864 4476 24806
rect 5552 24177 5580 27520
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 6104 24834 6132 27520
rect 6368 25900 6420 25906
rect 6368 25842 6420 25848
rect 6012 24806 6132 24834
rect 5538 24168 5594 24177
rect 5538 24103 5594 24112
rect 5264 24064 5316 24070
rect 5264 24006 5316 24012
rect 5276 23594 5304 24006
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5540 23656 5592 23662
rect 5446 23624 5502 23633
rect 5264 23588 5316 23594
rect 5540 23598 5592 23604
rect 5446 23559 5502 23568
rect 5264 23530 5316 23536
rect 5460 23526 5488 23559
rect 4620 23520 4672 23526
rect 5448 23520 5500 23526
rect 4620 23462 4672 23468
rect 5354 23488 5410 23497
rect 4528 22432 4580 22438
rect 4528 22374 4580 22380
rect 4540 18290 4568 22374
rect 4528 18284 4580 18290
rect 4528 18226 4580 18232
rect 4448 17836 4568 17864
rect 4436 17740 4488 17746
rect 4436 17682 4488 17688
rect 4448 17338 4476 17682
rect 4436 17332 4488 17338
rect 4436 17274 4488 17280
rect 4158 17232 4214 17241
rect 4158 17167 4214 17176
rect 4344 16992 4396 16998
rect 4344 16934 4396 16940
rect 4250 16824 4306 16833
rect 4250 16759 4306 16768
rect 4080 16510 4200 16538
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 4080 15638 4108 16390
rect 4068 15632 4120 15638
rect 4068 15574 4120 15580
rect 3988 15456 4108 15484
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 3988 13462 4016 14350
rect 3976 13456 4028 13462
rect 3976 13398 4028 13404
rect 3988 12986 4016 13398
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 3896 12838 4016 12866
rect 3884 12776 3936 12782
rect 3884 12718 3936 12724
rect 3896 12306 3924 12718
rect 3884 12300 3936 12306
rect 3884 12242 3936 12248
rect 3790 12200 3846 12209
rect 3790 12135 3846 12144
rect 3700 11212 3752 11218
rect 3700 11154 3752 11160
rect 3700 11076 3752 11082
rect 3700 11018 3752 11024
rect 3712 10606 3740 11018
rect 3700 10600 3752 10606
rect 3700 10542 3752 10548
rect 3608 10532 3660 10538
rect 3608 10474 3660 10480
rect 3516 10192 3568 10198
rect 3516 10134 3568 10140
rect 3516 9920 3568 9926
rect 3516 9862 3568 9868
rect 3528 8430 3556 9862
rect 3620 9382 3648 10474
rect 3698 10432 3754 10441
rect 3698 10367 3754 10376
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3620 8906 3648 9318
rect 3608 8900 3660 8906
rect 3608 8842 3660 8848
rect 3516 8424 3568 8430
rect 3516 8366 3568 8372
rect 3620 8090 3648 8842
rect 3712 8537 3740 10367
rect 3698 8528 3754 8537
rect 3698 8463 3754 8472
rect 3700 8288 3752 8294
rect 3700 8230 3752 8236
rect 3608 8084 3660 8090
rect 3608 8026 3660 8032
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 3344 7126 3464 7154
rect 3344 5098 3372 7126
rect 3620 6866 3648 7278
rect 3608 6860 3660 6866
rect 3608 6802 3660 6808
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3436 5370 3464 6598
rect 3620 6458 3648 6802
rect 3608 6452 3660 6458
rect 3608 6394 3660 6400
rect 3620 5846 3648 6394
rect 3608 5840 3660 5846
rect 3608 5782 3660 5788
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 3332 5092 3384 5098
rect 3332 5034 3384 5040
rect 3240 4820 3292 4826
rect 3240 4762 3292 4768
rect 3344 4758 3372 5034
rect 3332 4752 3384 4758
rect 3332 4694 3384 4700
rect 3332 4548 3384 4554
rect 3332 4490 3384 4496
rect 3344 2650 3372 4490
rect 3712 4049 3740 8230
rect 3804 5166 3832 12135
rect 3884 11620 3936 11626
rect 3884 11562 3936 11568
rect 3896 11354 3924 11562
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 3896 11150 3924 11290
rect 3884 11144 3936 11150
rect 3884 11086 3936 11092
rect 3988 10554 4016 12838
rect 4080 10713 4108 15456
rect 4172 12442 4200 16510
rect 4264 14074 4292 16759
rect 4252 14068 4304 14074
rect 4252 14010 4304 14016
rect 4356 13297 4384 16934
rect 4434 16824 4490 16833
rect 4434 16759 4490 16768
rect 4342 13288 4398 13297
rect 4342 13223 4398 13232
rect 4448 12764 4476 16759
rect 4540 15858 4568 17836
rect 4632 17270 4660 23462
rect 5448 23462 5500 23468
rect 5354 23423 5410 23432
rect 4896 23180 4948 23186
rect 4896 23122 4948 23128
rect 4804 22976 4856 22982
rect 4804 22918 4856 22924
rect 4712 21548 4764 21554
rect 4712 21490 4764 21496
rect 4724 20602 4752 21490
rect 4816 21185 4844 22918
rect 4908 21962 4936 23122
rect 4986 22808 5042 22817
rect 4986 22743 4988 22752
rect 5040 22743 5042 22752
rect 4988 22714 5040 22720
rect 5000 22506 5028 22714
rect 4988 22500 5040 22506
rect 4988 22442 5040 22448
rect 5080 22432 5132 22438
rect 5080 22374 5132 22380
rect 5092 22234 5120 22374
rect 5080 22228 5132 22234
rect 5080 22170 5132 22176
rect 4988 22092 5040 22098
rect 4988 22034 5040 22040
rect 4896 21956 4948 21962
rect 4896 21898 4948 21904
rect 5000 21486 5028 22034
rect 4988 21480 5040 21486
rect 4988 21422 5040 21428
rect 4802 21176 4858 21185
rect 4802 21111 4858 21120
rect 4712 20596 4764 20602
rect 4712 20538 4764 20544
rect 4816 20330 4844 21111
rect 4896 21004 4948 21010
rect 4896 20946 4948 20952
rect 4804 20324 4856 20330
rect 4804 20266 4856 20272
rect 4908 19836 4936 20946
rect 5000 20913 5028 21422
rect 4986 20904 5042 20913
rect 4986 20839 5042 20848
rect 5092 20466 5120 22170
rect 5172 22024 5224 22030
rect 5172 21966 5224 21972
rect 5184 21690 5212 21966
rect 5172 21684 5224 21690
rect 5172 21626 5224 21632
rect 5172 21548 5224 21554
rect 5172 21490 5224 21496
rect 5184 21078 5212 21490
rect 5172 21072 5224 21078
rect 5172 21014 5224 21020
rect 5080 20460 5132 20466
rect 5080 20402 5132 20408
rect 5184 20262 5212 21014
rect 5172 20256 5224 20262
rect 5172 20198 5224 20204
rect 5080 19848 5132 19854
rect 4908 19808 5080 19836
rect 5080 19790 5132 19796
rect 5092 19553 5120 19790
rect 5078 19544 5134 19553
rect 5078 19479 5134 19488
rect 4896 19168 4948 19174
rect 4896 19110 4948 19116
rect 4712 18828 4764 18834
rect 4712 18770 4764 18776
rect 4804 18828 4856 18834
rect 4804 18770 4856 18776
rect 4724 18222 4752 18770
rect 4712 18216 4764 18222
rect 4710 18184 4712 18193
rect 4764 18184 4766 18193
rect 4710 18119 4766 18128
rect 4816 18086 4844 18770
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 4620 17264 4672 17270
rect 4620 17206 4672 17212
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4724 16658 4752 16934
rect 4712 16652 4764 16658
rect 4712 16594 4764 16600
rect 4620 16584 4672 16590
rect 4620 16526 4672 16532
rect 4632 16046 4660 16526
rect 4712 16176 4764 16182
rect 4712 16118 4764 16124
rect 4620 16040 4672 16046
rect 4724 16017 4752 16118
rect 4620 15982 4672 15988
rect 4710 16008 4766 16017
rect 4710 15943 4766 15952
rect 4540 15830 4660 15858
rect 4448 12736 4568 12764
rect 4436 12640 4488 12646
rect 4250 12608 4306 12617
rect 4436 12582 4488 12588
rect 4250 12543 4306 12552
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 4264 12306 4292 12543
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 4160 11688 4212 11694
rect 4160 11630 4212 11636
rect 4172 11218 4200 11630
rect 4264 11558 4292 12242
rect 4252 11552 4304 11558
rect 4304 11512 4384 11540
rect 4252 11494 4304 11500
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 4172 11064 4200 11154
rect 4172 11036 4292 11064
rect 4066 10704 4122 10713
rect 4066 10639 4122 10648
rect 3988 10526 4108 10554
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3988 10062 4016 10406
rect 4080 10248 4108 10526
rect 4080 10220 4200 10248
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 3976 10056 4028 10062
rect 3882 10024 3938 10033
rect 3976 9998 4028 10004
rect 3882 9959 3884 9968
rect 3936 9959 3938 9968
rect 3884 9930 3936 9936
rect 3896 9178 3924 9930
rect 3884 9172 3936 9178
rect 3884 9114 3936 9120
rect 3988 9042 4016 9998
rect 4080 9178 4108 10066
rect 4172 9178 4200 10220
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 3974 8664 4030 8673
rect 3974 8599 4030 8608
rect 3988 8498 4016 8599
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 3988 7857 4016 8434
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 3974 7848 4030 7857
rect 3974 7783 4030 7792
rect 3974 7168 4030 7177
rect 3974 7103 4030 7112
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3896 6361 3924 6598
rect 3882 6352 3938 6361
rect 3882 6287 3938 6296
rect 3988 5710 4016 7103
rect 4080 6458 4108 8366
rect 4172 8362 4200 8910
rect 4264 8838 4292 11036
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4160 8356 4212 8362
rect 4160 8298 4212 8304
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 4172 5794 4200 8298
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4264 6662 4292 7142
rect 4252 6656 4304 6662
rect 4252 6598 4304 6604
rect 4264 5914 4292 6598
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 4172 5766 4292 5794
rect 4356 5778 4384 11512
rect 4448 10606 4476 12582
rect 4540 10985 4568 12736
rect 4526 10976 4582 10985
rect 4526 10911 4582 10920
rect 4632 10826 4660 15830
rect 4710 15736 4766 15745
rect 4908 15722 4936 19110
rect 4988 18284 5040 18290
rect 4988 18226 5040 18232
rect 5000 16153 5028 18226
rect 5092 17542 5120 19479
rect 5368 19242 5396 23423
rect 5552 23254 5580 23598
rect 5906 23352 5962 23361
rect 5906 23287 5908 23296
rect 5960 23287 5962 23296
rect 5908 23258 5960 23264
rect 5540 23248 5592 23254
rect 5540 23190 5592 23196
rect 5540 23044 5592 23050
rect 5540 22986 5592 22992
rect 5552 22642 5580 22986
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5540 22636 5592 22642
rect 5540 22578 5592 22584
rect 5538 22400 5594 22409
rect 5538 22335 5594 22344
rect 5448 22024 5500 22030
rect 5448 21966 5500 21972
rect 5460 21350 5488 21966
rect 5448 21344 5500 21350
rect 5448 21286 5500 21292
rect 5460 20806 5488 21286
rect 5448 20800 5500 20806
rect 5448 20742 5500 20748
rect 5448 20256 5500 20262
rect 5448 20198 5500 20204
rect 5460 19718 5488 20198
rect 5448 19712 5500 19718
rect 5446 19680 5448 19689
rect 5500 19680 5502 19689
rect 5446 19615 5502 19624
rect 5356 19236 5408 19242
rect 5356 19178 5408 19184
rect 5172 19168 5224 19174
rect 5172 19110 5224 19116
rect 5184 18737 5212 19110
rect 5552 18902 5580 22335
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5816 19372 5868 19378
rect 5816 19314 5868 19320
rect 5828 19174 5856 19314
rect 5816 19168 5868 19174
rect 5816 19110 5868 19116
rect 5540 18896 5592 18902
rect 5540 18838 5592 18844
rect 5828 18766 5856 19110
rect 5356 18760 5408 18766
rect 5170 18728 5226 18737
rect 5356 18702 5408 18708
rect 5816 18760 5868 18766
rect 5816 18702 5868 18708
rect 5170 18663 5226 18672
rect 5264 18624 5316 18630
rect 5264 18566 5316 18572
rect 5276 18329 5304 18566
rect 5262 18320 5318 18329
rect 5368 18290 5396 18702
rect 5448 18692 5500 18698
rect 5448 18634 5500 18640
rect 5262 18255 5318 18264
rect 5356 18284 5408 18290
rect 5356 18226 5408 18232
rect 5172 18080 5224 18086
rect 5172 18022 5224 18028
rect 5184 17785 5212 18022
rect 5460 17882 5488 18634
rect 5540 18624 5592 18630
rect 5540 18566 5592 18572
rect 5448 17876 5500 17882
rect 5448 17818 5500 17824
rect 5170 17776 5226 17785
rect 5170 17711 5226 17720
rect 5080 17536 5132 17542
rect 5080 17478 5132 17484
rect 5092 17202 5120 17478
rect 5080 17196 5132 17202
rect 5080 17138 5132 17144
rect 5264 17196 5316 17202
rect 5264 17138 5316 17144
rect 4986 16144 5042 16153
rect 4986 16079 5042 16088
rect 4710 15671 4766 15680
rect 4816 15694 4936 15722
rect 4724 15434 4752 15671
rect 4712 15428 4764 15434
rect 4712 15370 4764 15376
rect 4712 14816 4764 14822
rect 4712 14758 4764 14764
rect 4724 14482 4752 14758
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 4724 14006 4752 14418
rect 4712 14000 4764 14006
rect 4710 13968 4712 13977
rect 4764 13968 4766 13977
rect 4710 13903 4766 13912
rect 4712 13864 4764 13870
rect 4712 13806 4764 13812
rect 4724 13326 4752 13806
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4724 12646 4752 13262
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4816 11937 4844 15694
rect 4896 15632 4948 15638
rect 4896 15574 4948 15580
rect 4908 14550 4936 15574
rect 4896 14544 4948 14550
rect 4896 14486 4948 14492
rect 5000 13954 5028 16079
rect 5092 16046 5120 17138
rect 5276 16522 5304 17138
rect 5448 16720 5500 16726
rect 5448 16662 5500 16668
rect 5356 16652 5408 16658
rect 5356 16594 5408 16600
rect 5264 16516 5316 16522
rect 5264 16458 5316 16464
rect 5276 16250 5304 16458
rect 5264 16244 5316 16250
rect 5264 16186 5316 16192
rect 5080 16040 5132 16046
rect 5080 15982 5132 15988
rect 5080 15904 5132 15910
rect 5264 15904 5316 15910
rect 5080 15846 5132 15852
rect 5170 15872 5226 15881
rect 5092 15706 5120 15846
rect 5264 15846 5316 15852
rect 5170 15807 5226 15816
rect 5080 15700 5132 15706
rect 5080 15642 5132 15648
rect 5184 15570 5212 15807
rect 5276 15638 5304 15846
rect 5264 15632 5316 15638
rect 5264 15574 5316 15580
rect 5172 15564 5224 15570
rect 5172 15506 5224 15512
rect 5080 14816 5132 14822
rect 5078 14784 5080 14793
rect 5132 14784 5134 14793
rect 5078 14719 5134 14728
rect 5184 14074 5212 15506
rect 5264 15496 5316 15502
rect 5264 15438 5316 15444
rect 5276 15162 5304 15438
rect 5264 15156 5316 15162
rect 5264 15098 5316 15104
rect 5276 15065 5304 15098
rect 5262 15056 5318 15065
rect 5262 14991 5318 15000
rect 5368 14618 5396 16594
rect 5460 16046 5488 16662
rect 5448 16040 5500 16046
rect 5448 15982 5500 15988
rect 5448 15700 5500 15706
rect 5552 15688 5580 18566
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5816 18284 5868 18290
rect 5816 18226 5868 18232
rect 5828 17814 5856 18226
rect 5816 17808 5868 17814
rect 5816 17750 5868 17756
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5724 16176 5776 16182
rect 5724 16118 5776 16124
rect 5736 15706 5764 16118
rect 5500 15660 5580 15688
rect 5448 15642 5500 15648
rect 5446 15600 5502 15609
rect 5446 15535 5502 15544
rect 5460 15337 5488 15535
rect 5446 15328 5502 15337
rect 5446 15263 5502 15272
rect 5356 14612 5408 14618
rect 5356 14554 5408 14560
rect 5448 14544 5500 14550
rect 5448 14486 5500 14492
rect 5356 14272 5408 14278
rect 5356 14214 5408 14220
rect 5262 14104 5318 14113
rect 5172 14068 5224 14074
rect 5262 14039 5318 14048
rect 5172 14010 5224 14016
rect 5000 13926 5212 13954
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 4802 11928 4858 11937
rect 4802 11863 4858 11872
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4540 10798 4660 10826
rect 4436 10600 4488 10606
rect 4436 10542 4488 10548
rect 4436 10192 4488 10198
rect 4436 10134 4488 10140
rect 4448 9722 4476 10134
rect 4436 9716 4488 9722
rect 4436 9658 4488 9664
rect 4434 8392 4490 8401
rect 4434 8327 4436 8336
rect 4488 8327 4490 8336
rect 4436 8298 4488 8304
rect 4448 8090 4476 8298
rect 4436 8084 4488 8090
rect 4436 8026 4488 8032
rect 4540 7954 4568 10798
rect 4724 10538 4752 11154
rect 4908 10577 4936 12922
rect 4988 12708 5040 12714
rect 4988 12650 5040 12656
rect 5000 12102 5028 12650
rect 5078 12608 5134 12617
rect 5078 12543 5134 12552
rect 4988 12096 5040 12102
rect 4988 12038 5040 12044
rect 4894 10568 4950 10577
rect 4712 10532 4764 10538
rect 4894 10503 4950 10512
rect 4712 10474 4764 10480
rect 4724 10062 4752 10474
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 4632 9586 4660 9862
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4632 8974 4660 9522
rect 4816 9382 4844 10066
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 4632 8294 4660 8774
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4528 7948 4580 7954
rect 4528 7890 4580 7896
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4448 7410 4476 7686
rect 4436 7404 4488 7410
rect 4436 7346 4488 7352
rect 4448 7002 4476 7346
rect 4436 6996 4488 7002
rect 4436 6938 4488 6944
rect 4632 6798 4660 8230
rect 4724 8022 4752 9114
rect 4712 8016 4764 8022
rect 4712 7958 4764 7964
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4436 6384 4488 6390
rect 4436 6326 4488 6332
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 4080 5234 4108 5646
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 4080 4690 4108 5170
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 3698 4040 3754 4049
rect 3698 3975 3754 3984
rect 3424 3120 3476 3126
rect 3424 3062 3476 3068
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 3436 480 3464 3062
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 3528 2650 3556 2994
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 3528 2446 3556 2586
rect 3516 2440 3568 2446
rect 3516 2382 3568 2388
rect 3712 2009 3740 3975
rect 3988 3602 4016 4082
rect 4160 3664 4212 3670
rect 4160 3606 4212 3612
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3698 2000 3754 2009
rect 3698 1935 3754 1944
rect 3896 626 3924 3334
rect 4172 3058 4200 3606
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 4264 2990 4292 5766
rect 4344 5772 4396 5778
rect 4344 5714 4396 5720
rect 4356 5370 4384 5714
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 4448 4826 4476 6326
rect 4710 6216 4766 6225
rect 4710 6151 4766 6160
rect 4724 5914 4752 6151
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4724 5370 4752 5850
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4618 5264 4674 5273
rect 4618 5199 4674 5208
rect 4436 4820 4488 4826
rect 4356 4780 4436 4808
rect 4356 3194 4384 4780
rect 4436 4762 4488 4768
rect 4528 4616 4580 4622
rect 4528 4558 4580 4564
rect 4540 4457 4568 4558
rect 4526 4448 4582 4457
rect 4448 4406 4526 4434
rect 4344 3188 4396 3194
rect 4344 3130 4396 3136
rect 4252 2984 4304 2990
rect 3974 2952 4030 2961
rect 4252 2926 4304 2932
rect 3974 2887 3976 2896
rect 4028 2887 4030 2896
rect 3976 2858 4028 2864
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 4264 2281 4292 2790
rect 4448 2417 4476 4406
rect 4526 4383 4582 4392
rect 4632 2802 4660 5199
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4724 4078 4752 4558
rect 4712 4072 4764 4078
rect 4712 4014 4764 4020
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4540 2774 4660 2802
rect 4434 2408 4490 2417
rect 4434 2343 4490 2352
rect 4250 2272 4306 2281
rect 4250 2207 4306 2216
rect 3896 598 4016 626
rect 3988 480 4016 598
rect 4540 480 4568 2774
rect 4724 2582 4752 3538
rect 4816 3505 4844 9318
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 4908 6866 4936 8570
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 4908 6254 4936 6802
rect 4896 6248 4948 6254
rect 4896 6190 4948 6196
rect 5000 5409 5028 12038
rect 5092 9042 5120 12543
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 5080 7812 5132 7818
rect 5080 7754 5132 7760
rect 5092 7274 5120 7754
rect 5080 7268 5132 7274
rect 5080 7210 5132 7216
rect 5092 5914 5120 7210
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 5092 5710 5120 5850
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 4986 5400 5042 5409
rect 5092 5370 5120 5646
rect 4986 5335 5042 5344
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 5184 5234 5212 13926
rect 5276 10810 5304 14039
rect 5368 13394 5396 14214
rect 5460 13394 5488 14486
rect 5552 14346 5580 15660
rect 5724 15700 5776 15706
rect 5724 15642 5776 15648
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5540 14340 5592 14346
rect 5540 14282 5592 14288
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5722 13696 5778 13705
rect 5552 13530 5580 13670
rect 5722 13631 5778 13640
rect 5736 13530 5764 13631
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5552 13433 5580 13466
rect 5538 13424 5594 13433
rect 5356 13388 5408 13394
rect 5356 13330 5408 13336
rect 5448 13388 5500 13394
rect 5538 13359 5594 13368
rect 5448 13330 5500 13336
rect 5356 12844 5408 12850
rect 5356 12786 5408 12792
rect 5368 12102 5396 12786
rect 5460 12306 5488 13330
rect 5920 13297 5948 13806
rect 5906 13288 5962 13297
rect 5906 13223 5962 13232
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 6012 12968 6040 24806
rect 6380 24410 6408 25842
rect 6458 24440 6514 24449
rect 6368 24404 6420 24410
rect 6458 24375 6514 24384
rect 6368 24346 6420 24352
rect 6184 24268 6236 24274
rect 6184 24210 6236 24216
rect 6092 23724 6144 23730
rect 6092 23666 6144 23672
rect 6104 22710 6132 23666
rect 6196 23662 6224 24210
rect 6276 24064 6328 24070
rect 6276 24006 6328 24012
rect 6184 23656 6236 23662
rect 6184 23598 6236 23604
rect 6184 23248 6236 23254
rect 6184 23190 6236 23196
rect 6092 22704 6144 22710
rect 6196 22681 6224 23190
rect 6288 22982 6316 24006
rect 6368 23520 6420 23526
rect 6368 23462 6420 23468
rect 6276 22976 6328 22982
rect 6276 22918 6328 22924
rect 6092 22646 6144 22652
rect 6182 22672 6238 22681
rect 6182 22607 6184 22616
rect 6236 22607 6238 22616
rect 6184 22578 6236 22584
rect 6288 22522 6316 22918
rect 6104 22494 6316 22522
rect 6104 21554 6132 22494
rect 6184 22432 6236 22438
rect 6184 22374 6236 22380
rect 6092 21548 6144 21554
rect 6092 21490 6144 21496
rect 6092 20052 6144 20058
rect 6092 19994 6144 20000
rect 6104 18154 6132 19994
rect 6092 18148 6144 18154
rect 6092 18090 6144 18096
rect 6092 17672 6144 17678
rect 6092 17614 6144 17620
rect 6104 17202 6132 17614
rect 6092 17196 6144 17202
rect 6092 17138 6144 17144
rect 6092 16788 6144 16794
rect 6092 16730 6144 16736
rect 6104 15706 6132 16730
rect 6092 15700 6144 15706
rect 6092 15642 6144 15648
rect 6092 15564 6144 15570
rect 6092 15506 6144 15512
rect 6104 13802 6132 15506
rect 6092 13796 6144 13802
rect 6092 13738 6144 13744
rect 5920 12940 6040 12968
rect 5540 12368 5592 12374
rect 5540 12310 5592 12316
rect 5448 12300 5500 12306
rect 5448 12242 5500 12248
rect 5356 12096 5408 12102
rect 5356 12038 5408 12044
rect 5368 11286 5396 12038
rect 5552 11898 5580 12310
rect 5920 12209 5948 12940
rect 6196 12866 6224 22374
rect 6380 21593 6408 23462
rect 6366 21584 6422 21593
rect 6366 21519 6422 21528
rect 6276 20256 6328 20262
rect 6276 20198 6328 20204
rect 6288 18834 6316 20198
rect 6368 19712 6420 19718
rect 6368 19654 6420 19660
rect 6380 19242 6408 19654
rect 6368 19236 6420 19242
rect 6368 19178 6420 19184
rect 6276 18828 6328 18834
rect 6276 18770 6328 18776
rect 6288 17490 6316 18770
rect 6380 18222 6408 19178
rect 6368 18216 6420 18222
rect 6368 18158 6420 18164
rect 6472 17796 6500 24375
rect 6656 23769 6684 27520
rect 7104 25220 7156 25226
rect 7104 25162 7156 25168
rect 6734 25120 6790 25129
rect 6734 25055 6790 25064
rect 6642 23760 6698 23769
rect 6642 23695 6698 23704
rect 6552 23316 6604 23322
rect 6552 23258 6604 23264
rect 6564 22817 6592 23258
rect 6748 23202 6776 25055
rect 7116 24954 7144 25162
rect 7104 24948 7156 24954
rect 7104 24890 7156 24896
rect 7116 24342 7144 24890
rect 7104 24336 7156 24342
rect 7104 24278 7156 24284
rect 7196 24064 7248 24070
rect 7196 24006 7248 24012
rect 7208 23905 7236 24006
rect 7194 23896 7250 23905
rect 7194 23831 7250 23840
rect 7208 23662 7236 23831
rect 7196 23656 7248 23662
rect 7196 23598 7248 23604
rect 7300 23361 7328 27520
rect 7852 26194 7880 27520
rect 8300 26240 8352 26246
rect 7748 26172 7800 26178
rect 7852 26166 7972 26194
rect 8300 26182 8352 26188
rect 7748 26114 7800 26120
rect 7654 25936 7710 25945
rect 7654 25871 7710 25880
rect 7472 25764 7524 25770
rect 7472 25706 7524 25712
rect 7380 25152 7432 25158
rect 7380 25094 7432 25100
rect 7392 24274 7420 25094
rect 7380 24268 7432 24274
rect 7380 24210 7432 24216
rect 7392 23866 7420 24210
rect 7380 23860 7432 23866
rect 7380 23802 7432 23808
rect 7484 23798 7512 25706
rect 7668 24954 7696 25871
rect 7656 24948 7708 24954
rect 7656 24890 7708 24896
rect 7564 24744 7616 24750
rect 7564 24686 7616 24692
rect 7472 23792 7524 23798
rect 7472 23734 7524 23740
rect 7286 23352 7342 23361
rect 7286 23287 7342 23296
rect 6656 23174 6776 23202
rect 7104 23180 7156 23186
rect 6550 22808 6606 22817
rect 6550 22743 6552 22752
rect 6604 22743 6606 22752
rect 6552 22714 6604 22720
rect 6564 22683 6592 22714
rect 6552 22568 6604 22574
rect 6552 22510 6604 22516
rect 6564 21690 6592 22510
rect 6656 22438 6684 23174
rect 7104 23122 7156 23128
rect 7012 23112 7064 23118
rect 7012 23054 7064 23060
rect 6736 23044 6788 23050
rect 6736 22986 6788 22992
rect 6644 22432 6696 22438
rect 6644 22374 6696 22380
rect 6644 21956 6696 21962
rect 6644 21898 6696 21904
rect 6552 21684 6604 21690
rect 6552 21626 6604 21632
rect 6564 20534 6592 21626
rect 6656 21554 6684 21898
rect 6644 21548 6696 21554
rect 6644 21490 6696 21496
rect 6552 20528 6604 20534
rect 6552 20470 6604 20476
rect 6550 20360 6606 20369
rect 6550 20295 6552 20304
rect 6604 20295 6606 20304
rect 6552 20266 6604 20272
rect 6656 19854 6684 21490
rect 6748 20058 6776 22986
rect 6920 21888 6972 21894
rect 7024 21876 7052 23054
rect 7116 22506 7144 23122
rect 7194 23080 7250 23089
rect 7194 23015 7250 23024
rect 7208 22681 7236 23015
rect 7472 22976 7524 22982
rect 7472 22918 7524 22924
rect 7194 22672 7250 22681
rect 7194 22607 7250 22616
rect 7288 22636 7340 22642
rect 7104 22500 7156 22506
rect 7104 22442 7156 22448
rect 7208 22166 7236 22607
rect 7288 22578 7340 22584
rect 7300 22234 7328 22578
rect 7484 22574 7512 22918
rect 7472 22568 7524 22574
rect 7472 22510 7524 22516
rect 7380 22432 7432 22438
rect 7380 22374 7432 22380
rect 7392 22273 7420 22374
rect 7378 22264 7434 22273
rect 7288 22228 7340 22234
rect 7378 22199 7434 22208
rect 7288 22170 7340 22176
rect 7196 22160 7248 22166
rect 7196 22102 7248 22108
rect 7288 22092 7340 22098
rect 7288 22034 7340 22040
rect 7300 22001 7328 22034
rect 7286 21992 7342 22001
rect 7286 21927 7342 21936
rect 6972 21848 7052 21876
rect 6920 21830 6972 21836
rect 6932 21486 6960 21830
rect 6920 21480 6972 21486
rect 6920 21422 6972 21428
rect 6932 21146 6960 21422
rect 7300 21418 7328 21927
rect 7484 21457 7512 22510
rect 7470 21448 7526 21457
rect 7288 21412 7340 21418
rect 7470 21383 7526 21392
rect 7288 21354 7340 21360
rect 6920 21140 6972 21146
rect 6920 21082 6972 21088
rect 6828 20800 6880 20806
rect 6828 20742 6880 20748
rect 6736 20052 6788 20058
rect 6736 19994 6788 20000
rect 6840 19904 6868 20742
rect 7012 20528 7064 20534
rect 7010 20496 7012 20505
rect 7064 20496 7066 20505
rect 7010 20431 7066 20440
rect 7104 20392 7156 20398
rect 7104 20334 7156 20340
rect 6920 19916 6972 19922
rect 6840 19876 6920 19904
rect 6644 19848 6696 19854
rect 6644 19790 6696 19796
rect 6656 19553 6684 19790
rect 6642 19544 6698 19553
rect 6642 19479 6698 19488
rect 6644 19304 6696 19310
rect 6550 19272 6606 19281
rect 6644 19246 6696 19252
rect 6550 19207 6606 19216
rect 6564 19174 6592 19207
rect 6552 19168 6604 19174
rect 6552 19110 6604 19116
rect 6472 17768 6592 17796
rect 6288 17462 6500 17490
rect 6276 17196 6328 17202
rect 6276 17138 6328 17144
rect 6288 16590 6316 17138
rect 6366 16960 6422 16969
rect 6366 16895 6422 16904
rect 6276 16584 6328 16590
rect 6276 16526 6328 16532
rect 6276 16448 6328 16454
rect 6276 16390 6328 16396
rect 6288 16182 6316 16390
rect 6276 16176 6328 16182
rect 6276 16118 6328 16124
rect 6276 15632 6328 15638
rect 6276 15574 6328 15580
rect 6288 14822 6316 15574
rect 6380 15570 6408 16895
rect 6368 15564 6420 15570
rect 6368 15506 6420 15512
rect 6276 14816 6328 14822
rect 6276 14758 6328 14764
rect 6368 14816 6420 14822
rect 6368 14758 6420 14764
rect 6288 14414 6316 14758
rect 6276 14408 6328 14414
rect 6276 14350 6328 14356
rect 6288 13938 6316 14350
rect 6380 14278 6408 14758
rect 6368 14272 6420 14278
rect 6368 14214 6420 14220
rect 6276 13932 6328 13938
rect 6276 13874 6328 13880
rect 6380 13870 6408 14214
rect 6368 13864 6420 13870
rect 6368 13806 6420 13812
rect 6276 13796 6328 13802
rect 6276 13738 6328 13744
rect 6012 12838 6224 12866
rect 5906 12200 5962 12209
rect 5906 12135 5962 12144
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5448 11620 5500 11626
rect 5448 11562 5500 11568
rect 5356 11280 5408 11286
rect 5356 11222 5408 11228
rect 5460 11082 5488 11562
rect 5552 11354 5580 11834
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 5538 11248 5594 11257
rect 5538 11183 5594 11192
rect 5448 11076 5500 11082
rect 5448 11018 5500 11024
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5552 9466 5580 11183
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5724 10736 5776 10742
rect 5722 10704 5724 10713
rect 5776 10704 5778 10713
rect 5722 10639 5778 10648
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5632 9512 5684 9518
rect 5460 9438 5580 9466
rect 5630 9480 5632 9489
rect 5684 9480 5686 9489
rect 5460 8090 5488 9438
rect 5630 9415 5686 9424
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5552 8537 5580 9318
rect 5644 9178 5672 9415
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 5630 8936 5686 8945
rect 5630 8871 5632 8880
rect 5684 8871 5686 8880
rect 5632 8842 5684 8848
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5538 8528 5594 8537
rect 5538 8463 5594 8472
rect 5814 8120 5870 8129
rect 5448 8084 5500 8090
rect 5448 8026 5500 8032
rect 5540 8084 5592 8090
rect 5814 8055 5816 8064
rect 5540 8026 5592 8032
rect 5868 8055 5870 8064
rect 5816 8026 5868 8032
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 5276 7206 5304 7890
rect 5356 7880 5408 7886
rect 5354 7848 5356 7857
rect 5408 7848 5410 7857
rect 5354 7783 5410 7792
rect 5460 7546 5488 8026
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5552 7342 5580 8026
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 5276 6497 5304 7142
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5552 6746 5580 6802
rect 5460 6718 5580 6746
rect 5262 6488 5318 6497
rect 5262 6423 5318 6432
rect 5262 6352 5318 6361
rect 5262 6287 5318 6296
rect 5276 6254 5304 6287
rect 5264 6248 5316 6254
rect 5264 6190 5316 6196
rect 5356 6112 5408 6118
rect 5356 6054 5408 6060
rect 5368 5642 5396 6054
rect 5356 5636 5408 5642
rect 5356 5578 5408 5584
rect 5368 5370 5396 5578
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 5460 5114 5488 6718
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5552 6254 5580 6598
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 5540 5840 5592 5846
rect 5540 5782 5592 5788
rect 5184 5086 5488 5114
rect 4802 3496 4858 3505
rect 4802 3431 4858 3440
rect 5184 3194 5212 5086
rect 5552 4826 5580 5782
rect 5814 5672 5870 5681
rect 5814 5607 5816 5616
rect 5868 5607 5870 5616
rect 5816 5578 5868 5584
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5816 5160 5868 5166
rect 5814 5128 5816 5137
rect 5868 5128 5870 5137
rect 5814 5063 5870 5072
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5828 4758 5856 5063
rect 6012 4758 6040 12838
rect 6090 12744 6146 12753
rect 6090 12679 6146 12688
rect 6104 9450 6132 12679
rect 6288 12374 6316 13738
rect 6366 13560 6422 13569
rect 6366 13495 6422 13504
rect 6276 12368 6328 12374
rect 6276 12310 6328 12316
rect 6182 11928 6238 11937
rect 6182 11863 6238 11872
rect 6196 11665 6224 11863
rect 6182 11656 6238 11665
rect 6182 11591 6238 11600
rect 6184 11552 6236 11558
rect 6184 11494 6236 11500
rect 6196 9500 6224 11494
rect 6380 11354 6408 13495
rect 6368 11348 6420 11354
rect 6368 11290 6420 11296
rect 6276 11076 6328 11082
rect 6276 11018 6328 11024
rect 6288 10810 6316 11018
rect 6368 11008 6420 11014
rect 6368 10950 6420 10956
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 6276 10600 6328 10606
rect 6276 10542 6328 10548
rect 6288 10062 6316 10542
rect 6380 10266 6408 10950
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 6288 9654 6316 9998
rect 6380 9722 6408 10202
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6276 9648 6328 9654
rect 6276 9590 6328 9596
rect 6196 9472 6316 9500
rect 6092 9444 6144 9450
rect 6092 9386 6144 9392
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6196 8809 6224 8978
rect 6182 8800 6238 8809
rect 6182 8735 6238 8744
rect 6288 8650 6316 9472
rect 6368 9104 6420 9110
rect 6368 9046 6420 9052
rect 6196 8622 6316 8650
rect 6380 8634 6408 9046
rect 6368 8628 6420 8634
rect 6092 7744 6144 7750
rect 6092 7686 6144 7692
rect 6104 6905 6132 7686
rect 6090 6896 6146 6905
rect 6090 6831 6146 6840
rect 6092 6656 6144 6662
rect 6092 6598 6144 6604
rect 5816 4752 5868 4758
rect 5816 4694 5868 4700
rect 6000 4752 6052 4758
rect 6000 4694 6052 4700
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5262 4312 5318 4321
rect 5262 4247 5318 4256
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5276 2650 5304 4247
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5368 3670 5396 3878
rect 5356 3664 5408 3670
rect 5356 3606 5408 3612
rect 5460 3398 5488 4558
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 6012 4282 6040 4694
rect 6000 4276 6052 4282
rect 6000 4218 6052 4224
rect 6104 4185 6132 6598
rect 6090 4176 6146 4185
rect 6090 4111 6146 4120
rect 6104 4010 6132 4111
rect 6092 4004 6144 4010
rect 6092 3946 6144 3952
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 4712 2576 4764 2582
rect 4712 2518 4764 2524
rect 5080 2508 5132 2514
rect 5080 2450 5132 2456
rect 5092 480 5120 2450
rect 5460 1986 5488 3334
rect 5552 3194 5580 3674
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 6090 3224 6146 3233
rect 5540 3188 5592 3194
rect 6090 3159 6146 3168
rect 5540 3130 5592 3136
rect 6104 2990 6132 3159
rect 6092 2984 6144 2990
rect 6092 2926 6144 2932
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5460 1958 5672 1986
rect 5644 480 5672 1958
rect 6196 480 6224 8622
rect 6368 8570 6420 8576
rect 6472 7993 6500 17462
rect 6458 7984 6514 7993
rect 6458 7919 6514 7928
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6366 7304 6422 7313
rect 6366 7239 6422 7248
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 6288 5030 6316 7142
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6380 4808 6408 7239
rect 6472 7206 6500 7822
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6472 6769 6500 7142
rect 6458 6760 6514 6769
rect 6458 6695 6514 6704
rect 6458 6488 6514 6497
rect 6458 6423 6514 6432
rect 6472 6390 6500 6423
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6472 5302 6500 5646
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 6380 4780 6500 4808
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 6288 4146 6316 4558
rect 6276 4140 6328 4146
rect 6276 4082 6328 4088
rect 6288 3738 6316 4082
rect 6380 3942 6408 4626
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 6276 3732 6328 3738
rect 6276 3674 6328 3680
rect 6380 3369 6408 3878
rect 6366 3360 6422 3369
rect 6366 3295 6422 3304
rect 6380 3097 6408 3295
rect 6366 3088 6422 3097
rect 6366 3023 6422 3032
rect 6472 2854 6500 4780
rect 6564 3738 6592 17768
rect 6656 17746 6684 19246
rect 6840 18970 6868 19876
rect 6920 19858 6972 19864
rect 6828 18964 6880 18970
rect 7116 18952 7144 20334
rect 7484 19310 7512 21383
rect 7576 20398 7604 24686
rect 7760 24410 7788 26114
rect 7840 26036 7892 26042
rect 7840 25978 7892 25984
rect 7748 24404 7800 24410
rect 7748 24346 7800 24352
rect 7852 23882 7880 25978
rect 7668 23854 7880 23882
rect 7668 22250 7696 23854
rect 7944 23089 7972 26166
rect 8312 24410 8340 26182
rect 8404 24834 8432 27520
rect 8760 26104 8812 26110
rect 8760 26046 8812 26052
rect 8668 25356 8720 25362
rect 8668 25298 8720 25304
rect 8680 24886 8708 25298
rect 8772 24954 8800 26046
rect 8944 25968 8996 25974
rect 8944 25910 8996 25916
rect 8852 25832 8904 25838
rect 8852 25774 8904 25780
rect 8760 24948 8812 24954
rect 8760 24890 8812 24896
rect 8668 24880 8720 24886
rect 8666 24848 8668 24857
rect 8720 24848 8722 24857
rect 8404 24806 8616 24834
rect 8300 24404 8352 24410
rect 8300 24346 8352 24352
rect 8312 23662 8340 24346
rect 8484 24268 8536 24274
rect 8484 24210 8536 24216
rect 8496 23730 8524 24210
rect 8484 23724 8536 23730
rect 8484 23666 8536 23672
rect 8300 23656 8352 23662
rect 8300 23598 8352 23604
rect 8300 23520 8352 23526
rect 8300 23462 8352 23468
rect 8116 23180 8168 23186
rect 8116 23122 8168 23128
rect 8024 23112 8076 23118
rect 7930 23080 7986 23089
rect 8024 23054 8076 23060
rect 7930 23015 7986 23024
rect 7932 22636 7984 22642
rect 7932 22578 7984 22584
rect 7944 22386 7972 22578
rect 8036 22506 8064 23054
rect 8128 22778 8156 23122
rect 8312 23118 8340 23462
rect 8300 23112 8352 23118
rect 8352 23072 8432 23100
rect 8300 23054 8352 23060
rect 8300 22976 8352 22982
rect 8220 22936 8300 22964
rect 8116 22772 8168 22778
rect 8116 22714 8168 22720
rect 8024 22500 8076 22506
rect 8024 22442 8076 22448
rect 7944 22358 8064 22386
rect 7668 22222 7788 22250
rect 7656 22160 7708 22166
rect 7656 22102 7708 22108
rect 7564 20392 7616 20398
rect 7564 20334 7616 20340
rect 7564 20256 7616 20262
rect 7564 20198 7616 20204
rect 7576 20097 7604 20198
rect 7562 20088 7618 20097
rect 7562 20023 7618 20032
rect 7472 19304 7524 19310
rect 7472 19246 7524 19252
rect 7380 19236 7432 19242
rect 7380 19178 7432 19184
rect 7196 19168 7248 19174
rect 7392 19122 7420 19178
rect 7248 19116 7420 19122
rect 7196 19110 7420 19116
rect 7208 19094 7420 19110
rect 7116 18924 7236 18952
rect 6828 18906 6880 18912
rect 6920 18896 6972 18902
rect 6920 18838 6972 18844
rect 6828 18624 6880 18630
rect 6828 18566 6880 18572
rect 6736 18420 6788 18426
rect 6736 18362 6788 18368
rect 6644 17740 6696 17746
rect 6644 17682 6696 17688
rect 6644 17536 6696 17542
rect 6644 17478 6696 17484
rect 6656 16726 6684 17478
rect 6644 16720 6696 16726
rect 6644 16662 6696 16668
rect 6644 16584 6696 16590
rect 6644 16526 6696 16532
rect 6656 13297 6684 16526
rect 6748 13462 6776 18362
rect 6840 17882 6868 18566
rect 6828 17876 6880 17882
rect 6828 17818 6880 17824
rect 6828 17740 6880 17746
rect 6828 17682 6880 17688
rect 6840 16425 6868 17682
rect 6932 16590 6960 18838
rect 7104 18828 7156 18834
rect 7104 18770 7156 18776
rect 7116 18086 7144 18770
rect 7104 18080 7156 18086
rect 7104 18022 7156 18028
rect 7010 17776 7066 17785
rect 7010 17711 7012 17720
rect 7064 17711 7066 17720
rect 7012 17682 7064 17688
rect 7024 17338 7052 17682
rect 7012 17332 7064 17338
rect 7012 17274 7064 17280
rect 7116 17218 7144 18022
rect 7208 17513 7236 18924
rect 7668 18902 7696 22102
rect 7656 18896 7708 18902
rect 7656 18838 7708 18844
rect 7380 18760 7432 18766
rect 7380 18702 7432 18708
rect 7392 18426 7420 18702
rect 7380 18420 7432 18426
rect 7380 18362 7432 18368
rect 7668 18222 7696 18838
rect 7760 18834 7788 22222
rect 7932 22228 7984 22234
rect 7932 22170 7984 22176
rect 7840 20052 7892 20058
rect 7840 19994 7892 20000
rect 7748 18828 7800 18834
rect 7748 18770 7800 18776
rect 7852 18601 7880 19994
rect 7838 18592 7894 18601
rect 7838 18527 7894 18536
rect 7656 18216 7708 18222
rect 7656 18158 7708 18164
rect 7472 17672 7524 17678
rect 7472 17614 7524 17620
rect 7380 17604 7432 17610
rect 7380 17546 7432 17552
rect 7194 17504 7250 17513
rect 7194 17439 7250 17448
rect 7024 17190 7144 17218
rect 6920 16584 6972 16590
rect 6920 16526 6972 16532
rect 6920 16448 6972 16454
rect 6826 16416 6882 16425
rect 6920 16390 6972 16396
rect 6826 16351 6882 16360
rect 6826 16144 6882 16153
rect 6932 16114 6960 16390
rect 6826 16079 6882 16088
rect 6920 16108 6972 16114
rect 6840 16046 6868 16079
rect 6920 16050 6972 16056
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 6840 15337 6868 15846
rect 6826 15328 6882 15337
rect 6826 15263 6882 15272
rect 6826 15192 6882 15201
rect 6826 15127 6882 15136
rect 6840 14958 6868 15127
rect 6932 14958 6960 16050
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 6840 14385 6868 14894
rect 6932 14822 6960 14894
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 7024 14498 7052 17190
rect 7392 17134 7420 17546
rect 7380 17128 7432 17134
rect 7380 17070 7432 17076
rect 7104 16652 7156 16658
rect 7104 16594 7156 16600
rect 7116 16046 7144 16594
rect 7196 16448 7248 16454
rect 7196 16390 7248 16396
rect 7104 16040 7156 16046
rect 7104 15982 7156 15988
rect 7104 15904 7156 15910
rect 7104 15846 7156 15852
rect 7116 14618 7144 15846
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 7208 14550 7236 16390
rect 7378 16008 7434 16017
rect 7378 15943 7434 15952
rect 7288 15360 7340 15366
rect 7288 15302 7340 15308
rect 7300 15201 7328 15302
rect 7286 15192 7342 15201
rect 7286 15127 7342 15136
rect 7286 14784 7342 14793
rect 7286 14719 7342 14728
rect 7196 14544 7248 14550
rect 7024 14470 7144 14498
rect 7196 14486 7248 14492
rect 6826 14376 6882 14385
rect 6826 14311 6882 14320
rect 7012 14340 7064 14346
rect 7012 14282 7064 14288
rect 6828 14000 6880 14006
rect 6828 13942 6880 13948
rect 6920 14000 6972 14006
rect 6920 13942 6972 13948
rect 6840 13705 6868 13942
rect 6826 13696 6882 13705
rect 6826 13631 6882 13640
rect 6736 13456 6788 13462
rect 6736 13398 6788 13404
rect 6642 13288 6698 13297
rect 6642 13223 6698 13232
rect 6656 12986 6684 13223
rect 6644 12980 6696 12986
rect 6644 12922 6696 12928
rect 6748 12918 6776 13398
rect 6736 12912 6788 12918
rect 6736 12854 6788 12860
rect 6642 12744 6698 12753
rect 6642 12679 6644 12688
rect 6696 12679 6698 12688
rect 6644 12650 6696 12656
rect 6748 12442 6776 12854
rect 6736 12436 6788 12442
rect 6736 12378 6788 12384
rect 6932 12306 6960 13942
rect 6920 12300 6972 12306
rect 6920 12242 6972 12248
rect 6734 12064 6790 12073
rect 6734 11999 6790 12008
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 6656 9994 6684 11086
rect 6644 9988 6696 9994
rect 6644 9930 6696 9936
rect 6644 8356 6696 8362
rect 6644 8298 6696 8304
rect 6552 3732 6604 3738
rect 6552 3674 6604 3680
rect 6656 3670 6684 8298
rect 6644 3664 6696 3670
rect 6644 3606 6696 3612
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 6552 2304 6604 2310
rect 6550 2272 6552 2281
rect 6604 2272 6606 2281
rect 6550 2207 6606 2216
rect 6748 480 6776 11999
rect 7024 11558 7052 14282
rect 7116 12238 7144 14470
rect 7208 13530 7236 14486
rect 7300 13938 7328 14719
rect 7392 14550 7420 15943
rect 7380 14544 7432 14550
rect 7380 14486 7432 14492
rect 7288 13932 7340 13938
rect 7288 13874 7340 13880
rect 7378 13560 7434 13569
rect 7196 13524 7248 13530
rect 7484 13530 7512 17614
rect 7564 15904 7616 15910
rect 7564 15846 7616 15852
rect 7576 14890 7604 15846
rect 7668 15450 7696 18158
rect 7838 17912 7894 17921
rect 7838 17847 7894 17856
rect 7668 15422 7788 15450
rect 7656 15360 7708 15366
rect 7656 15302 7708 15308
rect 7668 15065 7696 15302
rect 7654 15056 7710 15065
rect 7654 14991 7710 15000
rect 7564 14884 7616 14890
rect 7564 14826 7616 14832
rect 7378 13495 7434 13504
rect 7472 13524 7524 13530
rect 7196 13466 7248 13472
rect 7392 12782 7420 13495
rect 7472 13466 7524 13472
rect 7576 12986 7604 14826
rect 7654 14104 7710 14113
rect 7654 14039 7710 14048
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7668 12850 7696 14039
rect 7656 12844 7708 12850
rect 7576 12804 7656 12832
rect 7380 12776 7432 12782
rect 7380 12718 7432 12724
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7116 11694 7144 12038
rect 7286 11928 7342 11937
rect 7286 11863 7342 11872
rect 7300 11762 7328 11863
rect 7288 11756 7340 11762
rect 7288 11698 7340 11704
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 6840 10690 6868 11494
rect 7012 11280 7064 11286
rect 7012 11222 7064 11228
rect 6840 10674 6960 10690
rect 6840 10668 6972 10674
rect 6840 10662 6920 10668
rect 6920 10610 6972 10616
rect 6828 10464 6880 10470
rect 6826 10432 6828 10441
rect 7024 10452 7052 11222
rect 6880 10432 7052 10452
rect 6882 10424 7052 10432
rect 6826 10367 6882 10376
rect 6826 10296 6882 10305
rect 6826 10231 6882 10240
rect 6840 8673 6868 10231
rect 7116 9722 7144 11630
rect 7194 10024 7250 10033
rect 7194 9959 7196 9968
rect 7248 9959 7250 9968
rect 7196 9930 7248 9936
rect 7288 9920 7340 9926
rect 7288 9862 7340 9868
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 7102 9072 7158 9081
rect 7102 9007 7158 9016
rect 6826 8664 6882 8673
rect 6826 8599 6882 8608
rect 7116 8430 7144 9007
rect 7300 8838 7328 9862
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 7300 8634 7328 8774
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7196 8560 7248 8566
rect 7196 8502 7248 8508
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 6840 6866 6868 7822
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6932 6866 6960 7686
rect 7012 7472 7064 7478
rect 7012 7414 7064 7420
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6932 5914 6960 6802
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 7024 5846 7052 7414
rect 7116 7274 7144 7822
rect 7104 7268 7156 7274
rect 7104 7210 7156 7216
rect 7104 6180 7156 6186
rect 7104 6122 7156 6128
rect 7012 5840 7064 5846
rect 7012 5782 7064 5788
rect 6828 5772 6880 5778
rect 6880 5732 6960 5760
rect 6828 5714 6880 5720
rect 6932 5370 6960 5732
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6840 2145 6868 4966
rect 7024 4826 7052 5510
rect 7116 5166 7144 6122
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 7024 4690 7052 4762
rect 7012 4684 7064 4690
rect 7012 4626 7064 4632
rect 7012 4004 7064 4010
rect 7012 3946 7064 3952
rect 7024 3058 7052 3946
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 7024 2514 7052 2994
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 6826 2136 6882 2145
rect 6826 2071 6882 2080
rect 7208 2009 7236 8502
rect 7300 8401 7328 8570
rect 7286 8392 7342 8401
rect 7286 8327 7342 8336
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7300 7206 7328 7890
rect 7288 7200 7340 7206
rect 7286 7168 7288 7177
rect 7340 7168 7342 7177
rect 7286 7103 7342 7112
rect 7288 5772 7340 5778
rect 7288 5714 7340 5720
rect 7300 5098 7328 5714
rect 7392 5409 7420 12718
rect 7463 12436 7515 12442
rect 7576 12424 7604 12804
rect 7656 12786 7708 12792
rect 7515 12396 7604 12424
rect 7463 12378 7515 12384
rect 7760 12322 7788 15422
rect 7852 14278 7880 17847
rect 7944 14346 7972 22170
rect 8036 20058 8064 22358
rect 8116 22024 8168 22030
rect 8116 21966 8168 21972
rect 8024 20052 8076 20058
rect 8024 19994 8076 20000
rect 8128 19378 8156 21966
rect 8220 21146 8248 22936
rect 8300 22918 8352 22924
rect 8404 22030 8432 23072
rect 8482 22944 8538 22953
rect 8482 22879 8538 22888
rect 8392 22024 8444 22030
rect 8392 21966 8444 21972
rect 8392 21888 8444 21894
rect 8392 21830 8444 21836
rect 8404 21486 8432 21830
rect 8392 21480 8444 21486
rect 8392 21422 8444 21428
rect 8208 21140 8260 21146
rect 8208 21082 8260 21088
rect 8300 21004 8352 21010
rect 8300 20946 8352 20952
rect 8312 20602 8340 20946
rect 8390 20904 8446 20913
rect 8390 20839 8446 20848
rect 8300 20596 8352 20602
rect 8300 20538 8352 20544
rect 8116 19372 8168 19378
rect 8116 19314 8168 19320
rect 8022 19272 8078 19281
rect 8022 19207 8024 19216
rect 8076 19207 8078 19216
rect 8024 19178 8076 19184
rect 8404 18970 8432 20839
rect 8496 19836 8524 22879
rect 8588 21457 8616 24806
rect 8666 24783 8722 24792
rect 8760 24744 8812 24750
rect 8760 24686 8812 24692
rect 8668 23792 8720 23798
rect 8668 23734 8720 23740
rect 8680 22234 8708 23734
rect 8668 22228 8720 22234
rect 8668 22170 8720 22176
rect 8668 22092 8720 22098
rect 8668 22034 8720 22040
rect 8680 21593 8708 22034
rect 8666 21584 8722 21593
rect 8666 21519 8722 21528
rect 8574 21448 8630 21457
rect 8680 21418 8708 21519
rect 8574 21383 8630 21392
rect 8668 21412 8720 21418
rect 8668 21354 8720 21360
rect 8496 19808 8616 19836
rect 8392 18964 8444 18970
rect 8392 18906 8444 18912
rect 8484 18828 8536 18834
rect 8484 18770 8536 18776
rect 8024 18624 8076 18630
rect 8300 18624 8352 18630
rect 8024 18566 8076 18572
rect 8128 18584 8300 18612
rect 8036 18154 8064 18566
rect 8024 18148 8076 18154
rect 8024 18090 8076 18096
rect 8036 17814 8064 18090
rect 8024 17808 8076 17814
rect 8024 17750 8076 17756
rect 8036 17377 8064 17750
rect 8128 17746 8156 18584
rect 8300 18566 8352 18572
rect 8496 18086 8524 18770
rect 8484 18080 8536 18086
rect 8484 18022 8536 18028
rect 8116 17740 8168 17746
rect 8116 17682 8168 17688
rect 8022 17368 8078 17377
rect 8022 17303 8024 17312
rect 8076 17303 8078 17312
rect 8024 17274 8076 17280
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 8036 14550 8064 16730
rect 8128 15745 8156 17682
rect 8208 17536 8260 17542
rect 8208 17478 8260 17484
rect 8220 16658 8248 17478
rect 8392 17060 8444 17066
rect 8392 17002 8444 17008
rect 8404 16833 8432 17002
rect 8390 16824 8446 16833
rect 8390 16759 8446 16768
rect 8298 16688 8354 16697
rect 8208 16652 8260 16658
rect 8298 16623 8300 16632
rect 8208 16594 8260 16600
rect 8352 16623 8354 16632
rect 8300 16594 8352 16600
rect 8220 16250 8248 16594
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 8392 16176 8444 16182
rect 8392 16118 8444 16124
rect 8114 15736 8170 15745
rect 8114 15671 8170 15680
rect 8300 15632 8352 15638
rect 8298 15600 8300 15609
rect 8352 15600 8354 15609
rect 8298 15535 8354 15544
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 8116 14816 8168 14822
rect 8116 14758 8168 14764
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8024 14544 8076 14550
rect 8024 14486 8076 14492
rect 8128 14482 8156 14758
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 7932 14340 7984 14346
rect 7932 14282 7984 14288
rect 8024 14340 8076 14346
rect 8024 14282 8076 14288
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7930 13832 7986 13841
rect 7930 13767 7986 13776
rect 7944 13326 7972 13767
rect 7932 13320 7984 13326
rect 7932 13262 7984 13268
rect 7484 12294 7788 12322
rect 7840 12300 7892 12306
rect 7484 9761 7512 12294
rect 7840 12242 7892 12248
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 7576 9874 7604 12174
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 7668 10146 7696 11494
rect 7760 11354 7788 12174
rect 7852 11558 7880 12242
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7748 11348 7800 11354
rect 7748 11290 7800 11296
rect 7852 11150 7880 11494
rect 7840 11144 7892 11150
rect 7840 11086 7892 11092
rect 7668 10118 7788 10146
rect 7656 10056 7708 10062
rect 7654 10024 7656 10033
rect 7708 10024 7710 10033
rect 7654 9959 7710 9968
rect 7576 9846 7696 9874
rect 7470 9752 7526 9761
rect 7470 9687 7526 9696
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 7564 9376 7616 9382
rect 7564 9318 7616 9324
rect 7484 7002 7512 9318
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7484 6118 7512 6734
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 7378 5400 7434 5409
rect 7378 5335 7434 5344
rect 7484 5234 7512 6054
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7378 5128 7434 5137
rect 7288 5092 7340 5098
rect 7378 5063 7434 5072
rect 7288 5034 7340 5040
rect 7300 4826 7328 5034
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 7392 4706 7420 5063
rect 7470 4992 7526 5001
rect 7470 4927 7526 4936
rect 7300 4678 7420 4706
rect 7194 2000 7250 2009
rect 7194 1935 7250 1944
rect 7300 480 7328 4678
rect 7484 4457 7512 4927
rect 7470 4448 7526 4457
rect 7470 4383 7526 4392
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 7484 3738 7512 4014
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7484 2922 7512 3334
rect 7472 2916 7524 2922
rect 7472 2858 7524 2864
rect 7470 2680 7526 2689
rect 7470 2615 7526 2624
rect 7484 2582 7512 2615
rect 7472 2576 7524 2582
rect 7472 2518 7524 2524
rect 7576 1601 7604 9318
rect 7668 8265 7696 9846
rect 7654 8256 7710 8265
rect 7654 8191 7710 8200
rect 7760 3534 7788 10118
rect 7838 9752 7894 9761
rect 7838 9687 7894 9696
rect 7852 5250 7880 9687
rect 7944 9518 7972 13262
rect 8036 12442 8064 14282
rect 8128 13852 8156 14418
rect 8220 14414 8248 14758
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 8312 14006 8340 15302
rect 8300 14000 8352 14006
rect 8300 13942 8352 13948
rect 8128 13824 8340 13852
rect 8312 13462 8340 13824
rect 8300 13456 8352 13462
rect 8300 13398 8352 13404
rect 8404 13394 8432 16118
rect 8496 15910 8524 18022
rect 8484 15904 8536 15910
rect 8484 15846 8536 15852
rect 8482 14512 8538 14521
rect 8482 14447 8538 14456
rect 8496 14074 8524 14447
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8482 13832 8538 13841
rect 8482 13767 8538 13776
rect 8392 13388 8444 13394
rect 8392 13330 8444 13336
rect 8496 13274 8524 13767
rect 8404 13258 8524 13274
rect 8392 13252 8524 13258
rect 8444 13246 8524 13252
rect 8392 13194 8444 13200
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 8114 12880 8170 12889
rect 8114 12815 8170 12824
rect 8024 12436 8076 12442
rect 8024 12378 8076 12384
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 8036 10266 8064 12038
rect 8128 11626 8156 12815
rect 8312 12782 8340 13126
rect 8300 12776 8352 12782
rect 8298 12744 8300 12753
rect 8352 12744 8354 12753
rect 8298 12679 8354 12688
rect 8206 11792 8262 11801
rect 8206 11727 8262 11736
rect 8116 11620 8168 11626
rect 8116 11562 8168 11568
rect 8220 11558 8248 11727
rect 8208 11552 8260 11558
rect 8206 11520 8208 11529
rect 8300 11552 8352 11558
rect 8260 11520 8262 11529
rect 8300 11494 8352 11500
rect 8206 11455 8262 11464
rect 8116 10804 8168 10810
rect 8312 10792 8340 11494
rect 8168 10764 8340 10792
rect 8116 10746 8168 10752
rect 8024 10260 8076 10266
rect 8024 10202 8076 10208
rect 8128 10198 8156 10746
rect 8298 10296 8354 10305
rect 8298 10231 8354 10240
rect 8116 10192 8168 10198
rect 8116 10134 8168 10140
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 8024 8288 8076 8294
rect 8024 8230 8076 8236
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 7944 7342 7972 7686
rect 8036 7410 8064 8230
rect 8116 7812 8168 7818
rect 8116 7754 8168 7760
rect 8128 7410 8156 7754
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 8116 7404 8168 7410
rect 8116 7346 8168 7352
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 8036 6934 8064 7346
rect 8024 6928 8076 6934
rect 8024 6870 8076 6876
rect 8128 6798 8156 7346
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 7932 6724 7984 6730
rect 7932 6666 7984 6672
rect 7944 5914 7972 6666
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 7932 5908 7984 5914
rect 7932 5850 7984 5856
rect 8036 5710 8064 6054
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 8036 5302 8064 5646
rect 8024 5296 8076 5302
rect 7852 5222 7972 5250
rect 8024 5238 8076 5244
rect 7840 5160 7892 5166
rect 7840 5102 7892 5108
rect 7852 3738 7880 5102
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 7760 3210 7788 3470
rect 7944 3233 7972 5222
rect 8024 5024 8076 5030
rect 8022 4992 8024 5001
rect 8076 4992 8078 5001
rect 8022 4927 8078 4936
rect 8128 4010 8156 6190
rect 8220 5370 8248 8774
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 8220 4622 8248 5170
rect 8312 5137 8340 10231
rect 8404 8090 8432 13194
rect 8482 12744 8538 12753
rect 8482 12679 8538 12688
rect 8496 12238 8524 12679
rect 8484 12232 8536 12238
rect 8484 12174 8536 12180
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 8496 11286 8524 11494
rect 8588 11354 8616 19808
rect 8680 19530 8708 21354
rect 8772 21078 8800 24686
rect 8864 24410 8892 25774
rect 8956 25498 8984 25910
rect 8944 25492 8996 25498
rect 8944 25434 8996 25440
rect 8852 24404 8904 24410
rect 8852 24346 8904 24352
rect 8944 23724 8996 23730
rect 8944 23666 8996 23672
rect 8852 22432 8904 22438
rect 8852 22374 8904 22380
rect 8864 21350 8892 22374
rect 8852 21344 8904 21350
rect 8852 21286 8904 21292
rect 8760 21072 8812 21078
rect 8760 21014 8812 21020
rect 8760 20936 8812 20942
rect 8760 20878 8812 20884
rect 8772 20058 8800 20878
rect 8864 20641 8892 21286
rect 8850 20632 8906 20641
rect 8850 20567 8906 20576
rect 8852 20324 8904 20330
rect 8852 20266 8904 20272
rect 8760 20052 8812 20058
rect 8760 19994 8812 20000
rect 8680 19502 8800 19530
rect 8666 19408 8722 19417
rect 8666 19343 8722 19352
rect 8680 19310 8708 19343
rect 8668 19304 8720 19310
rect 8668 19246 8720 19252
rect 8668 16992 8720 16998
rect 8668 16934 8720 16940
rect 8680 12617 8708 16934
rect 8772 16182 8800 19502
rect 8864 19378 8892 20266
rect 8956 19990 8984 23666
rect 9048 21593 9076 27520
rect 9600 26160 9628 27520
rect 9324 26132 9628 26160
rect 9128 25696 9180 25702
rect 9128 25638 9180 25644
rect 9140 23866 9168 25638
rect 9324 25362 9352 26132
rect 9954 26072 10010 26081
rect 9954 26007 10010 26016
rect 9312 25356 9364 25362
rect 9312 25298 9364 25304
rect 9588 25356 9640 25362
rect 9588 25298 9640 25304
rect 9312 24948 9364 24954
rect 9312 24890 9364 24896
rect 9324 23866 9352 24890
rect 9496 24812 9548 24818
rect 9496 24754 9548 24760
rect 9404 24064 9456 24070
rect 9404 24006 9456 24012
rect 9128 23860 9180 23866
rect 9128 23802 9180 23808
rect 9312 23860 9364 23866
rect 9312 23802 9364 23808
rect 9310 23760 9366 23769
rect 9416 23730 9444 24006
rect 9310 23695 9366 23704
rect 9404 23724 9456 23730
rect 9128 22976 9180 22982
rect 9128 22918 9180 22924
rect 9140 22574 9168 22918
rect 9324 22658 9352 23695
rect 9404 23666 9456 23672
rect 9416 22778 9444 23666
rect 9404 22772 9456 22778
rect 9404 22714 9456 22720
rect 9220 22636 9272 22642
rect 9324 22630 9444 22658
rect 9220 22578 9272 22584
rect 9128 22568 9180 22574
rect 9128 22510 9180 22516
rect 9128 22228 9180 22234
rect 9128 22170 9180 22176
rect 9034 21584 9090 21593
rect 9034 21519 9090 21528
rect 9036 21480 9088 21486
rect 9036 21422 9088 21428
rect 9048 20942 9076 21422
rect 9036 20936 9088 20942
rect 9034 20904 9036 20913
rect 9088 20904 9090 20913
rect 9034 20839 9090 20848
rect 9034 20360 9090 20369
rect 9034 20295 9090 20304
rect 9048 20262 9076 20295
rect 9036 20256 9088 20262
rect 9036 20198 9088 20204
rect 8944 19984 8996 19990
rect 8944 19926 8996 19932
rect 8956 19514 8984 19926
rect 8944 19508 8996 19514
rect 8944 19450 8996 19456
rect 8852 19372 8904 19378
rect 8852 19314 8904 19320
rect 8852 19168 8904 19174
rect 8852 19110 8904 19116
rect 8864 17610 8892 19110
rect 8956 18902 8984 19450
rect 9140 18952 9168 22170
rect 9232 21894 9260 22578
rect 9312 22500 9364 22506
rect 9312 22442 9364 22448
rect 9220 21888 9272 21894
rect 9220 21830 9272 21836
rect 9232 21486 9260 21830
rect 9220 21480 9272 21486
rect 9220 21422 9272 21428
rect 9220 21072 9272 21078
rect 9220 21014 9272 21020
rect 9048 18924 9168 18952
rect 8944 18896 8996 18902
rect 8944 18838 8996 18844
rect 8852 17604 8904 17610
rect 8852 17546 8904 17552
rect 8864 16250 8892 17546
rect 8944 17536 8996 17542
rect 8944 17478 8996 17484
rect 8852 16244 8904 16250
rect 8852 16186 8904 16192
rect 8760 16176 8812 16182
rect 8760 16118 8812 16124
rect 8760 16040 8812 16046
rect 8760 15982 8812 15988
rect 8772 15337 8800 15982
rect 8852 15972 8904 15978
rect 8852 15914 8904 15920
rect 8758 15328 8814 15337
rect 8758 15263 8814 15272
rect 8760 15156 8812 15162
rect 8760 15098 8812 15104
rect 8772 14414 8800 15098
rect 8760 14408 8812 14414
rect 8760 14350 8812 14356
rect 8760 14272 8812 14278
rect 8760 14214 8812 14220
rect 8772 13734 8800 14214
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 8760 13388 8812 13394
rect 8760 13330 8812 13336
rect 8666 12608 8722 12617
rect 8666 12543 8722 12552
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8484 11280 8536 11286
rect 8484 11222 8536 11228
rect 8680 11150 8708 12174
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 8496 10146 8524 11086
rect 8668 11008 8720 11014
rect 8668 10950 8720 10956
rect 8576 10532 8628 10538
rect 8576 10474 8628 10480
rect 8588 10266 8616 10474
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8496 10118 8616 10146
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 8496 9382 8524 9522
rect 8588 9382 8616 10118
rect 8680 9926 8708 10950
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8576 9376 8628 9382
rect 8576 9318 8628 9324
rect 8496 9042 8524 9318
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8496 8498 8524 8978
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8404 7546 8432 8026
rect 8496 7886 8524 8434
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8392 7268 8444 7274
rect 8496 7256 8524 7822
rect 8588 7313 8616 8910
rect 8680 8809 8708 9862
rect 8666 8800 8722 8809
rect 8666 8735 8722 8744
rect 8680 7342 8708 8735
rect 8668 7336 8720 7342
rect 8444 7228 8524 7256
rect 8574 7304 8630 7313
rect 8668 7278 8720 7284
rect 8574 7239 8630 7248
rect 8392 7210 8444 7216
rect 8404 6662 8432 7210
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8390 5672 8446 5681
rect 8390 5607 8446 5616
rect 8298 5128 8354 5137
rect 8298 5063 8354 5072
rect 8404 4758 8432 5607
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8496 5001 8524 5510
rect 8576 5296 8628 5302
rect 8576 5238 8628 5244
rect 8482 4992 8538 5001
rect 8482 4927 8538 4936
rect 8392 4752 8444 4758
rect 8392 4694 8444 4700
rect 8484 4752 8536 4758
rect 8484 4694 8536 4700
rect 8208 4616 8260 4622
rect 8260 4576 8340 4604
rect 8496 4593 8524 4694
rect 8208 4558 8260 4564
rect 8116 4004 8168 4010
rect 8116 3946 8168 3952
rect 8312 3942 8340 4576
rect 8482 4584 8538 4593
rect 8588 4554 8616 5238
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 8680 4593 8708 4966
rect 8666 4584 8722 4593
rect 8482 4519 8538 4528
rect 8576 4548 8628 4554
rect 8666 4519 8722 4528
rect 8576 4490 8628 4496
rect 8772 4162 8800 13330
rect 8864 9602 8892 15914
rect 8956 15881 8984 17478
rect 9048 16046 9076 18924
rect 9128 18828 9180 18834
rect 9128 18770 9180 18776
rect 9140 18630 9168 18770
rect 9128 18624 9180 18630
rect 9128 18566 9180 18572
rect 9140 18086 9168 18566
rect 9128 18080 9180 18086
rect 9126 18048 9128 18057
rect 9180 18048 9182 18057
rect 9126 17983 9182 17992
rect 9128 17740 9180 17746
rect 9128 17682 9180 17688
rect 9140 16998 9168 17682
rect 9232 17338 9260 21014
rect 9324 18465 9352 22442
rect 9416 21865 9444 22630
rect 9508 22234 9536 24754
rect 9496 22228 9548 22234
rect 9496 22170 9548 22176
rect 9402 21856 9458 21865
rect 9402 21791 9458 21800
rect 9600 21706 9628 25298
rect 9772 25220 9824 25226
rect 9772 25162 9824 25168
rect 9678 24440 9734 24449
rect 9678 24375 9734 24384
rect 9692 24138 9720 24375
rect 9680 24132 9732 24138
rect 9680 24074 9732 24080
rect 9784 24070 9812 25162
rect 9968 24886 9996 26007
rect 9956 24880 10008 24886
rect 10152 24834 10180 27520
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10230 25256 10286 25265
rect 10230 25191 10286 25200
rect 9956 24822 10008 24828
rect 10060 24806 10180 24834
rect 9772 24064 9824 24070
rect 9772 24006 9824 24012
rect 9680 23520 9732 23526
rect 9680 23462 9732 23468
rect 9692 23050 9720 23462
rect 9680 23044 9732 23050
rect 9680 22986 9732 22992
rect 9784 22658 9812 24006
rect 9864 23860 9916 23866
rect 9864 23802 9916 23808
rect 9876 23497 9904 23802
rect 9956 23724 10008 23730
rect 9956 23666 10008 23672
rect 9862 23488 9918 23497
rect 9862 23423 9918 23432
rect 9692 22630 9812 22658
rect 9692 22030 9720 22630
rect 9770 22536 9826 22545
rect 9770 22471 9826 22480
rect 9680 22024 9732 22030
rect 9680 21966 9732 21972
rect 9416 21678 9628 21706
rect 9692 21690 9720 21966
rect 9680 21684 9732 21690
rect 9310 18456 9366 18465
rect 9310 18391 9366 18400
rect 9310 17640 9366 17649
rect 9310 17575 9312 17584
rect 9364 17575 9366 17584
rect 9312 17546 9364 17552
rect 9220 17332 9272 17338
rect 9220 17274 9272 17280
rect 9324 17134 9352 17546
rect 9312 17128 9364 17134
rect 9218 17096 9274 17105
rect 9312 17070 9364 17076
rect 9218 17031 9274 17040
rect 9232 16998 9260 17031
rect 9128 16992 9180 16998
rect 9128 16934 9180 16940
rect 9220 16992 9272 16998
rect 9220 16934 9272 16940
rect 9310 16824 9366 16833
rect 9310 16759 9366 16768
rect 9324 16726 9352 16759
rect 9312 16720 9364 16726
rect 9312 16662 9364 16668
rect 9128 16448 9180 16454
rect 9128 16390 9180 16396
rect 9140 16266 9168 16390
rect 9218 16280 9274 16289
rect 9140 16238 9218 16266
rect 9140 16114 9168 16238
rect 9218 16215 9274 16224
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 9220 16108 9272 16114
rect 9220 16050 9272 16056
rect 9036 16040 9088 16046
rect 9036 15982 9088 15988
rect 9126 16008 9182 16017
rect 9126 15943 9182 15952
rect 9036 15904 9088 15910
rect 8942 15872 8998 15881
rect 9036 15846 9088 15852
rect 8942 15807 8998 15816
rect 8944 15700 8996 15706
rect 8944 15642 8996 15648
rect 8956 14113 8984 15642
rect 8942 14104 8998 14113
rect 8942 14039 8998 14048
rect 8942 13968 8998 13977
rect 8942 13903 8944 13912
rect 8996 13903 8998 13912
rect 8944 13874 8996 13880
rect 8956 13530 8984 13874
rect 8944 13524 8996 13530
rect 8944 13466 8996 13472
rect 9048 12617 9076 15846
rect 9140 15570 9168 15943
rect 9232 15706 9260 16050
rect 9220 15700 9272 15706
rect 9220 15642 9272 15648
rect 9128 15564 9180 15570
rect 9128 15506 9180 15512
rect 9140 15178 9168 15506
rect 9140 15150 9260 15178
rect 9128 15088 9180 15094
rect 9126 15056 9128 15065
rect 9180 15056 9182 15065
rect 9126 14991 9182 15000
rect 9232 14618 9260 15150
rect 9220 14612 9272 14618
rect 9140 14572 9220 14600
rect 9034 12608 9090 12617
rect 9034 12543 9090 12552
rect 9140 12442 9168 14572
rect 9220 14554 9272 14560
rect 9312 14476 9364 14482
rect 9312 14418 9364 14424
rect 9218 13696 9274 13705
rect 9218 13631 9274 13640
rect 9232 13530 9260 13631
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 9220 13388 9272 13394
rect 9220 13330 9272 13336
rect 9232 12782 9260 13330
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 9128 12436 9180 12442
rect 9128 12378 9180 12384
rect 9036 12368 9088 12374
rect 9036 12310 9088 12316
rect 9048 10305 9076 12310
rect 9128 12300 9180 12306
rect 9128 12242 9180 12248
rect 9140 11898 9168 12242
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 9324 11354 9352 14418
rect 9416 13802 9444 21678
rect 9680 21626 9732 21632
rect 9692 21128 9720 21626
rect 9508 21100 9720 21128
rect 9508 20788 9536 21100
rect 9692 21010 9720 21100
rect 9588 21004 9640 21010
rect 9588 20946 9640 20952
rect 9680 21004 9732 21010
rect 9680 20946 9732 20952
rect 9600 20890 9628 20946
rect 9600 20862 9720 20890
rect 9508 20760 9628 20788
rect 9494 19816 9550 19825
rect 9494 19751 9550 19760
rect 9508 16697 9536 19751
rect 9600 19394 9628 20760
rect 9692 20602 9720 20862
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 9784 19854 9812 22471
rect 9968 22001 9996 23666
rect 9954 21992 10010 22001
rect 9954 21927 10010 21936
rect 9968 21690 9996 21927
rect 9956 21684 10008 21690
rect 9956 21626 10008 21632
rect 9956 21004 10008 21010
rect 9956 20946 10008 20952
rect 9968 20466 9996 20946
rect 10060 20584 10088 24806
rect 10244 24596 10272 25191
rect 10692 24880 10744 24886
rect 10692 24822 10744 24828
rect 10152 24568 10272 24596
rect 10152 22098 10180 24568
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10508 24268 10560 24274
rect 10704 24256 10732 24822
rect 10796 24313 10824 27520
rect 10874 25392 10930 25401
rect 10980 25362 11100 25378
rect 10874 25327 10930 25336
rect 10968 25356 11100 25362
rect 10888 25129 10916 25327
rect 11020 25350 11100 25356
rect 10968 25298 11020 25304
rect 10874 25120 10930 25129
rect 10874 25055 10930 25064
rect 10968 24608 11020 24614
rect 10968 24550 11020 24556
rect 10508 24210 10560 24216
rect 10612 24228 10732 24256
rect 10782 24304 10838 24313
rect 10782 24239 10838 24248
rect 10876 24268 10928 24274
rect 10520 23662 10548 24210
rect 10508 23656 10560 23662
rect 10508 23598 10560 23604
rect 10612 23610 10640 24228
rect 10876 24210 10928 24216
rect 10784 24200 10836 24206
rect 10784 24142 10836 24148
rect 10612 23582 10732 23610
rect 10796 23594 10824 24142
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10704 23066 10732 23582
rect 10784 23588 10836 23594
rect 10784 23530 10836 23536
rect 10612 23038 10732 23066
rect 10506 22536 10562 22545
rect 10506 22471 10508 22480
rect 10560 22471 10562 22480
rect 10508 22442 10560 22448
rect 10612 22420 10640 23038
rect 10692 22976 10744 22982
rect 10692 22918 10744 22924
rect 10704 22574 10732 22918
rect 10692 22568 10744 22574
rect 10692 22510 10744 22516
rect 10612 22392 10732 22420
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10598 22128 10654 22137
rect 10140 22092 10192 22098
rect 10598 22063 10654 22072
rect 10140 22034 10192 22040
rect 10612 21418 10640 22063
rect 10704 21962 10732 22392
rect 10692 21956 10744 21962
rect 10692 21898 10744 21904
rect 10690 21448 10746 21457
rect 10600 21412 10652 21418
rect 10690 21383 10746 21392
rect 10600 21354 10652 21360
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10704 20602 10732 21383
rect 10692 20596 10744 20602
rect 10060 20556 10180 20584
rect 9956 20460 10008 20466
rect 9956 20402 10008 20408
rect 10048 20392 10100 20398
rect 10048 20334 10100 20340
rect 9956 20256 10008 20262
rect 9862 20224 9918 20233
rect 9956 20198 10008 20204
rect 9862 20159 9918 20168
rect 9772 19848 9824 19854
rect 9772 19790 9824 19796
rect 9784 19514 9812 19790
rect 9772 19508 9824 19514
rect 9772 19450 9824 19456
rect 9580 19366 9628 19394
rect 9580 19242 9608 19366
rect 9580 19236 9640 19242
rect 9580 19196 9588 19236
rect 9588 19178 9640 19184
rect 9600 18766 9628 19178
rect 9588 18760 9640 18766
rect 9588 18702 9640 18708
rect 9600 18222 9628 18702
rect 9588 18216 9640 18222
rect 9588 18158 9640 18164
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 9494 16688 9550 16697
rect 9494 16623 9550 16632
rect 9496 15904 9548 15910
rect 9496 15846 9548 15852
rect 9508 15366 9536 15846
rect 9496 15360 9548 15366
rect 9496 15302 9548 15308
rect 9600 14618 9628 17138
rect 9692 16561 9720 17478
rect 9772 17264 9824 17270
rect 9772 17206 9824 17212
rect 9678 16552 9734 16561
rect 9678 16487 9734 16496
rect 9678 16416 9734 16425
rect 9678 16351 9734 16360
rect 9692 15706 9720 16351
rect 9784 16130 9812 17206
rect 9876 16946 9904 20159
rect 9968 20097 9996 20198
rect 9954 20088 10010 20097
rect 9954 20023 10010 20032
rect 10060 19258 10088 20334
rect 10152 19938 10180 20556
rect 10692 20538 10744 20544
rect 10796 20398 10824 23530
rect 10888 23050 10916 24210
rect 10980 23361 11008 24550
rect 11072 24410 11100 25350
rect 11152 24744 11204 24750
rect 11150 24712 11152 24721
rect 11204 24712 11206 24721
rect 11150 24647 11206 24656
rect 11244 24608 11296 24614
rect 11242 24576 11244 24585
rect 11296 24576 11298 24585
rect 11242 24511 11298 24520
rect 11242 24440 11298 24449
rect 11060 24404 11112 24410
rect 11242 24375 11298 24384
rect 11060 24346 11112 24352
rect 11256 23866 11284 24375
rect 11244 23860 11296 23866
rect 11244 23802 11296 23808
rect 11242 23760 11298 23769
rect 11242 23695 11298 23704
rect 11256 23662 11284 23695
rect 11060 23656 11112 23662
rect 11058 23624 11060 23633
rect 11244 23656 11296 23662
rect 11112 23624 11114 23633
rect 11244 23598 11296 23604
rect 11058 23559 11114 23568
rect 11060 23520 11112 23526
rect 11060 23462 11112 23468
rect 10966 23352 11022 23361
rect 11072 23322 11100 23462
rect 10966 23287 11022 23296
rect 11060 23316 11112 23322
rect 11060 23258 11112 23264
rect 10876 23044 10928 23050
rect 10876 22986 10928 22992
rect 10888 20777 10916 22986
rect 11072 22778 11100 23258
rect 11152 23112 11204 23118
rect 11152 23054 11204 23060
rect 11060 22772 11112 22778
rect 11060 22714 11112 22720
rect 11060 22432 11112 22438
rect 11060 22374 11112 22380
rect 10968 21888 11020 21894
rect 11072 21842 11100 22374
rect 11164 22166 11192 23054
rect 11244 22636 11296 22642
rect 11244 22578 11296 22584
rect 11152 22160 11204 22166
rect 11152 22102 11204 22108
rect 11256 22098 11284 22578
rect 11244 22092 11296 22098
rect 11244 22034 11296 22040
rect 11150 21992 11206 22001
rect 11150 21927 11206 21936
rect 11020 21836 11100 21842
rect 10968 21830 11100 21836
rect 10980 21814 11100 21830
rect 11072 21729 11100 21814
rect 11058 21720 11114 21729
rect 11058 21655 11114 21664
rect 10968 21412 11020 21418
rect 10968 21354 11020 21360
rect 10874 20768 10930 20777
rect 10874 20703 10930 20712
rect 10876 20596 10928 20602
rect 10876 20538 10928 20544
rect 10784 20392 10836 20398
rect 10784 20334 10836 20340
rect 10692 20324 10744 20330
rect 10692 20266 10744 20272
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10416 19984 10468 19990
rect 10152 19910 10272 19938
rect 10416 19926 10468 19932
rect 10060 19230 10171 19258
rect 10244 19242 10272 19910
rect 10428 19281 10456 19926
rect 10414 19272 10470 19281
rect 9956 19168 10008 19174
rect 9956 19110 10008 19116
rect 10048 19168 10100 19174
rect 10048 19110 10100 19116
rect 9959 18986 9987 19110
rect 9959 18958 9996 18986
rect 10060 18970 10088 19110
rect 9968 17270 9996 18958
rect 10048 18964 10100 18970
rect 10048 18906 10100 18912
rect 10143 18680 10171 19230
rect 10232 19236 10284 19242
rect 10414 19207 10470 19216
rect 10232 19178 10284 19184
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10232 18896 10284 18902
rect 10232 18838 10284 18844
rect 10060 18652 10171 18680
rect 9956 17264 10008 17270
rect 9956 17206 10008 17212
rect 9876 16918 9996 16946
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 9876 16250 9904 16730
rect 9968 16250 9996 16918
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 9956 16244 10008 16250
rect 9956 16186 10008 16192
rect 9784 16102 9996 16130
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9864 15700 9916 15706
rect 9864 15642 9916 15648
rect 9772 15428 9824 15434
rect 9772 15370 9824 15376
rect 9784 14890 9812 15370
rect 9772 14884 9824 14890
rect 9772 14826 9824 14832
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9600 14006 9628 14554
rect 9784 14414 9812 14826
rect 9772 14408 9824 14414
rect 9678 14376 9734 14385
rect 9734 14356 9772 14362
rect 9734 14350 9824 14356
rect 9734 14334 9812 14350
rect 9678 14311 9734 14320
rect 9588 14000 9640 14006
rect 9588 13942 9640 13948
rect 9692 13818 9720 14311
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 9404 13796 9456 13802
rect 9404 13738 9456 13744
rect 9600 13790 9720 13818
rect 9600 13394 9628 13790
rect 9680 13728 9732 13734
rect 9680 13670 9732 13676
rect 9588 13388 9640 13394
rect 9588 13330 9640 13336
rect 9588 13252 9640 13258
rect 9588 13194 9640 13200
rect 9600 13161 9628 13194
rect 9586 13152 9642 13161
rect 9586 13087 9642 13096
rect 9588 12980 9640 12986
rect 9588 12922 9640 12928
rect 9496 11688 9548 11694
rect 9496 11630 9548 11636
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9128 10532 9180 10538
rect 9128 10474 9180 10480
rect 9034 10296 9090 10305
rect 9034 10231 9090 10240
rect 9140 10010 9168 10474
rect 9218 10432 9274 10441
rect 9218 10367 9274 10376
rect 9232 10198 9260 10367
rect 9220 10192 9272 10198
rect 9220 10134 9272 10140
rect 9324 10130 9352 11290
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9312 10124 9364 10130
rect 9312 10066 9364 10072
rect 9140 9982 9260 10010
rect 9126 9888 9182 9897
rect 9126 9823 9182 9832
rect 8864 9574 9076 9602
rect 8944 9512 8996 9518
rect 8942 9480 8944 9489
rect 8996 9480 8998 9489
rect 8942 9415 8998 9424
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 8852 8424 8904 8430
rect 8850 8392 8852 8401
rect 8904 8392 8906 8401
rect 8850 8327 8906 8336
rect 8850 7848 8906 7857
rect 8850 7783 8906 7792
rect 8864 7274 8892 7783
rect 8852 7268 8904 7274
rect 8852 7210 8904 7216
rect 8852 5024 8904 5030
rect 8852 4966 8904 4972
rect 8864 4486 8892 4966
rect 8852 4480 8904 4486
rect 8852 4422 8904 4428
rect 8956 4321 8984 9318
rect 8942 4312 8998 4321
rect 8942 4247 8998 4256
rect 8772 4134 8984 4162
rect 8392 4004 8444 4010
rect 8392 3946 8444 3952
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8220 3466 8248 3674
rect 8298 3632 8354 3641
rect 8298 3567 8354 3576
rect 8208 3460 8260 3466
rect 8208 3402 8260 3408
rect 7930 3224 7986 3233
rect 7760 3194 7880 3210
rect 7760 3188 7892 3194
rect 7760 3182 7840 3188
rect 7930 3159 7986 3168
rect 7840 3130 7892 3136
rect 7932 2916 7984 2922
rect 7932 2858 7984 2864
rect 7944 2650 7972 2858
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 7562 1592 7618 1601
rect 7562 1527 7618 1536
rect 7746 1456 7802 1465
rect 7746 1391 7802 1400
rect 7760 610 7788 1391
rect 8312 1034 8340 3567
rect 8404 2553 8432 3946
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 8666 3496 8722 3505
rect 8496 3194 8524 3470
rect 8666 3431 8722 3440
rect 8680 3194 8708 3431
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8668 3188 8720 3194
rect 8668 3130 8720 3136
rect 8390 2544 8446 2553
rect 8390 2479 8446 2488
rect 8312 1006 8432 1034
rect 7748 604 7800 610
rect 7748 546 7800 552
rect 7840 604 7892 610
rect 7840 546 7892 552
rect 7852 480 7880 546
rect 8404 480 8432 1006
rect 8956 480 8984 4134
rect 9048 2514 9076 9574
rect 9140 8362 9168 9823
rect 9232 9450 9260 9982
rect 9220 9444 9272 9450
rect 9220 9386 9272 9392
rect 9128 8356 9180 8362
rect 9128 8298 9180 8304
rect 9126 8256 9182 8265
rect 9126 8191 9182 8200
rect 9140 5166 9168 8191
rect 9232 7206 9260 9386
rect 9416 9382 9444 11018
rect 9508 9994 9536 11630
rect 9600 10606 9628 12922
rect 9692 12442 9720 13670
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9784 12322 9812 14214
rect 9876 12986 9904 15642
rect 9968 14278 9996 16102
rect 10060 16096 10088 18652
rect 10244 18612 10272 18838
rect 10152 18584 10272 18612
rect 10152 17785 10180 18584
rect 10704 18426 10732 20266
rect 10782 20224 10838 20233
rect 10782 20159 10838 20168
rect 10796 20058 10824 20159
rect 10784 20052 10836 20058
rect 10784 19994 10836 20000
rect 10782 18864 10838 18873
rect 10782 18799 10838 18808
rect 10692 18420 10744 18426
rect 10692 18362 10744 18368
rect 10692 18284 10744 18290
rect 10692 18226 10744 18232
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10704 17882 10732 18226
rect 10692 17876 10744 17882
rect 10692 17818 10744 17824
rect 10138 17776 10194 17785
rect 10138 17711 10194 17720
rect 10416 17740 10468 17746
rect 10416 17682 10468 17688
rect 10232 17672 10284 17678
rect 10232 17614 10284 17620
rect 10244 17202 10272 17614
rect 10428 17270 10456 17682
rect 10416 17264 10468 17270
rect 10414 17232 10416 17241
rect 10468 17232 10470 17241
rect 10232 17196 10284 17202
rect 10414 17167 10470 17176
rect 10232 17138 10284 17144
rect 10796 16998 10824 18799
rect 10888 17921 10916 20538
rect 10980 18086 11008 21354
rect 11072 21185 11100 21655
rect 11058 21176 11114 21185
rect 11058 21111 11114 21120
rect 11058 20904 11114 20913
rect 11058 20839 11060 20848
rect 11112 20839 11114 20848
rect 11060 20810 11112 20816
rect 11164 19786 11192 21927
rect 11256 21350 11284 22034
rect 11244 21344 11296 21350
rect 11244 21286 11296 21292
rect 11242 21176 11298 21185
rect 11242 21111 11298 21120
rect 11256 20097 11284 21111
rect 11242 20088 11298 20097
rect 11242 20023 11298 20032
rect 11152 19780 11204 19786
rect 11152 19722 11204 19728
rect 11060 19712 11112 19718
rect 11060 19654 11112 19660
rect 11072 19553 11100 19654
rect 11058 19544 11114 19553
rect 11058 19479 11114 19488
rect 11152 19168 11204 19174
rect 11204 19128 11284 19156
rect 11152 19110 11204 19116
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 10968 18080 11020 18086
rect 10968 18022 11020 18028
rect 10874 17912 10930 17921
rect 10874 17847 10930 17856
rect 10876 17808 10928 17814
rect 10876 17750 10928 17756
rect 10888 17134 10916 17750
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10784 16992 10836 16998
rect 10980 16980 11008 18022
rect 11072 17678 11100 18770
rect 11150 18592 11206 18601
rect 11150 18527 11206 18536
rect 11164 18057 11192 18527
rect 11150 18048 11206 18057
rect 11150 17983 11206 17992
rect 11060 17672 11112 17678
rect 11060 17614 11112 17620
rect 11072 17338 11100 17614
rect 11060 17332 11112 17338
rect 11060 17274 11112 17280
rect 11060 17196 11112 17202
rect 11060 17138 11112 17144
rect 10784 16934 10836 16940
rect 10888 16952 11008 16980
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10690 16824 10746 16833
rect 10690 16759 10692 16768
rect 10744 16759 10746 16768
rect 10692 16730 10744 16736
rect 10232 16652 10284 16658
rect 10232 16594 10284 16600
rect 10060 16068 10180 16096
rect 10048 15972 10100 15978
rect 10048 15914 10100 15920
rect 10060 14958 10088 15914
rect 10048 14952 10100 14958
rect 10048 14894 10100 14900
rect 9956 14272 10008 14278
rect 9956 14214 10008 14220
rect 10046 14240 10102 14249
rect 10046 14175 10102 14184
rect 10060 14074 10088 14175
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 9956 14000 10008 14006
rect 9956 13942 10008 13948
rect 9968 13462 9996 13942
rect 9956 13456 10008 13462
rect 9956 13398 10008 13404
rect 9968 12986 9996 13398
rect 9864 12980 9916 12986
rect 9864 12922 9916 12928
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 9956 12844 10008 12850
rect 9956 12786 10008 12792
rect 9968 12374 9996 12786
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 9864 12368 9916 12374
rect 9692 12294 9812 12322
rect 9862 12336 9864 12345
rect 9956 12368 10008 12374
rect 9916 12336 9918 12345
rect 9692 11937 9720 12294
rect 9956 12310 10008 12316
rect 9862 12271 9918 12280
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 9772 12096 9824 12102
rect 9772 12038 9824 12044
rect 9678 11928 9734 11937
rect 9784 11898 9812 12038
rect 9678 11863 9734 11872
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 9692 11393 9720 11698
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 9678 11384 9734 11393
rect 9678 11319 9734 11328
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 9586 10296 9642 10305
rect 9586 10231 9642 10240
rect 9496 9988 9548 9994
rect 9496 9930 9548 9936
rect 9404 9376 9456 9382
rect 9324 9324 9404 9330
rect 9324 9318 9456 9324
rect 9324 9302 9444 9318
rect 9324 9110 9352 9302
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 9312 9104 9364 9110
rect 9312 9046 9364 9052
rect 9310 8664 9366 8673
rect 9310 8599 9366 8608
rect 9324 8090 9352 8599
rect 9312 8084 9364 8090
rect 9312 8026 9364 8032
rect 9220 7200 9272 7206
rect 9220 7142 9272 7148
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9232 5574 9260 6598
rect 9220 5568 9272 5574
rect 9220 5510 9272 5516
rect 9232 5234 9260 5510
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 9128 5160 9180 5166
rect 9128 5102 9180 5108
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9140 4826 9168 4966
rect 9128 4820 9180 4826
rect 9128 4762 9180 4768
rect 9232 4214 9260 5170
rect 9220 4208 9272 4214
rect 9220 4150 9272 4156
rect 9128 3936 9180 3942
rect 9126 3904 9128 3913
rect 9180 3904 9182 3913
rect 9126 3839 9182 3848
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 9140 3346 9168 3674
rect 9232 3534 9260 4150
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9140 3318 9260 3346
rect 9232 3126 9260 3318
rect 9220 3120 9272 3126
rect 9218 3088 9220 3097
rect 9272 3088 9274 3097
rect 9218 3023 9274 3032
rect 9324 2553 9352 6598
rect 9416 4622 9444 9114
rect 9508 9110 9536 9930
rect 9600 9897 9628 10231
rect 9586 9888 9642 9897
rect 9586 9823 9642 9832
rect 9588 9512 9640 9518
rect 9692 9500 9720 10746
rect 9784 10130 9812 11630
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9640 9472 9720 9500
rect 9588 9454 9640 9460
rect 9600 9178 9628 9454
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9496 9104 9548 9110
rect 9496 9046 9548 9052
rect 9772 8968 9824 8974
rect 9678 8936 9734 8945
rect 9772 8910 9824 8916
rect 9678 8871 9680 8880
rect 9732 8871 9734 8880
rect 9680 8842 9732 8848
rect 9784 8673 9812 8910
rect 9770 8664 9826 8673
rect 9770 8599 9826 8608
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 9600 8242 9628 8366
rect 9772 8356 9824 8362
rect 9772 8298 9824 8304
rect 9600 8214 9720 8242
rect 9588 7336 9640 7342
rect 9588 7278 9640 7284
rect 9600 7206 9628 7278
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 9600 6798 9628 7142
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9692 5914 9720 8214
rect 9784 8129 9812 8298
rect 9770 8120 9826 8129
rect 9770 8055 9826 8064
rect 9772 7812 9824 7818
rect 9772 7754 9824 7760
rect 9784 7546 9812 7754
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9784 6458 9812 6802
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9680 5908 9732 5914
rect 9680 5850 9732 5856
rect 9678 5808 9734 5817
rect 9678 5743 9734 5752
rect 9494 5128 9550 5137
rect 9692 5114 9720 5743
rect 9770 5264 9826 5273
rect 9770 5199 9826 5208
rect 9494 5063 9496 5072
rect 9548 5063 9550 5072
rect 9600 5086 9720 5114
rect 9496 5034 9548 5040
rect 9508 4826 9536 5034
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 9404 4616 9456 4622
rect 9404 4558 9456 4564
rect 9600 4162 9628 5086
rect 9678 4992 9734 5001
rect 9678 4927 9734 4936
rect 9692 4282 9720 4927
rect 9784 4826 9812 5199
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9876 4554 9904 12174
rect 9954 10568 10010 10577
rect 9954 10503 10010 10512
rect 9968 9178 9996 10503
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 10060 8673 10088 12718
rect 10152 12238 10180 16068
rect 10244 15978 10272 16594
rect 10324 16584 10376 16590
rect 10324 16526 10376 16532
rect 10336 16250 10364 16526
rect 10600 16516 10652 16522
rect 10600 16458 10652 16464
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 10612 16046 10640 16458
rect 10692 16448 10744 16454
rect 10692 16390 10744 16396
rect 10600 16040 10652 16046
rect 10600 15982 10652 15988
rect 10232 15972 10284 15978
rect 10232 15914 10284 15920
rect 10704 15910 10732 16390
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10692 15904 10744 15910
rect 10690 15872 10692 15881
rect 10744 15872 10746 15881
rect 10289 15804 10585 15824
rect 10690 15807 10746 15816
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10796 15706 10824 16050
rect 10784 15700 10836 15706
rect 10784 15642 10836 15648
rect 10784 14952 10836 14958
rect 10784 14894 10836 14900
rect 10692 14816 10744 14822
rect 10692 14758 10744 14764
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10704 14550 10732 14758
rect 10692 14544 10744 14550
rect 10692 14486 10744 14492
rect 10704 14074 10732 14486
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10692 13728 10744 13734
rect 10692 13670 10744 13676
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10600 13456 10652 13462
rect 10600 13398 10652 13404
rect 10612 12782 10640 13398
rect 10704 12850 10732 13670
rect 10796 13462 10824 14894
rect 10784 13456 10836 13462
rect 10784 13398 10836 13404
rect 10784 13252 10836 13258
rect 10784 13194 10836 13200
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10600 12776 10652 12782
rect 10600 12718 10652 12724
rect 10692 12708 10744 12714
rect 10692 12650 10744 12656
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10232 12368 10284 12374
rect 10232 12310 10284 12316
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 10244 11778 10272 12310
rect 10324 11892 10376 11898
rect 10324 11834 10376 11840
rect 10152 11750 10272 11778
rect 10046 8664 10102 8673
rect 10046 8599 10102 8608
rect 9956 7744 10008 7750
rect 9956 7686 10008 7692
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 9968 7342 9996 7686
rect 9956 7336 10008 7342
rect 9956 7278 10008 7284
rect 9968 6118 9996 7278
rect 10060 6361 10088 7686
rect 10046 6352 10102 6361
rect 10046 6287 10102 6296
rect 9956 6112 10008 6118
rect 9956 6054 10008 6060
rect 9968 5642 9996 6054
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 10060 5681 10088 5714
rect 10046 5672 10102 5681
rect 9956 5636 10008 5642
rect 10046 5607 10102 5616
rect 9956 5578 10008 5584
rect 9968 5370 9996 5578
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 10060 5250 10088 5510
rect 9968 5222 10088 5250
rect 9864 4548 9916 4554
rect 9864 4490 9916 4496
rect 9680 4276 9732 4282
rect 9680 4218 9732 4224
rect 9862 4176 9918 4185
rect 9600 4134 9720 4162
rect 9586 3768 9642 3777
rect 9692 3738 9720 4134
rect 9968 4162 9996 5222
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 9918 4134 9996 4162
rect 9862 4111 9918 4120
rect 9586 3703 9642 3712
rect 9680 3732 9732 3738
rect 9600 2650 9628 3703
rect 9680 3674 9732 3680
rect 9692 2961 9720 3674
rect 9876 3602 9904 4111
rect 9956 4072 10008 4078
rect 9956 4014 10008 4020
rect 9968 3942 9996 4014
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 9954 3768 10010 3777
rect 9954 3703 9956 3712
rect 10008 3703 10010 3712
rect 9956 3674 10008 3680
rect 9864 3596 9916 3602
rect 9864 3538 9916 3544
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 9678 2952 9734 2961
rect 9876 2922 9904 3334
rect 9968 3194 9996 3470
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 9678 2887 9734 2896
rect 9864 2916 9916 2922
rect 9864 2858 9916 2864
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9310 2544 9366 2553
rect 9036 2508 9088 2514
rect 9692 2514 9720 2790
rect 9310 2479 9366 2488
rect 9496 2508 9548 2514
rect 9036 2450 9088 2456
rect 9324 1737 9352 2479
rect 9496 2450 9548 2456
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 9310 1728 9366 1737
rect 9310 1663 9366 1672
rect 9508 480 9536 2450
rect 10060 480 10088 5102
rect 10152 4706 10180 11750
rect 10336 11665 10364 11834
rect 10322 11656 10378 11665
rect 10322 11591 10378 11600
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10704 11336 10732 12650
rect 10796 12646 10824 13194
rect 10784 12640 10836 12646
rect 10784 12582 10836 12588
rect 10796 12374 10824 12582
rect 10784 12368 10836 12374
rect 10784 12310 10836 12316
rect 10888 11898 10916 16952
rect 11072 16182 11100 17138
rect 11060 16176 11112 16182
rect 11060 16118 11112 16124
rect 11072 15162 11100 16118
rect 11164 15638 11192 17983
rect 11152 15632 11204 15638
rect 11152 15574 11204 15580
rect 11164 15162 11192 15574
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 11152 15156 11204 15162
rect 11152 15098 11204 15104
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 10980 13530 11008 13806
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 11072 13190 11100 14894
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 10966 13016 11022 13025
rect 10966 12951 11022 12960
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 10888 11626 10916 11698
rect 10876 11620 10928 11626
rect 10876 11562 10928 11568
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10520 11308 10732 11336
rect 10232 11076 10284 11082
rect 10232 11018 10284 11024
rect 10244 10849 10272 11018
rect 10230 10840 10286 10849
rect 10520 10810 10548 11308
rect 10796 11257 10824 11494
rect 10782 11248 10838 11257
rect 10600 11212 10652 11218
rect 10782 11183 10838 11192
rect 10600 11154 10652 11160
rect 10612 11121 10640 11154
rect 10888 11150 10916 11562
rect 10876 11144 10928 11150
rect 10598 11112 10654 11121
rect 10654 11070 10732 11098
rect 10876 11086 10928 11092
rect 10598 11047 10654 11056
rect 10230 10775 10286 10784
rect 10508 10804 10560 10810
rect 10508 10746 10560 10752
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10704 10266 10732 11070
rect 10782 10296 10838 10305
rect 10692 10260 10744 10266
rect 10782 10231 10838 10240
rect 10876 10260 10928 10266
rect 10692 10202 10744 10208
rect 10796 10198 10824 10231
rect 10876 10202 10928 10208
rect 10784 10192 10836 10198
rect 10784 10134 10836 10140
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 10336 9489 10364 10066
rect 10322 9480 10378 9489
rect 10322 9415 10378 9424
rect 10692 9376 10744 9382
rect 10690 9344 10692 9353
rect 10744 9344 10746 9353
rect 10289 9276 10585 9296
rect 10690 9279 10746 9288
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10244 8634 10272 8910
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10598 8392 10654 8401
rect 10598 8327 10600 8336
rect 10652 8327 10654 8336
rect 10600 8298 10652 8304
rect 10690 8256 10746 8265
rect 10289 8188 10585 8208
rect 10690 8191 10746 8200
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10704 8090 10732 8191
rect 10692 8084 10744 8090
rect 10888 8072 10916 10202
rect 10692 8026 10744 8032
rect 10796 8044 10916 8072
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10704 7002 10732 8026
rect 10692 6996 10744 7002
rect 10692 6938 10744 6944
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10690 6624 10746 6633
rect 10428 6254 10456 6598
rect 10690 6559 10746 6568
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10704 5817 10732 6559
rect 10690 5808 10746 5817
rect 10690 5743 10746 5752
rect 10600 5568 10652 5574
rect 10600 5510 10652 5516
rect 10612 5234 10640 5510
rect 10796 5302 10824 8044
rect 10980 5760 11008 12951
rect 11164 12170 11192 13126
rect 11256 12442 11284 19128
rect 11348 16833 11376 27520
rect 11900 26382 11928 27520
rect 11888 26376 11940 26382
rect 11888 26318 11940 26324
rect 11518 25936 11574 25945
rect 11518 25871 11574 25880
rect 11428 24812 11480 24818
rect 11428 24754 11480 24760
rect 11440 24138 11468 24754
rect 11428 24132 11480 24138
rect 11428 24074 11480 24080
rect 11532 23866 11560 25871
rect 11612 25356 11664 25362
rect 11612 25298 11664 25304
rect 11796 25356 11848 25362
rect 11796 25298 11848 25304
rect 11624 24818 11652 25298
rect 11808 25226 11836 25298
rect 11796 25220 11848 25226
rect 11796 25162 11848 25168
rect 11612 24812 11664 24818
rect 11612 24754 11664 24760
rect 11980 24812 12032 24818
rect 11980 24754 12032 24760
rect 11612 24404 11664 24410
rect 11612 24346 11664 24352
rect 11520 23860 11572 23866
rect 11520 23802 11572 23808
rect 11520 23588 11572 23594
rect 11520 23530 11572 23536
rect 11426 22808 11482 22817
rect 11426 22743 11428 22752
rect 11480 22743 11482 22752
rect 11428 22714 11480 22720
rect 11426 21720 11482 21729
rect 11426 21655 11482 21664
rect 11440 21457 11468 21655
rect 11426 21448 11482 21457
rect 11426 21383 11482 21392
rect 11428 21344 11480 21350
rect 11428 21286 11480 21292
rect 11440 19854 11468 21286
rect 11532 20534 11560 23530
rect 11520 20528 11572 20534
rect 11520 20470 11572 20476
rect 11520 20324 11572 20330
rect 11520 20266 11572 20272
rect 11532 20058 11560 20266
rect 11520 20052 11572 20058
rect 11520 19994 11572 20000
rect 11428 19848 11480 19854
rect 11428 19790 11480 19796
rect 11440 19174 11468 19790
rect 11518 19544 11574 19553
rect 11518 19479 11574 19488
rect 11428 19168 11480 19174
rect 11428 19110 11480 19116
rect 11440 18630 11468 19110
rect 11532 18902 11560 19479
rect 11520 18896 11572 18902
rect 11520 18838 11572 18844
rect 11518 18728 11574 18737
rect 11518 18663 11574 18672
rect 11428 18624 11480 18630
rect 11428 18566 11480 18572
rect 11440 18290 11468 18566
rect 11532 18426 11560 18663
rect 11520 18420 11572 18426
rect 11520 18362 11572 18368
rect 11428 18284 11480 18290
rect 11428 18226 11480 18232
rect 11426 17912 11482 17921
rect 11426 17847 11482 17856
rect 11334 16824 11390 16833
rect 11334 16759 11390 16768
rect 11440 16658 11468 17847
rect 11532 17814 11560 18362
rect 11520 17808 11572 17814
rect 11520 17750 11572 17756
rect 11624 16726 11652 24346
rect 11704 24064 11756 24070
rect 11704 24006 11756 24012
rect 11716 21321 11744 24006
rect 11796 23248 11848 23254
rect 11796 23190 11848 23196
rect 11808 22982 11836 23190
rect 11796 22976 11848 22982
rect 11796 22918 11848 22924
rect 11808 22012 11836 22918
rect 11992 22098 12020 24754
rect 12256 24744 12308 24750
rect 12256 24686 12308 24692
rect 12164 24608 12216 24614
rect 12164 24550 12216 24556
rect 12176 24410 12204 24550
rect 12164 24404 12216 24410
rect 12164 24346 12216 24352
rect 12072 24200 12124 24206
rect 12072 24142 12124 24148
rect 12084 23254 12112 24142
rect 12176 23322 12204 24346
rect 12268 24041 12296 24686
rect 12440 24404 12492 24410
rect 12440 24346 12492 24352
rect 12348 24268 12400 24274
rect 12348 24210 12400 24216
rect 12254 24032 12310 24041
rect 12254 23967 12310 23976
rect 12164 23316 12216 23322
rect 12164 23258 12216 23264
rect 12072 23248 12124 23254
rect 12072 23190 12124 23196
rect 12072 23112 12124 23118
rect 12072 23054 12124 23060
rect 11980 22092 12032 22098
rect 11980 22034 12032 22040
rect 11808 21984 11928 22012
rect 11702 21312 11758 21321
rect 11702 21247 11758 21256
rect 11900 21026 11928 21984
rect 12084 21978 12112 23054
rect 12164 22976 12216 22982
rect 12164 22918 12216 22924
rect 12176 22681 12204 22918
rect 12360 22710 12388 24210
rect 12452 24041 12480 24346
rect 12438 24032 12494 24041
rect 12438 23967 12494 23976
rect 12438 23760 12494 23769
rect 12438 23695 12494 23704
rect 12452 23662 12480 23695
rect 12440 23656 12492 23662
rect 12440 23598 12492 23604
rect 12440 23180 12492 23186
rect 12440 23122 12492 23128
rect 12452 22778 12480 23122
rect 12440 22772 12492 22778
rect 12440 22714 12492 22720
rect 12348 22704 12400 22710
rect 12162 22672 12218 22681
rect 12348 22646 12400 22652
rect 12162 22607 12218 22616
rect 12256 22636 12308 22642
rect 12256 22578 12308 22584
rect 12162 22536 12218 22545
rect 12162 22471 12218 22480
rect 11992 21950 12112 21978
rect 11992 21894 12020 21950
rect 11980 21888 12032 21894
rect 11980 21830 12032 21836
rect 11808 20998 11928 21026
rect 11704 20528 11756 20534
rect 11704 20470 11756 20476
rect 11716 18601 11744 20470
rect 11808 18834 11836 20998
rect 11992 20466 12020 21830
rect 12176 21026 12204 22471
rect 12268 21690 12296 22578
rect 12440 22432 12492 22438
rect 12440 22374 12492 22380
rect 12452 22166 12480 22374
rect 12348 22160 12400 22166
rect 12348 22102 12400 22108
rect 12440 22160 12492 22166
rect 12440 22102 12492 22108
rect 12360 21690 12388 22102
rect 12256 21684 12308 21690
rect 12256 21626 12308 21632
rect 12348 21684 12400 21690
rect 12348 21626 12400 21632
rect 12346 21448 12402 21457
rect 12346 21383 12402 21392
rect 12084 20998 12204 21026
rect 11980 20460 12032 20466
rect 11980 20402 12032 20408
rect 11980 19984 12032 19990
rect 11980 19926 12032 19932
rect 11888 19780 11940 19786
rect 11888 19722 11940 19728
rect 11900 19174 11928 19722
rect 11992 19174 12020 19926
rect 11888 19168 11940 19174
rect 11886 19136 11888 19145
rect 11980 19168 12032 19174
rect 11940 19136 11942 19145
rect 11980 19110 12032 19116
rect 11886 19071 11942 19080
rect 11992 18952 12020 19110
rect 11900 18924 12020 18952
rect 11796 18828 11848 18834
rect 11796 18770 11848 18776
rect 11796 18692 11848 18698
rect 11796 18634 11848 18640
rect 11702 18592 11758 18601
rect 11702 18527 11758 18536
rect 11702 18320 11758 18329
rect 11702 18255 11758 18264
rect 11716 17814 11744 18255
rect 11704 17808 11756 17814
rect 11704 17750 11756 17756
rect 11716 16794 11744 17750
rect 11704 16788 11756 16794
rect 11704 16730 11756 16736
rect 11612 16720 11664 16726
rect 11612 16662 11664 16668
rect 11808 16658 11836 18634
rect 11428 16652 11480 16658
rect 11428 16594 11480 16600
rect 11796 16652 11848 16658
rect 11796 16594 11848 16600
rect 11426 16144 11482 16153
rect 11426 16079 11482 16088
rect 11610 16144 11666 16153
rect 11610 16079 11666 16088
rect 11440 15910 11468 16079
rect 11428 15904 11480 15910
rect 11428 15846 11480 15852
rect 11518 14104 11574 14113
rect 11518 14039 11574 14048
rect 11428 13864 11480 13870
rect 11334 13832 11390 13841
rect 11428 13806 11480 13812
rect 11334 13767 11390 13776
rect 11348 12850 11376 13767
rect 11440 13433 11468 13806
rect 11426 13424 11482 13433
rect 11426 13359 11482 13368
rect 11336 12844 11388 12850
rect 11336 12786 11388 12792
rect 11244 12436 11296 12442
rect 11244 12378 11296 12384
rect 11428 12368 11480 12374
rect 11428 12310 11480 12316
rect 11244 12300 11296 12306
rect 11244 12242 11296 12248
rect 11152 12164 11204 12170
rect 11152 12106 11204 12112
rect 11058 11656 11114 11665
rect 11058 11591 11060 11600
rect 11112 11591 11114 11600
rect 11060 11562 11112 11568
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 11072 10810 11100 11290
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 11060 10192 11112 10198
rect 11060 10134 11112 10140
rect 11072 9382 11100 10134
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 11164 8242 11192 11494
rect 11256 11082 11284 12242
rect 11440 12209 11468 12310
rect 11426 12200 11482 12209
rect 11426 12135 11482 12144
rect 11532 11354 11560 14039
rect 11624 11694 11652 16079
rect 11808 15570 11836 16594
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 11808 14521 11836 14758
rect 11794 14512 11850 14521
rect 11704 14476 11756 14482
rect 11794 14447 11850 14456
rect 11704 14418 11756 14424
rect 11716 13938 11744 14418
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11704 13932 11756 13938
rect 11704 13874 11756 13880
rect 11808 13462 11836 14010
rect 11796 13456 11848 13462
rect 11796 13398 11848 13404
rect 11702 13288 11758 13297
rect 11808 13258 11836 13398
rect 11702 13223 11758 13232
rect 11796 13252 11848 13258
rect 11716 13138 11744 13223
rect 11796 13194 11848 13200
rect 11716 13110 11836 13138
rect 11702 13016 11758 13025
rect 11702 12951 11704 12960
rect 11756 12951 11758 12960
rect 11704 12922 11756 12928
rect 11702 12472 11758 12481
rect 11702 12407 11758 12416
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 11520 11348 11572 11354
rect 11520 11290 11572 11296
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11336 11144 11388 11150
rect 11336 11086 11388 11092
rect 11244 11076 11296 11082
rect 11244 11018 11296 11024
rect 11256 10538 11284 11018
rect 11348 10810 11376 11086
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 11244 10532 11296 10538
rect 11244 10474 11296 10480
rect 11348 10198 11376 10746
rect 11336 10192 11388 10198
rect 11336 10134 11388 10140
rect 11348 9722 11376 10134
rect 11532 10130 11560 11154
rect 11610 10704 11666 10713
rect 11610 10639 11666 10648
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11336 9716 11388 9722
rect 11336 9658 11388 9664
rect 11244 9172 11296 9178
rect 11244 9114 11296 9120
rect 11256 8430 11284 9114
rect 11336 9036 11388 9042
rect 11336 8978 11388 8984
rect 11348 8498 11376 8978
rect 11532 8974 11560 10066
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11072 7993 11100 8230
rect 11164 8214 11284 8242
rect 11058 7984 11114 7993
rect 11058 7919 11114 7928
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 11072 7274 11100 7822
rect 11060 7268 11112 7274
rect 11060 7210 11112 7216
rect 11152 7268 11204 7274
rect 11152 7210 11204 7216
rect 11072 6662 11100 7210
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11164 6474 11192 7210
rect 10888 5732 11008 5760
rect 11072 6446 11192 6474
rect 10784 5296 10836 5302
rect 10784 5238 10836 5244
rect 10600 5228 10652 5234
rect 10600 5170 10652 5176
rect 10888 5166 10916 5732
rect 10968 5296 11020 5302
rect 10968 5238 11020 5244
rect 10876 5160 10928 5166
rect 10876 5102 10928 5108
rect 10784 5024 10836 5030
rect 10690 4992 10746 5001
rect 10289 4924 10585 4944
rect 10784 4966 10836 4972
rect 10690 4927 10746 4936
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10704 4826 10732 4927
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10152 4678 10732 4706
rect 10140 4548 10192 4554
rect 10140 4490 10192 4496
rect 10152 3233 10180 4490
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10138 3224 10194 3233
rect 10138 3159 10194 3168
rect 10152 2689 10180 3159
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10138 2680 10194 2689
rect 10289 2672 10585 2692
rect 10138 2615 10194 2624
rect 10704 1442 10732 4678
rect 10796 4554 10824 4966
rect 10980 4758 11008 5238
rect 11072 5030 11100 6446
rect 11152 5840 11204 5846
rect 11152 5782 11204 5788
rect 11164 5574 11192 5782
rect 11152 5568 11204 5574
rect 11256 5545 11284 8214
rect 11348 8090 11376 8434
rect 11336 8084 11388 8090
rect 11336 8026 11388 8032
rect 11348 7546 11376 8026
rect 11336 7540 11388 7546
rect 11336 7482 11388 7488
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11152 5510 11204 5516
rect 11242 5536 11298 5545
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 10968 4752 11020 4758
rect 10968 4694 11020 4700
rect 10784 4548 10836 4554
rect 10784 4490 10836 4496
rect 10796 4298 10824 4490
rect 10796 4270 10916 4298
rect 10782 2680 10838 2689
rect 10782 2615 10838 2624
rect 10796 2582 10824 2615
rect 10888 2582 10916 4270
rect 10980 4214 11008 4694
rect 11164 4622 11192 5510
rect 11242 5471 11298 5480
rect 11348 5234 11376 6802
rect 11532 6254 11560 8910
rect 11520 6248 11572 6254
rect 11520 6190 11572 6196
rect 11518 5944 11574 5953
rect 11518 5879 11520 5888
rect 11572 5879 11574 5888
rect 11520 5850 11572 5856
rect 11244 5228 11296 5234
rect 11244 5170 11296 5176
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 11256 4758 11284 5170
rect 11532 5030 11560 5850
rect 11624 5098 11652 10639
rect 11612 5092 11664 5098
rect 11612 5034 11664 5040
rect 11520 5024 11572 5030
rect 11426 4992 11482 5001
rect 11520 4966 11572 4972
rect 11426 4927 11482 4936
rect 11244 4752 11296 4758
rect 11244 4694 11296 4700
rect 11334 4720 11390 4729
rect 11334 4655 11336 4664
rect 11388 4655 11390 4664
rect 11336 4626 11388 4632
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 10968 4208 11020 4214
rect 10968 4150 11020 4156
rect 11348 4078 11376 4626
rect 11440 4146 11468 4927
rect 11716 4604 11744 12407
rect 11808 9178 11836 13110
rect 11900 12356 11928 18924
rect 11980 16652 12032 16658
rect 11980 16594 12032 16600
rect 11992 15706 12020 16594
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 12084 15144 12112 20998
rect 12164 20936 12216 20942
rect 12162 20904 12164 20913
rect 12216 20904 12218 20913
rect 12162 20839 12218 20848
rect 12360 20058 12388 21383
rect 12440 21344 12492 21350
rect 12440 21286 12492 21292
rect 12452 21049 12480 21286
rect 12438 21040 12494 21049
rect 12438 20975 12494 20984
rect 12452 20806 12480 20975
rect 12440 20800 12492 20806
rect 12440 20742 12492 20748
rect 12438 20632 12494 20641
rect 12438 20567 12440 20576
rect 12492 20567 12494 20576
rect 12440 20538 12492 20544
rect 12348 20052 12400 20058
rect 12348 19994 12400 20000
rect 12440 19916 12492 19922
rect 12440 19858 12492 19864
rect 12164 19780 12216 19786
rect 12164 19722 12216 19728
rect 11992 15116 12112 15144
rect 11992 12458 12020 15116
rect 12176 13705 12204 19722
rect 12452 19700 12480 19858
rect 12360 19672 12480 19700
rect 12256 18828 12308 18834
rect 12256 18770 12308 18776
rect 12268 18358 12296 18770
rect 12256 18352 12308 18358
rect 12256 18294 12308 18300
rect 12360 17882 12388 19672
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 12452 18737 12480 18770
rect 12438 18728 12494 18737
rect 12438 18663 12494 18672
rect 12440 18624 12492 18630
rect 12440 18566 12492 18572
rect 12348 17876 12400 17882
rect 12348 17818 12400 17824
rect 12452 17814 12480 18566
rect 12440 17808 12492 17814
rect 12440 17750 12492 17756
rect 12254 17368 12310 17377
rect 12254 17303 12310 17312
rect 12268 17202 12296 17303
rect 12544 17270 12572 27520
rect 13096 26042 13124 27520
rect 13084 26036 13136 26042
rect 13084 25978 13136 25984
rect 13176 26036 13228 26042
rect 13176 25978 13228 25984
rect 12992 25356 13044 25362
rect 12992 25298 13044 25304
rect 12898 24712 12954 24721
rect 12898 24647 12954 24656
rect 12808 24064 12860 24070
rect 12714 24032 12770 24041
rect 12808 24006 12860 24012
rect 12714 23967 12770 23976
rect 12728 23798 12756 23967
rect 12716 23792 12768 23798
rect 12716 23734 12768 23740
rect 12820 23526 12848 24006
rect 12912 23730 12940 24647
rect 13004 24614 13032 25298
rect 13188 25158 13216 25978
rect 13176 25152 13228 25158
rect 13176 25094 13228 25100
rect 13544 25152 13596 25158
rect 13544 25094 13596 25100
rect 13556 24750 13584 25094
rect 13648 24936 13676 27520
rect 13912 25356 13964 25362
rect 13912 25298 13964 25304
rect 13820 25288 13872 25294
rect 13820 25230 13872 25236
rect 13648 24908 13768 24936
rect 13634 24848 13690 24857
rect 13634 24783 13636 24792
rect 13688 24783 13690 24792
rect 13636 24754 13688 24760
rect 13084 24744 13136 24750
rect 13084 24686 13136 24692
rect 13544 24744 13596 24750
rect 13544 24686 13596 24692
rect 12992 24608 13044 24614
rect 12992 24550 13044 24556
rect 12900 23724 12952 23730
rect 12900 23666 12952 23672
rect 12808 23520 12860 23526
rect 12808 23462 12860 23468
rect 12716 23112 12768 23118
rect 12716 23054 12768 23060
rect 12622 21992 12678 22001
rect 12622 21927 12678 21936
rect 12532 17264 12584 17270
rect 12532 17206 12584 17212
rect 12256 17196 12308 17202
rect 12256 17138 12308 17144
rect 12438 17096 12494 17105
rect 12348 17060 12400 17066
rect 12438 17031 12494 17040
rect 12348 17002 12400 17008
rect 12360 16250 12388 17002
rect 12452 16998 12480 17031
rect 12440 16992 12492 16998
rect 12440 16934 12492 16940
rect 12348 16244 12400 16250
rect 12348 16186 12400 16192
rect 12346 15872 12402 15881
rect 12346 15807 12402 15816
rect 12360 15162 12388 15807
rect 12348 15156 12400 15162
rect 12348 15098 12400 15104
rect 12532 15088 12584 15094
rect 12532 15030 12584 15036
rect 12544 14929 12572 15030
rect 12530 14920 12586 14929
rect 12530 14855 12586 14864
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12452 14414 12480 14758
rect 12532 14476 12584 14482
rect 12532 14418 12584 14424
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 12452 14249 12480 14350
rect 12438 14240 12494 14249
rect 12438 14175 12494 14184
rect 12256 13932 12308 13938
rect 12256 13874 12308 13880
rect 12162 13696 12218 13705
rect 12162 13631 12218 13640
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 12176 12986 12204 13330
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 11992 12430 12112 12458
rect 11900 12328 12020 12356
rect 11900 12238 11928 12269
rect 11888 12232 11940 12238
rect 11886 12200 11888 12209
rect 11940 12200 11942 12209
rect 11886 12135 11942 12144
rect 11900 11898 11928 12135
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11992 11801 12020 12328
rect 11978 11792 12034 11801
rect 11978 11727 12034 11736
rect 11888 11688 11940 11694
rect 11888 11630 11940 11636
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 11794 8664 11850 8673
rect 11794 8599 11796 8608
rect 11848 8599 11850 8608
rect 11796 8570 11848 8576
rect 11808 8430 11836 8570
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 11900 8362 11928 11630
rect 11992 8673 12020 11727
rect 12084 11694 12112 12430
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 12176 11626 12204 12242
rect 12268 12170 12296 13874
rect 12544 13802 12572 14418
rect 12532 13796 12584 13802
rect 12532 13738 12584 13744
rect 12530 13696 12586 13705
rect 12530 13631 12586 13640
rect 12544 13530 12572 13631
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 12544 12986 12572 13466
rect 12636 13161 12664 21927
rect 12728 21672 12756 23054
rect 12820 22114 12848 23462
rect 12900 22500 12952 22506
rect 12900 22442 12952 22448
rect 12912 22234 12940 22442
rect 13004 22273 13032 24550
rect 12990 22264 13046 22273
rect 12900 22228 12952 22234
rect 12990 22199 13046 22208
rect 12900 22170 12952 22176
rect 12820 22086 12940 22114
rect 12728 21644 12848 21672
rect 12714 21584 12770 21593
rect 12714 21519 12770 21528
rect 12728 17678 12756 21519
rect 12820 20913 12848 21644
rect 12806 20904 12862 20913
rect 12806 20839 12862 20848
rect 12808 20392 12860 20398
rect 12808 20334 12860 20340
rect 12820 20233 12848 20334
rect 12806 20224 12862 20233
rect 12806 20159 12862 20168
rect 12808 19848 12860 19854
rect 12808 19790 12860 19796
rect 12820 19514 12848 19790
rect 12808 19508 12860 19514
rect 12808 19450 12860 19456
rect 12820 18970 12848 19450
rect 12808 18964 12860 18970
rect 12808 18906 12860 18912
rect 12806 18864 12862 18873
rect 12806 18799 12862 18808
rect 12820 18426 12848 18799
rect 12912 18442 12940 22086
rect 12990 20224 13046 20233
rect 12990 20159 13046 20168
rect 13004 19990 13032 20159
rect 13096 20058 13124 24686
rect 13268 24676 13320 24682
rect 13268 24618 13320 24624
rect 13176 24064 13228 24070
rect 13176 24006 13228 24012
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 12992 19984 13044 19990
rect 12992 19926 13044 19932
rect 13004 19310 13032 19926
rect 12992 19304 13044 19310
rect 12992 19246 13044 19252
rect 13004 18970 13032 19246
rect 12992 18964 13044 18970
rect 12992 18906 13044 18912
rect 12808 18420 12860 18426
rect 12912 18414 13124 18442
rect 12808 18362 12860 18368
rect 12900 18352 12952 18358
rect 12900 18294 12952 18300
rect 12716 17672 12768 17678
rect 12716 17614 12768 17620
rect 12806 17640 12862 17649
rect 12806 17575 12862 17584
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12728 17134 12756 17478
rect 12820 17377 12848 17575
rect 12806 17368 12862 17377
rect 12806 17303 12862 17312
rect 12808 17264 12860 17270
rect 12808 17206 12860 17212
rect 12716 17128 12768 17134
rect 12716 17070 12768 17076
rect 12728 15706 12756 17070
rect 12716 15700 12768 15706
rect 12716 15642 12768 15648
rect 12820 15586 12848 17206
rect 12912 16794 12940 18294
rect 12992 18080 13044 18086
rect 12992 18022 13044 18028
rect 13004 17921 13032 18022
rect 12990 17912 13046 17921
rect 12990 17847 13046 17856
rect 12992 17672 13044 17678
rect 12992 17614 13044 17620
rect 12900 16788 12952 16794
rect 12900 16730 12952 16736
rect 12900 16108 12952 16114
rect 12900 16050 12952 16056
rect 12728 15558 12848 15586
rect 12622 13152 12678 13161
rect 12728 13138 12756 15558
rect 12912 15450 12940 16050
rect 12820 15422 12940 15450
rect 12820 15366 12848 15422
rect 12808 15360 12860 15366
rect 12806 15328 12808 15337
rect 12860 15328 12862 15337
rect 12806 15263 12862 15272
rect 12820 14770 12848 15263
rect 13004 14929 13032 17614
rect 13096 17542 13124 18414
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 13084 17264 13136 17270
rect 13084 17206 13136 17212
rect 12990 14920 13046 14929
rect 12990 14855 13046 14864
rect 12820 14742 13032 14770
rect 12808 14340 12860 14346
rect 12808 14282 12860 14288
rect 12820 13326 12848 14282
rect 12900 14272 12952 14278
rect 12900 14214 12952 14220
rect 12912 13977 12940 14214
rect 12898 13968 12954 13977
rect 12898 13903 12954 13912
rect 13004 13852 13032 14742
rect 12912 13824 13032 13852
rect 12808 13320 12860 13326
rect 12808 13262 12860 13268
rect 12728 13110 12848 13138
rect 12622 13087 12678 13096
rect 12714 13016 12770 13025
rect 12532 12980 12584 12986
rect 12714 12951 12770 12960
rect 12532 12922 12584 12928
rect 12728 12850 12756 12951
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12452 12442 12480 12718
rect 12624 12708 12676 12714
rect 12544 12668 12624 12696
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12256 12164 12308 12170
rect 12256 12106 12308 12112
rect 12256 11688 12308 11694
rect 12256 11630 12308 11636
rect 12164 11620 12216 11626
rect 12164 11562 12216 11568
rect 12268 11286 12296 11630
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12256 11280 12308 11286
rect 12256 11222 12308 11228
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 12084 10742 12112 11154
rect 12164 11008 12216 11014
rect 12164 10950 12216 10956
rect 12254 10976 12310 10985
rect 12176 10810 12204 10950
rect 12254 10911 12310 10920
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12072 10736 12124 10742
rect 12072 10678 12124 10684
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 11978 8664 12034 8673
rect 11978 8599 12034 8608
rect 11888 8356 11940 8362
rect 11888 8298 11940 8304
rect 11888 7744 11940 7750
rect 11888 7686 11940 7692
rect 11900 6225 11928 7686
rect 11980 6248 12032 6254
rect 11886 6216 11942 6225
rect 11980 6190 12032 6196
rect 11886 6151 11942 6160
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 11900 5370 11928 5714
rect 11992 5710 12020 6190
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 11888 5364 11940 5370
rect 11888 5306 11940 5312
rect 11888 5092 11940 5098
rect 11888 5034 11940 5040
rect 11532 4576 11744 4604
rect 11900 4593 11928 5034
rect 11886 4584 11942 4593
rect 11428 4140 11480 4146
rect 11428 4082 11480 4088
rect 11336 4072 11388 4078
rect 11336 4014 11388 4020
rect 11428 3936 11480 3942
rect 11426 3904 11428 3913
rect 11480 3904 11482 3913
rect 11426 3839 11482 3848
rect 11532 3754 11560 4576
rect 11886 4519 11942 4528
rect 11900 4486 11928 4519
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 11886 4312 11942 4321
rect 11886 4247 11942 4256
rect 11610 4040 11666 4049
rect 11610 3975 11666 3984
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 11164 3726 11560 3754
rect 10784 2576 10836 2582
rect 10784 2518 10836 2524
rect 10876 2576 10928 2582
rect 10876 2518 10928 2524
rect 10980 2417 11008 3674
rect 11058 3224 11114 3233
rect 11058 3159 11060 3168
rect 11112 3159 11114 3168
rect 11060 3130 11112 3136
rect 11060 2916 11112 2922
rect 11060 2858 11112 2864
rect 11072 2650 11100 2858
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 10966 2408 11022 2417
rect 10966 2343 11022 2352
rect 10612 1414 10732 1442
rect 10612 480 10640 1414
rect 11164 480 11192 3726
rect 11624 3670 11652 3975
rect 11612 3664 11664 3670
rect 11612 3606 11664 3612
rect 11624 3194 11652 3606
rect 11704 3528 11756 3534
rect 11704 3470 11756 3476
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 11716 3126 11744 3470
rect 11704 3120 11756 3126
rect 11704 3062 11756 3068
rect 11704 2576 11756 2582
rect 11704 2518 11756 2524
rect 11716 480 11744 2518
rect 11900 610 11928 4247
rect 11992 2990 12020 5646
rect 12084 3641 12112 9318
rect 12268 9217 12296 10911
rect 12452 10554 12480 11290
rect 12360 10526 12480 10554
rect 12360 10282 12388 10526
rect 12360 10254 12480 10282
rect 12452 9602 12480 10254
rect 12544 9738 12572 12668
rect 12624 12650 12676 12656
rect 12622 12608 12678 12617
rect 12622 12543 12678 12552
rect 12636 10130 12664 12543
rect 12728 12442 12756 12786
rect 12716 12436 12768 12442
rect 12716 12378 12768 12384
rect 12820 11354 12848 13110
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 12808 10736 12860 10742
rect 12808 10678 12860 10684
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12728 10305 12756 10406
rect 12714 10296 12770 10305
rect 12714 10231 12770 10240
rect 12624 10124 12676 10130
rect 12624 10066 12676 10072
rect 12820 9994 12848 10678
rect 12912 10554 12940 13824
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 13004 11150 13032 12038
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 12912 10526 13032 10554
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 12912 10266 12940 10406
rect 12900 10260 12952 10266
rect 12900 10202 12952 10208
rect 12900 10124 12952 10130
rect 12900 10066 12952 10072
rect 12808 9988 12860 9994
rect 12808 9930 12860 9936
rect 12544 9710 12756 9738
rect 12820 9722 12848 9930
rect 12728 9625 12756 9710
rect 12808 9716 12860 9722
rect 12808 9658 12860 9664
rect 12714 9616 12770 9625
rect 12452 9574 12572 9602
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 12452 9330 12480 9454
rect 12360 9302 12480 9330
rect 12254 9208 12310 9217
rect 12254 9143 12310 9152
rect 12268 7954 12296 9143
rect 12360 8090 12388 9302
rect 12544 8537 12572 9574
rect 12912 9602 12940 10066
rect 12714 9551 12770 9560
rect 12820 9574 12940 9602
rect 12820 8566 12848 9574
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12912 8974 12940 9318
rect 12900 8968 12952 8974
rect 12900 8910 12952 8916
rect 12912 8634 12940 8910
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 12808 8560 12860 8566
rect 12530 8528 12586 8537
rect 12808 8502 12860 8508
rect 12530 8463 12586 8472
rect 12820 8362 12848 8502
rect 12808 8356 12860 8362
rect 12808 8298 12860 8304
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12256 7948 12308 7954
rect 12256 7890 12308 7896
rect 12164 7472 12216 7478
rect 12162 7440 12164 7449
rect 12216 7440 12218 7449
rect 12162 7375 12218 7384
rect 12268 7002 12296 7890
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 12360 7585 12388 7822
rect 12346 7576 12402 7585
rect 12346 7511 12348 7520
rect 12400 7511 12402 7520
rect 12624 7540 12676 7546
rect 12348 7482 12400 7488
rect 12624 7482 12676 7488
rect 12360 7451 12388 7482
rect 12452 7342 12480 7373
rect 12440 7336 12492 7342
rect 12438 7304 12440 7313
rect 12492 7304 12494 7313
rect 12438 7239 12494 7248
rect 12452 7002 12480 7239
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 12440 6996 12492 7002
rect 12440 6938 12492 6944
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12176 5574 12204 6054
rect 12348 5840 12400 5846
rect 12348 5782 12400 5788
rect 12360 5624 12388 5782
rect 12544 5624 12572 7142
rect 12360 5596 12572 5624
rect 12164 5568 12216 5574
rect 12164 5510 12216 5516
rect 12176 4622 12204 5510
rect 12438 5128 12494 5137
rect 12438 5063 12494 5072
rect 12452 5030 12480 5063
rect 12348 5024 12400 5030
rect 12348 4966 12400 4972
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12360 4826 12388 4966
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12164 4616 12216 4622
rect 12164 4558 12216 4564
rect 12176 4282 12204 4558
rect 12256 4548 12308 4554
rect 12256 4490 12308 4496
rect 12164 4276 12216 4282
rect 12164 4218 12216 4224
rect 12070 3632 12126 3641
rect 12268 3602 12296 4490
rect 12636 4146 12664 7482
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12728 5778 12756 7346
rect 12716 5772 12768 5778
rect 12716 5714 12768 5720
rect 12728 4826 12756 5714
rect 12820 4978 12848 8298
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12912 7478 12940 8230
rect 12900 7472 12952 7478
rect 12900 7414 12952 7420
rect 12912 7206 12940 7414
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12900 6656 12952 6662
rect 12900 6598 12952 6604
rect 12912 5302 12940 6598
rect 13004 5370 13032 10526
rect 13096 9738 13124 17206
rect 13188 12458 13216 24006
rect 13280 22574 13308 24618
rect 13544 24336 13596 24342
rect 13542 24304 13544 24313
rect 13596 24304 13598 24313
rect 13452 24268 13504 24274
rect 13598 24262 13676 24290
rect 13542 24239 13598 24248
rect 13452 24210 13504 24216
rect 13360 24200 13412 24206
rect 13464 24177 13492 24210
rect 13360 24142 13412 24148
rect 13450 24168 13506 24177
rect 13372 23730 13400 24142
rect 13450 24103 13506 24112
rect 13544 24132 13596 24138
rect 13464 23798 13492 24103
rect 13544 24074 13596 24080
rect 13452 23792 13504 23798
rect 13452 23734 13504 23740
rect 13360 23724 13412 23730
rect 13360 23666 13412 23672
rect 13372 23118 13400 23666
rect 13556 23254 13584 24074
rect 13648 23798 13676 24262
rect 13636 23792 13688 23798
rect 13636 23734 13688 23740
rect 13634 23352 13690 23361
rect 13634 23287 13636 23296
rect 13688 23287 13690 23296
rect 13636 23258 13688 23264
rect 13544 23248 13596 23254
rect 13544 23190 13596 23196
rect 13360 23112 13412 23118
rect 13360 23054 13412 23060
rect 13268 22568 13320 22574
rect 13268 22510 13320 22516
rect 13372 22506 13400 23054
rect 13556 22794 13584 23190
rect 13636 23112 13688 23118
rect 13636 23054 13688 23060
rect 13464 22766 13584 22794
rect 13648 22778 13676 23054
rect 13636 22772 13688 22778
rect 13360 22500 13412 22506
rect 13360 22442 13412 22448
rect 13268 22228 13320 22234
rect 13268 22170 13320 22176
rect 13280 17270 13308 22170
rect 13372 21350 13400 22442
rect 13464 22234 13492 22766
rect 13636 22714 13688 22720
rect 13544 22636 13596 22642
rect 13544 22578 13596 22584
rect 13556 22438 13584 22578
rect 13544 22432 13596 22438
rect 13544 22374 13596 22380
rect 13452 22228 13504 22234
rect 13452 22170 13504 22176
rect 13450 22128 13506 22137
rect 13450 22063 13506 22072
rect 13360 21344 13412 21350
rect 13360 21286 13412 21292
rect 13360 20800 13412 20806
rect 13360 20742 13412 20748
rect 13372 19417 13400 20742
rect 13358 19408 13414 19417
rect 13358 19343 13414 19352
rect 13358 18456 13414 18465
rect 13358 18391 13360 18400
rect 13412 18391 13414 18400
rect 13360 18362 13412 18368
rect 13360 17536 13412 17542
rect 13360 17478 13412 17484
rect 13268 17264 13320 17270
rect 13268 17206 13320 17212
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 13280 14074 13308 14554
rect 13268 14068 13320 14074
rect 13268 14010 13320 14016
rect 13266 13968 13322 13977
rect 13266 13903 13322 13912
rect 13280 13682 13308 13903
rect 13372 13841 13400 17478
rect 13358 13832 13414 13841
rect 13358 13767 13414 13776
rect 13280 13654 13400 13682
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 13280 12850 13308 13466
rect 13268 12844 13320 12850
rect 13268 12786 13320 12792
rect 13266 12744 13322 12753
rect 13266 12679 13322 12688
rect 13280 12646 13308 12679
rect 13268 12640 13320 12646
rect 13268 12582 13320 12588
rect 13188 12430 13308 12458
rect 13176 11620 13228 11626
rect 13176 11562 13228 11568
rect 13188 11354 13216 11562
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 13188 11014 13216 11290
rect 13176 11008 13228 11014
rect 13176 10950 13228 10956
rect 13188 10674 13216 10950
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 13096 9710 13216 9738
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 13096 8838 13124 9522
rect 13188 8945 13216 9710
rect 13174 8936 13230 8945
rect 13174 8871 13230 8880
rect 13084 8832 13136 8838
rect 13084 8774 13136 8780
rect 13084 8492 13136 8498
rect 13084 8434 13136 8440
rect 13096 8090 13124 8434
rect 13084 8084 13136 8090
rect 13084 8026 13136 8032
rect 13188 8022 13216 8871
rect 13176 8016 13228 8022
rect 13176 7958 13228 7964
rect 13084 7812 13136 7818
rect 13084 7754 13136 7760
rect 13096 7290 13124 7754
rect 13188 7410 13216 7958
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 13096 7262 13216 7290
rect 13084 6996 13136 7002
rect 13084 6938 13136 6944
rect 13096 5914 13124 6938
rect 13188 6882 13216 7262
rect 13280 7002 13308 12430
rect 13372 10169 13400 13654
rect 13464 12458 13492 22063
rect 13556 21010 13584 22374
rect 13648 22137 13676 22714
rect 13740 22273 13768 24908
rect 13726 22264 13782 22273
rect 13726 22199 13782 22208
rect 13634 22128 13690 22137
rect 13634 22063 13690 22072
rect 13728 22092 13780 22098
rect 13728 22034 13780 22040
rect 13636 21888 13688 21894
rect 13636 21830 13688 21836
rect 13544 21004 13596 21010
rect 13544 20946 13596 20952
rect 13556 20602 13584 20946
rect 13544 20596 13596 20602
rect 13544 20538 13596 20544
rect 13556 20074 13584 20538
rect 13648 20505 13676 21830
rect 13740 21690 13768 22034
rect 13728 21684 13780 21690
rect 13728 21626 13780 21632
rect 13832 21554 13860 25230
rect 13924 25158 13952 25298
rect 13912 25152 13964 25158
rect 13912 25094 13964 25100
rect 13924 24954 13952 25094
rect 13912 24948 13964 24954
rect 13912 24890 13964 24896
rect 14292 23905 14320 27520
rect 14648 25424 14700 25430
rect 14648 25366 14700 25372
rect 14660 24954 14688 25366
rect 14740 25152 14792 25158
rect 14740 25094 14792 25100
rect 14752 24993 14780 25094
rect 14738 24984 14794 24993
rect 14648 24948 14700 24954
rect 14738 24919 14794 24928
rect 14648 24890 14700 24896
rect 14844 24834 14872 27520
rect 15292 25152 15344 25158
rect 15292 25094 15344 25100
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14384 24806 14872 24834
rect 14924 24880 14976 24886
rect 14924 24822 14976 24828
rect 15106 24848 15162 24857
rect 14094 23896 14150 23905
rect 14094 23831 14150 23840
rect 14278 23896 14334 23905
rect 14278 23831 14334 23840
rect 13912 23520 13964 23526
rect 13912 23462 13964 23468
rect 13820 21548 13872 21554
rect 13740 21508 13820 21536
rect 13740 21146 13768 21508
rect 13820 21490 13872 21496
rect 13820 21344 13872 21350
rect 13820 21286 13872 21292
rect 13728 21140 13780 21146
rect 13728 21082 13780 21088
rect 13634 20496 13690 20505
rect 13634 20431 13690 20440
rect 13740 20262 13768 21082
rect 13728 20256 13780 20262
rect 13728 20198 13780 20204
rect 13832 20210 13860 21286
rect 13924 20369 13952 23462
rect 14108 23254 14136 23831
rect 14280 23792 14332 23798
rect 14280 23734 14332 23740
rect 14096 23248 14148 23254
rect 14096 23190 14148 23196
rect 14188 23180 14240 23186
rect 14188 23122 14240 23128
rect 14096 22024 14148 22030
rect 14096 21966 14148 21972
rect 14002 21856 14058 21865
rect 14002 21791 14058 21800
rect 13910 20360 13966 20369
rect 13910 20295 13966 20304
rect 13832 20182 13952 20210
rect 13556 20046 13768 20074
rect 13542 19952 13598 19961
rect 13542 19887 13544 19896
rect 13596 19887 13598 19896
rect 13544 19858 13596 19864
rect 13740 19394 13768 20046
rect 13740 19366 13860 19394
rect 13542 19272 13598 19281
rect 13542 19207 13598 19216
rect 13636 19236 13688 19242
rect 13556 18222 13584 19207
rect 13636 19178 13688 19184
rect 13544 18216 13596 18222
rect 13544 18158 13596 18164
rect 13544 18080 13596 18086
rect 13544 18022 13596 18028
rect 13556 17882 13584 18022
rect 13544 17876 13596 17882
rect 13544 17818 13596 17824
rect 13556 16794 13584 17818
rect 13648 17746 13676 19178
rect 13832 19174 13860 19366
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 13818 19000 13874 19009
rect 13924 18986 13952 20182
rect 13874 18958 13952 18986
rect 13818 18935 13874 18944
rect 13728 18692 13780 18698
rect 13728 18634 13780 18640
rect 13740 17814 13768 18634
rect 13728 17808 13780 17814
rect 13728 17750 13780 17756
rect 13636 17740 13688 17746
rect 13636 17682 13688 17688
rect 13832 17660 13860 18935
rect 14016 17898 14044 21791
rect 14108 21690 14136 21966
rect 14096 21684 14148 21690
rect 14096 21626 14148 21632
rect 14096 21412 14148 21418
rect 14096 21354 14148 21360
rect 14108 21146 14136 21354
rect 14096 21140 14148 21146
rect 14096 21082 14148 21088
rect 14200 21078 14228 23122
rect 14188 21072 14240 21078
rect 14188 21014 14240 21020
rect 14096 21004 14148 21010
rect 14096 20946 14148 20952
rect 13634 17640 13690 17649
rect 13634 17575 13636 17584
rect 13688 17575 13690 17584
rect 13740 17632 13860 17660
rect 13924 17870 14044 17898
rect 13636 17546 13688 17552
rect 13634 17368 13690 17377
rect 13634 17303 13690 17312
rect 13648 16969 13676 17303
rect 13634 16960 13690 16969
rect 13634 16895 13690 16904
rect 13544 16788 13596 16794
rect 13544 16730 13596 16736
rect 13740 16590 13768 17632
rect 13820 17536 13872 17542
rect 13820 17478 13872 17484
rect 13832 17202 13860 17478
rect 13820 17196 13872 17202
rect 13820 17138 13872 17144
rect 13728 16584 13780 16590
rect 13728 16526 13780 16532
rect 13740 16250 13768 16526
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13832 16182 13860 17138
rect 13820 16176 13872 16182
rect 13820 16118 13872 16124
rect 13820 16040 13872 16046
rect 13818 16008 13820 16017
rect 13872 16008 13874 16017
rect 13818 15943 13874 15952
rect 13924 15892 13952 17870
rect 14004 17808 14056 17814
rect 14004 17750 14056 17756
rect 14016 16794 14044 17750
rect 14004 16788 14056 16794
rect 14004 16730 14056 16736
rect 14108 16425 14136 20946
rect 14200 20874 14228 21014
rect 14188 20868 14240 20874
rect 14188 20810 14240 20816
rect 14186 20496 14242 20505
rect 14186 20431 14242 20440
rect 14200 20330 14228 20431
rect 14188 20324 14240 20330
rect 14188 20266 14240 20272
rect 14200 20058 14228 20266
rect 14188 20052 14240 20058
rect 14188 19994 14240 20000
rect 14186 19680 14242 19689
rect 14186 19615 14242 19624
rect 14200 18766 14228 19615
rect 14188 18760 14240 18766
rect 14188 18702 14240 18708
rect 14186 17504 14242 17513
rect 14186 17439 14242 17448
rect 14200 17338 14228 17439
rect 14188 17332 14240 17338
rect 14188 17274 14240 17280
rect 14186 17096 14242 17105
rect 14186 17031 14242 17040
rect 14200 16794 14228 17031
rect 14188 16788 14240 16794
rect 14188 16730 14240 16736
rect 14094 16416 14150 16425
rect 14094 16351 14150 16360
rect 14096 16176 14148 16182
rect 14096 16118 14148 16124
rect 14186 16144 14242 16153
rect 13832 15864 13952 15892
rect 13728 15632 13780 15638
rect 13728 15574 13780 15580
rect 13636 15496 13688 15502
rect 13636 15438 13688 15444
rect 13542 14920 13598 14929
rect 13542 14855 13598 14864
rect 13556 14618 13584 14855
rect 13648 14822 13676 15438
rect 13740 14822 13768 15574
rect 13832 15094 13860 15864
rect 13820 15088 13872 15094
rect 13820 15030 13872 15036
rect 13636 14816 13688 14822
rect 13636 14758 13688 14764
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13544 14340 13596 14346
rect 13544 14282 13596 14288
rect 13556 13462 13584 14282
rect 13544 13456 13596 13462
rect 13544 13398 13596 13404
rect 13556 12782 13584 13398
rect 13544 12776 13596 12782
rect 13544 12718 13596 12724
rect 13556 12617 13584 12718
rect 13542 12608 13598 12617
rect 13542 12543 13598 12552
rect 13464 12430 13584 12458
rect 13450 10840 13506 10849
rect 13450 10775 13452 10784
rect 13504 10775 13506 10784
rect 13452 10746 13504 10752
rect 13464 10538 13492 10746
rect 13452 10532 13504 10538
rect 13452 10474 13504 10480
rect 13358 10160 13414 10169
rect 13358 10095 13414 10104
rect 13452 9920 13504 9926
rect 13452 9862 13504 9868
rect 13464 9518 13492 9862
rect 13452 9512 13504 9518
rect 13358 9480 13414 9489
rect 13452 9454 13504 9460
rect 13358 9415 13414 9424
rect 13268 6996 13320 7002
rect 13268 6938 13320 6944
rect 13188 6854 13308 6882
rect 13176 6792 13228 6798
rect 13176 6734 13228 6740
rect 13188 6254 13216 6734
rect 13176 6248 13228 6254
rect 13176 6190 13228 6196
rect 13280 5914 13308 6854
rect 13084 5908 13136 5914
rect 13084 5850 13136 5856
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13372 5817 13400 9415
rect 13452 8424 13504 8430
rect 13452 8366 13504 8372
rect 13464 7177 13492 8366
rect 13450 7168 13506 7177
rect 13450 7103 13506 7112
rect 13452 6112 13504 6118
rect 13452 6054 13504 6060
rect 13358 5808 13414 5817
rect 13176 5772 13228 5778
rect 13358 5743 13414 5752
rect 13176 5714 13228 5720
rect 12992 5364 13044 5370
rect 13044 5324 13124 5352
rect 12992 5306 13044 5312
rect 12900 5296 12952 5302
rect 12900 5238 12952 5244
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 13004 5098 13032 5170
rect 12992 5092 13044 5098
rect 12992 5034 13044 5040
rect 12820 4950 13032 4978
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12900 4752 12952 4758
rect 12900 4694 12952 4700
rect 12912 4214 12940 4694
rect 12900 4208 12952 4214
rect 12900 4150 12952 4156
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12532 4072 12584 4078
rect 12532 4014 12584 4020
rect 12544 3738 12572 4014
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 12070 3567 12126 3576
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 12532 3460 12584 3466
rect 12532 3402 12584 3408
rect 12544 3346 12572 3402
rect 12360 3318 12572 3346
rect 11980 2984 12032 2990
rect 11980 2926 12032 2932
rect 12360 2650 12388 3318
rect 12348 2644 12400 2650
rect 12348 2586 12400 2592
rect 12636 2553 12664 3878
rect 12806 3768 12862 3777
rect 12806 3703 12808 3712
rect 12860 3703 12862 3712
rect 12808 3674 12860 3680
rect 12808 3392 12860 3398
rect 12808 3334 12860 3340
rect 12716 2916 12768 2922
rect 12716 2858 12768 2864
rect 12622 2544 12678 2553
rect 12622 2479 12678 2488
rect 12072 2440 12124 2446
rect 12070 2408 12072 2417
rect 12728 2417 12756 2858
rect 12124 2408 12126 2417
rect 12070 2343 12126 2352
rect 12714 2408 12770 2417
rect 12714 2343 12770 2352
rect 11888 604 11940 610
rect 11888 546 11940 552
rect 12256 604 12308 610
rect 12256 546 12308 552
rect 12268 480 12296 546
rect 12820 480 12848 3334
rect 13004 1465 13032 4950
rect 13096 2281 13124 5324
rect 13188 3738 13216 5714
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 13268 3596 13320 3602
rect 13268 3538 13320 3544
rect 13280 3505 13308 3538
rect 13266 3496 13322 3505
rect 13266 3431 13322 3440
rect 13082 2272 13138 2281
rect 13082 2207 13138 2216
rect 12990 1456 13046 1465
rect 12990 1391 13046 1400
rect 13372 480 13400 5743
rect 13464 5098 13492 6054
rect 13452 5092 13504 5098
rect 13452 5034 13504 5040
rect 13556 4078 13584 12430
rect 13648 11898 13676 14758
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13740 12594 13768 14010
rect 13832 13462 13860 15030
rect 14108 14958 14136 16118
rect 14186 16079 14242 16088
rect 13912 14952 13964 14958
rect 13912 14894 13964 14900
rect 14096 14952 14148 14958
rect 14096 14894 14148 14900
rect 13924 13841 13952 14894
rect 14096 14816 14148 14822
rect 14094 14784 14096 14793
rect 14148 14784 14150 14793
rect 14094 14719 14150 14728
rect 14004 14272 14056 14278
rect 14004 14214 14056 14220
rect 14096 14272 14148 14278
rect 14096 14214 14148 14220
rect 13910 13832 13966 13841
rect 14016 13802 14044 14214
rect 13910 13767 13912 13776
rect 13964 13767 13966 13776
rect 14004 13796 14056 13802
rect 13912 13738 13964 13744
rect 14004 13738 14056 13744
rect 13924 13707 13952 13738
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 13924 12617 13952 13330
rect 13910 12608 13966 12617
rect 13740 12566 13860 12594
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13740 12073 13768 12106
rect 13726 12064 13782 12073
rect 13726 11999 13782 12008
rect 13636 11892 13688 11898
rect 13636 11834 13688 11840
rect 13634 11792 13690 11801
rect 13634 11727 13690 11736
rect 13648 8430 13676 11727
rect 13832 10826 13860 12566
rect 13910 12543 13966 12552
rect 13910 12472 13966 12481
rect 13910 12407 13966 12416
rect 13924 11694 13952 12407
rect 14016 12306 14044 13738
rect 14108 12753 14136 14214
rect 14200 13734 14228 16079
rect 14292 14385 14320 23734
rect 14384 16697 14412 24806
rect 14740 24608 14792 24614
rect 14646 24576 14702 24585
rect 14740 24550 14792 24556
rect 14646 24511 14702 24520
rect 14554 23760 14610 23769
rect 14660 23746 14688 24511
rect 14752 23769 14780 24550
rect 14936 24052 14964 24822
rect 15106 24783 15162 24792
rect 15120 24750 15148 24783
rect 15108 24744 15160 24750
rect 15108 24686 15160 24692
rect 15304 24154 15332 25094
rect 15396 24698 15424 27520
rect 15672 25486 15976 25514
rect 15672 25430 15700 25486
rect 15948 25430 15976 25486
rect 15660 25424 15712 25430
rect 15660 25366 15712 25372
rect 15936 25424 15988 25430
rect 15936 25366 15988 25372
rect 15752 25356 15804 25362
rect 15804 25316 15884 25344
rect 15752 25298 15804 25304
rect 15476 25152 15528 25158
rect 15476 25094 15528 25100
rect 15488 24886 15516 25094
rect 15476 24880 15528 24886
rect 15476 24822 15528 24828
rect 15752 24744 15804 24750
rect 15396 24670 15700 24698
rect 15752 24686 15804 24692
rect 15476 24268 15528 24274
rect 15476 24210 15528 24216
rect 15304 24126 15424 24154
rect 14844 24024 14964 24052
rect 15292 24064 15344 24070
rect 14610 23718 14688 23746
rect 14554 23695 14610 23704
rect 14556 23656 14608 23662
rect 14556 23598 14608 23604
rect 14568 22982 14596 23598
rect 14556 22976 14608 22982
rect 14554 22944 14556 22953
rect 14608 22944 14610 22953
rect 14554 22879 14610 22888
rect 14660 22642 14688 23718
rect 14738 23760 14794 23769
rect 14738 23695 14794 23704
rect 14740 23044 14792 23050
rect 14740 22986 14792 22992
rect 14648 22636 14700 22642
rect 14648 22578 14700 22584
rect 14464 22568 14516 22574
rect 14464 22510 14516 22516
rect 14476 20505 14504 22510
rect 14554 22400 14610 22409
rect 14554 22335 14610 22344
rect 14462 20496 14518 20505
rect 14462 20431 14518 20440
rect 14464 17672 14516 17678
rect 14464 17614 14516 17620
rect 14476 17066 14504 17614
rect 14464 17060 14516 17066
rect 14464 17002 14516 17008
rect 14370 16688 14426 16697
rect 14370 16623 14426 16632
rect 14370 16552 14426 16561
rect 14370 16487 14426 16496
rect 14384 15706 14412 16487
rect 14372 15700 14424 15706
rect 14372 15642 14424 15648
rect 14384 14890 14412 15642
rect 14372 14884 14424 14890
rect 14372 14826 14424 14832
rect 14278 14376 14334 14385
rect 14278 14311 14334 14320
rect 14384 14074 14412 14826
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 14568 13954 14596 22335
rect 14648 22092 14700 22098
rect 14648 22034 14700 22040
rect 14660 21350 14688 22034
rect 14648 21344 14700 21350
rect 14648 21286 14700 21292
rect 14660 19514 14688 21286
rect 14752 21146 14780 22986
rect 14844 22778 14872 24024
rect 15292 24006 15344 24012
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15106 23624 15162 23633
rect 15106 23559 15162 23568
rect 15120 23526 15148 23559
rect 15108 23520 15160 23526
rect 15304 23497 15332 24006
rect 15108 23462 15160 23468
rect 15290 23488 15346 23497
rect 15290 23423 15346 23432
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 14832 22772 14884 22778
rect 14832 22714 14884 22720
rect 15396 22642 15424 24126
rect 15488 23866 15516 24210
rect 15568 24200 15620 24206
rect 15568 24142 15620 24148
rect 15476 23860 15528 23866
rect 15476 23802 15528 23808
rect 15580 23361 15608 24142
rect 15566 23352 15622 23361
rect 15566 23287 15622 23296
rect 15568 23180 15620 23186
rect 15568 23122 15620 23128
rect 15476 23112 15528 23118
rect 15476 23054 15528 23060
rect 14924 22636 14976 22642
rect 15384 22636 15436 22642
rect 14924 22578 14976 22584
rect 15304 22596 15384 22624
rect 14936 21876 14964 22578
rect 14844 21848 14964 21876
rect 14740 21140 14792 21146
rect 14740 21082 14792 21088
rect 14752 20398 14780 21082
rect 14740 20392 14792 20398
rect 14740 20334 14792 20340
rect 14648 19508 14700 19514
rect 14648 19450 14700 19456
rect 14648 18760 14700 18766
rect 14648 18702 14700 18708
rect 14660 18086 14688 18702
rect 14740 18692 14792 18698
rect 14740 18634 14792 18640
rect 14752 18290 14780 18634
rect 14740 18284 14792 18290
rect 14740 18226 14792 18232
rect 14648 18080 14700 18086
rect 14648 18022 14700 18028
rect 14660 15858 14688 18022
rect 14752 17882 14780 18226
rect 14740 17876 14792 17882
rect 14740 17818 14792 17824
rect 14752 16522 14780 17818
rect 14740 16516 14792 16522
rect 14740 16458 14792 16464
rect 14752 16250 14780 16458
rect 14740 16244 14792 16250
rect 14740 16186 14792 16192
rect 14752 15978 14780 16186
rect 14740 15972 14792 15978
rect 14740 15914 14792 15920
rect 14660 15830 14780 15858
rect 14648 15360 14700 15366
rect 14648 15302 14700 15308
rect 14660 14278 14688 15302
rect 14648 14272 14700 14278
rect 14648 14214 14700 14220
rect 14752 14090 14780 15830
rect 14476 13926 14596 13954
rect 14660 14062 14780 14090
rect 14188 13728 14240 13734
rect 14476 13682 14504 13926
rect 14188 13670 14240 13676
rect 14384 13654 14504 13682
rect 14188 13320 14240 13326
rect 14188 13262 14240 13268
rect 14094 12744 14150 12753
rect 14094 12679 14150 12688
rect 14094 12608 14150 12617
rect 14094 12543 14150 12552
rect 14004 12300 14056 12306
rect 14004 12242 14056 12248
rect 14108 12186 14136 12543
rect 14016 12158 14136 12186
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 14016 11370 14044 12158
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 14108 11830 14136 12038
rect 14096 11824 14148 11830
rect 14096 11766 14148 11772
rect 14016 11342 14136 11370
rect 14004 11280 14056 11286
rect 14002 11248 14004 11257
rect 14056 11248 14058 11257
rect 14002 11183 14058 11192
rect 13832 10798 13952 10826
rect 13924 10554 13952 10798
rect 14016 10656 14044 11183
rect 14108 10996 14136 11342
rect 14200 11257 14228 13262
rect 14384 12288 14412 13654
rect 14464 13456 14516 13462
rect 14464 13398 14516 13404
rect 14292 12260 14412 12288
rect 14186 11248 14242 11257
rect 14186 11183 14242 11192
rect 14188 11008 14240 11014
rect 14108 10968 14188 10996
rect 14188 10950 14240 10956
rect 14096 10668 14148 10674
rect 14016 10628 14096 10656
rect 14096 10610 14148 10616
rect 13924 10526 14136 10554
rect 13726 10432 13782 10441
rect 13726 10367 13782 10376
rect 13740 9897 13768 10367
rect 14004 10260 14056 10266
rect 14004 10202 14056 10208
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13726 9888 13782 9897
rect 13726 9823 13782 9832
rect 13832 9761 13860 10066
rect 13910 9888 13966 9897
rect 13910 9823 13966 9832
rect 13818 9752 13874 9761
rect 13818 9687 13820 9696
rect 13872 9687 13874 9696
rect 13820 9658 13872 9664
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 13740 9178 13768 9590
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 13636 8424 13688 8430
rect 13636 8366 13688 8372
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 13648 7546 13676 7890
rect 13740 7886 13768 8774
rect 13832 8090 13860 9318
rect 13924 9160 13952 9823
rect 14016 9722 14044 10202
rect 14004 9716 14056 9722
rect 14004 9658 14056 9664
rect 13924 9132 14044 9160
rect 13912 9036 13964 9042
rect 13912 8978 13964 8984
rect 13924 8634 13952 8978
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 13912 8424 13964 8430
rect 13910 8392 13912 8401
rect 13964 8392 13966 8401
rect 13910 8327 13966 8336
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13910 7984 13966 7993
rect 13910 7919 13912 7928
rect 13964 7919 13966 7928
rect 13912 7890 13964 7896
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13820 7812 13872 7818
rect 13820 7754 13872 7760
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13832 7478 13860 7754
rect 13924 7546 13952 7890
rect 13912 7540 13964 7546
rect 13912 7482 13964 7488
rect 13820 7472 13872 7478
rect 13820 7414 13872 7420
rect 13832 6934 13860 7414
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 13728 6928 13780 6934
rect 13728 6870 13780 6876
rect 13820 6928 13872 6934
rect 13820 6870 13872 6876
rect 13740 6474 13768 6870
rect 13648 6458 13860 6474
rect 13648 6452 13872 6458
rect 13648 6446 13820 6452
rect 13648 4826 13676 6446
rect 13820 6394 13872 6400
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13740 5234 13768 5850
rect 13818 5536 13874 5545
rect 13818 5471 13874 5480
rect 13832 5370 13860 5471
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 13452 3936 13504 3942
rect 13740 3890 13768 5170
rect 13832 5166 13860 5306
rect 13924 5273 13952 7346
rect 13910 5264 13966 5273
rect 13910 5199 13966 5208
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 14016 4826 14044 9132
rect 14108 8022 14136 10526
rect 14200 10062 14228 10950
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14200 8974 14228 9998
rect 14292 9058 14320 12260
rect 14476 12220 14504 13398
rect 14384 12192 14504 12220
rect 14384 9466 14412 12192
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14476 9722 14504 12038
rect 14556 11688 14608 11694
rect 14556 11630 14608 11636
rect 14568 11286 14596 11630
rect 14556 11280 14608 11286
rect 14556 11222 14608 11228
rect 14556 10804 14608 10810
rect 14556 10746 14608 10752
rect 14568 10674 14596 10746
rect 14556 10668 14608 10674
rect 14556 10610 14608 10616
rect 14464 9716 14516 9722
rect 14464 9658 14516 9664
rect 14568 9586 14596 10610
rect 14660 10198 14688 14062
rect 14738 13424 14794 13433
rect 14738 13359 14794 13368
rect 14752 12986 14780 13359
rect 14740 12980 14792 12986
rect 14740 12922 14792 12928
rect 14740 12300 14792 12306
rect 14740 12242 14792 12248
rect 14752 11558 14780 12242
rect 14740 11552 14792 11558
rect 14740 11494 14792 11500
rect 14648 10192 14700 10198
rect 14646 10160 14648 10169
rect 14700 10160 14702 10169
rect 14646 10095 14702 10104
rect 14648 9920 14700 9926
rect 14648 9862 14700 9868
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 14384 9438 14596 9466
rect 14292 9030 14412 9058
rect 14188 8968 14240 8974
rect 14188 8910 14240 8916
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 14188 8832 14240 8838
rect 14188 8774 14240 8780
rect 14096 8016 14148 8022
rect 14096 7958 14148 7964
rect 14096 7880 14148 7886
rect 14096 7822 14148 7828
rect 14108 7002 14136 7822
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 14004 4820 14056 4826
rect 14004 4762 14056 4768
rect 13820 4684 13872 4690
rect 13820 4626 13872 4632
rect 13832 3942 13860 4626
rect 13912 4480 13964 4486
rect 13912 4422 13964 4428
rect 13452 3878 13504 3884
rect 13464 3233 13492 3878
rect 13648 3862 13768 3890
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13648 3398 13676 3862
rect 13924 3754 13952 4422
rect 14016 4282 14044 4762
rect 14108 4593 14136 6734
rect 14094 4584 14150 4593
rect 14094 4519 14150 4528
rect 14004 4276 14056 4282
rect 14004 4218 14056 4224
rect 14002 4040 14058 4049
rect 14002 3975 14058 3984
rect 14096 4004 14148 4010
rect 14016 3942 14044 3975
rect 14096 3946 14148 3952
rect 14004 3936 14056 3942
rect 14108 3913 14136 3946
rect 14004 3878 14056 3884
rect 14094 3904 14150 3913
rect 14094 3839 14150 3848
rect 13740 3738 13952 3754
rect 13728 3732 13952 3738
rect 13780 3726 13952 3732
rect 13728 3674 13780 3680
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13450 3224 13506 3233
rect 13450 3159 13506 3168
rect 14002 3224 14058 3233
rect 14002 3159 14058 3168
rect 13912 3120 13964 3126
rect 13450 3088 13506 3097
rect 13912 3062 13964 3068
rect 13450 3023 13506 3032
rect 13464 1193 13492 3023
rect 13924 2961 13952 3062
rect 13910 2952 13966 2961
rect 13910 2887 13966 2896
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 13450 1184 13506 1193
rect 13450 1119 13506 1128
rect 13924 480 13952 2790
rect 14016 1737 14044 3159
rect 14002 1728 14058 1737
rect 14002 1663 14058 1672
rect 3146 368 3202 377
rect 3146 303 3202 312
rect 3422 0 3478 480
rect 3974 0 4030 480
rect 4526 0 4582 480
rect 5078 0 5134 480
rect 5630 0 5686 480
rect 6182 0 6238 480
rect 6734 0 6790 480
rect 7286 0 7342 480
rect 7838 0 7894 480
rect 8390 0 8446 480
rect 8942 0 8998 480
rect 9494 0 9550 480
rect 10046 0 10102 480
rect 10598 0 10654 480
rect 11150 0 11206 480
rect 11702 0 11758 480
rect 12254 0 12310 480
rect 12806 0 12862 480
rect 13358 0 13414 480
rect 13910 0 13966 480
rect 14200 105 14228 8774
rect 14292 7410 14320 8910
rect 14384 8242 14412 9030
rect 14464 8900 14516 8906
rect 14464 8842 14516 8848
rect 14476 8362 14504 8842
rect 14464 8356 14516 8362
rect 14464 8298 14516 8304
rect 14384 8214 14504 8242
rect 14370 8120 14426 8129
rect 14476 8090 14504 8214
rect 14370 8055 14426 8064
rect 14464 8084 14516 8090
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14278 7304 14334 7313
rect 14278 7239 14334 7248
rect 14292 7206 14320 7239
rect 14280 7200 14332 7206
rect 14280 7142 14332 7148
rect 14384 7018 14412 8055
rect 14464 8026 14516 8032
rect 14464 7744 14516 7750
rect 14464 7686 14516 7692
rect 14476 7449 14504 7686
rect 14462 7440 14518 7449
rect 14462 7375 14464 7384
rect 14516 7375 14518 7384
rect 14464 7346 14516 7352
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 14292 6990 14412 7018
rect 14292 5370 14320 6990
rect 14372 6112 14424 6118
rect 14372 6054 14424 6060
rect 14280 5364 14332 5370
rect 14280 5306 14332 5312
rect 14280 5092 14332 5098
rect 14280 5034 14332 5040
rect 14292 2854 14320 5034
rect 14384 4078 14412 6054
rect 14476 4214 14504 7142
rect 14568 4978 14596 9438
rect 14660 9382 14688 9862
rect 14648 9376 14700 9382
rect 14648 9318 14700 9324
rect 14752 9194 14780 11494
rect 14660 9166 14780 9194
rect 14660 7732 14688 9166
rect 14740 9104 14792 9110
rect 14740 9046 14792 9052
rect 14752 8809 14780 9046
rect 14738 8800 14794 8809
rect 14738 8735 14794 8744
rect 14738 8664 14794 8673
rect 14738 8599 14794 8608
rect 14752 7857 14780 8599
rect 14738 7848 14794 7857
rect 14738 7783 14794 7792
rect 14660 7704 14780 7732
rect 14648 6928 14700 6934
rect 14648 6870 14700 6876
rect 14660 5098 14688 6870
rect 14752 6225 14780 7704
rect 14844 6934 14872 21848
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14924 21548 14976 21554
rect 14924 21490 14976 21496
rect 14936 20942 14964 21490
rect 14924 20936 14976 20942
rect 14924 20878 14976 20884
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15304 20602 15332 22596
rect 15384 22578 15436 22584
rect 15488 21962 15516 23054
rect 15580 22778 15608 23122
rect 15568 22772 15620 22778
rect 15568 22714 15620 22720
rect 15566 22672 15622 22681
rect 15566 22607 15622 22616
rect 15580 22574 15608 22607
rect 15568 22568 15620 22574
rect 15568 22510 15620 22516
rect 15580 22234 15608 22510
rect 15568 22228 15620 22234
rect 15568 22170 15620 22176
rect 15568 22024 15620 22030
rect 15568 21966 15620 21972
rect 15476 21956 15528 21962
rect 15476 21898 15528 21904
rect 15384 21888 15436 21894
rect 15384 21830 15436 21836
rect 15396 21418 15424 21830
rect 15384 21412 15436 21418
rect 15384 21354 15436 21360
rect 15384 21072 15436 21078
rect 15384 21014 15436 21020
rect 15292 20596 15344 20602
rect 15292 20538 15344 20544
rect 15396 20466 15424 21014
rect 15488 20602 15516 21898
rect 15580 20806 15608 21966
rect 15568 20800 15620 20806
rect 15568 20742 15620 20748
rect 15580 20641 15608 20742
rect 15566 20632 15622 20641
rect 15476 20596 15528 20602
rect 15566 20567 15622 20576
rect 15476 20538 15528 20544
rect 14924 20460 14976 20466
rect 14924 20402 14976 20408
rect 15384 20460 15436 20466
rect 15384 20402 15436 20408
rect 14936 20058 14964 20402
rect 15292 20324 15344 20330
rect 15292 20266 15344 20272
rect 15200 20256 15252 20262
rect 15200 20198 15252 20204
rect 14924 20052 14976 20058
rect 14924 19994 14976 20000
rect 15212 19922 15240 20198
rect 15200 19916 15252 19922
rect 15200 19858 15252 19864
rect 15304 19786 15332 20266
rect 15384 20256 15436 20262
rect 15384 20198 15436 20204
rect 15292 19780 15344 19786
rect 15292 19722 15344 19728
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15106 19272 15162 19281
rect 15106 19207 15162 19216
rect 15120 18970 15148 19207
rect 15108 18964 15160 18970
rect 15108 18906 15160 18912
rect 15292 18624 15344 18630
rect 15292 18566 15344 18572
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15304 18034 15332 18566
rect 15120 18006 15332 18034
rect 15120 17814 15148 18006
rect 15290 17912 15346 17921
rect 15290 17847 15292 17856
rect 15344 17847 15346 17856
rect 15292 17818 15344 17824
rect 15108 17808 15160 17814
rect 15108 17750 15160 17756
rect 15292 17740 15344 17746
rect 15292 17682 15344 17688
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15198 17232 15254 17241
rect 15304 17218 15332 17682
rect 15254 17190 15332 17218
rect 15198 17167 15254 17176
rect 15108 17060 15160 17066
rect 15108 17002 15160 17008
rect 15120 16726 15148 17002
rect 15108 16720 15160 16726
rect 15108 16662 15160 16668
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15304 15858 15332 17190
rect 15396 16153 15424 20198
rect 15476 19916 15528 19922
rect 15476 19858 15528 19864
rect 15488 18290 15516 19858
rect 15672 19394 15700 24670
rect 15580 19366 15700 19394
rect 15476 18284 15528 18290
rect 15476 18226 15528 18232
rect 15476 17740 15528 17746
rect 15476 17682 15528 17688
rect 15488 17338 15516 17682
rect 15476 17332 15528 17338
rect 15476 17274 15528 17280
rect 15382 16144 15438 16153
rect 15382 16079 15438 16088
rect 15304 15830 15424 15858
rect 15292 15360 15344 15366
rect 15292 15302 15344 15308
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15304 14793 15332 15302
rect 15290 14784 15346 14793
rect 15290 14719 15346 14728
rect 15292 14272 15344 14278
rect 15292 14214 15344 14220
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15198 13832 15254 13841
rect 15198 13767 15254 13776
rect 15212 13394 15240 13767
rect 15200 13388 15252 13394
rect 15200 13330 15252 13336
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15304 12986 15332 14214
rect 15396 14006 15424 15830
rect 15488 14550 15516 17274
rect 15580 14958 15608 19366
rect 15660 19236 15712 19242
rect 15660 19178 15712 19184
rect 15672 18193 15700 19178
rect 15764 19174 15792 24686
rect 15856 24614 15884 25316
rect 15936 25288 15988 25294
rect 15936 25230 15988 25236
rect 15948 24750 15976 25230
rect 16040 24857 16068 27520
rect 16592 25974 16620 27520
rect 17144 26178 17172 27520
rect 17132 26172 17184 26178
rect 17132 26114 17184 26120
rect 16580 25968 16632 25974
rect 16580 25910 16632 25916
rect 17224 25968 17276 25974
rect 17224 25910 17276 25916
rect 17236 25498 17264 25910
rect 17788 25906 17816 27520
rect 17960 26376 18012 26382
rect 17960 26318 18012 26324
rect 17776 25900 17828 25906
rect 17776 25842 17828 25848
rect 17224 25492 17276 25498
rect 17224 25434 17276 25440
rect 16946 25392 17002 25401
rect 17314 25392 17370 25401
rect 16946 25327 17002 25336
rect 17132 25356 17184 25362
rect 16120 25288 16172 25294
rect 16120 25230 16172 25236
rect 16488 25288 16540 25294
rect 16488 25230 16540 25236
rect 16026 24848 16082 24857
rect 16026 24783 16082 24792
rect 15936 24744 15988 24750
rect 16132 24698 16160 25230
rect 16304 24880 16356 24886
rect 16304 24822 16356 24828
rect 15936 24686 15988 24692
rect 16040 24682 16160 24698
rect 16028 24676 16160 24682
rect 16080 24670 16160 24676
rect 16028 24618 16080 24624
rect 15844 24608 15896 24614
rect 15844 24550 15896 24556
rect 15936 24608 15988 24614
rect 15936 24550 15988 24556
rect 15856 22545 15884 24550
rect 15948 23254 15976 24550
rect 16040 24274 16068 24618
rect 16028 24268 16080 24274
rect 16028 24210 16080 24216
rect 16040 23866 16068 24210
rect 16212 24200 16264 24206
rect 16212 24142 16264 24148
rect 16028 23860 16080 23866
rect 16028 23802 16080 23808
rect 16120 23724 16172 23730
rect 16120 23666 16172 23672
rect 15936 23248 15988 23254
rect 15936 23190 15988 23196
rect 15936 23112 15988 23118
rect 15936 23054 15988 23060
rect 15842 22536 15898 22545
rect 15842 22471 15898 22480
rect 15948 21978 15976 23054
rect 16028 22772 16080 22778
rect 16028 22714 16080 22720
rect 15856 21962 15976 21978
rect 15844 21956 15976 21962
rect 15896 21950 15976 21956
rect 15844 21898 15896 21904
rect 15936 21888 15988 21894
rect 15936 21830 15988 21836
rect 15948 21706 15976 21830
rect 15856 21678 15976 21706
rect 15752 19168 15804 19174
rect 15752 19110 15804 19116
rect 15764 18601 15792 19110
rect 15856 18834 15884 21678
rect 16040 21570 16068 22714
rect 15948 21542 16068 21570
rect 16132 21554 16160 23666
rect 16224 23662 16252 24142
rect 16212 23656 16264 23662
rect 16212 23598 16264 23604
rect 16224 22982 16252 23598
rect 16212 22976 16264 22982
rect 16212 22918 16264 22924
rect 16120 21548 16172 21554
rect 15844 18828 15896 18834
rect 15844 18770 15896 18776
rect 15750 18592 15806 18601
rect 15750 18527 15806 18536
rect 15658 18184 15714 18193
rect 15658 18119 15714 18128
rect 15568 14952 15620 14958
rect 15568 14894 15620 14900
rect 15568 14816 15620 14822
rect 15568 14758 15620 14764
rect 15476 14544 15528 14550
rect 15476 14486 15528 14492
rect 15476 14340 15528 14346
rect 15476 14282 15528 14288
rect 15384 14000 15436 14006
rect 15384 13942 15436 13948
rect 15384 13456 15436 13462
rect 15384 13398 15436 13404
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15396 12850 15424 13398
rect 15384 12844 15436 12850
rect 15384 12786 15436 12792
rect 15488 12782 15516 14282
rect 15580 13569 15608 14758
rect 15566 13560 15622 13569
rect 15566 13495 15622 13504
rect 15580 13394 15608 13495
rect 15568 13388 15620 13394
rect 15568 13330 15620 13336
rect 15580 12918 15608 13330
rect 15672 12918 15700 18119
rect 15856 18086 15884 18770
rect 15844 18080 15896 18086
rect 15844 18022 15896 18028
rect 15948 17882 15976 21542
rect 16120 21490 16172 21496
rect 16224 21434 16252 22918
rect 16316 22438 16344 24822
rect 16500 23730 16528 25230
rect 16764 25152 16816 25158
rect 16764 25094 16816 25100
rect 16856 25152 16908 25158
rect 16856 25094 16908 25100
rect 16578 24848 16634 24857
rect 16578 24783 16634 24792
rect 16592 24018 16620 24783
rect 16776 24614 16804 25094
rect 16868 24954 16896 25094
rect 16856 24948 16908 24954
rect 16856 24890 16908 24896
rect 16856 24812 16908 24818
rect 16856 24754 16908 24760
rect 16672 24608 16724 24614
rect 16672 24550 16724 24556
rect 16764 24608 16816 24614
rect 16764 24550 16816 24556
rect 16684 24138 16712 24550
rect 16672 24132 16724 24138
rect 16672 24074 16724 24080
rect 16592 23990 16712 24018
rect 16488 23724 16540 23730
rect 16488 23666 16540 23672
rect 16396 23520 16448 23526
rect 16394 23488 16396 23497
rect 16448 23488 16450 23497
rect 16394 23423 16450 23432
rect 16394 23216 16450 23225
rect 16394 23151 16450 23160
rect 16408 22794 16436 23151
rect 16580 23112 16632 23118
rect 16580 23054 16632 23060
rect 16592 22794 16620 23054
rect 16408 22778 16620 22794
rect 16408 22772 16632 22778
rect 16408 22766 16580 22772
rect 16304 22432 16356 22438
rect 16304 22374 16356 22380
rect 16304 22024 16356 22030
rect 16304 21966 16356 21972
rect 16040 21406 16252 21434
rect 16040 18834 16068 21406
rect 16316 21350 16344 21966
rect 16408 21894 16436 22766
rect 16580 22714 16632 22720
rect 16488 22636 16540 22642
rect 16488 22578 16540 22584
rect 16396 21888 16448 21894
rect 16396 21830 16448 21836
rect 16394 21720 16450 21729
rect 16394 21655 16450 21664
rect 16120 21344 16172 21350
rect 16304 21344 16356 21350
rect 16120 21286 16172 21292
rect 16210 21312 16266 21321
rect 16028 18828 16080 18834
rect 16028 18770 16080 18776
rect 15936 17876 15988 17882
rect 15936 17818 15988 17824
rect 15752 17672 15804 17678
rect 15752 17614 15804 17620
rect 16028 17672 16080 17678
rect 16028 17614 16080 17620
rect 15764 16794 15792 17614
rect 16040 17241 16068 17614
rect 16026 17232 16082 17241
rect 16026 17167 16082 17176
rect 15752 16788 15804 16794
rect 15752 16730 15804 16736
rect 16040 16726 16068 17167
rect 16028 16720 16080 16726
rect 16028 16662 16080 16668
rect 15844 16652 15896 16658
rect 15844 16594 15896 16600
rect 15856 15638 15884 16594
rect 15936 16584 15988 16590
rect 15936 16526 15988 16532
rect 15948 16289 15976 16526
rect 15934 16280 15990 16289
rect 16040 16250 16068 16662
rect 15934 16215 15990 16224
rect 16028 16244 16080 16250
rect 15844 15632 15896 15638
rect 15844 15574 15896 15580
rect 15752 14544 15804 14550
rect 15752 14486 15804 14492
rect 15568 12912 15620 12918
rect 15568 12854 15620 12860
rect 15660 12912 15712 12918
rect 15660 12854 15712 12860
rect 15108 12776 15160 12782
rect 15476 12776 15528 12782
rect 15108 12718 15160 12724
rect 15290 12744 15346 12753
rect 15120 12442 15148 12718
rect 15476 12718 15528 12724
rect 15290 12679 15346 12688
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 15212 12442 15240 12582
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15304 11150 15332 12679
rect 15384 12300 15436 12306
rect 15384 12242 15436 12248
rect 15396 11150 15424 12242
rect 15660 11620 15712 11626
rect 15660 11562 15712 11568
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15304 10742 15332 11086
rect 15292 10736 15344 10742
rect 15292 10678 15344 10684
rect 15396 10588 15424 11086
rect 15304 10560 15424 10588
rect 15304 10062 15332 10560
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14924 9648 14976 9654
rect 14924 9590 14976 9596
rect 14936 9178 14964 9590
rect 15014 9480 15070 9489
rect 15304 9450 15332 9998
rect 15014 9415 15016 9424
rect 15068 9415 15070 9424
rect 15292 9444 15344 9450
rect 15016 9386 15068 9392
rect 15292 9386 15344 9392
rect 14924 9172 14976 9178
rect 14924 9114 14976 9120
rect 14924 8900 14976 8906
rect 15028 8888 15056 9386
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 15212 8974 15240 9318
rect 15396 9092 15424 10202
rect 15304 9064 15424 9092
rect 15200 8968 15252 8974
rect 15200 8910 15252 8916
rect 14976 8860 15056 8888
rect 14924 8842 14976 8848
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15200 8560 15252 8566
rect 15014 8528 15070 8537
rect 15200 8502 15252 8508
rect 15014 8463 15016 8472
rect 15068 8463 15070 8472
rect 15016 8434 15068 8440
rect 15016 8356 15068 8362
rect 15016 8298 15068 8304
rect 15028 8022 15056 8298
rect 15016 8016 15068 8022
rect 14922 7984 14978 7993
rect 15016 7958 15068 7964
rect 14922 7919 14978 7928
rect 14936 7886 14964 7919
rect 14924 7880 14976 7886
rect 14924 7822 14976 7828
rect 15212 7732 15240 8502
rect 15304 8242 15332 9064
rect 15382 8936 15438 8945
rect 15382 8871 15438 8880
rect 15396 8634 15424 8871
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15304 8214 15424 8242
rect 15290 8120 15346 8129
rect 15290 8055 15292 8064
rect 15344 8055 15346 8064
rect 15292 8026 15344 8032
rect 15212 7704 15332 7732
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14832 6928 14884 6934
rect 14832 6870 14884 6876
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14738 6216 14794 6225
rect 14738 6151 14794 6160
rect 14844 5778 14872 6598
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15200 6180 15252 6186
rect 15200 6122 15252 6128
rect 15212 6089 15240 6122
rect 15198 6080 15254 6089
rect 15198 6015 15254 6024
rect 15212 5794 15240 6015
rect 15304 5914 15332 7704
rect 15396 6089 15424 8214
rect 15488 6882 15516 11494
rect 15580 11393 15608 11494
rect 15566 11384 15622 11393
rect 15566 11319 15622 11328
rect 15568 11212 15620 11218
rect 15568 11154 15620 11160
rect 15580 10810 15608 11154
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 15566 10024 15622 10033
rect 15566 9959 15622 9968
rect 15580 9654 15608 9959
rect 15672 9897 15700 11562
rect 15658 9888 15714 9897
rect 15658 9823 15714 9832
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 15568 9648 15620 9654
rect 15568 9590 15620 9596
rect 15568 9036 15620 9042
rect 15568 8978 15620 8984
rect 15580 8498 15608 8978
rect 15568 8492 15620 8498
rect 15568 8434 15620 8440
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 15580 7546 15608 7890
rect 15672 7818 15700 9658
rect 15660 7812 15712 7818
rect 15660 7754 15712 7760
rect 15568 7540 15620 7546
rect 15568 7482 15620 7488
rect 15658 7032 15714 7041
rect 15658 6967 15714 6976
rect 15488 6854 15608 6882
rect 15476 6792 15528 6798
rect 15474 6760 15476 6769
rect 15528 6760 15530 6769
rect 15474 6695 15530 6704
rect 15382 6080 15438 6089
rect 15382 6015 15438 6024
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 14832 5772 14884 5778
rect 15212 5766 15332 5794
rect 14832 5714 14884 5720
rect 14740 5568 14792 5574
rect 14740 5510 14792 5516
rect 14648 5092 14700 5098
rect 14648 5034 14700 5040
rect 14568 4950 14688 4978
rect 14660 4214 14688 4950
rect 14464 4208 14516 4214
rect 14464 4150 14516 4156
rect 14648 4208 14700 4214
rect 14648 4150 14700 4156
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14372 3392 14424 3398
rect 14372 3334 14424 3340
rect 14384 3194 14412 3334
rect 14372 3188 14424 3194
rect 14372 3130 14424 3136
rect 14280 2848 14332 2854
rect 14280 2790 14332 2796
rect 14278 2408 14334 2417
rect 14278 2343 14280 2352
rect 14332 2343 14334 2352
rect 14280 2314 14332 2320
rect 14384 480 14412 3130
rect 14476 2553 14504 4150
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 14568 3534 14596 4082
rect 14648 4072 14700 4078
rect 14648 4014 14700 4020
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 14660 2689 14688 4014
rect 14752 3942 14780 5510
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15304 4758 15332 5766
rect 15580 5624 15608 6854
rect 15672 6118 15700 6967
rect 15660 6112 15712 6118
rect 15660 6054 15712 6060
rect 15658 5944 15714 5953
rect 15658 5879 15660 5888
rect 15712 5879 15714 5888
rect 15660 5850 15712 5856
rect 15488 5596 15608 5624
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 15396 5166 15424 5510
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 15292 4752 15344 4758
rect 15292 4694 15344 4700
rect 15304 4622 15332 4694
rect 15292 4616 15344 4622
rect 15292 4558 15344 4564
rect 14832 4480 14884 4486
rect 14832 4422 14884 4428
rect 14844 4049 14872 4422
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14924 4140 14976 4146
rect 14924 4082 14976 4088
rect 14830 4040 14886 4049
rect 14830 3975 14886 3984
rect 14740 3936 14792 3942
rect 14738 3904 14740 3913
rect 14792 3904 14794 3913
rect 14936 3890 14964 4082
rect 14738 3839 14794 3848
rect 14844 3862 14964 3890
rect 14646 2680 14702 2689
rect 14646 2615 14702 2624
rect 14462 2544 14518 2553
rect 14462 2479 14518 2488
rect 14844 1986 14872 3862
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15108 2984 15160 2990
rect 15304 2972 15332 4558
rect 15488 3720 15516 5596
rect 15566 5536 15622 5545
rect 15566 5471 15622 5480
rect 15580 5302 15608 5471
rect 15672 5370 15700 5850
rect 15660 5364 15712 5370
rect 15660 5306 15712 5312
rect 15568 5296 15620 5302
rect 15568 5238 15620 5244
rect 15658 5264 15714 5273
rect 15658 5199 15714 5208
rect 15672 4570 15700 5199
rect 15580 4542 15700 4570
rect 15580 4146 15608 4542
rect 15658 4448 15714 4457
rect 15658 4383 15714 4392
rect 15568 4140 15620 4146
rect 15568 4082 15620 4088
rect 15580 4010 15608 4082
rect 15568 4004 15620 4010
rect 15568 3946 15620 3952
rect 15672 3738 15700 4383
rect 15764 4282 15792 14486
rect 15856 14414 15884 15574
rect 15948 15366 15976 16215
rect 16028 16186 16080 16192
rect 15936 15360 15988 15366
rect 15936 15302 15988 15308
rect 16026 15328 16082 15337
rect 16026 15263 16082 15272
rect 15936 14952 15988 14958
rect 15936 14894 15988 14900
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 15856 14006 15884 14350
rect 15844 14000 15896 14006
rect 15844 13942 15896 13948
rect 15844 13728 15896 13734
rect 15844 13670 15896 13676
rect 15856 13002 15884 13670
rect 15948 13161 15976 14894
rect 16040 13530 16068 15263
rect 16028 13524 16080 13530
rect 16028 13466 16080 13472
rect 15934 13152 15990 13161
rect 15934 13087 15990 13096
rect 15856 12974 16068 13002
rect 15844 12912 15896 12918
rect 15844 12854 15896 12860
rect 15856 11642 15884 12854
rect 15934 12336 15990 12345
rect 15934 12271 15990 12280
rect 15948 12238 15976 12271
rect 15936 12232 15988 12238
rect 15936 12174 15988 12180
rect 15936 12096 15988 12102
rect 15936 12038 15988 12044
rect 15948 11762 15976 12038
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 15856 11614 15976 11642
rect 15844 11552 15896 11558
rect 15844 11494 15896 11500
rect 15856 9722 15884 11494
rect 15948 10470 15976 11614
rect 15936 10464 15988 10470
rect 15936 10406 15988 10412
rect 15948 9761 15976 10406
rect 15934 9752 15990 9761
rect 15844 9716 15896 9722
rect 15934 9687 15990 9696
rect 15844 9658 15896 9664
rect 15842 9616 15898 9625
rect 15842 9551 15898 9560
rect 15936 9580 15988 9586
rect 15856 9518 15884 9551
rect 15936 9522 15988 9528
rect 15844 9512 15896 9518
rect 15844 9454 15896 9460
rect 15948 9353 15976 9522
rect 15934 9344 15990 9353
rect 15934 9279 15990 9288
rect 15844 9172 15896 9178
rect 15844 9114 15896 9120
rect 15856 8809 15884 9114
rect 15934 9072 15990 9081
rect 15934 9007 15990 9016
rect 15842 8800 15898 8809
rect 15842 8735 15898 8744
rect 15948 8673 15976 9007
rect 15934 8664 15990 8673
rect 15934 8599 15990 8608
rect 15842 8256 15898 8265
rect 15842 8191 15898 8200
rect 15856 7546 15884 8191
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 15856 7342 15884 7482
rect 15844 7336 15896 7342
rect 15844 7278 15896 7284
rect 15844 6860 15896 6866
rect 15844 6802 15896 6808
rect 15856 5710 15884 6802
rect 15948 5914 15976 8599
rect 16040 6610 16068 12974
rect 16132 6730 16160 21286
rect 16304 21286 16356 21292
rect 16210 21247 16266 21256
rect 16224 18970 16252 21247
rect 16316 21078 16344 21286
rect 16304 21072 16356 21078
rect 16304 21014 16356 21020
rect 16408 20924 16436 21655
rect 16316 20896 16436 20924
rect 16500 21162 16528 22578
rect 16500 21146 16620 21162
rect 16500 21140 16632 21146
rect 16500 21134 16580 21140
rect 16212 18964 16264 18970
rect 16212 18906 16264 18912
rect 16212 18828 16264 18834
rect 16212 18770 16264 18776
rect 16224 13920 16252 18770
rect 16316 18154 16344 20896
rect 16500 19990 16528 21134
rect 16580 21082 16632 21088
rect 16488 19984 16540 19990
rect 16488 19926 16540 19932
rect 16500 19514 16528 19926
rect 16580 19712 16632 19718
rect 16580 19654 16632 19660
rect 16488 19508 16540 19514
rect 16488 19450 16540 19456
rect 16592 18952 16620 19654
rect 16684 19145 16712 23990
rect 16776 23866 16804 24550
rect 16868 24342 16896 24754
rect 16856 24336 16908 24342
rect 16856 24278 16908 24284
rect 16856 24064 16908 24070
rect 16856 24006 16908 24012
rect 16764 23860 16816 23866
rect 16764 23802 16816 23808
rect 16762 23352 16818 23361
rect 16762 23287 16764 23296
rect 16816 23287 16818 23296
rect 16764 23258 16816 23264
rect 16764 22976 16816 22982
rect 16868 22964 16896 24006
rect 16960 23322 16988 25327
rect 17314 25327 17370 25336
rect 17132 25298 17184 25304
rect 17144 24818 17172 25298
rect 17224 25220 17276 25226
rect 17224 25162 17276 25168
rect 17236 24954 17264 25162
rect 17224 24948 17276 24954
rect 17224 24890 17276 24896
rect 17132 24812 17184 24818
rect 17132 24754 17184 24760
rect 17132 24676 17184 24682
rect 17132 24618 17184 24624
rect 17040 24132 17092 24138
rect 17040 24074 17092 24080
rect 16948 23316 17000 23322
rect 16948 23258 17000 23264
rect 16948 23044 17000 23050
rect 16948 22986 17000 22992
rect 16816 22936 16896 22964
rect 16764 22918 16816 22924
rect 16776 22642 16804 22918
rect 16960 22794 16988 22986
rect 17052 22953 17080 24074
rect 17038 22944 17094 22953
rect 17038 22879 17094 22888
rect 16868 22766 16988 22794
rect 16764 22636 16816 22642
rect 16764 22578 16816 22584
rect 16868 21962 16896 22766
rect 17038 22536 17094 22545
rect 17038 22471 17094 22480
rect 17052 22438 17080 22471
rect 17040 22432 17092 22438
rect 17040 22374 17092 22380
rect 16948 22024 17000 22030
rect 16948 21966 17000 21972
rect 16856 21956 16908 21962
rect 16856 21898 16908 21904
rect 16764 20460 16816 20466
rect 16764 20402 16816 20408
rect 16776 19378 16804 20402
rect 16764 19372 16816 19378
rect 16764 19314 16816 19320
rect 16670 19136 16726 19145
rect 16670 19071 16726 19080
rect 16500 18924 16620 18952
rect 16500 18766 16528 18924
rect 16868 18816 16896 21898
rect 16960 21865 16988 21966
rect 16946 21856 17002 21865
rect 16946 21791 17002 21800
rect 16960 21350 16988 21791
rect 17040 21616 17092 21622
rect 17040 21558 17092 21564
rect 16948 21344 17000 21350
rect 16948 21286 17000 21292
rect 16960 21010 16988 21286
rect 16948 21004 17000 21010
rect 16948 20946 17000 20952
rect 16946 20768 17002 20777
rect 16946 20703 17002 20712
rect 16960 19310 16988 20703
rect 16948 19304 17000 19310
rect 16948 19246 17000 19252
rect 16592 18788 16896 18816
rect 16948 18828 17000 18834
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 16488 18216 16540 18222
rect 16488 18158 16540 18164
rect 16304 18148 16356 18154
rect 16304 18090 16356 18096
rect 16316 17542 16344 18090
rect 16396 18080 16448 18086
rect 16396 18022 16448 18028
rect 16304 17536 16356 17542
rect 16304 17478 16356 17484
rect 16316 17338 16344 17478
rect 16304 17332 16356 17338
rect 16304 17274 16356 17280
rect 16408 17218 16436 18022
rect 16500 17746 16528 18158
rect 16488 17740 16540 17746
rect 16488 17682 16540 17688
rect 16486 17504 16542 17513
rect 16486 17439 16542 17448
rect 16316 17190 16436 17218
rect 16316 15337 16344 17190
rect 16396 16516 16448 16522
rect 16396 16458 16448 16464
rect 16408 16250 16436 16458
rect 16396 16244 16448 16250
rect 16396 16186 16448 16192
rect 16500 15706 16528 17439
rect 16488 15700 16540 15706
rect 16408 15660 16488 15688
rect 16408 15473 16436 15660
rect 16488 15642 16540 15648
rect 16488 15564 16540 15570
rect 16488 15506 16540 15512
rect 16394 15464 16450 15473
rect 16394 15399 16450 15408
rect 16302 15328 16358 15337
rect 16302 15263 16358 15272
rect 16408 15162 16436 15399
rect 16396 15156 16448 15162
rect 16396 15098 16448 15104
rect 16396 14952 16448 14958
rect 16396 14894 16448 14900
rect 16408 14482 16436 14894
rect 16500 14822 16528 15506
rect 16488 14816 16540 14822
rect 16488 14758 16540 14764
rect 16500 14618 16528 14758
rect 16488 14612 16540 14618
rect 16488 14554 16540 14560
rect 16396 14476 16448 14482
rect 16396 14418 16448 14424
rect 16224 13892 16528 13920
rect 16302 13832 16358 13841
rect 16302 13767 16358 13776
rect 16316 12986 16344 13767
rect 16396 13728 16448 13734
rect 16396 13670 16448 13676
rect 16304 12980 16356 12986
rect 16304 12922 16356 12928
rect 16210 12880 16266 12889
rect 16210 12815 16212 12824
rect 16264 12815 16266 12824
rect 16212 12786 16264 12792
rect 16304 12708 16356 12714
rect 16304 12650 16356 12656
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16224 10554 16252 11834
rect 16316 10674 16344 12650
rect 16408 12442 16436 13670
rect 16396 12436 16448 12442
rect 16396 12378 16448 12384
rect 16394 11928 16450 11937
rect 16394 11863 16396 11872
rect 16448 11863 16450 11872
rect 16396 11834 16448 11840
rect 16500 11354 16528 13892
rect 16592 12186 16620 18788
rect 16948 18770 17000 18776
rect 16764 18692 16816 18698
rect 16764 18634 16816 18640
rect 16672 18624 16724 18630
rect 16672 18566 16724 18572
rect 16684 18057 16712 18566
rect 16670 18048 16726 18057
rect 16670 17983 16726 17992
rect 16672 17604 16724 17610
rect 16672 17546 16724 17552
rect 16684 17377 16712 17546
rect 16776 17542 16804 18634
rect 16960 18358 16988 18770
rect 16856 18352 16908 18358
rect 16854 18320 16856 18329
rect 16948 18352 17000 18358
rect 16908 18320 16910 18329
rect 16948 18294 17000 18300
rect 16854 18255 16910 18264
rect 16868 17814 16896 18255
rect 16856 17808 16908 17814
rect 16856 17750 16908 17756
rect 16764 17536 16816 17542
rect 16764 17478 16816 17484
rect 16670 17368 16726 17377
rect 16670 17303 16726 17312
rect 16684 16794 16712 17303
rect 16672 16788 16724 16794
rect 16672 16730 16724 16736
rect 16684 16454 16712 16730
rect 16672 16448 16724 16454
rect 16672 16390 16724 16396
rect 16672 15496 16724 15502
rect 16672 15438 16724 15444
rect 16684 14346 16712 15438
rect 16672 14340 16724 14346
rect 16672 14282 16724 14288
rect 16684 13938 16712 14282
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 16672 13184 16724 13190
rect 16672 13126 16724 13132
rect 16684 12442 16712 13126
rect 16776 12481 16804 17478
rect 16868 17338 16896 17750
rect 16856 17332 16908 17338
rect 16856 17274 16908 17280
rect 17052 16776 17080 21558
rect 16960 16748 17080 16776
rect 16960 16130 16988 16748
rect 17038 16688 17094 16697
rect 17038 16623 17040 16632
rect 17092 16623 17094 16632
rect 17040 16594 17092 16600
rect 17052 16250 17080 16594
rect 17040 16244 17092 16250
rect 17040 16186 17092 16192
rect 16960 16102 17080 16130
rect 16948 16040 17000 16046
rect 16948 15982 17000 15988
rect 16856 14476 16908 14482
rect 16856 14418 16908 14424
rect 16868 14385 16896 14418
rect 16854 14376 16910 14385
rect 16854 14311 16910 14320
rect 16868 14074 16896 14311
rect 16856 14068 16908 14074
rect 16856 14010 16908 14016
rect 16856 13864 16908 13870
rect 16854 13832 16856 13841
rect 16908 13832 16910 13841
rect 16854 13767 16910 13776
rect 16762 12472 16818 12481
rect 16672 12436 16724 12442
rect 16762 12407 16818 12416
rect 16672 12378 16724 12384
rect 16856 12300 16908 12306
rect 16856 12242 16908 12248
rect 16592 12158 16712 12186
rect 16684 12102 16712 12158
rect 16672 12096 16724 12102
rect 16672 12038 16724 12044
rect 16580 11824 16632 11830
rect 16580 11766 16632 11772
rect 16670 11792 16726 11801
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16394 10840 16450 10849
rect 16394 10775 16396 10784
rect 16448 10775 16450 10784
rect 16396 10746 16448 10752
rect 16304 10668 16356 10674
rect 16304 10610 16356 10616
rect 16224 10526 16436 10554
rect 16212 10464 16264 10470
rect 16210 10432 16212 10441
rect 16264 10432 16266 10441
rect 16210 10367 16266 10376
rect 16304 10192 16356 10198
rect 16304 10134 16356 10140
rect 16210 9752 16266 9761
rect 16210 9687 16266 9696
rect 16224 6866 16252 9687
rect 16316 9654 16344 10134
rect 16304 9648 16356 9654
rect 16304 9590 16356 9596
rect 16302 9344 16358 9353
rect 16302 9279 16358 9288
rect 16316 9110 16344 9279
rect 16304 9104 16356 9110
rect 16304 9046 16356 9052
rect 16304 8832 16356 8838
rect 16304 8774 16356 8780
rect 16316 8537 16344 8774
rect 16302 8528 16358 8537
rect 16302 8463 16358 8472
rect 16408 8106 16436 10526
rect 16500 10198 16528 11290
rect 16488 10192 16540 10198
rect 16488 10134 16540 10140
rect 16592 10112 16620 11766
rect 16868 11762 16896 12242
rect 16960 12209 16988 15982
rect 17052 15026 17080 16102
rect 17040 15020 17092 15026
rect 17040 14962 17092 14968
rect 17040 14816 17092 14822
rect 17040 14758 17092 14764
rect 17052 13841 17080 14758
rect 17038 13832 17094 13841
rect 17038 13767 17094 13776
rect 16946 12200 17002 12209
rect 16946 12135 17002 12144
rect 16670 11727 16726 11736
rect 16856 11756 16908 11762
rect 16684 11626 16712 11727
rect 16856 11698 16908 11704
rect 16764 11688 16816 11694
rect 16764 11630 16816 11636
rect 16672 11620 16724 11626
rect 16672 11562 16724 11568
rect 16776 11506 16804 11630
rect 16572 10084 16620 10112
rect 16684 11478 16804 11506
rect 16572 10044 16600 10084
rect 16500 10016 16600 10044
rect 16500 9722 16528 10016
rect 16684 9908 16712 11478
rect 16868 10674 16896 11698
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 16856 10464 16908 10470
rect 16856 10406 16908 10412
rect 16592 9880 16712 9908
rect 16764 9920 16816 9926
rect 16488 9716 16540 9722
rect 16488 9658 16540 9664
rect 16486 9616 16542 9625
rect 16486 9551 16542 9560
rect 16500 9081 16528 9551
rect 16486 9072 16542 9081
rect 16486 9007 16542 9016
rect 16592 8566 16620 9880
rect 16868 9897 16896 10406
rect 16960 10266 16988 12135
rect 17038 11112 17094 11121
rect 17038 11047 17094 11056
rect 16948 10260 17000 10266
rect 16948 10202 17000 10208
rect 16946 10024 17002 10033
rect 16946 9959 17002 9968
rect 16764 9862 16816 9868
rect 16854 9888 16910 9897
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 16580 8560 16632 8566
rect 16580 8502 16632 8508
rect 16304 8084 16356 8090
rect 16408 8078 16528 8106
rect 16304 8026 16356 8032
rect 16212 6860 16264 6866
rect 16212 6802 16264 6808
rect 16120 6724 16172 6730
rect 16120 6666 16172 6672
rect 16040 6582 16160 6610
rect 15936 5908 15988 5914
rect 15936 5850 15988 5856
rect 15844 5704 15896 5710
rect 15844 5646 15896 5652
rect 16026 5672 16082 5681
rect 15856 5302 15884 5646
rect 16026 5607 16028 5616
rect 16080 5607 16082 5616
rect 16028 5578 16080 5584
rect 15936 5568 15988 5574
rect 15936 5510 15988 5516
rect 15844 5296 15896 5302
rect 15844 5238 15896 5244
rect 15844 5160 15896 5166
rect 15844 5102 15896 5108
rect 15752 4276 15804 4282
rect 15752 4218 15804 4224
rect 15856 4214 15884 5102
rect 15948 5001 15976 5510
rect 16026 5400 16082 5409
rect 16026 5335 16082 5344
rect 16040 5234 16068 5335
rect 16028 5228 16080 5234
rect 16028 5170 16080 5176
rect 15934 4992 15990 5001
rect 15934 4927 15990 4936
rect 16040 4826 16068 5170
rect 16028 4820 16080 4826
rect 16028 4762 16080 4768
rect 16028 4276 16080 4282
rect 16028 4218 16080 4224
rect 15844 4208 15896 4214
rect 15844 4150 15896 4156
rect 15660 3732 15712 3738
rect 15488 3692 15608 3720
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 15160 2944 15332 2972
rect 15108 2926 15160 2932
rect 14924 2848 14976 2854
rect 14924 2790 14976 2796
rect 14936 2582 14964 2790
rect 14924 2576 14976 2582
rect 14924 2518 14976 2524
rect 15120 2514 15148 2926
rect 15384 2916 15436 2922
rect 15384 2858 15436 2864
rect 15108 2508 15160 2514
rect 15108 2450 15160 2456
rect 15396 2378 15424 2858
rect 15488 2650 15516 3538
rect 15580 2825 15608 3692
rect 15660 3674 15712 3680
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 15856 2922 15884 3470
rect 15844 2916 15896 2922
rect 15844 2858 15896 2864
rect 15566 2816 15622 2825
rect 15566 2751 15622 2760
rect 15476 2644 15528 2650
rect 15476 2586 15528 2592
rect 15384 2372 15436 2378
rect 15384 2314 15436 2320
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14844 1958 14964 1986
rect 14936 480 14964 1958
rect 15488 480 15516 2246
rect 16040 480 16068 4218
rect 16132 2310 16160 6582
rect 16316 6322 16344 8026
rect 16396 8016 16448 8022
rect 16396 7958 16448 7964
rect 16408 7857 16436 7958
rect 16394 7848 16450 7857
rect 16394 7783 16450 7792
rect 16396 7200 16448 7206
rect 16396 7142 16448 7148
rect 16408 6934 16436 7142
rect 16396 6928 16448 6934
rect 16396 6870 16448 6876
rect 16396 6656 16448 6662
rect 16396 6598 16448 6604
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 16224 4282 16252 6054
rect 16408 5760 16436 6598
rect 16316 5732 16436 5760
rect 16212 4276 16264 4282
rect 16212 4218 16264 4224
rect 16316 4146 16344 5732
rect 16500 5658 16528 8078
rect 16578 7712 16634 7721
rect 16578 7647 16634 7656
rect 16592 6905 16620 7647
rect 16578 6896 16634 6905
rect 16578 6831 16634 6840
rect 16684 6798 16712 9590
rect 16776 8498 16804 9862
rect 16854 9823 16910 9832
rect 16856 9716 16908 9722
rect 16856 9658 16908 9664
rect 16868 8945 16896 9658
rect 16854 8936 16910 8945
rect 16854 8871 16910 8880
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16764 8356 16816 8362
rect 16764 8298 16816 8304
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16684 5914 16712 6734
rect 16672 5908 16724 5914
rect 16672 5850 16724 5856
rect 16580 5840 16632 5846
rect 16580 5782 16632 5788
rect 16408 5630 16528 5658
rect 16408 5001 16436 5630
rect 16488 5568 16540 5574
rect 16488 5510 16540 5516
rect 16500 5250 16528 5510
rect 16592 5370 16620 5782
rect 16580 5364 16632 5370
rect 16580 5306 16632 5312
rect 16500 5222 16712 5250
rect 16394 4992 16450 5001
rect 16394 4927 16450 4936
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16316 3670 16344 4082
rect 16408 4078 16436 4927
rect 16488 4684 16540 4690
rect 16488 4626 16540 4632
rect 16500 4214 16528 4626
rect 16684 4593 16712 5222
rect 16776 4729 16804 8298
rect 16868 6730 16896 8871
rect 16856 6724 16908 6730
rect 16856 6666 16908 6672
rect 16854 6624 16910 6633
rect 16854 6559 16910 6568
rect 16868 5914 16896 6559
rect 16960 6458 16988 9959
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 16948 6112 17000 6118
rect 16948 6054 17000 6060
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 16762 4720 16818 4729
rect 16762 4655 16818 4664
rect 16670 4584 16726 4593
rect 16670 4519 16726 4528
rect 16856 4480 16908 4486
rect 16856 4422 16908 4428
rect 16488 4208 16540 4214
rect 16488 4150 16540 4156
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16762 3768 16818 3777
rect 16762 3703 16818 3712
rect 16776 3670 16804 3703
rect 16304 3664 16356 3670
rect 16304 3606 16356 3612
rect 16764 3664 16816 3670
rect 16764 3606 16816 3612
rect 16868 3534 16896 4422
rect 16960 4078 16988 6054
rect 16948 4072 17000 4078
rect 16948 4014 17000 4020
rect 16948 3936 17000 3942
rect 16948 3878 17000 3884
rect 16960 3738 16988 3878
rect 16948 3732 17000 3738
rect 16948 3674 17000 3680
rect 16856 3528 16908 3534
rect 16856 3470 16908 3476
rect 16868 3194 16896 3470
rect 16580 3188 16632 3194
rect 16580 3130 16632 3136
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 16592 2802 16620 3130
rect 16500 2774 16620 2802
rect 16500 2446 16528 2774
rect 17052 2650 17080 11047
rect 17144 3738 17172 24618
rect 17328 24449 17356 25327
rect 17776 24608 17828 24614
rect 17776 24550 17828 24556
rect 17314 24440 17370 24449
rect 17314 24375 17370 24384
rect 17408 24336 17460 24342
rect 17788 24313 17816 24550
rect 17972 24392 18000 26318
rect 18236 26240 18288 26246
rect 18236 26182 18288 26188
rect 18052 25152 18104 25158
rect 18052 25094 18104 25100
rect 18064 24886 18092 25094
rect 18052 24880 18104 24886
rect 18052 24822 18104 24828
rect 18248 24818 18276 26182
rect 18340 26110 18368 27520
rect 18328 26104 18380 26110
rect 18328 26046 18380 26052
rect 18892 25770 18920 27520
rect 19536 25838 19564 27520
rect 20088 26602 20116 27520
rect 19996 26574 20116 26602
rect 19524 25832 19576 25838
rect 19524 25774 19576 25780
rect 18880 25764 18932 25770
rect 18880 25706 18932 25712
rect 18972 25764 19024 25770
rect 18972 25706 19024 25712
rect 18880 25356 18932 25362
rect 18880 25298 18932 25304
rect 18510 25120 18566 25129
rect 18510 25055 18566 25064
rect 18418 24984 18474 24993
rect 18418 24919 18474 24928
rect 18236 24812 18288 24818
rect 18236 24754 18288 24760
rect 18236 24404 18288 24410
rect 17972 24364 18092 24392
rect 17408 24278 17460 24284
rect 17774 24304 17830 24313
rect 17316 24200 17368 24206
rect 17316 24142 17368 24148
rect 17328 23798 17356 24142
rect 17316 23792 17368 23798
rect 17316 23734 17368 23740
rect 17420 23644 17448 24278
rect 17500 24268 17552 24274
rect 17774 24239 17830 24248
rect 17960 24268 18012 24274
rect 17500 24210 17552 24216
rect 17328 23616 17448 23644
rect 17224 23316 17276 23322
rect 17224 23258 17276 23264
rect 17236 22778 17264 23258
rect 17224 22772 17276 22778
rect 17224 22714 17276 22720
rect 17328 22574 17356 23616
rect 17512 23526 17540 24210
rect 17788 23594 17816 24239
rect 17960 24210 18012 24216
rect 17776 23588 17828 23594
rect 17776 23530 17828 23536
rect 17500 23520 17552 23526
rect 17500 23462 17552 23468
rect 17406 23352 17462 23361
rect 17406 23287 17462 23296
rect 17316 22568 17368 22574
rect 17316 22510 17368 22516
rect 17222 22128 17278 22137
rect 17222 22063 17224 22072
rect 17276 22063 17278 22072
rect 17224 22034 17276 22040
rect 17236 21690 17264 22034
rect 17224 21684 17276 21690
rect 17224 21626 17276 21632
rect 17222 18864 17278 18873
rect 17222 18799 17278 18808
rect 17236 16794 17264 18799
rect 17224 16788 17276 16794
rect 17224 16730 17276 16736
rect 17224 15904 17276 15910
rect 17224 15846 17276 15852
rect 17236 15337 17264 15846
rect 17222 15328 17278 15337
rect 17222 15263 17278 15272
rect 17224 14544 17276 14550
rect 17224 14486 17276 14492
rect 17236 14414 17264 14486
rect 17224 14408 17276 14414
rect 17224 14350 17276 14356
rect 17236 14074 17264 14350
rect 17224 14068 17276 14074
rect 17224 14010 17276 14016
rect 17222 13968 17278 13977
rect 17222 13903 17278 13912
rect 17236 13870 17264 13903
rect 17224 13864 17276 13870
rect 17224 13806 17276 13812
rect 17328 11626 17356 22510
rect 17420 20398 17448 23287
rect 17512 21185 17540 23462
rect 17972 23338 18000 24210
rect 18064 23526 18092 24364
rect 18236 24346 18288 24352
rect 18144 24064 18196 24070
rect 18144 24006 18196 24012
rect 18156 23594 18184 24006
rect 18144 23588 18196 23594
rect 18144 23530 18196 23536
rect 18052 23520 18104 23526
rect 18052 23462 18104 23468
rect 17604 23310 18000 23338
rect 18064 23322 18092 23462
rect 18052 23316 18104 23322
rect 17498 21176 17554 21185
rect 17498 21111 17554 21120
rect 17408 20392 17460 20398
rect 17408 20334 17460 20340
rect 17498 19952 17554 19961
rect 17498 19887 17554 19896
rect 17408 19712 17460 19718
rect 17408 19654 17460 19660
rect 17420 19417 17448 19654
rect 17406 19408 17462 19417
rect 17406 19343 17462 19352
rect 17512 19310 17540 19887
rect 17500 19304 17552 19310
rect 17500 19246 17552 19252
rect 17500 18828 17552 18834
rect 17500 18770 17552 18776
rect 17512 18193 17540 18770
rect 17498 18184 17554 18193
rect 17498 18119 17500 18128
rect 17552 18119 17554 18128
rect 17500 18090 17552 18096
rect 17408 17876 17460 17882
rect 17408 17818 17460 17824
rect 17420 17785 17448 17818
rect 17406 17776 17462 17785
rect 17406 17711 17462 17720
rect 17500 17740 17552 17746
rect 17500 17682 17552 17688
rect 17512 17270 17540 17682
rect 17500 17264 17552 17270
rect 17500 17206 17552 17212
rect 17408 17128 17460 17134
rect 17408 17070 17460 17076
rect 17420 16522 17448 17070
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17408 16516 17460 16522
rect 17408 16458 17460 16464
rect 17420 15910 17448 16458
rect 17512 16250 17540 16526
rect 17500 16244 17552 16250
rect 17500 16186 17552 16192
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 17500 15428 17552 15434
rect 17500 15370 17552 15376
rect 17408 15020 17460 15026
rect 17408 14962 17460 14968
rect 17420 13410 17448 14962
rect 17512 14618 17540 15370
rect 17500 14612 17552 14618
rect 17500 14554 17552 14560
rect 17512 13530 17540 14554
rect 17604 13530 17632 23310
rect 18052 23258 18104 23264
rect 17776 23180 17828 23186
rect 17776 23122 17828 23128
rect 17684 23044 17736 23050
rect 17684 22986 17736 22992
rect 17696 17252 17724 22986
rect 17788 22438 17816 23122
rect 17776 22432 17828 22438
rect 17774 22400 17776 22409
rect 18144 22432 18196 22438
rect 17828 22400 17830 22409
rect 18248 22409 18276 24346
rect 18432 23322 18460 24919
rect 18420 23316 18472 23322
rect 18420 23258 18472 23264
rect 18328 22500 18380 22506
rect 18380 22460 18460 22488
rect 18328 22442 18380 22448
rect 18144 22374 18196 22380
rect 18234 22400 18290 22409
rect 17774 22335 17830 22344
rect 17868 22024 17920 22030
rect 17868 21966 17920 21972
rect 17880 20534 17908 21966
rect 18156 21894 18184 22374
rect 18234 22335 18290 22344
rect 18144 21888 18196 21894
rect 18144 21830 18196 21836
rect 17960 21412 18012 21418
rect 17960 21354 18012 21360
rect 17868 20528 17920 20534
rect 17868 20470 17920 20476
rect 17776 20256 17828 20262
rect 17776 20198 17828 20204
rect 17788 19825 17816 20198
rect 17972 20074 18000 21354
rect 18052 21344 18104 21350
rect 18052 21286 18104 21292
rect 18064 21049 18092 21286
rect 18050 21040 18106 21049
rect 18050 20975 18106 20984
rect 18050 20632 18106 20641
rect 18050 20567 18052 20576
rect 18104 20567 18106 20576
rect 18052 20538 18104 20544
rect 17880 20058 18000 20074
rect 17868 20052 18000 20058
rect 17920 20046 18000 20052
rect 17868 19994 17920 20000
rect 17774 19816 17830 19825
rect 17774 19751 17830 19760
rect 17868 18080 17920 18086
rect 17868 18022 17920 18028
rect 17696 17224 17816 17252
rect 17684 16448 17736 16454
rect 17684 16390 17736 16396
rect 17696 16046 17724 16390
rect 17684 16040 17736 16046
rect 17684 15982 17736 15988
rect 17684 15904 17736 15910
rect 17684 15846 17736 15852
rect 17696 15473 17724 15846
rect 17682 15464 17738 15473
rect 17682 15399 17738 15408
rect 17684 14952 17736 14958
rect 17684 14894 17736 14900
rect 17696 14521 17724 14894
rect 17682 14512 17738 14521
rect 17682 14447 17738 14456
rect 17684 13932 17736 13938
rect 17684 13874 17736 13880
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17592 13524 17644 13530
rect 17592 13466 17644 13472
rect 17696 13462 17724 13874
rect 17684 13456 17736 13462
rect 17420 13382 17632 13410
rect 17684 13398 17736 13404
rect 17498 13016 17554 13025
rect 17498 12951 17500 12960
rect 17552 12951 17554 12960
rect 17500 12922 17552 12928
rect 17498 12744 17554 12753
rect 17498 12679 17554 12688
rect 17512 12442 17540 12679
rect 17500 12436 17552 12442
rect 17500 12378 17552 12384
rect 17408 12096 17460 12102
rect 17408 12038 17460 12044
rect 17224 11620 17276 11626
rect 17224 11562 17276 11568
rect 17316 11620 17368 11626
rect 17316 11562 17368 11568
rect 17236 11529 17264 11562
rect 17222 11520 17278 11529
rect 17222 11455 17278 11464
rect 17420 11218 17448 12038
rect 17512 11898 17540 12378
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17500 11620 17552 11626
rect 17500 11562 17552 11568
rect 17408 11212 17460 11218
rect 17408 11154 17460 11160
rect 17224 9920 17276 9926
rect 17224 9862 17276 9868
rect 17316 9920 17368 9926
rect 17316 9862 17368 9868
rect 17236 7857 17264 9862
rect 17328 9518 17356 9862
rect 17420 9761 17448 11154
rect 17406 9752 17462 9761
rect 17406 9687 17462 9696
rect 17512 9636 17540 11562
rect 17420 9608 17540 9636
rect 17316 9512 17368 9518
rect 17316 9454 17368 9460
rect 17328 9110 17356 9454
rect 17316 9104 17368 9110
rect 17316 9046 17368 9052
rect 17316 8968 17368 8974
rect 17316 8910 17368 8916
rect 17328 8634 17356 8910
rect 17316 8628 17368 8634
rect 17316 8570 17368 8576
rect 17316 8492 17368 8498
rect 17316 8434 17368 8440
rect 17222 7848 17278 7857
rect 17222 7783 17278 7792
rect 17328 3777 17356 8434
rect 17420 7426 17448 9608
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17512 9042 17540 9318
rect 17500 9036 17552 9042
rect 17500 8978 17552 8984
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 17512 7546 17540 8570
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 17420 7398 17540 7426
rect 17408 7336 17460 7342
rect 17408 7278 17460 7284
rect 17420 5522 17448 7278
rect 17512 6118 17540 7398
rect 17604 7274 17632 13382
rect 17682 10976 17738 10985
rect 17682 10911 17738 10920
rect 17696 9217 17724 10911
rect 17682 9208 17738 9217
rect 17682 9143 17738 9152
rect 17696 8537 17724 9143
rect 17682 8528 17738 8537
rect 17682 8463 17738 8472
rect 17684 8424 17736 8430
rect 17684 8366 17736 8372
rect 17696 7970 17724 8366
rect 17788 8090 17816 17224
rect 17880 16028 17908 18022
rect 17972 17338 18000 20046
rect 18052 19984 18104 19990
rect 18052 19926 18104 19932
rect 18064 19174 18092 19926
rect 18052 19168 18104 19174
rect 18052 19110 18104 19116
rect 18052 18896 18104 18902
rect 18052 18838 18104 18844
rect 17960 17332 18012 17338
rect 17960 17274 18012 17280
rect 18064 16794 18092 18838
rect 18156 16810 18184 21830
rect 18248 18970 18276 22335
rect 18328 22024 18380 22030
rect 18328 21966 18380 21972
rect 18340 21622 18368 21966
rect 18328 21616 18380 21622
rect 18328 21558 18380 21564
rect 18328 21344 18380 21350
rect 18328 21286 18380 21292
rect 18340 19417 18368 21286
rect 18326 19408 18382 19417
rect 18326 19343 18382 19352
rect 18328 19168 18380 19174
rect 18328 19110 18380 19116
rect 18236 18964 18288 18970
rect 18236 18906 18288 18912
rect 18248 18222 18276 18906
rect 18340 18850 18368 19110
rect 18432 18970 18460 22460
rect 18524 21457 18552 25055
rect 18602 24984 18658 24993
rect 18602 24919 18658 24928
rect 18616 24585 18644 24919
rect 18892 24614 18920 25298
rect 18984 25226 19012 25706
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19996 25498 20024 26574
rect 20076 26444 20128 26450
rect 20076 26386 20128 26392
rect 19984 25492 20036 25498
rect 19984 25434 20036 25440
rect 18972 25220 19024 25226
rect 18972 25162 19024 25168
rect 19984 24880 20036 24886
rect 19984 24822 20036 24828
rect 19800 24744 19852 24750
rect 19798 24712 19800 24721
rect 19852 24712 19854 24721
rect 19248 24676 19300 24682
rect 19798 24647 19854 24656
rect 19248 24618 19300 24624
rect 18880 24608 18932 24614
rect 18602 24576 18658 24585
rect 18880 24550 18932 24556
rect 18602 24511 18658 24520
rect 18696 24200 18748 24206
rect 18696 24142 18748 24148
rect 18604 24132 18656 24138
rect 18604 24074 18656 24080
rect 18616 23730 18644 24074
rect 18708 23769 18736 24142
rect 18694 23760 18750 23769
rect 18604 23724 18656 23730
rect 18694 23695 18750 23704
rect 18604 23666 18656 23672
rect 18788 23520 18840 23526
rect 18788 23462 18840 23468
rect 18800 23236 18828 23462
rect 18892 23361 18920 24550
rect 18972 23724 19024 23730
rect 18972 23666 19024 23672
rect 18878 23352 18934 23361
rect 18878 23287 18934 23296
rect 18800 23208 18920 23236
rect 18696 22704 18748 22710
rect 18696 22646 18748 22652
rect 18602 21720 18658 21729
rect 18602 21655 18658 21664
rect 18616 21554 18644 21655
rect 18604 21548 18656 21554
rect 18604 21490 18656 21496
rect 18510 21448 18566 21457
rect 18510 21383 18566 21392
rect 18602 21312 18658 21321
rect 18602 21247 18658 21256
rect 18616 21146 18644 21247
rect 18604 21140 18656 21146
rect 18604 21082 18656 21088
rect 18604 21004 18656 21010
rect 18604 20946 18656 20952
rect 18512 20800 18564 20806
rect 18512 20742 18564 20748
rect 18524 20466 18552 20742
rect 18512 20460 18564 20466
rect 18512 20402 18564 20408
rect 18524 20058 18552 20402
rect 18512 20052 18564 20058
rect 18512 19994 18564 20000
rect 18510 19544 18566 19553
rect 18510 19479 18566 19488
rect 18524 18970 18552 19479
rect 18616 19281 18644 20946
rect 18602 19272 18658 19281
rect 18602 19207 18658 19216
rect 18602 19000 18658 19009
rect 18420 18964 18472 18970
rect 18420 18906 18472 18912
rect 18512 18964 18564 18970
rect 18602 18935 18658 18944
rect 18512 18906 18564 18912
rect 18340 18822 18460 18850
rect 18236 18216 18288 18222
rect 18236 18158 18288 18164
rect 18432 17882 18460 18822
rect 18616 18766 18644 18935
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18604 18624 18656 18630
rect 18604 18566 18656 18572
rect 18510 18456 18566 18465
rect 18510 18391 18566 18400
rect 18420 17876 18472 17882
rect 18420 17818 18472 17824
rect 18524 17082 18552 18391
rect 18616 18290 18644 18566
rect 18604 18284 18656 18290
rect 18604 18226 18656 18232
rect 18604 18148 18656 18154
rect 18604 18090 18656 18096
rect 18432 17054 18552 17082
rect 18052 16788 18104 16794
rect 18156 16782 18368 16810
rect 18052 16730 18104 16736
rect 18144 16720 18196 16726
rect 18144 16662 18196 16668
rect 18156 16590 18184 16662
rect 18144 16584 18196 16590
rect 18144 16526 18196 16532
rect 18156 16046 18184 16526
rect 18144 16040 18196 16046
rect 17880 16000 18092 16028
rect 17960 15496 18012 15502
rect 17960 15438 18012 15444
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 17880 13546 17908 15302
rect 17972 14618 18000 15438
rect 18064 15065 18092 16000
rect 18144 15982 18196 15988
rect 18156 15144 18184 15982
rect 18236 15156 18288 15162
rect 18156 15116 18236 15144
rect 18236 15098 18288 15104
rect 18050 15056 18106 15065
rect 18050 14991 18106 15000
rect 18248 14822 18276 15098
rect 18236 14816 18288 14822
rect 18236 14758 18288 14764
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 18144 14544 18196 14550
rect 18144 14486 18196 14492
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 17972 14006 18000 14418
rect 18052 14068 18104 14074
rect 18052 14010 18104 14016
rect 17960 14000 18012 14006
rect 17960 13942 18012 13948
rect 18064 13870 18092 14010
rect 18156 13870 18184 14486
rect 18248 14074 18276 14758
rect 18236 14068 18288 14074
rect 18236 14010 18288 14016
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 18144 13864 18196 13870
rect 18144 13806 18196 13812
rect 17880 13530 18000 13546
rect 17880 13524 18012 13530
rect 17880 13518 17960 13524
rect 17960 13466 18012 13472
rect 18234 13424 18290 13433
rect 18234 13359 18236 13368
rect 18288 13359 18290 13368
rect 18236 13330 18288 13336
rect 17866 13152 17922 13161
rect 17866 13087 17922 13096
rect 18050 13152 18106 13161
rect 18050 13087 18106 13096
rect 17880 12889 17908 13087
rect 17866 12880 17922 12889
rect 17866 12815 17922 12824
rect 17880 12374 17908 12815
rect 18064 12646 18092 13087
rect 18236 12776 18288 12782
rect 18236 12718 18288 12724
rect 18052 12640 18104 12646
rect 18104 12600 18184 12628
rect 18052 12582 18104 12588
rect 17868 12368 17920 12374
rect 17868 12310 17920 12316
rect 17960 11620 18012 11626
rect 17960 11562 18012 11568
rect 17972 11082 18000 11562
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 17960 11076 18012 11082
rect 17960 11018 18012 11024
rect 17868 9444 17920 9450
rect 17868 9386 17920 9392
rect 17880 8974 17908 9386
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 17776 8084 17828 8090
rect 17776 8026 17828 8032
rect 17696 7942 17816 7970
rect 17684 7880 17736 7886
rect 17684 7822 17736 7828
rect 17592 7268 17644 7274
rect 17592 7210 17644 7216
rect 17592 6996 17644 7002
rect 17696 6984 17724 7822
rect 17788 7546 17816 7942
rect 17776 7540 17828 7546
rect 17776 7482 17828 7488
rect 17644 6956 17724 6984
rect 17592 6938 17644 6944
rect 17500 6112 17552 6118
rect 17500 6054 17552 6060
rect 17500 5704 17552 5710
rect 17498 5672 17500 5681
rect 17552 5672 17554 5681
rect 17498 5607 17554 5616
rect 17420 5494 17540 5522
rect 17314 3768 17370 3777
rect 17132 3732 17184 3738
rect 17314 3703 17370 3712
rect 17132 3674 17184 3680
rect 17144 3058 17172 3674
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 17040 2644 17092 2650
rect 17040 2586 17092 2592
rect 16948 2508 17000 2514
rect 16948 2450 17000 2456
rect 16488 2440 16540 2446
rect 16488 2382 16540 2388
rect 16960 2310 16988 2450
rect 17512 2428 17540 5494
rect 17604 4593 17632 6938
rect 17774 6488 17830 6497
rect 17774 6423 17776 6432
rect 17828 6423 17830 6432
rect 17776 6394 17828 6400
rect 17880 6361 17908 8774
rect 17682 6352 17738 6361
rect 17682 6287 17738 6296
rect 17866 6352 17922 6361
rect 17866 6287 17922 6296
rect 17696 5914 17724 6287
rect 17684 5908 17736 5914
rect 17684 5850 17736 5856
rect 17972 4706 18000 11018
rect 18064 10266 18092 11494
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 18156 10130 18184 12600
rect 18248 11354 18276 12718
rect 18340 12345 18368 16782
rect 18432 16017 18460 17054
rect 18512 16992 18564 16998
rect 18512 16934 18564 16940
rect 18418 16008 18474 16017
rect 18418 15943 18474 15952
rect 18420 15496 18472 15502
rect 18420 15438 18472 15444
rect 18432 15162 18460 15438
rect 18420 15156 18472 15162
rect 18420 15098 18472 15104
rect 18432 14550 18460 15098
rect 18420 14544 18472 14550
rect 18420 14486 18472 14492
rect 18420 13728 18472 13734
rect 18420 13670 18472 13676
rect 18432 13326 18460 13670
rect 18420 13320 18472 13326
rect 18420 13262 18472 13268
rect 18432 12986 18460 13262
rect 18420 12980 18472 12986
rect 18420 12922 18472 12928
rect 18420 12368 18472 12374
rect 18326 12336 18382 12345
rect 18420 12310 18472 12316
rect 18326 12271 18382 12280
rect 18236 11348 18288 11354
rect 18236 11290 18288 11296
rect 18248 11150 18276 11290
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 18144 10124 18196 10130
rect 18144 10066 18196 10072
rect 18052 9920 18104 9926
rect 18052 9862 18104 9868
rect 17696 4678 18000 4706
rect 17590 4584 17646 4593
rect 17590 4519 17646 4528
rect 17696 3398 17724 4678
rect 18064 4672 18092 9862
rect 18156 9722 18184 10066
rect 18144 9716 18196 9722
rect 18144 9658 18196 9664
rect 18340 9654 18368 12271
rect 18328 9648 18380 9654
rect 18328 9590 18380 9596
rect 18236 9512 18288 9518
rect 18236 9454 18288 9460
rect 18144 9376 18196 9382
rect 18248 9353 18276 9454
rect 18144 9318 18196 9324
rect 18234 9344 18290 9353
rect 18156 5681 18184 9318
rect 18234 9279 18290 9288
rect 18236 8832 18288 8838
rect 18236 8774 18288 8780
rect 18248 8362 18276 8774
rect 18236 8356 18288 8362
rect 18236 8298 18288 8304
rect 18248 7342 18276 8298
rect 18328 8016 18380 8022
rect 18326 7984 18328 7993
rect 18380 7984 18382 7993
rect 18326 7919 18382 7928
rect 18236 7336 18288 7342
rect 18236 7278 18288 7284
rect 18340 7206 18368 7919
rect 18432 7886 18460 12310
rect 18524 10690 18552 16934
rect 18616 16726 18644 18090
rect 18604 16720 18656 16726
rect 18604 16662 18656 16668
rect 18604 15972 18656 15978
rect 18604 15914 18656 15920
rect 18616 15366 18644 15914
rect 18604 15360 18656 15366
rect 18604 15302 18656 15308
rect 18604 14952 18656 14958
rect 18604 14894 18656 14900
rect 18616 14414 18644 14894
rect 18604 14408 18656 14414
rect 18604 14350 18656 14356
rect 18616 13462 18644 14350
rect 18604 13456 18656 13462
rect 18604 13398 18656 13404
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 18616 11286 18644 11698
rect 18604 11280 18656 11286
rect 18604 11222 18656 11228
rect 18708 11121 18736 22646
rect 18786 21992 18842 22001
rect 18786 21927 18842 21936
rect 18694 11112 18750 11121
rect 18694 11047 18750 11056
rect 18696 10804 18748 10810
rect 18696 10746 18748 10752
rect 18524 10662 18644 10690
rect 18512 10600 18564 10606
rect 18512 10542 18564 10548
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 18328 7200 18380 7206
rect 18328 7142 18380 7148
rect 18328 6384 18380 6390
rect 18328 6326 18380 6332
rect 18340 6118 18368 6326
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18328 6112 18380 6118
rect 18328 6054 18380 6060
rect 18234 5944 18290 5953
rect 18290 5902 18368 5930
rect 18234 5879 18236 5888
rect 18288 5879 18290 5888
rect 18236 5850 18288 5856
rect 18236 5772 18288 5778
rect 18236 5714 18288 5720
rect 18142 5672 18198 5681
rect 18142 5607 18198 5616
rect 18248 5370 18276 5714
rect 18340 5370 18368 5902
rect 18432 5710 18460 6190
rect 18420 5704 18472 5710
rect 18420 5646 18472 5652
rect 18236 5364 18288 5370
rect 18236 5306 18288 5312
rect 18328 5364 18380 5370
rect 18328 5306 18380 5312
rect 18064 4644 18184 4672
rect 17960 4616 18012 4622
rect 17866 4584 17922 4593
rect 18012 4576 18092 4604
rect 17960 4558 18012 4564
rect 17866 4519 17868 4528
rect 17920 4519 17922 4528
rect 17868 4490 17920 4496
rect 17960 4480 18012 4486
rect 17960 4422 18012 4428
rect 17684 3392 17736 3398
rect 17684 3334 17736 3340
rect 17776 3392 17828 3398
rect 17776 3334 17828 3340
rect 17788 2990 17816 3334
rect 17972 2990 18000 4422
rect 18064 3738 18092 4576
rect 18052 3732 18104 3738
rect 18052 3674 18104 3680
rect 18050 3496 18106 3505
rect 18050 3431 18106 3440
rect 18064 3194 18092 3431
rect 18052 3188 18104 3194
rect 18052 3130 18104 3136
rect 18156 3097 18184 4644
rect 18248 4185 18276 5306
rect 18432 5114 18460 5646
rect 18340 5098 18460 5114
rect 18328 5092 18460 5098
rect 18380 5086 18460 5092
rect 18328 5034 18380 5040
rect 18340 4690 18368 5034
rect 18418 4720 18474 4729
rect 18328 4684 18380 4690
rect 18418 4655 18474 4664
rect 18328 4626 18380 4632
rect 18340 4593 18368 4626
rect 18326 4584 18382 4593
rect 18326 4519 18382 4528
rect 18340 4214 18368 4519
rect 18432 4282 18460 4655
rect 18420 4276 18472 4282
rect 18420 4218 18472 4224
rect 18328 4208 18380 4214
rect 18234 4176 18290 4185
rect 18328 4150 18380 4156
rect 18234 4111 18290 4120
rect 18418 3904 18474 3913
rect 18418 3839 18474 3848
rect 18432 3466 18460 3839
rect 18420 3460 18472 3466
rect 18420 3402 18472 3408
rect 18142 3088 18198 3097
rect 18142 3023 18198 3032
rect 17776 2984 17828 2990
rect 17774 2952 17776 2961
rect 17960 2984 18012 2990
rect 17828 2952 17830 2961
rect 17960 2926 18012 2932
rect 18420 2984 18472 2990
rect 18420 2926 18472 2932
rect 17774 2887 17830 2896
rect 18326 2680 18382 2689
rect 18326 2615 18328 2624
rect 18380 2615 18382 2624
rect 18328 2586 18380 2592
rect 18432 2553 18460 2926
rect 18234 2544 18290 2553
rect 18234 2479 18290 2488
rect 18418 2544 18474 2553
rect 18418 2479 18474 2488
rect 17052 2400 17540 2428
rect 18248 2428 18276 2479
rect 18248 2400 18460 2428
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 16672 2304 16724 2310
rect 16948 2304 17000 2310
rect 16672 2246 16724 2252
rect 16762 2272 16818 2281
rect 16684 2145 16712 2246
rect 16762 2207 16818 2216
rect 16946 2272 16948 2281
rect 17000 2272 17002 2281
rect 16946 2207 17002 2216
rect 16670 2136 16726 2145
rect 16670 2071 16726 2080
rect 16776 1601 16804 2207
rect 16762 1592 16818 1601
rect 16762 1527 16818 1536
rect 17052 1442 17080 2400
rect 17132 2304 17184 2310
rect 17132 2246 17184 2252
rect 17592 2304 17644 2310
rect 17592 2246 17644 2252
rect 16592 1414 17080 1442
rect 16592 480 16620 1414
rect 17144 480 17172 2246
rect 17604 1329 17632 2246
rect 18432 2009 18460 2400
rect 18234 2000 18290 2009
rect 18234 1935 18290 1944
rect 18418 2000 18474 2009
rect 18418 1935 18474 1944
rect 17682 1864 17738 1873
rect 17682 1799 17738 1808
rect 17590 1320 17646 1329
rect 17590 1255 17646 1264
rect 17696 480 17724 1799
rect 18248 480 18276 1935
rect 18524 1873 18552 10542
rect 18616 8514 18644 10662
rect 18708 8673 18736 10746
rect 18694 8664 18750 8673
rect 18694 8599 18750 8608
rect 18616 8486 18736 8514
rect 18604 7744 18656 7750
rect 18604 7686 18656 7692
rect 18616 7274 18644 7686
rect 18604 7268 18656 7274
rect 18604 7210 18656 7216
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 18616 6458 18644 6734
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 18708 5953 18736 8486
rect 18800 8090 18828 21927
rect 18892 11529 18920 23208
rect 18984 23118 19012 23666
rect 19156 23588 19208 23594
rect 19156 23530 19208 23536
rect 19064 23248 19116 23254
rect 19064 23190 19116 23196
rect 18972 23112 19024 23118
rect 18972 23054 19024 23060
rect 19076 22778 19104 23190
rect 19064 22772 19116 22778
rect 19064 22714 19116 22720
rect 18970 22264 19026 22273
rect 18970 22199 19026 22208
rect 18984 21729 19012 22199
rect 19064 22160 19116 22166
rect 19064 22102 19116 22108
rect 18970 21720 19026 21729
rect 18970 21655 19026 21664
rect 19076 21350 19104 22102
rect 19064 21344 19116 21350
rect 19064 21286 19116 21292
rect 19076 21185 19104 21286
rect 19062 21176 19118 21185
rect 19062 21111 19118 21120
rect 18972 20936 19024 20942
rect 18972 20878 19024 20884
rect 19062 20904 19118 20913
rect 18984 20602 19012 20878
rect 19062 20839 19118 20848
rect 18972 20596 19024 20602
rect 18972 20538 19024 20544
rect 18984 20233 19012 20538
rect 18970 20224 19026 20233
rect 18970 20159 19026 20168
rect 18972 20052 19024 20058
rect 18972 19994 19024 20000
rect 18984 18170 19012 19994
rect 19076 18426 19104 20839
rect 19064 18420 19116 18426
rect 19064 18362 19116 18368
rect 18984 18142 19104 18170
rect 18972 17536 19024 17542
rect 18972 17478 19024 17484
rect 18984 17241 19012 17478
rect 18970 17232 19026 17241
rect 18970 17167 18972 17176
rect 19024 17167 19026 17176
rect 18972 17138 19024 17144
rect 18984 17107 19012 17138
rect 18972 16992 19024 16998
rect 18972 16934 19024 16940
rect 18984 14482 19012 16934
rect 19076 16425 19104 18142
rect 19062 16416 19118 16425
rect 19062 16351 19118 16360
rect 18972 14476 19024 14482
rect 18972 14418 19024 14424
rect 18972 12096 19024 12102
rect 18972 12038 19024 12044
rect 18984 11937 19012 12038
rect 18970 11928 19026 11937
rect 18970 11863 19026 11872
rect 18970 11792 19026 11801
rect 18970 11727 19026 11736
rect 18878 11520 18934 11529
rect 18878 11455 18934 11464
rect 18880 11212 18932 11218
rect 18880 11154 18932 11160
rect 18892 11121 18920 11154
rect 18878 11112 18934 11121
rect 18878 11047 18934 11056
rect 18984 10554 19012 11727
rect 19076 10810 19104 16351
rect 19168 11801 19196 23530
rect 19260 23225 19288 24618
rect 19340 24608 19392 24614
rect 19340 24550 19392 24556
rect 19246 23216 19302 23225
rect 19246 23151 19302 23160
rect 19248 22432 19300 22438
rect 19246 22400 19248 22409
rect 19300 22400 19302 22409
rect 19246 22335 19302 22344
rect 19248 21888 19300 21894
rect 19248 21830 19300 21836
rect 19260 20448 19288 21830
rect 19352 20618 19380 24550
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19996 24410 20024 24822
rect 20088 24614 20116 26386
rect 20640 26081 20668 27520
rect 21088 26852 21140 26858
rect 21088 26794 21140 26800
rect 20626 26072 20682 26081
rect 20626 26007 20682 26016
rect 20628 25356 20680 25362
rect 20628 25298 20680 25304
rect 20076 24608 20128 24614
rect 20076 24550 20128 24556
rect 20536 24608 20588 24614
rect 20640 24596 20668 25298
rect 20996 25152 21048 25158
rect 20996 25094 21048 25100
rect 21008 24750 21036 25094
rect 20996 24744 21048 24750
rect 20996 24686 21048 24692
rect 21100 24614 21128 26794
rect 21284 25702 21312 27520
rect 21272 25696 21324 25702
rect 21272 25638 21324 25644
rect 21180 25356 21232 25362
rect 21180 25298 21232 25304
rect 21192 24857 21220 25298
rect 21362 25256 21418 25265
rect 21836 25226 21864 27520
rect 22388 25974 22416 27520
rect 23032 26194 23060 27520
rect 22664 26166 23060 26194
rect 22376 25968 22428 25974
rect 22376 25910 22428 25916
rect 22468 25832 22520 25838
rect 22468 25774 22520 25780
rect 22192 25696 22244 25702
rect 22192 25638 22244 25644
rect 21362 25191 21418 25200
rect 21824 25220 21876 25226
rect 21270 25120 21326 25129
rect 21270 25055 21326 25064
rect 21178 24848 21234 24857
rect 21178 24783 21180 24792
rect 21232 24783 21234 24792
rect 21180 24754 21232 24760
rect 20720 24608 20772 24614
rect 20640 24576 20720 24596
rect 21088 24608 21140 24614
rect 20772 24576 20774 24585
rect 20640 24568 20718 24576
rect 20536 24550 20588 24556
rect 19984 24404 20036 24410
rect 19984 24346 20036 24352
rect 19982 24304 20038 24313
rect 19982 24239 20038 24248
rect 20352 24268 20404 24274
rect 19432 23520 19484 23526
rect 19430 23488 19432 23497
rect 19484 23488 19486 23497
rect 19430 23423 19486 23432
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19800 23112 19852 23118
rect 19800 23054 19852 23060
rect 19614 22944 19670 22953
rect 19614 22879 19670 22888
rect 19628 22778 19656 22879
rect 19616 22772 19668 22778
rect 19616 22714 19668 22720
rect 19812 22642 19840 23054
rect 19996 22692 20024 24239
rect 20352 24210 20404 24216
rect 20364 24070 20392 24210
rect 20352 24064 20404 24070
rect 20352 24006 20404 24012
rect 20168 23792 20220 23798
rect 20168 23734 20220 23740
rect 20180 23633 20208 23734
rect 20166 23624 20222 23633
rect 20076 23588 20128 23594
rect 20166 23559 20222 23568
rect 20076 23530 20128 23536
rect 20088 23497 20116 23530
rect 20260 23520 20312 23526
rect 20074 23488 20130 23497
rect 20260 23462 20312 23468
rect 20074 23423 20130 23432
rect 20168 22976 20220 22982
rect 20272 22964 20300 23462
rect 20364 23361 20392 24006
rect 20442 23896 20498 23905
rect 20442 23831 20498 23840
rect 20350 23352 20406 23361
rect 20350 23287 20406 23296
rect 20220 22936 20300 22964
rect 20168 22918 20220 22924
rect 20180 22817 20208 22918
rect 20166 22808 20222 22817
rect 20166 22743 20222 22752
rect 19996 22664 20300 22692
rect 19800 22636 19852 22642
rect 19800 22578 19852 22584
rect 19524 22500 19576 22506
rect 19524 22442 19576 22448
rect 19536 22098 19564 22442
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19524 22092 19576 22098
rect 19524 22034 19576 22040
rect 19432 21548 19484 21554
rect 19432 21490 19484 21496
rect 19444 21146 19472 21490
rect 19536 21457 19564 22034
rect 19984 21616 20036 21622
rect 19984 21558 20036 21564
rect 19522 21448 19578 21457
rect 19522 21383 19578 21392
rect 19524 21344 19576 21350
rect 19524 21286 19576 21292
rect 19432 21140 19484 21146
rect 19432 21082 19484 21088
rect 19536 20788 19564 21286
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19616 20800 19668 20806
rect 19536 20768 19616 20788
rect 19708 20800 19760 20806
rect 19668 20768 19670 20777
rect 19536 20760 19614 20768
rect 19708 20742 19760 20748
rect 19614 20703 19670 20712
rect 19352 20590 19472 20618
rect 19340 20460 19392 20466
rect 19260 20420 19340 20448
rect 19340 20402 19392 20408
rect 19248 19712 19300 19718
rect 19248 19654 19300 19660
rect 19260 19242 19288 19654
rect 19248 19236 19300 19242
rect 19248 19178 19300 19184
rect 19352 18970 19380 20402
rect 19444 19310 19472 20590
rect 19720 20346 19748 20742
rect 19536 20318 19748 20346
rect 19432 19304 19484 19310
rect 19432 19246 19484 19252
rect 19248 18964 19300 18970
rect 19248 18906 19300 18912
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 19260 18034 19288 18906
rect 19444 18850 19472 19246
rect 19352 18822 19472 18850
rect 19536 18850 19564 20318
rect 19996 20262 20024 21558
rect 20074 21312 20130 21321
rect 20074 21247 20130 21256
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19996 19961 20024 20198
rect 19982 19952 20038 19961
rect 19982 19887 20038 19896
rect 19984 19168 20036 19174
rect 19984 19110 20036 19116
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19536 18822 19840 18850
rect 19352 18154 19380 18822
rect 19616 18760 19668 18766
rect 19616 18702 19668 18708
rect 19432 18624 19484 18630
rect 19432 18566 19484 18572
rect 19340 18148 19392 18154
rect 19340 18090 19392 18096
rect 19260 18006 19380 18034
rect 19352 17882 19380 18006
rect 19444 17921 19472 18566
rect 19628 18068 19656 18702
rect 19536 18040 19656 18068
rect 19812 18068 19840 18822
rect 19996 18222 20024 19110
rect 19984 18216 20036 18222
rect 19984 18158 20036 18164
rect 19812 18040 20024 18068
rect 19430 17912 19486 17921
rect 19340 17876 19392 17882
rect 19430 17847 19486 17856
rect 19536 17864 19564 18040
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19536 17836 19656 17864
rect 19340 17818 19392 17824
rect 19248 17808 19300 17814
rect 19248 17750 19300 17756
rect 19260 17134 19288 17750
rect 19524 17740 19576 17746
rect 19524 17682 19576 17688
rect 19248 17128 19300 17134
rect 19248 17070 19300 17076
rect 19430 16824 19486 16833
rect 19536 16794 19564 17682
rect 19628 17610 19656 17836
rect 19708 17672 19760 17678
rect 19708 17614 19760 17620
rect 19616 17604 19668 17610
rect 19616 17546 19668 17552
rect 19720 17338 19748 17614
rect 19708 17332 19760 17338
rect 19708 17274 19760 17280
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19430 16759 19486 16768
rect 19524 16788 19576 16794
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 19260 16114 19288 16594
rect 19248 16108 19300 16114
rect 19248 16050 19300 16056
rect 19340 15904 19392 15910
rect 19340 15846 19392 15852
rect 19248 15020 19300 15026
rect 19352 15008 19380 15846
rect 19444 15706 19472 16759
rect 19524 16730 19576 16736
rect 19524 16448 19576 16454
rect 19524 16390 19576 16396
rect 19432 15700 19484 15706
rect 19432 15642 19484 15648
rect 19444 15026 19472 15642
rect 19536 15366 19564 16390
rect 19996 16096 20024 18040
rect 20088 17338 20116 21247
rect 20168 20460 20220 20466
rect 20168 20402 20220 20408
rect 20180 19718 20208 20402
rect 20168 19712 20220 19718
rect 20168 19654 20220 19660
rect 20166 19136 20222 19145
rect 20166 19071 20222 19080
rect 20180 18601 20208 19071
rect 20166 18592 20222 18601
rect 20166 18527 20222 18536
rect 20166 17368 20222 17377
rect 20076 17332 20128 17338
rect 20166 17303 20222 17312
rect 20076 17274 20128 17280
rect 19996 16068 20116 16096
rect 19982 16008 20038 16017
rect 19982 15943 20038 15952
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19708 15496 19760 15502
rect 19708 15438 19760 15444
rect 19524 15360 19576 15366
rect 19524 15302 19576 15308
rect 19300 14980 19380 15008
rect 19432 15020 19484 15026
rect 19248 14962 19300 14968
rect 19432 14962 19484 14968
rect 19340 14884 19392 14890
rect 19340 14826 19392 14832
rect 19352 14618 19380 14826
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 19246 14104 19302 14113
rect 19246 14039 19302 14048
rect 19154 11792 19210 11801
rect 19154 11727 19210 11736
rect 19260 11665 19288 14039
rect 19352 13161 19380 14554
rect 19338 13152 19394 13161
rect 19338 13087 19394 13096
rect 19536 13025 19564 15302
rect 19720 14890 19748 15438
rect 19708 14884 19760 14890
rect 19708 14826 19760 14832
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19996 14618 20024 15943
rect 20088 15337 20116 16068
rect 20074 15328 20130 15337
rect 20074 15263 20130 15272
rect 20088 14770 20116 15263
rect 20180 15201 20208 17303
rect 20166 15192 20222 15201
rect 20166 15127 20222 15136
rect 20088 14742 20208 14770
rect 20074 14648 20130 14657
rect 19984 14612 20036 14618
rect 20074 14583 20130 14592
rect 19984 14554 20036 14560
rect 20088 14482 20116 14583
rect 20076 14476 20128 14482
rect 20076 14418 20128 14424
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 20088 13462 20116 14418
rect 20076 13456 20128 13462
rect 20076 13398 20128 13404
rect 20180 13274 20208 14742
rect 19996 13246 20208 13274
rect 19522 13016 19578 13025
rect 19522 12951 19578 12960
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19524 12300 19576 12306
rect 19524 12242 19576 12248
rect 19246 11656 19302 11665
rect 19246 11591 19302 11600
rect 19246 10976 19302 10985
rect 19246 10911 19302 10920
rect 19064 10804 19116 10810
rect 19064 10746 19116 10752
rect 18892 10526 19012 10554
rect 18892 10033 18920 10526
rect 18972 10464 19024 10470
rect 19024 10424 19104 10452
rect 18972 10406 19024 10412
rect 18878 10024 18934 10033
rect 18878 9959 18934 9968
rect 18972 9104 19024 9110
rect 18972 9046 19024 9052
rect 18984 8634 19012 9046
rect 18972 8628 19024 8634
rect 18972 8570 19024 8576
rect 18984 8090 19012 8570
rect 18788 8084 18840 8090
rect 18788 8026 18840 8032
rect 18972 8084 19024 8090
rect 18972 8026 19024 8032
rect 18880 7948 18932 7954
rect 18880 7890 18932 7896
rect 18788 7336 18840 7342
rect 18788 7278 18840 7284
rect 18800 6798 18828 7278
rect 18892 7002 18920 7890
rect 18972 7540 19024 7546
rect 18972 7482 19024 7488
rect 18880 6996 18932 7002
rect 18880 6938 18932 6944
rect 18788 6792 18840 6798
rect 18788 6734 18840 6740
rect 18694 5944 18750 5953
rect 18694 5879 18750 5888
rect 18984 5817 19012 7482
rect 18970 5808 19026 5817
rect 18970 5743 19026 5752
rect 18788 5636 18840 5642
rect 18788 5578 18840 5584
rect 18696 5160 18748 5166
rect 18696 5102 18748 5108
rect 18708 4758 18736 5102
rect 18696 4752 18748 4758
rect 18696 4694 18748 4700
rect 18800 4146 18828 5578
rect 18788 4140 18840 4146
rect 18788 4082 18840 4088
rect 18696 4004 18748 4010
rect 18696 3946 18748 3952
rect 18708 3369 18736 3946
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18800 3670 18828 3878
rect 18880 3732 18932 3738
rect 18880 3674 18932 3680
rect 18788 3664 18840 3670
rect 18788 3606 18840 3612
rect 18694 3360 18750 3369
rect 18694 3295 18750 3304
rect 18708 2990 18736 3295
rect 18800 3194 18828 3606
rect 18892 3233 18920 3674
rect 18970 3496 19026 3505
rect 18970 3431 19026 3440
rect 18878 3224 18934 3233
rect 18788 3188 18840 3194
rect 18878 3159 18934 3168
rect 18788 3130 18840 3136
rect 18880 3052 18932 3058
rect 18880 2994 18932 3000
rect 18696 2984 18748 2990
rect 18696 2926 18748 2932
rect 18892 2446 18920 2994
rect 18880 2440 18932 2446
rect 18880 2382 18932 2388
rect 18984 2258 19012 3431
rect 19076 2961 19104 10424
rect 19260 10266 19288 10911
rect 19536 10810 19564 12242
rect 19996 11801 20024 13246
rect 20076 12912 20128 12918
rect 20074 12880 20076 12889
rect 20128 12880 20130 12889
rect 20074 12815 20130 12824
rect 20272 12782 20300 22664
rect 20352 22568 20404 22574
rect 20352 22510 20404 22516
rect 20364 20806 20392 22510
rect 20352 20800 20404 20806
rect 20352 20742 20404 20748
rect 20350 20496 20406 20505
rect 20350 20431 20406 20440
rect 20364 20233 20392 20431
rect 20350 20224 20406 20233
rect 20350 20159 20406 20168
rect 20350 17776 20406 17785
rect 20350 17711 20406 17720
rect 20364 17377 20392 17711
rect 20350 17368 20406 17377
rect 20350 17303 20406 17312
rect 20456 17082 20484 23831
rect 20548 23497 20576 24550
rect 21088 24550 21140 24556
rect 20718 24511 20774 24520
rect 21284 24274 21312 25055
rect 21376 24410 21404 25191
rect 21824 25162 21876 25168
rect 22204 24886 22232 25638
rect 22480 25294 22508 25774
rect 22468 25288 22520 25294
rect 22468 25230 22520 25236
rect 22466 24984 22522 24993
rect 22664 24954 22692 26166
rect 23584 25378 23612 27520
rect 23938 25392 23994 25401
rect 22744 25356 22796 25362
rect 22744 25298 22796 25304
rect 22928 25356 22980 25362
rect 23584 25350 23704 25378
rect 22928 25298 22980 25304
rect 22466 24919 22522 24928
rect 22652 24948 22704 24954
rect 22192 24880 22244 24886
rect 22192 24822 22244 24828
rect 22480 24818 22508 24919
rect 22652 24890 22704 24896
rect 22468 24812 22520 24818
rect 22468 24754 22520 24760
rect 22652 24812 22704 24818
rect 22652 24754 22704 24760
rect 21456 24744 21508 24750
rect 21456 24686 21508 24692
rect 21364 24404 21416 24410
rect 21364 24346 21416 24352
rect 21272 24268 21324 24274
rect 21272 24210 21324 24216
rect 20720 24200 20772 24206
rect 20720 24142 20772 24148
rect 21086 24168 21142 24177
rect 20534 23488 20590 23497
rect 20534 23423 20590 23432
rect 20732 23322 20760 24142
rect 21086 24103 21142 24112
rect 20904 24064 20956 24070
rect 20904 24006 20956 24012
rect 20916 23662 20944 24006
rect 20904 23656 20956 23662
rect 20904 23598 20956 23604
rect 20720 23316 20772 23322
rect 20720 23258 20772 23264
rect 20720 22976 20772 22982
rect 20720 22918 20772 22924
rect 20732 22574 20760 22918
rect 20916 22778 20944 23598
rect 20904 22772 20956 22778
rect 20904 22714 20956 22720
rect 20720 22568 20772 22574
rect 20720 22510 20772 22516
rect 20904 22160 20956 22166
rect 20902 22128 20904 22137
rect 20956 22128 20958 22137
rect 20902 22063 20958 22072
rect 20536 21888 20588 21894
rect 20536 21830 20588 21836
rect 20548 21554 20576 21830
rect 20718 21584 20774 21593
rect 20536 21548 20588 21554
rect 20718 21519 20720 21528
rect 20536 21490 20588 21496
rect 20772 21519 20774 21528
rect 20720 21490 20772 21496
rect 20548 20806 20576 21490
rect 20902 21448 20958 21457
rect 20902 21383 20958 21392
rect 20916 21350 20944 21383
rect 20904 21344 20956 21350
rect 20904 21286 20956 21292
rect 20812 21140 20864 21146
rect 20812 21082 20864 21088
rect 20720 21004 20772 21010
rect 20720 20946 20772 20952
rect 20536 20800 20588 20806
rect 20536 20742 20588 20748
rect 20548 19990 20576 20742
rect 20732 20602 20760 20946
rect 20720 20596 20772 20602
rect 20720 20538 20772 20544
rect 20732 20505 20760 20538
rect 20718 20496 20774 20505
rect 20718 20431 20774 20440
rect 20536 19984 20588 19990
rect 20536 19926 20588 19932
rect 20536 19712 20588 19718
rect 20536 19654 20588 19660
rect 20364 17054 20484 17082
rect 20364 13530 20392 17054
rect 20444 16992 20496 16998
rect 20444 16934 20496 16940
rect 20456 16726 20484 16934
rect 20444 16720 20496 16726
rect 20444 16662 20496 16668
rect 20444 15156 20496 15162
rect 20444 15098 20496 15104
rect 20456 14929 20484 15098
rect 20442 14920 20498 14929
rect 20442 14855 20498 14864
rect 20352 13524 20404 13530
rect 20352 13466 20404 13472
rect 20548 12832 20576 19654
rect 20824 19446 20852 21082
rect 20996 20936 21048 20942
rect 20902 20904 20958 20913
rect 20996 20878 21048 20884
rect 20902 20839 20904 20848
rect 20956 20839 20958 20848
rect 20904 20810 20956 20816
rect 21008 20602 21036 20878
rect 20996 20596 21048 20602
rect 20996 20538 21048 20544
rect 20812 19440 20864 19446
rect 20812 19382 20864 19388
rect 21008 19378 21036 20538
rect 20996 19372 21048 19378
rect 20996 19314 21048 19320
rect 20902 19272 20958 19281
rect 20902 19207 20958 19216
rect 20996 19236 21048 19242
rect 20916 18630 20944 19207
rect 20996 19178 21048 19184
rect 20904 18624 20956 18630
rect 20904 18566 20956 18572
rect 20718 18456 20774 18465
rect 20718 18391 20774 18400
rect 20732 18086 20760 18391
rect 20904 18148 20956 18154
rect 20904 18090 20956 18096
rect 20720 18080 20772 18086
rect 20720 18022 20772 18028
rect 20916 17134 20944 18090
rect 21008 17649 21036 19178
rect 21100 18834 21128 24103
rect 21284 23594 21312 24210
rect 21376 23866 21404 24346
rect 21364 23860 21416 23866
rect 21364 23802 21416 23808
rect 21272 23588 21324 23594
rect 21272 23530 21324 23536
rect 21364 23180 21416 23186
rect 21364 23122 21416 23128
rect 21376 22438 21404 23122
rect 21364 22432 21416 22438
rect 21364 22374 21416 22380
rect 21180 22228 21232 22234
rect 21180 22170 21232 22176
rect 21192 21690 21220 22170
rect 21468 22114 21496 24686
rect 21824 24676 21876 24682
rect 21824 24618 21876 24624
rect 21836 24585 21864 24618
rect 21916 24608 21968 24614
rect 21822 24576 21878 24585
rect 21916 24550 21968 24556
rect 21822 24511 21878 24520
rect 21824 24064 21876 24070
rect 21824 24006 21876 24012
rect 21732 22568 21784 22574
rect 21732 22510 21784 22516
rect 21548 22432 21600 22438
rect 21548 22374 21600 22380
rect 21560 22234 21588 22374
rect 21744 22234 21772 22510
rect 21548 22228 21600 22234
rect 21548 22170 21600 22176
rect 21732 22228 21784 22234
rect 21732 22170 21784 22176
rect 21468 22086 21588 22114
rect 21180 21684 21232 21690
rect 21180 21626 21232 21632
rect 21456 21616 21508 21622
rect 21456 21558 21508 21564
rect 21180 21072 21232 21078
rect 21180 21014 21232 21020
rect 21192 20602 21220 21014
rect 21180 20596 21232 20602
rect 21180 20538 21232 20544
rect 21270 20360 21326 20369
rect 21270 20295 21326 20304
rect 21284 19990 21312 20295
rect 21272 19984 21324 19990
rect 21272 19926 21324 19932
rect 21180 19168 21232 19174
rect 21180 19110 21232 19116
rect 21192 18902 21220 19110
rect 21284 18970 21312 19926
rect 21364 19848 21416 19854
rect 21364 19790 21416 19796
rect 21376 19689 21404 19790
rect 21468 19718 21496 21558
rect 21456 19712 21508 19718
rect 21362 19680 21418 19689
rect 21456 19654 21508 19660
rect 21362 19615 21418 19624
rect 21376 19514 21404 19615
rect 21364 19508 21416 19514
rect 21364 19450 21416 19456
rect 21456 19168 21508 19174
rect 21456 19110 21508 19116
rect 21272 18964 21324 18970
rect 21272 18906 21324 18912
rect 21180 18896 21232 18902
rect 21180 18838 21232 18844
rect 21088 18828 21140 18834
rect 21088 18770 21140 18776
rect 21364 18760 21416 18766
rect 21364 18702 21416 18708
rect 21086 18184 21142 18193
rect 21086 18119 21142 18128
rect 20994 17640 21050 17649
rect 20994 17575 21050 17584
rect 20996 17536 21048 17542
rect 20996 17478 21048 17484
rect 20904 17128 20956 17134
rect 20904 17070 20956 17076
rect 20720 16788 20772 16794
rect 20720 16730 20772 16736
rect 20626 16416 20682 16425
rect 20626 16351 20682 16360
rect 20640 15910 20668 16351
rect 20732 16250 20760 16730
rect 20916 16590 20944 17070
rect 20904 16584 20956 16590
rect 20904 16526 20956 16532
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 21008 16046 21036 17478
rect 20996 16040 21048 16046
rect 20996 15982 21048 15988
rect 20628 15904 20680 15910
rect 20628 15846 20680 15852
rect 21008 15706 21036 15982
rect 20996 15700 21048 15706
rect 20996 15642 21048 15648
rect 20720 15632 20772 15638
rect 20720 15574 20772 15580
rect 20626 15464 20682 15473
rect 20626 15399 20682 15408
rect 20640 14958 20668 15399
rect 20732 15162 20760 15574
rect 20904 15360 20956 15366
rect 20810 15328 20866 15337
rect 20904 15302 20956 15308
rect 20810 15263 20866 15272
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20628 14952 20680 14958
rect 20628 14894 20680 14900
rect 20640 14618 20668 14894
rect 20628 14612 20680 14618
rect 20628 14554 20680 14560
rect 20824 14074 20852 15263
rect 20916 15065 20944 15302
rect 20902 15056 20958 15065
rect 20902 14991 20958 15000
rect 20994 14376 21050 14385
rect 20994 14311 21050 14320
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20718 13968 20774 13977
rect 20718 13903 20720 13912
rect 20772 13903 20774 13912
rect 20720 13874 20772 13880
rect 20812 13388 20864 13394
rect 20812 13330 20864 13336
rect 20548 12804 20760 12832
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 20536 12640 20588 12646
rect 20536 12582 20588 12588
rect 20076 12232 20128 12238
rect 20076 12174 20128 12180
rect 19982 11792 20038 11801
rect 19982 11727 20038 11736
rect 19984 11688 20036 11694
rect 19984 11630 20036 11636
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19890 11248 19946 11257
rect 19890 11183 19892 11192
rect 19944 11183 19946 11192
rect 19892 11154 19944 11160
rect 19524 10804 19576 10810
rect 19524 10746 19576 10752
rect 19904 10742 19932 11154
rect 19800 10736 19852 10742
rect 19800 10678 19852 10684
rect 19892 10736 19944 10742
rect 19892 10678 19944 10684
rect 19812 10606 19840 10678
rect 19800 10600 19852 10606
rect 19800 10542 19852 10548
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19338 10296 19394 10305
rect 19248 10260 19300 10266
rect 19622 10288 19918 10308
rect 19338 10231 19394 10240
rect 19432 10260 19484 10266
rect 19248 10202 19300 10208
rect 19248 10124 19300 10130
rect 19248 10066 19300 10072
rect 19156 10056 19208 10062
rect 19156 9998 19208 10004
rect 19168 9722 19196 9998
rect 19260 9722 19288 10066
rect 19156 9716 19208 9722
rect 19156 9658 19208 9664
rect 19248 9716 19300 9722
rect 19248 9658 19300 9664
rect 19352 8650 19380 10231
rect 19432 10202 19484 10208
rect 19444 9450 19472 10202
rect 19996 10062 20024 11630
rect 20088 11626 20116 12174
rect 20444 12096 20496 12102
rect 20444 12038 20496 12044
rect 20456 11762 20484 12038
rect 20260 11756 20312 11762
rect 20260 11698 20312 11704
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 20272 11665 20300 11698
rect 20258 11656 20314 11665
rect 20076 11620 20128 11626
rect 20258 11591 20314 11600
rect 20076 11562 20128 11568
rect 20088 11150 20116 11562
rect 20168 11348 20220 11354
rect 20168 11290 20220 11296
rect 20076 11144 20128 11150
rect 20076 11086 20128 11092
rect 20180 10062 20208 11290
rect 20444 11280 20496 11286
rect 20444 11222 20496 11228
rect 20352 11076 20404 11082
rect 20352 11018 20404 11024
rect 20258 10704 20314 10713
rect 20258 10639 20260 10648
rect 20312 10639 20314 10648
rect 20260 10610 20312 10616
rect 20272 10198 20300 10610
rect 20364 10266 20392 11018
rect 20352 10260 20404 10266
rect 20352 10202 20404 10208
rect 20260 10192 20312 10198
rect 20260 10134 20312 10140
rect 19984 10056 20036 10062
rect 19984 9998 20036 10004
rect 20168 10056 20220 10062
rect 20168 9998 20220 10004
rect 19522 9616 19578 9625
rect 19522 9551 19578 9560
rect 19432 9444 19484 9450
rect 19432 9386 19484 9392
rect 19536 8974 19564 9551
rect 19996 9450 20024 9998
rect 20456 9704 20484 11222
rect 20548 10266 20576 12582
rect 20628 11620 20680 11626
rect 20628 11562 20680 11568
rect 20640 11354 20668 11562
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 20732 11286 20760 12804
rect 20824 12646 20852 13330
rect 21008 12986 21036 14311
rect 21100 13530 21128 18119
rect 21272 18080 21324 18086
rect 21376 18057 21404 18702
rect 21468 18698 21496 19110
rect 21560 19009 21588 22086
rect 21836 22080 21864 24006
rect 21744 22052 21864 22080
rect 21640 20256 21692 20262
rect 21640 20198 21692 20204
rect 21652 20058 21680 20198
rect 21640 20052 21692 20058
rect 21640 19994 21692 20000
rect 21744 19786 21772 22052
rect 21824 21956 21876 21962
rect 21824 21898 21876 21904
rect 21836 21554 21864 21898
rect 21824 21548 21876 21554
rect 21824 21490 21876 21496
rect 21836 21010 21864 21490
rect 21824 21004 21876 21010
rect 21824 20946 21876 20952
rect 21928 20097 21956 24550
rect 22480 24410 22508 24754
rect 22560 24608 22612 24614
rect 22560 24550 22612 24556
rect 22468 24404 22520 24410
rect 22468 24346 22520 24352
rect 22374 24304 22430 24313
rect 22374 24239 22430 24248
rect 22284 23724 22336 23730
rect 22284 23666 22336 23672
rect 22100 23520 22152 23526
rect 22020 23480 22100 23508
rect 22020 23322 22048 23480
rect 22100 23462 22152 23468
rect 22008 23316 22060 23322
rect 22008 23258 22060 23264
rect 22296 23118 22324 23666
rect 22100 23112 22152 23118
rect 22100 23054 22152 23060
rect 22284 23112 22336 23118
rect 22284 23054 22336 23060
rect 22112 22642 22140 23054
rect 22100 22636 22152 22642
rect 22100 22578 22152 22584
rect 22112 22166 22140 22578
rect 22100 22160 22152 22166
rect 22100 22102 22152 22108
rect 22284 22092 22336 22098
rect 22284 22034 22336 22040
rect 22192 22024 22244 22030
rect 22192 21966 22244 21972
rect 22204 21729 22232 21966
rect 22190 21720 22246 21729
rect 22190 21655 22192 21664
rect 22244 21655 22246 21664
rect 22192 21626 22244 21632
rect 22296 21350 22324 22034
rect 22284 21344 22336 21350
rect 22284 21286 22336 21292
rect 22190 21040 22246 21049
rect 22190 20975 22246 20984
rect 22100 20800 22152 20806
rect 22100 20742 22152 20748
rect 22112 20482 22140 20742
rect 22020 20454 22140 20482
rect 22020 20398 22048 20454
rect 22008 20392 22060 20398
rect 22008 20334 22060 20340
rect 21914 20088 21970 20097
rect 21914 20023 21970 20032
rect 21824 19984 21876 19990
rect 21824 19926 21876 19932
rect 21732 19780 21784 19786
rect 21732 19722 21784 19728
rect 21732 19372 21784 19378
rect 21732 19314 21784 19320
rect 21546 19000 21602 19009
rect 21744 18970 21772 19314
rect 21546 18935 21602 18944
rect 21732 18964 21784 18970
rect 21732 18906 21784 18912
rect 21640 18828 21692 18834
rect 21640 18770 21692 18776
rect 21548 18760 21600 18766
rect 21546 18728 21548 18737
rect 21600 18728 21602 18737
rect 21456 18692 21508 18698
rect 21546 18663 21602 18672
rect 21456 18634 21508 18640
rect 21560 18426 21588 18663
rect 21548 18420 21600 18426
rect 21548 18362 21600 18368
rect 21456 18080 21508 18086
rect 21272 18022 21324 18028
rect 21362 18048 21418 18057
rect 21180 17604 21232 17610
rect 21180 17546 21232 17552
rect 21192 16289 21220 17546
rect 21178 16280 21234 16289
rect 21178 16215 21234 16224
rect 21180 15428 21232 15434
rect 21180 15370 21232 15376
rect 21192 14890 21220 15370
rect 21180 14884 21232 14890
rect 21180 14826 21232 14832
rect 21192 14618 21220 14826
rect 21180 14612 21232 14618
rect 21180 14554 21232 14560
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 20996 12980 21048 12986
rect 20996 12922 21048 12928
rect 20996 12776 21048 12782
rect 20996 12718 21048 12724
rect 20812 12640 20864 12646
rect 20812 12582 20864 12588
rect 20824 12481 20852 12582
rect 20810 12472 20866 12481
rect 20810 12407 20866 12416
rect 20904 12232 20956 12238
rect 20904 12174 20956 12180
rect 20916 11694 20944 12174
rect 20904 11688 20956 11694
rect 20904 11630 20956 11636
rect 20812 11552 20864 11558
rect 20812 11494 20864 11500
rect 20720 11280 20772 11286
rect 20720 11222 20772 11228
rect 20720 11008 20772 11014
rect 20718 10976 20720 10985
rect 20772 10976 20774 10985
rect 20718 10911 20774 10920
rect 20732 10606 20760 10911
rect 20824 10674 20852 11494
rect 20916 10849 20944 11630
rect 20902 10840 20958 10849
rect 20902 10775 20958 10784
rect 20812 10668 20864 10674
rect 20812 10610 20864 10616
rect 20720 10600 20772 10606
rect 20720 10542 20772 10548
rect 20536 10260 20588 10266
rect 20536 10202 20588 10208
rect 21008 10130 21036 12718
rect 21180 12640 21232 12646
rect 21180 12582 21232 12588
rect 21192 12238 21220 12582
rect 21284 12424 21312 18022
rect 21456 18022 21508 18028
rect 21362 17983 21418 17992
rect 21468 17814 21496 18022
rect 21456 17808 21508 17814
rect 21456 17750 21508 17756
rect 21548 17740 21600 17746
rect 21548 17682 21600 17688
rect 21456 17672 21508 17678
rect 21456 17614 21508 17620
rect 21364 16992 21416 16998
rect 21364 16934 21416 16940
rect 21376 14929 21404 16934
rect 21468 16658 21496 17614
rect 21560 16658 21588 17682
rect 21456 16652 21508 16658
rect 21456 16594 21508 16600
rect 21548 16652 21600 16658
rect 21548 16594 21600 16600
rect 21652 15706 21680 18770
rect 21836 18306 21864 19926
rect 22008 19916 22060 19922
rect 22060 19876 22140 19904
rect 22008 19858 22060 19864
rect 21916 19848 21968 19854
rect 21968 19796 22048 19802
rect 21916 19790 22048 19796
rect 21928 19774 22048 19790
rect 21916 19712 21968 19718
rect 21916 19654 21968 19660
rect 21928 19242 21956 19654
rect 22020 19446 22048 19774
rect 22008 19440 22060 19446
rect 22008 19382 22060 19388
rect 22006 19272 22062 19281
rect 21916 19236 21968 19242
rect 22006 19207 22062 19216
rect 21916 19178 21968 19184
rect 21914 19000 21970 19009
rect 21914 18935 21970 18944
rect 21744 18278 21864 18306
rect 21640 15700 21692 15706
rect 21640 15642 21692 15648
rect 21548 15564 21600 15570
rect 21548 15506 21600 15512
rect 21362 14920 21418 14929
rect 21362 14855 21418 14864
rect 21364 14544 21416 14550
rect 21364 14486 21416 14492
rect 21454 14512 21510 14521
rect 21376 13938 21404 14486
rect 21560 14498 21588 15506
rect 21510 14470 21588 14498
rect 21454 14447 21510 14456
rect 21560 14278 21588 14470
rect 21640 14476 21692 14482
rect 21640 14418 21692 14424
rect 21548 14272 21600 14278
rect 21548 14214 21600 14220
rect 21364 13932 21416 13938
rect 21364 13874 21416 13880
rect 21376 13462 21404 13874
rect 21364 13456 21416 13462
rect 21364 13398 21416 13404
rect 21364 12436 21416 12442
rect 21284 12396 21364 12424
rect 21180 12232 21232 12238
rect 21086 12200 21142 12209
rect 21180 12174 21232 12180
rect 21086 12135 21142 12144
rect 21100 10742 21128 12135
rect 21192 11558 21220 12174
rect 21284 11830 21312 12396
rect 21364 12378 21416 12384
rect 21456 12164 21508 12170
rect 21456 12106 21508 12112
rect 21272 11824 21324 11830
rect 21272 11766 21324 11772
rect 21180 11552 21232 11558
rect 21180 11494 21232 11500
rect 21192 11082 21220 11494
rect 21180 11076 21232 11082
rect 21180 11018 21232 11024
rect 21178 10840 21234 10849
rect 21178 10775 21234 10784
rect 21088 10736 21140 10742
rect 21088 10678 21140 10684
rect 21192 10169 21220 10775
rect 21284 10713 21312 11766
rect 21468 11762 21496 12106
rect 21456 11756 21508 11762
rect 21456 11698 21508 11704
rect 21364 11212 21416 11218
rect 21364 11154 21416 11160
rect 21376 10810 21404 11154
rect 21364 10804 21416 10810
rect 21364 10746 21416 10752
rect 21270 10704 21326 10713
rect 21270 10639 21326 10648
rect 21560 10441 21588 14214
rect 21652 13530 21680 14418
rect 21744 13870 21772 18278
rect 21824 18148 21876 18154
rect 21824 18090 21876 18096
rect 21732 13864 21784 13870
rect 21730 13832 21732 13841
rect 21784 13832 21786 13841
rect 21730 13767 21786 13776
rect 21744 13741 21772 13767
rect 21640 13524 21692 13530
rect 21640 13466 21692 13472
rect 21652 13376 21680 13466
rect 21652 13348 21772 13376
rect 21638 13016 21694 13025
rect 21638 12951 21694 12960
rect 21652 12850 21680 12951
rect 21640 12844 21692 12850
rect 21640 12786 21692 12792
rect 21640 10668 21692 10674
rect 21640 10610 21692 10616
rect 21546 10432 21602 10441
rect 21546 10367 21602 10376
rect 21652 10266 21680 10610
rect 21456 10260 21508 10266
rect 21456 10202 21508 10208
rect 21640 10260 21692 10266
rect 21640 10202 21692 10208
rect 21178 10160 21234 10169
rect 20628 10124 20680 10130
rect 20628 10066 20680 10072
rect 20996 10124 21048 10130
rect 21178 10095 21234 10104
rect 20996 10066 21048 10072
rect 20456 9676 20576 9704
rect 19984 9444 20036 9450
rect 19984 9386 20036 9392
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19996 9178 20024 9386
rect 20350 9344 20406 9353
rect 20350 9279 20406 9288
rect 19984 9172 20036 9178
rect 19984 9114 20036 9120
rect 19524 8968 19576 8974
rect 19524 8910 19576 8916
rect 19352 8622 19472 8650
rect 19536 8634 19564 8910
rect 19614 8664 19670 8673
rect 19340 8560 19392 8566
rect 19340 8502 19392 8508
rect 19352 8378 19380 8502
rect 19260 8350 19380 8378
rect 19260 7970 19288 8350
rect 19340 8288 19392 8294
rect 19340 8230 19392 8236
rect 19168 7942 19288 7970
rect 19168 6934 19196 7942
rect 19352 7886 19380 8230
rect 19248 7880 19300 7886
rect 19248 7822 19300 7828
rect 19340 7880 19392 7886
rect 19340 7822 19392 7828
rect 19260 7478 19288 7822
rect 19352 7546 19380 7822
rect 19340 7540 19392 7546
rect 19340 7482 19392 7488
rect 19248 7472 19300 7478
rect 19248 7414 19300 7420
rect 19260 7002 19288 7414
rect 19340 7200 19392 7206
rect 19340 7142 19392 7148
rect 19248 6996 19300 7002
rect 19248 6938 19300 6944
rect 19156 6928 19208 6934
rect 19156 6870 19208 6876
rect 19352 6186 19380 7142
rect 19444 6866 19472 8622
rect 19524 8628 19576 8634
rect 19614 8599 19670 8608
rect 19524 8570 19576 8576
rect 19628 8430 19656 8599
rect 19616 8424 19668 8430
rect 19616 8366 19668 8372
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 20076 8016 20128 8022
rect 20076 7958 20128 7964
rect 20088 7546 20116 7958
rect 20076 7540 20128 7546
rect 20076 7482 20128 7488
rect 20260 7404 20312 7410
rect 20260 7346 20312 7352
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 20272 7002 20300 7346
rect 20260 6996 20312 7002
rect 20260 6938 20312 6944
rect 19432 6860 19484 6866
rect 19432 6802 19484 6808
rect 19444 6322 19472 6802
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 19432 6316 19484 6322
rect 19432 6258 19484 6264
rect 19628 6225 19656 6734
rect 19614 6216 19670 6225
rect 19340 6180 19392 6186
rect 19614 6151 19670 6160
rect 20168 6180 20220 6186
rect 19340 6122 19392 6128
rect 20168 6122 20220 6128
rect 20076 6112 20128 6118
rect 19154 6080 19210 6089
rect 20076 6054 20128 6060
rect 19154 6015 19210 6024
rect 19168 4185 19196 6015
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19246 5944 19302 5953
rect 19622 5936 19918 5956
rect 20088 5953 20116 6054
rect 20074 5944 20130 5953
rect 19246 5879 19302 5888
rect 20074 5879 20130 5888
rect 19260 5846 19288 5879
rect 19248 5840 19300 5846
rect 19248 5782 19300 5788
rect 19984 5772 20036 5778
rect 19984 5714 20036 5720
rect 19524 5704 19576 5710
rect 19524 5646 19576 5652
rect 19432 5636 19484 5642
rect 19432 5578 19484 5584
rect 19248 5568 19300 5574
rect 19248 5510 19300 5516
rect 19260 5098 19288 5510
rect 19444 5216 19472 5578
rect 19352 5188 19472 5216
rect 19248 5092 19300 5098
rect 19248 5034 19300 5040
rect 19352 5001 19380 5188
rect 19432 5092 19484 5098
rect 19432 5034 19484 5040
rect 19338 4992 19394 5001
rect 19338 4927 19394 4936
rect 19246 4856 19302 4865
rect 19444 4826 19472 5034
rect 19246 4791 19302 4800
rect 19432 4820 19484 4826
rect 19154 4176 19210 4185
rect 19154 4111 19210 4120
rect 19154 3768 19210 3777
rect 19154 3703 19210 3712
rect 19168 3602 19196 3703
rect 19156 3596 19208 3602
rect 19156 3538 19208 3544
rect 19260 3074 19288 4791
rect 19432 4762 19484 4768
rect 19444 4282 19472 4762
rect 19432 4276 19484 4282
rect 19432 4218 19484 4224
rect 19338 4040 19394 4049
rect 19338 3975 19394 3984
rect 19352 3194 19380 3975
rect 19444 3738 19472 4218
rect 19432 3732 19484 3738
rect 19432 3674 19484 3680
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19260 3046 19380 3074
rect 19062 2952 19118 2961
rect 19062 2887 19118 2896
rect 18800 2230 19012 2258
rect 18510 1864 18566 1873
rect 18510 1799 18566 1808
rect 18800 480 18828 2230
rect 19352 480 19380 3046
rect 19430 2816 19486 2825
rect 19430 2751 19486 2760
rect 19444 2582 19472 2751
rect 19432 2576 19484 2582
rect 19432 2518 19484 2524
rect 19536 2281 19564 5646
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19996 4486 20024 5714
rect 20180 5574 20208 6122
rect 20168 5568 20220 5574
rect 20168 5510 20220 5516
rect 20180 5030 20208 5510
rect 20168 5024 20220 5030
rect 20168 4966 20220 4972
rect 19984 4480 20036 4486
rect 19982 4448 19984 4457
rect 20036 4448 20038 4457
rect 19982 4383 20038 4392
rect 20180 4214 20208 4966
rect 20272 4826 20300 6938
rect 20364 5545 20392 9279
rect 20444 8628 20496 8634
rect 20548 8616 20576 9676
rect 20640 9654 20668 10066
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20628 9648 20680 9654
rect 20628 9590 20680 9596
rect 20732 9518 20760 9998
rect 20720 9512 20772 9518
rect 20772 9472 20852 9500
rect 20720 9454 20772 9460
rect 20824 9382 20852 9472
rect 21362 9480 21418 9489
rect 21362 9415 21418 9424
rect 20812 9376 20864 9382
rect 20812 9318 20864 9324
rect 20994 9344 21050 9353
rect 20824 8906 20852 9318
rect 20994 9279 21050 9288
rect 20812 8900 20864 8906
rect 20812 8842 20864 8848
rect 20496 8588 20576 8616
rect 20444 8570 20496 8576
rect 20456 8362 20484 8570
rect 20548 8378 20576 8588
rect 20720 8424 20772 8430
rect 20718 8392 20720 8401
rect 20772 8392 20774 8401
rect 20444 8356 20496 8362
rect 20548 8350 20668 8378
rect 20444 8298 20496 8304
rect 20536 8288 20588 8294
rect 20640 8276 20668 8350
rect 20718 8327 20774 8336
rect 20720 8288 20772 8294
rect 20640 8248 20720 8276
rect 20536 8230 20588 8236
rect 20720 8230 20772 8236
rect 20548 7750 20576 8230
rect 20824 7886 20852 8842
rect 20904 8832 20956 8838
rect 20904 8774 20956 8780
rect 20916 7993 20944 8774
rect 20902 7984 20958 7993
rect 20902 7919 20958 7928
rect 20812 7880 20864 7886
rect 20812 7822 20864 7828
rect 20536 7744 20588 7750
rect 20536 7686 20588 7692
rect 20444 7200 20496 7206
rect 20444 7142 20496 7148
rect 20456 6730 20484 7142
rect 20444 6724 20496 6730
rect 20444 6666 20496 6672
rect 20350 5536 20406 5545
rect 20350 5471 20406 5480
rect 20260 4820 20312 4826
rect 20260 4762 20312 4768
rect 20168 4208 20220 4214
rect 20168 4150 20220 4156
rect 20456 4146 20484 6666
rect 20548 6633 20576 7686
rect 20628 7200 20680 7206
rect 20628 7142 20680 7148
rect 20640 6662 20668 7142
rect 20720 6792 20772 6798
rect 20720 6734 20772 6740
rect 20628 6656 20680 6662
rect 20534 6624 20590 6633
rect 20628 6598 20680 6604
rect 20534 6559 20590 6568
rect 20536 6248 20588 6254
rect 20536 6190 20588 6196
rect 20548 5778 20576 6190
rect 20536 5772 20588 5778
rect 20536 5714 20588 5720
rect 20640 5545 20668 6598
rect 20626 5536 20682 5545
rect 20626 5471 20682 5480
rect 20732 5386 20760 6734
rect 20824 5778 20852 7822
rect 21008 6730 21036 9279
rect 21376 9178 21404 9415
rect 21364 9172 21416 9178
rect 21364 9114 21416 9120
rect 21376 8634 21404 9114
rect 21468 8974 21496 10202
rect 21546 9480 21602 9489
rect 21546 9415 21602 9424
rect 21560 9081 21588 9415
rect 21744 9081 21772 13348
rect 21836 13326 21864 18090
rect 21928 17513 21956 18935
rect 22020 18601 22048 19207
rect 22006 18592 22062 18601
rect 22006 18527 22062 18536
rect 22112 18426 22140 19876
rect 22204 18834 22232 20975
rect 22296 19922 22324 21286
rect 22388 19990 22416 24239
rect 22468 23044 22520 23050
rect 22468 22986 22520 22992
rect 22480 20058 22508 22986
rect 22468 20052 22520 20058
rect 22468 19994 22520 20000
rect 22376 19984 22428 19990
rect 22376 19926 22428 19932
rect 22284 19916 22336 19922
rect 22284 19858 22336 19864
rect 22572 19802 22600 24550
rect 22664 24138 22692 24754
rect 22756 24274 22784 25298
rect 22940 24954 22968 25298
rect 23020 25288 23072 25294
rect 23020 25230 23072 25236
rect 23572 25288 23624 25294
rect 23572 25230 23624 25236
rect 22928 24948 22980 24954
rect 22928 24890 22980 24896
rect 23032 24818 23060 25230
rect 23480 25152 23532 25158
rect 23480 25094 23532 25100
rect 23020 24812 23072 24818
rect 23020 24754 23072 24760
rect 22928 24744 22980 24750
rect 22928 24686 22980 24692
rect 22744 24268 22796 24274
rect 22744 24210 22796 24216
rect 22652 24132 22704 24138
rect 22652 24074 22704 24080
rect 22664 23508 22692 24074
rect 22756 24041 22784 24210
rect 22836 24132 22888 24138
rect 22836 24074 22888 24080
rect 22742 24032 22798 24041
rect 22742 23967 22798 23976
rect 22744 23520 22796 23526
rect 22664 23480 22744 23508
rect 22744 23462 22796 23468
rect 22756 22817 22784 23462
rect 22742 22808 22798 22817
rect 22742 22743 22798 22752
rect 22848 20806 22876 24074
rect 22836 20800 22888 20806
rect 22836 20742 22888 20748
rect 22742 20632 22798 20641
rect 22742 20567 22744 20576
rect 22796 20567 22798 20576
rect 22744 20538 22796 20544
rect 22836 19916 22888 19922
rect 22836 19858 22888 19864
rect 22296 19774 22600 19802
rect 22744 19848 22796 19854
rect 22744 19790 22796 19796
rect 22192 18828 22244 18834
rect 22192 18770 22244 18776
rect 22100 18420 22152 18426
rect 22100 18362 22152 18368
rect 22006 17912 22062 17921
rect 22204 17882 22232 18770
rect 22006 17847 22062 17856
rect 22192 17876 22244 17882
rect 22020 17814 22048 17847
rect 22192 17818 22244 17824
rect 22008 17808 22060 17814
rect 22008 17750 22060 17756
rect 22008 17672 22060 17678
rect 22008 17614 22060 17620
rect 21914 17504 21970 17513
rect 21914 17439 21970 17448
rect 21928 17270 21956 17439
rect 21916 17264 21968 17270
rect 21916 17206 21968 17212
rect 22020 16998 22048 17614
rect 22008 16992 22060 16998
rect 22008 16934 22060 16940
rect 21916 16788 21968 16794
rect 21916 16730 21968 16736
rect 21928 16114 21956 16730
rect 22020 16726 22048 16934
rect 22008 16720 22060 16726
rect 22008 16662 22060 16668
rect 21916 16108 21968 16114
rect 21916 16050 21968 16056
rect 22020 16046 22048 16662
rect 22190 16552 22246 16561
rect 22190 16487 22246 16496
rect 22204 16114 22232 16487
rect 22192 16108 22244 16114
rect 22192 16050 22244 16056
rect 22008 16040 22060 16046
rect 22008 15982 22060 15988
rect 22020 15502 22048 15982
rect 22192 15972 22244 15978
rect 22192 15914 22244 15920
rect 22204 15706 22232 15914
rect 22192 15700 22244 15706
rect 22192 15642 22244 15648
rect 22296 15586 22324 19774
rect 22376 19712 22428 19718
rect 22376 19654 22428 19660
rect 22468 19712 22520 19718
rect 22468 19654 22520 19660
rect 22388 18970 22416 19654
rect 22376 18964 22428 18970
rect 22376 18906 22428 18912
rect 22388 18222 22416 18906
rect 22376 18216 22428 18222
rect 22376 18158 22428 18164
rect 22480 17921 22508 19654
rect 22560 19372 22612 19378
rect 22612 19332 22692 19360
rect 22560 19314 22612 19320
rect 22560 18896 22612 18902
rect 22560 18838 22612 18844
rect 22466 17912 22522 17921
rect 22572 17882 22600 18838
rect 22466 17847 22522 17856
rect 22560 17876 22612 17882
rect 22560 17818 22612 17824
rect 22468 17740 22520 17746
rect 22468 17682 22520 17688
rect 22376 17060 22428 17066
rect 22376 17002 22428 17008
rect 22204 15558 22324 15586
rect 22008 15496 22060 15502
rect 22008 15438 22060 15444
rect 22008 14952 22060 14958
rect 22008 14894 22060 14900
rect 21916 14612 21968 14618
rect 21916 14554 21968 14560
rect 21928 13870 21956 14554
rect 21916 13864 21968 13870
rect 21916 13806 21968 13812
rect 21824 13320 21876 13326
rect 21824 13262 21876 13268
rect 21822 13152 21878 13161
rect 21822 13087 21878 13096
rect 21546 9072 21602 9081
rect 21546 9007 21602 9016
rect 21730 9072 21786 9081
rect 21730 9007 21786 9016
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 21364 8628 21416 8634
rect 21364 8570 21416 8576
rect 21468 8498 21496 8910
rect 21456 8492 21508 8498
rect 21456 8434 21508 8440
rect 21468 8090 21496 8434
rect 21456 8084 21508 8090
rect 21456 8026 21508 8032
rect 21468 7410 21496 8026
rect 21456 7404 21508 7410
rect 21456 7346 21508 7352
rect 21836 6882 21864 13087
rect 21928 12481 21956 13806
rect 22020 13394 22048 14894
rect 22098 14104 22154 14113
rect 22098 14039 22154 14048
rect 22112 13870 22140 14039
rect 22100 13864 22152 13870
rect 22100 13806 22152 13812
rect 22008 13388 22060 13394
rect 22008 13330 22060 13336
rect 21914 12472 21970 12481
rect 21914 12407 21970 12416
rect 22008 12096 22060 12102
rect 22008 12038 22060 12044
rect 21916 11824 21968 11830
rect 21916 11766 21968 11772
rect 21928 11354 21956 11766
rect 22020 11762 22048 12038
rect 22008 11756 22060 11762
rect 22008 11698 22060 11704
rect 22020 11354 22048 11698
rect 21916 11348 21968 11354
rect 21916 11290 21968 11296
rect 22008 11348 22060 11354
rect 22008 11290 22060 11296
rect 21928 11150 21956 11290
rect 21916 11144 21968 11150
rect 21916 11086 21968 11092
rect 21928 10198 21956 11086
rect 22100 10668 22152 10674
rect 22100 10610 22152 10616
rect 21916 10192 21968 10198
rect 21916 10134 21968 10140
rect 22008 9920 22060 9926
rect 22008 9862 22060 9868
rect 22020 9450 22048 9862
rect 22112 9722 22140 10610
rect 22100 9716 22152 9722
rect 22100 9658 22152 9664
rect 22008 9444 22060 9450
rect 22008 9386 22060 9392
rect 22112 9160 22140 9658
rect 22020 9132 22140 9160
rect 22020 8022 22048 9132
rect 22008 8016 22060 8022
rect 22008 7958 22060 7964
rect 22006 7848 22062 7857
rect 22062 7806 22140 7834
rect 22006 7783 22062 7792
rect 21916 7404 21968 7410
rect 21916 7346 21968 7352
rect 21928 7002 21956 7346
rect 22008 7336 22060 7342
rect 22008 7278 22060 7284
rect 22020 7206 22048 7278
rect 22008 7200 22060 7206
rect 22008 7142 22060 7148
rect 21916 6996 21968 7002
rect 21916 6938 21968 6944
rect 21272 6860 21324 6866
rect 21272 6802 21324 6808
rect 21652 6854 21864 6882
rect 20996 6724 21048 6730
rect 20996 6666 21048 6672
rect 21284 5914 21312 6802
rect 21364 6656 21416 6662
rect 21364 6598 21416 6604
rect 21272 5908 21324 5914
rect 21272 5850 21324 5856
rect 20904 5840 20956 5846
rect 20904 5782 20956 5788
rect 20812 5772 20864 5778
rect 20812 5714 20864 5720
rect 20640 5358 20760 5386
rect 20444 4140 20496 4146
rect 20444 4082 20496 4088
rect 20442 4040 20498 4049
rect 20640 4010 20668 5358
rect 20720 5024 20772 5030
rect 20720 4966 20772 4972
rect 20442 3975 20498 3984
rect 20628 4004 20680 4010
rect 20352 3936 20404 3942
rect 20352 3878 20404 3884
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 20364 3466 20392 3878
rect 20076 3460 20128 3466
rect 20076 3402 20128 3408
rect 20352 3460 20404 3466
rect 20352 3402 20404 3408
rect 20088 3097 20116 3402
rect 20260 3392 20312 3398
rect 20260 3334 20312 3340
rect 20272 3126 20300 3334
rect 20260 3120 20312 3126
rect 19890 3088 19946 3097
rect 20074 3088 20130 3097
rect 19946 3046 20024 3074
rect 19890 3023 19946 3032
rect 19996 2938 20024 3046
rect 20260 3062 20312 3068
rect 20074 3023 20076 3032
rect 20128 3023 20130 3032
rect 20076 2994 20128 3000
rect 19996 2910 20116 2938
rect 20088 2825 20116 2910
rect 20074 2816 20130 2825
rect 19622 2748 19918 2768
rect 20074 2751 20130 2760
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19892 2576 19944 2582
rect 19892 2518 19944 2524
rect 19800 2508 19852 2514
rect 19800 2450 19852 2456
rect 19812 2310 19840 2450
rect 19800 2304 19852 2310
rect 19522 2272 19578 2281
rect 19800 2246 19852 2252
rect 19522 2207 19578 2216
rect 19812 1465 19840 2246
rect 19798 1456 19854 1465
rect 19798 1391 19854 1400
rect 19904 480 19932 2518
rect 20168 2304 20220 2310
rect 20168 2246 20220 2252
rect 20180 1465 20208 2246
rect 20272 1601 20300 3062
rect 20258 1592 20314 1601
rect 20258 1527 20314 1536
rect 20166 1456 20222 1465
rect 20166 1391 20222 1400
rect 20456 480 20484 3975
rect 20628 3946 20680 3952
rect 20732 3913 20760 4966
rect 20812 4276 20864 4282
rect 20812 4218 20864 4224
rect 20718 3904 20774 3913
rect 20718 3839 20774 3848
rect 20732 2922 20760 3839
rect 20720 2916 20772 2922
rect 20720 2858 20772 2864
rect 20824 2650 20852 4218
rect 20916 3194 20944 5782
rect 21284 5370 21312 5850
rect 21376 5658 21404 6598
rect 21376 5630 21496 5658
rect 21272 5364 21324 5370
rect 21272 5306 21324 5312
rect 21468 5030 21496 5630
rect 21456 5024 21508 5030
rect 21456 4966 21508 4972
rect 21468 4729 21496 4966
rect 21454 4720 21510 4729
rect 21272 4684 21324 4690
rect 21454 4655 21510 4664
rect 21272 4626 21324 4632
rect 20996 4548 21048 4554
rect 20996 4490 21048 4496
rect 21008 4049 21036 4490
rect 20994 4040 21050 4049
rect 20994 3975 21050 3984
rect 21284 3398 21312 4626
rect 21456 4616 21508 4622
rect 21456 4558 21508 4564
rect 21364 3936 21416 3942
rect 21364 3878 21416 3884
rect 21376 3641 21404 3878
rect 21362 3632 21418 3641
rect 21362 3567 21418 3576
rect 21468 3534 21496 4558
rect 21652 4554 21680 6854
rect 21824 6792 21876 6798
rect 21824 6734 21876 6740
rect 21732 6724 21784 6730
rect 21732 6666 21784 6672
rect 21744 5166 21772 6666
rect 21836 6458 21864 6734
rect 21824 6452 21876 6458
rect 21824 6394 21876 6400
rect 21836 5846 21864 6394
rect 22020 5914 22048 7142
rect 22112 6202 22140 7806
rect 22204 7206 22232 15558
rect 22282 15192 22338 15201
rect 22388 15162 22416 17002
rect 22282 15127 22338 15136
rect 22376 15156 22428 15162
rect 22296 14498 22324 15127
rect 22376 15098 22428 15104
rect 22296 14470 22416 14498
rect 22284 14408 22336 14414
rect 22284 14350 22336 14356
rect 22296 14006 22324 14350
rect 22284 14000 22336 14006
rect 22282 13968 22284 13977
rect 22336 13968 22338 13977
rect 22282 13903 22338 13912
rect 22284 13456 22336 13462
rect 22284 13398 22336 13404
rect 22296 12782 22324 13398
rect 22284 12776 22336 12782
rect 22284 12718 22336 12724
rect 22296 12442 22324 12718
rect 22284 12436 22336 12442
rect 22284 12378 22336 12384
rect 22282 12336 22338 12345
rect 22282 12271 22338 12280
rect 22296 9217 22324 12271
rect 22388 12238 22416 14470
rect 22376 12232 22428 12238
rect 22376 12174 22428 12180
rect 22480 11694 22508 17682
rect 22560 17128 22612 17134
rect 22558 17096 22560 17105
rect 22612 17096 22614 17105
rect 22558 17031 22614 17040
rect 22560 16992 22612 16998
rect 22560 16934 22612 16940
rect 22572 15910 22600 16934
rect 22560 15904 22612 15910
rect 22560 15846 22612 15852
rect 22558 15736 22614 15745
rect 22558 15671 22614 15680
rect 22572 13462 22600 15671
rect 22560 13456 22612 13462
rect 22560 13398 22612 13404
rect 22664 12084 22692 19332
rect 22756 19310 22784 19790
rect 22848 19514 22876 19858
rect 22940 19854 22968 24686
rect 23296 24200 23348 24206
rect 23296 24142 23348 24148
rect 23308 23322 23336 24142
rect 23492 23746 23520 25094
rect 23584 24614 23612 25230
rect 23572 24608 23624 24614
rect 23572 24550 23624 24556
rect 23400 23718 23520 23746
rect 23296 23316 23348 23322
rect 23296 23258 23348 23264
rect 23294 23216 23350 23225
rect 23294 23151 23350 23160
rect 23204 23044 23256 23050
rect 23204 22986 23256 22992
rect 23020 22976 23072 22982
rect 23018 22944 23020 22953
rect 23072 22944 23074 22953
rect 23018 22879 23074 22888
rect 23216 22438 23244 22986
rect 23204 22432 23256 22438
rect 23204 22374 23256 22380
rect 23308 22030 23336 23151
rect 23400 22574 23428 23718
rect 23480 23588 23532 23594
rect 23480 23530 23532 23536
rect 23492 23322 23520 23530
rect 23480 23316 23532 23322
rect 23480 23258 23532 23264
rect 23584 22710 23612 24550
rect 23676 23905 23704 25350
rect 23938 25327 23994 25336
rect 24032 25356 24084 25362
rect 23952 24342 23980 25327
rect 24032 25298 24084 25304
rect 24044 24682 24072 25298
rect 24136 25242 24164 27520
rect 24582 27160 24638 27169
rect 24582 27095 24638 27104
rect 24596 25430 24624 27095
rect 24688 26858 24716 27639
rect 24766 27520 24822 28000
rect 25318 27520 25374 28000
rect 25870 27520 25926 28000
rect 26514 27520 26570 28000
rect 27066 27520 27122 28000
rect 27618 27520 27674 28000
rect 24676 26852 24728 26858
rect 24676 26794 24728 26800
rect 24780 26738 24808 27520
rect 24688 26710 24808 26738
rect 24688 26042 24716 26710
rect 24766 26616 24822 26625
rect 24766 26551 24822 26560
rect 24780 26450 24808 26551
rect 24768 26444 24820 26450
rect 24768 26386 24820 26392
rect 24676 26036 24728 26042
rect 24676 25978 24728 25984
rect 25332 25945 25360 27520
rect 25318 25936 25374 25945
rect 25318 25871 25374 25880
rect 24766 25800 24822 25809
rect 25884 25770 25912 27520
rect 26528 25838 26556 27520
rect 26516 25832 26568 25838
rect 26516 25774 26568 25780
rect 24766 25735 24822 25744
rect 25872 25764 25924 25770
rect 24780 25702 24808 25735
rect 25872 25706 25924 25712
rect 24768 25696 24820 25702
rect 24768 25638 24820 25644
rect 24768 25492 24820 25498
rect 24768 25434 24820 25440
rect 24584 25424 24636 25430
rect 24780 25401 24808 25434
rect 24584 25366 24636 25372
rect 24766 25392 24822 25401
rect 24766 25327 24822 25336
rect 24136 25214 24256 25242
rect 24124 25152 24176 25158
rect 24124 25094 24176 25100
rect 24032 24676 24084 24682
rect 24032 24618 24084 24624
rect 23940 24336 23992 24342
rect 23940 24278 23992 24284
rect 23756 24268 23808 24274
rect 23756 24210 23808 24216
rect 23848 24268 23900 24274
rect 23848 24210 23900 24216
rect 23662 23896 23718 23905
rect 23662 23831 23718 23840
rect 23664 23520 23716 23526
rect 23664 23462 23716 23468
rect 23572 22704 23624 22710
rect 23572 22646 23624 22652
rect 23388 22568 23440 22574
rect 23388 22510 23440 22516
rect 23572 22568 23624 22574
rect 23572 22510 23624 22516
rect 23388 22432 23440 22438
rect 23388 22374 23440 22380
rect 23296 22024 23348 22030
rect 23296 21966 23348 21972
rect 23202 21856 23258 21865
rect 23202 21791 23258 21800
rect 23018 21448 23074 21457
rect 23018 21383 23074 21392
rect 22928 19848 22980 19854
rect 22928 19790 22980 19796
rect 22836 19508 22888 19514
rect 22836 19450 22888 19456
rect 22744 19304 22796 19310
rect 22848 19281 22876 19450
rect 22744 19246 22796 19252
rect 22834 19272 22890 19281
rect 22756 12170 22784 19246
rect 22834 19207 22890 19216
rect 23032 18850 23060 21383
rect 23112 21004 23164 21010
rect 23112 20946 23164 20952
rect 23124 19854 23152 20946
rect 23112 19848 23164 19854
rect 23112 19790 23164 19796
rect 22848 18822 23060 18850
rect 22848 16998 22876 18822
rect 23020 18760 23072 18766
rect 23020 18702 23072 18708
rect 23032 18442 23060 18702
rect 23124 18630 23152 19790
rect 23112 18624 23164 18630
rect 23112 18566 23164 18572
rect 22940 18414 23060 18442
rect 22940 18358 22968 18414
rect 22928 18352 22980 18358
rect 22926 18320 22928 18329
rect 22980 18320 22982 18329
rect 22926 18255 22982 18264
rect 23124 17814 23152 18566
rect 23112 17808 23164 17814
rect 23112 17750 23164 17756
rect 22928 17740 22980 17746
rect 22928 17682 22980 17688
rect 22940 16998 22968 17682
rect 23020 17672 23072 17678
rect 23020 17614 23072 17620
rect 23112 17672 23164 17678
rect 23112 17614 23164 17620
rect 23032 17377 23060 17614
rect 23018 17368 23074 17377
rect 23018 17303 23074 17312
rect 22836 16992 22888 16998
rect 22836 16934 22888 16940
rect 22928 16992 22980 16998
rect 22928 16934 22980 16940
rect 22834 16824 22890 16833
rect 22834 16759 22890 16768
rect 22848 12442 22876 16759
rect 22940 16046 22968 16934
rect 23032 16794 23060 17303
rect 23124 17066 23152 17614
rect 23112 17060 23164 17066
rect 23112 17002 23164 17008
rect 23124 16794 23152 17002
rect 23020 16788 23072 16794
rect 23020 16730 23072 16736
rect 23112 16788 23164 16794
rect 23112 16730 23164 16736
rect 23124 16674 23152 16730
rect 23032 16646 23152 16674
rect 23032 16561 23060 16646
rect 23018 16552 23074 16561
rect 23018 16487 23074 16496
rect 23112 16516 23164 16522
rect 23112 16458 23164 16464
rect 23124 16250 23152 16458
rect 23112 16244 23164 16250
rect 23112 16186 23164 16192
rect 22928 16040 22980 16046
rect 22928 15982 22980 15988
rect 22928 15564 22980 15570
rect 22928 15506 22980 15512
rect 22940 14822 22968 15506
rect 23020 15496 23072 15502
rect 23020 15438 23072 15444
rect 23032 15162 23060 15438
rect 23112 15360 23164 15366
rect 23112 15302 23164 15308
rect 23020 15156 23072 15162
rect 23020 15098 23072 15104
rect 23018 14920 23074 14929
rect 23018 14855 23020 14864
rect 23072 14855 23074 14864
rect 23020 14826 23072 14832
rect 22928 14816 22980 14822
rect 22928 14758 22980 14764
rect 22940 14618 22968 14758
rect 22928 14612 22980 14618
rect 22928 14554 22980 14560
rect 23124 14074 23152 15302
rect 23112 14068 23164 14074
rect 23112 14010 23164 14016
rect 22926 13832 22982 13841
rect 22926 13767 22982 13776
rect 22836 12436 22888 12442
rect 22836 12378 22888 12384
rect 22744 12164 22796 12170
rect 22744 12106 22796 12112
rect 22572 12056 22692 12084
rect 22468 11688 22520 11694
rect 22374 11656 22430 11665
rect 22468 11630 22520 11636
rect 22374 11591 22430 11600
rect 22388 11218 22416 11591
rect 22376 11212 22428 11218
rect 22376 11154 22428 11160
rect 22388 10810 22416 11154
rect 22468 11076 22520 11082
rect 22468 11018 22520 11024
rect 22376 10804 22428 10810
rect 22376 10746 22428 10752
rect 22480 10062 22508 11018
rect 22572 10538 22600 12056
rect 22650 11384 22706 11393
rect 22650 11319 22652 11328
rect 22704 11319 22706 11328
rect 22652 11290 22704 11296
rect 22560 10532 22612 10538
rect 22560 10474 22612 10480
rect 22468 10056 22520 10062
rect 22468 9998 22520 10004
rect 22572 9738 22600 10474
rect 22388 9710 22600 9738
rect 22282 9208 22338 9217
rect 22282 9143 22338 9152
rect 22388 9058 22416 9710
rect 22652 9512 22704 9518
rect 22652 9454 22704 9460
rect 22560 9444 22612 9450
rect 22560 9386 22612 9392
rect 22296 9030 22416 9058
rect 22296 7206 22324 9030
rect 22468 8832 22520 8838
rect 22468 8774 22520 8780
rect 22376 8492 22428 8498
rect 22376 8434 22428 8440
rect 22192 7200 22244 7206
rect 22192 7142 22244 7148
rect 22284 7200 22336 7206
rect 22284 7142 22336 7148
rect 22388 6225 22416 8434
rect 22480 7449 22508 8774
rect 22466 7440 22522 7449
rect 22466 7375 22522 7384
rect 22374 6216 22430 6225
rect 22112 6174 22324 6202
rect 22192 6112 22244 6118
rect 22192 6054 22244 6060
rect 22008 5908 22060 5914
rect 22008 5850 22060 5856
rect 21824 5840 21876 5846
rect 21876 5800 21956 5828
rect 21824 5782 21876 5788
rect 21928 5794 21956 5800
rect 21928 5766 22140 5794
rect 22112 5370 22140 5766
rect 22100 5364 22152 5370
rect 22100 5306 22152 5312
rect 21732 5160 21784 5166
rect 21732 5102 21784 5108
rect 21744 4826 21772 5102
rect 21824 5092 21876 5098
rect 21824 5034 21876 5040
rect 21732 4820 21784 4826
rect 21732 4762 21784 4768
rect 21730 4584 21786 4593
rect 21640 4548 21692 4554
rect 21730 4519 21732 4528
rect 21640 4490 21692 4496
rect 21784 4519 21786 4528
rect 21732 4490 21784 4496
rect 21652 4282 21680 4490
rect 21640 4276 21692 4282
rect 21640 4218 21692 4224
rect 21744 4214 21772 4490
rect 21732 4208 21784 4214
rect 21732 4150 21784 4156
rect 21836 3942 21864 5034
rect 22100 4480 22152 4486
rect 22020 4428 22100 4434
rect 22020 4422 22152 4428
rect 22020 4406 22140 4422
rect 21824 3936 21876 3942
rect 21824 3878 21876 3884
rect 21836 3670 21864 3878
rect 22020 3738 22048 4406
rect 22008 3732 22060 3738
rect 22008 3674 22060 3680
rect 21824 3664 21876 3670
rect 21824 3606 21876 3612
rect 21456 3528 21508 3534
rect 21456 3470 21508 3476
rect 21732 3528 21784 3534
rect 22204 3482 22232 6054
rect 22296 4826 22324 6174
rect 22374 6151 22430 6160
rect 22376 5908 22428 5914
rect 22376 5850 22428 5856
rect 22284 4820 22336 4826
rect 22284 4762 22336 4768
rect 22282 4448 22338 4457
rect 22388 4434 22416 5850
rect 22572 4758 22600 9386
rect 22664 8498 22692 9454
rect 22652 8492 22704 8498
rect 22652 8434 22704 8440
rect 22652 8288 22704 8294
rect 22652 8230 22704 8236
rect 22560 4752 22612 4758
rect 22560 4694 22612 4700
rect 22338 4406 22416 4434
rect 22282 4383 22338 4392
rect 22296 4010 22324 4383
rect 22376 4208 22428 4214
rect 22376 4150 22428 4156
rect 22284 4004 22336 4010
rect 22284 3946 22336 3952
rect 22296 3670 22324 3946
rect 22388 3738 22416 4150
rect 22572 4146 22600 4694
rect 22560 4140 22612 4146
rect 22560 4082 22612 4088
rect 22376 3732 22428 3738
rect 22376 3674 22428 3680
rect 22284 3664 22336 3670
rect 22284 3606 22336 3612
rect 22572 3505 22600 4082
rect 22664 3777 22692 8230
rect 22756 5001 22784 12106
rect 22834 10976 22890 10985
rect 22834 10911 22890 10920
rect 22848 10810 22876 10911
rect 22836 10804 22888 10810
rect 22836 10746 22888 10752
rect 22940 9450 22968 13767
rect 23018 13696 23074 13705
rect 23018 13631 23074 13640
rect 22928 9444 22980 9450
rect 22928 9386 22980 9392
rect 23032 9178 23060 13631
rect 23216 12850 23244 21791
rect 23308 21690 23336 21966
rect 23296 21684 23348 21690
rect 23296 21626 23348 21632
rect 23400 21570 23428 22374
rect 23584 21962 23612 22510
rect 23572 21956 23624 21962
rect 23572 21898 23624 21904
rect 23676 21729 23704 23462
rect 23768 22953 23796 24210
rect 23860 24177 23888 24210
rect 23846 24168 23902 24177
rect 23846 24103 23902 24112
rect 23846 23488 23902 23497
rect 23846 23423 23902 23432
rect 23754 22944 23810 22953
rect 23754 22879 23810 22888
rect 23860 22778 23888 23423
rect 24032 23248 24084 23254
rect 24032 23190 24084 23196
rect 23940 23112 23992 23118
rect 23940 23054 23992 23060
rect 23848 22772 23900 22778
rect 23848 22714 23900 22720
rect 23756 22704 23808 22710
rect 23756 22646 23808 22652
rect 23662 21720 23718 21729
rect 23768 21690 23796 22646
rect 23848 22568 23900 22574
rect 23848 22510 23900 22516
rect 23860 21865 23888 22510
rect 23952 22234 23980 23054
rect 24044 22438 24072 23190
rect 24032 22432 24084 22438
rect 24032 22374 24084 22380
rect 23940 22228 23992 22234
rect 23940 22170 23992 22176
rect 24044 22166 24072 22374
rect 24032 22160 24084 22166
rect 24032 22102 24084 22108
rect 24032 21956 24084 21962
rect 24032 21898 24084 21904
rect 23940 21888 23992 21894
rect 23846 21856 23902 21865
rect 23940 21830 23992 21836
rect 23846 21791 23902 21800
rect 23662 21655 23718 21664
rect 23756 21684 23808 21690
rect 23756 21626 23808 21632
rect 23400 21542 23888 21570
rect 23952 21554 23980 21830
rect 23572 21480 23624 21486
rect 23572 21422 23624 21428
rect 23296 21412 23348 21418
rect 23296 21354 23348 21360
rect 23308 21146 23336 21354
rect 23296 21140 23348 21146
rect 23296 21082 23348 21088
rect 23388 21140 23440 21146
rect 23388 21082 23440 21088
rect 23296 20800 23348 20806
rect 23296 20742 23348 20748
rect 23308 20466 23336 20742
rect 23296 20460 23348 20466
rect 23296 20402 23348 20408
rect 23400 20346 23428 21082
rect 23480 20936 23532 20942
rect 23480 20878 23532 20884
rect 23492 20641 23520 20878
rect 23478 20632 23534 20641
rect 23584 20602 23612 21422
rect 23664 21344 23716 21350
rect 23664 21286 23716 21292
rect 23676 21185 23704 21286
rect 23662 21176 23718 21185
rect 23662 21111 23718 21120
rect 23664 21004 23716 21010
rect 23664 20946 23716 20952
rect 23478 20567 23534 20576
rect 23572 20596 23624 20602
rect 23308 20318 23428 20346
rect 23308 17377 23336 20318
rect 23388 20256 23440 20262
rect 23388 20198 23440 20204
rect 23400 19718 23428 20198
rect 23388 19712 23440 19718
rect 23388 19654 23440 19660
rect 23492 19174 23520 20567
rect 23572 20538 23624 20544
rect 23676 20058 23704 20946
rect 23756 20800 23808 20806
rect 23756 20742 23808 20748
rect 23664 20052 23716 20058
rect 23664 19994 23716 20000
rect 23572 19848 23624 19854
rect 23572 19790 23624 19796
rect 23584 19514 23612 19790
rect 23572 19508 23624 19514
rect 23572 19450 23624 19456
rect 23664 19508 23716 19514
rect 23664 19450 23716 19456
rect 23570 19408 23626 19417
rect 23570 19343 23626 19352
rect 23480 19168 23532 19174
rect 23480 19110 23532 19116
rect 23480 18760 23532 18766
rect 23480 18702 23532 18708
rect 23388 18624 23440 18630
rect 23388 18566 23440 18572
rect 23294 17368 23350 17377
rect 23294 17303 23350 17312
rect 23296 16448 23348 16454
rect 23296 16390 23348 16396
rect 23308 14550 23336 16390
rect 23400 15366 23428 18566
rect 23492 18222 23520 18702
rect 23480 18216 23532 18222
rect 23480 18158 23532 18164
rect 23492 18086 23520 18158
rect 23480 18080 23532 18086
rect 23480 18022 23532 18028
rect 23584 17338 23612 19343
rect 23676 18630 23704 19450
rect 23664 18624 23716 18630
rect 23664 18566 23716 18572
rect 23664 18284 23716 18290
rect 23664 18226 23716 18232
rect 23676 17814 23704 18226
rect 23768 18086 23796 20742
rect 23756 18080 23808 18086
rect 23756 18022 23808 18028
rect 23664 17808 23716 17814
rect 23664 17750 23716 17756
rect 23572 17332 23624 17338
rect 23572 17274 23624 17280
rect 23570 17232 23626 17241
rect 23570 17167 23626 17176
rect 23584 16538 23612 17167
rect 23492 16510 23612 16538
rect 23388 15360 23440 15366
rect 23388 15302 23440 15308
rect 23386 15192 23442 15201
rect 23386 15127 23442 15136
rect 23296 14544 23348 14550
rect 23400 14521 23428 15127
rect 23296 14486 23348 14492
rect 23386 14512 23442 14521
rect 23386 14447 23442 14456
rect 23204 12844 23256 12850
rect 23204 12786 23256 12792
rect 23112 12776 23164 12782
rect 23112 12718 23164 12724
rect 23124 12345 23152 12718
rect 23388 12640 23440 12646
rect 23388 12582 23440 12588
rect 23400 12481 23428 12582
rect 23386 12472 23442 12481
rect 23296 12436 23348 12442
rect 23386 12407 23442 12416
rect 23296 12378 23348 12384
rect 23204 12368 23256 12374
rect 23110 12336 23166 12345
rect 23204 12310 23256 12316
rect 23110 12271 23166 12280
rect 23216 11354 23244 12310
rect 23308 12073 23336 12378
rect 23294 12064 23350 12073
rect 23294 11999 23350 12008
rect 23204 11348 23256 11354
rect 23204 11290 23256 11296
rect 23112 11008 23164 11014
rect 23308 10962 23336 11999
rect 23386 11112 23442 11121
rect 23386 11047 23442 11056
rect 23400 11014 23428 11047
rect 23112 10950 23164 10956
rect 23124 10266 23152 10950
rect 23216 10934 23336 10962
rect 23388 11008 23440 11014
rect 23388 10950 23440 10956
rect 23112 10260 23164 10266
rect 23112 10202 23164 10208
rect 23124 9518 23152 10202
rect 23112 9512 23164 9518
rect 23112 9454 23164 9460
rect 23110 9208 23166 9217
rect 23020 9172 23072 9178
rect 23110 9143 23166 9152
rect 23020 9114 23072 9120
rect 22836 9036 22888 9042
rect 22836 8978 22888 8984
rect 22848 8362 22876 8978
rect 22928 8968 22980 8974
rect 22926 8936 22928 8945
rect 22980 8936 22982 8945
rect 22926 8871 22982 8880
rect 22836 8356 22888 8362
rect 22836 8298 22888 8304
rect 22742 4992 22798 5001
rect 22742 4927 22798 4936
rect 22848 4593 22876 8298
rect 22940 8090 22968 8871
rect 23032 8634 23060 9114
rect 23020 8628 23072 8634
rect 23020 8570 23072 8576
rect 22928 8084 22980 8090
rect 22928 8026 22980 8032
rect 22928 7472 22980 7478
rect 22928 7414 22980 7420
rect 22940 4622 22968 7414
rect 23124 7018 23152 9143
rect 23032 6990 23152 7018
rect 22928 4616 22980 4622
rect 22834 4584 22890 4593
rect 22928 4558 22980 4564
rect 22834 4519 22890 4528
rect 22650 3768 22706 3777
rect 22848 3738 22876 4519
rect 22940 4282 22968 4558
rect 22928 4276 22980 4282
rect 22928 4218 22980 4224
rect 23032 4162 23060 6990
rect 23112 6928 23164 6934
rect 23112 6870 23164 6876
rect 23124 6458 23152 6870
rect 23112 6452 23164 6458
rect 23112 6394 23164 6400
rect 23216 5794 23244 10934
rect 23294 10840 23350 10849
rect 23294 10775 23350 10784
rect 23308 10146 23336 10775
rect 23492 10577 23520 16510
rect 23572 15904 23624 15910
rect 23572 15846 23624 15852
rect 23584 15609 23612 15846
rect 23570 15600 23626 15609
rect 23570 15535 23626 15544
rect 23572 15088 23624 15094
rect 23572 15030 23624 15036
rect 23584 14550 23612 15030
rect 23572 14544 23624 14550
rect 23572 14486 23624 14492
rect 23572 13796 23624 13802
rect 23572 13738 23624 13744
rect 23584 13394 23612 13738
rect 23572 13388 23624 13394
rect 23572 13330 23624 13336
rect 23570 12744 23626 12753
rect 23570 12679 23572 12688
rect 23624 12679 23626 12688
rect 23572 12650 23624 12656
rect 23570 12472 23626 12481
rect 23570 12407 23626 12416
rect 23584 11898 23612 12407
rect 23572 11892 23624 11898
rect 23572 11834 23624 11840
rect 23572 11552 23624 11558
rect 23572 11494 23624 11500
rect 23478 10568 23534 10577
rect 23478 10503 23534 10512
rect 23308 10130 23428 10146
rect 23308 10124 23440 10130
rect 23308 10118 23388 10124
rect 23388 10066 23440 10072
rect 23400 9654 23428 10066
rect 23480 9988 23532 9994
rect 23480 9930 23532 9936
rect 23492 9897 23520 9930
rect 23478 9888 23534 9897
rect 23478 9823 23534 9832
rect 23388 9648 23440 9654
rect 23388 9590 23440 9596
rect 23294 9480 23350 9489
rect 23294 9415 23350 9424
rect 23308 9110 23336 9415
rect 23492 9178 23520 9823
rect 23480 9172 23532 9178
rect 23480 9114 23532 9120
rect 23296 9104 23348 9110
rect 23584 9058 23612 11494
rect 23676 10996 23704 17750
rect 23756 17332 23808 17338
rect 23756 17274 23808 17280
rect 23768 16794 23796 17274
rect 23756 16788 23808 16794
rect 23756 16730 23808 16736
rect 23756 16652 23808 16658
rect 23756 16594 23808 16600
rect 23768 16454 23796 16594
rect 23756 16448 23808 16454
rect 23756 16390 23808 16396
rect 23860 16402 23888 21542
rect 23940 21548 23992 21554
rect 23940 21490 23992 21496
rect 23952 18850 23980 21490
rect 24044 19922 24072 21898
rect 24032 19916 24084 19922
rect 24032 19858 24084 19864
rect 24044 19825 24072 19858
rect 24030 19816 24086 19825
rect 24030 19751 24086 19760
rect 24032 19712 24084 19718
rect 24032 19654 24084 19660
rect 24044 19310 24072 19654
rect 24136 19310 24164 25094
rect 24228 24721 24256 25214
rect 25044 25220 25096 25226
rect 25044 25162 25096 25168
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 25056 24818 25084 25162
rect 26238 24848 26294 24857
rect 25044 24812 25096 24818
rect 26238 24783 26294 24792
rect 25044 24754 25096 24760
rect 24214 24712 24270 24721
rect 25778 24712 25834 24721
rect 24584 24676 24636 24682
rect 24214 24647 24270 24656
rect 24504 24636 24584 24664
rect 24504 24313 24532 24636
rect 25778 24647 25834 24656
rect 24584 24618 24636 24624
rect 24676 24608 24728 24614
rect 24676 24550 24728 24556
rect 24490 24304 24546 24313
rect 24490 24239 24492 24248
rect 24544 24239 24546 24248
rect 24492 24210 24544 24216
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24308 23724 24360 23730
rect 24308 23666 24360 23672
rect 24320 23497 24348 23666
rect 24306 23488 24362 23497
rect 24306 23423 24362 23432
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24216 21684 24268 21690
rect 24216 21626 24268 21632
rect 24032 19304 24084 19310
rect 24032 19246 24084 19252
rect 24124 19304 24176 19310
rect 24124 19246 24176 19252
rect 24044 18970 24072 19246
rect 24228 18986 24256 21626
rect 24688 21162 24716 24550
rect 24952 24268 25004 24274
rect 24952 24210 25004 24216
rect 24964 23866 24992 24210
rect 25134 24168 25190 24177
rect 25134 24103 25136 24112
rect 25188 24103 25190 24112
rect 25136 24074 25188 24080
rect 24952 23860 25004 23866
rect 24952 23802 25004 23808
rect 25226 23760 25282 23769
rect 25226 23695 25282 23704
rect 25240 23662 25268 23695
rect 24860 23656 24912 23662
rect 24860 23598 24912 23604
rect 25228 23656 25280 23662
rect 25228 23598 25280 23604
rect 25410 23624 25466 23633
rect 24872 23322 24900 23598
rect 25410 23559 25466 23568
rect 25424 23526 25452 23559
rect 25412 23520 25464 23526
rect 25412 23462 25464 23468
rect 25318 23352 25374 23361
rect 24860 23316 24912 23322
rect 25318 23287 25374 23296
rect 24860 23258 24912 23264
rect 25332 23254 25360 23287
rect 25320 23248 25372 23254
rect 25320 23190 25372 23196
rect 25044 23180 25096 23186
rect 25044 23122 25096 23128
rect 24860 22976 24912 22982
rect 24860 22918 24912 22924
rect 24872 22642 24900 22918
rect 25056 22710 25084 23122
rect 25320 23112 25372 23118
rect 25320 23054 25372 23060
rect 25410 23080 25466 23089
rect 25044 22704 25096 22710
rect 25042 22672 25044 22681
rect 25096 22672 25098 22681
rect 24860 22636 24912 22642
rect 25042 22607 25098 22616
rect 24860 22578 24912 22584
rect 24872 22234 24900 22578
rect 24860 22228 24912 22234
rect 24860 22170 24912 22176
rect 24768 22092 24820 22098
rect 24768 22034 24820 22040
rect 24780 21350 24808 22034
rect 24952 22024 25004 22030
rect 24952 21966 25004 21972
rect 24768 21344 24820 21350
rect 24768 21286 24820 21292
rect 24688 21146 24900 21162
rect 24688 21140 24912 21146
rect 24688 21134 24860 21140
rect 24860 21082 24912 21088
rect 24964 21078 24992 21966
rect 25332 21078 25360 23054
rect 25410 23015 25466 23024
rect 25424 21690 25452 23015
rect 25502 22536 25558 22545
rect 25502 22471 25558 22480
rect 25412 21684 25464 21690
rect 25412 21626 25464 21632
rect 25412 21140 25464 21146
rect 25412 21082 25464 21088
rect 24952 21072 25004 21078
rect 24952 21014 25004 21020
rect 25320 21072 25372 21078
rect 25320 21014 25372 21020
rect 24676 20936 24728 20942
rect 24676 20878 24728 20884
rect 25044 20936 25096 20942
rect 25044 20878 25096 20884
rect 25226 20904 25282 20913
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24688 20534 24716 20878
rect 24860 20800 24912 20806
rect 24860 20742 24912 20748
rect 24676 20528 24728 20534
rect 24676 20470 24728 20476
rect 24584 20460 24636 20466
rect 24584 20402 24636 20408
rect 24490 20088 24546 20097
rect 24490 20023 24492 20032
rect 24544 20023 24546 20032
rect 24492 19994 24544 20000
rect 24596 19854 24624 20402
rect 24768 20392 24820 20398
rect 24872 20380 24900 20742
rect 24820 20352 24900 20380
rect 24768 20334 24820 20340
rect 24952 20324 25004 20330
rect 24952 20266 25004 20272
rect 24964 20233 24992 20266
rect 24950 20224 25006 20233
rect 24950 20159 25006 20168
rect 24860 20052 24912 20058
rect 24860 19994 24912 20000
rect 24584 19848 24636 19854
rect 24584 19790 24636 19796
rect 24768 19712 24820 19718
rect 24674 19680 24730 19689
rect 24289 19612 24585 19632
rect 24768 19654 24820 19660
rect 24674 19615 24730 19624
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24584 19372 24636 19378
rect 24584 19314 24636 19320
rect 24032 18964 24084 18970
rect 24228 18958 24348 18986
rect 24032 18906 24084 18912
rect 24216 18896 24268 18902
rect 23952 18822 24072 18850
rect 24216 18838 24268 18844
rect 23940 18692 23992 18698
rect 23940 18634 23992 18640
rect 23952 18465 23980 18634
rect 23938 18456 23994 18465
rect 23938 18391 23994 18400
rect 24044 18306 24072 18822
rect 24124 18828 24176 18834
rect 24124 18770 24176 18776
rect 23952 18278 24072 18306
rect 23952 16674 23980 18278
rect 24136 18086 24164 18770
rect 24228 18154 24256 18838
rect 24320 18737 24348 18958
rect 24596 18873 24624 19314
rect 24582 18864 24638 18873
rect 24582 18799 24638 18808
rect 24306 18728 24362 18737
rect 24306 18663 24362 18672
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24216 18148 24268 18154
rect 24216 18090 24268 18096
rect 24124 18080 24176 18086
rect 24124 18022 24176 18028
rect 24032 17876 24084 17882
rect 24032 17818 24084 17824
rect 24044 17338 24072 17818
rect 24032 17332 24084 17338
rect 24032 17274 24084 17280
rect 24136 17134 24164 18022
rect 24688 17814 24716 19615
rect 24780 17898 24808 19654
rect 24872 18902 24900 19994
rect 25056 19718 25084 20878
rect 25226 20839 25282 20848
rect 25136 20596 25188 20602
rect 25136 20538 25188 20544
rect 25044 19712 25096 19718
rect 25044 19654 25096 19660
rect 25044 19440 25096 19446
rect 25044 19382 25096 19388
rect 24860 18896 24912 18902
rect 24860 18838 24912 18844
rect 24952 18692 25004 18698
rect 24952 18634 25004 18640
rect 24964 18426 24992 18634
rect 24952 18420 25004 18426
rect 24952 18362 25004 18368
rect 24780 17870 24900 17898
rect 24676 17808 24728 17814
rect 24676 17750 24728 17756
rect 24768 17740 24820 17746
rect 24768 17682 24820 17688
rect 24676 17672 24728 17678
rect 24676 17614 24728 17620
rect 24216 17536 24268 17542
rect 24216 17478 24268 17484
rect 24228 17202 24256 17478
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24216 17196 24268 17202
rect 24216 17138 24268 17144
rect 24124 17128 24176 17134
rect 24228 17105 24256 17138
rect 24124 17070 24176 17076
rect 24214 17096 24270 17105
rect 24214 17031 24270 17040
rect 24400 17060 24452 17066
rect 24400 17002 24452 17008
rect 24308 16992 24360 16998
rect 24308 16934 24360 16940
rect 23952 16646 24256 16674
rect 24032 16584 24084 16590
rect 24030 16552 24032 16561
rect 24084 16552 24086 16561
rect 24030 16487 24086 16496
rect 24124 16516 24176 16522
rect 24124 16458 24176 16464
rect 23768 16250 23796 16390
rect 23860 16374 23980 16402
rect 23846 16280 23902 16289
rect 23756 16244 23808 16250
rect 23846 16215 23902 16224
rect 23756 16186 23808 16192
rect 23754 16144 23810 16153
rect 23860 16114 23888 16215
rect 23754 16079 23810 16088
rect 23848 16108 23900 16114
rect 23768 15638 23796 16079
rect 23848 16050 23900 16056
rect 23848 15904 23900 15910
rect 23846 15872 23848 15881
rect 23900 15872 23902 15881
rect 23846 15807 23902 15816
rect 23756 15632 23808 15638
rect 23756 15574 23808 15580
rect 23860 15502 23888 15807
rect 23848 15496 23900 15502
rect 23768 15456 23848 15484
rect 23768 13734 23796 15456
rect 23848 15438 23900 15444
rect 23848 14408 23900 14414
rect 23848 14350 23900 14356
rect 23860 13802 23888 14350
rect 23952 13870 23980 16374
rect 24032 15496 24084 15502
rect 24032 15438 24084 15444
rect 24044 15337 24072 15438
rect 24030 15328 24086 15337
rect 24030 15263 24086 15272
rect 24136 15144 24164 16458
rect 24044 15116 24164 15144
rect 24044 14906 24072 15116
rect 24122 15056 24178 15065
rect 24122 14991 24124 15000
rect 24176 14991 24178 15000
rect 24124 14962 24176 14968
rect 24044 14878 24164 14906
rect 24032 14816 24084 14822
rect 24032 14758 24084 14764
rect 24044 14618 24072 14758
rect 24032 14612 24084 14618
rect 24032 14554 24084 14560
rect 24136 14550 24164 14878
rect 24124 14544 24176 14550
rect 24124 14486 24176 14492
rect 24122 14376 24178 14385
rect 24122 14311 24178 14320
rect 23940 13864 23992 13870
rect 23940 13806 23992 13812
rect 23848 13796 23900 13802
rect 23848 13738 23900 13744
rect 23756 13728 23808 13734
rect 23756 13670 23808 13676
rect 23952 13530 23980 13806
rect 24136 13705 24164 14311
rect 24122 13696 24178 13705
rect 24122 13631 24178 13640
rect 24228 13546 24256 16646
rect 24320 16522 24348 16934
rect 24412 16794 24440 17002
rect 24400 16788 24452 16794
rect 24400 16730 24452 16736
rect 24308 16516 24360 16522
rect 24308 16458 24360 16464
rect 24688 16454 24716 17614
rect 24780 17377 24808 17682
rect 24766 17368 24822 17377
rect 24766 17303 24768 17312
rect 24820 17303 24822 17312
rect 24768 17274 24820 17280
rect 24780 17243 24808 17274
rect 24872 17082 24900 17870
rect 24952 17604 25004 17610
rect 24952 17546 25004 17552
rect 24780 17054 24900 17082
rect 24676 16448 24728 16454
rect 24676 16390 24728 16396
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24688 16046 24716 16390
rect 24676 16040 24728 16046
rect 24676 15982 24728 15988
rect 24676 15632 24728 15638
rect 24676 15574 24728 15580
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24688 15162 24716 15574
rect 24676 15156 24728 15162
rect 24676 15098 24728 15104
rect 24306 15056 24362 15065
rect 24780 15042 24808 17054
rect 24860 16584 24912 16590
rect 24860 16526 24912 16532
rect 24872 16250 24900 16526
rect 24860 16244 24912 16250
rect 24860 16186 24912 16192
rect 24860 15972 24912 15978
rect 24860 15914 24912 15920
rect 24306 14991 24362 15000
rect 24688 15014 24808 15042
rect 24320 14385 24348 14991
rect 24584 14612 24636 14618
rect 24584 14554 24636 14560
rect 24596 14521 24624 14554
rect 24582 14512 24638 14521
rect 24582 14447 24638 14456
rect 24306 14376 24362 14385
rect 24306 14311 24362 14320
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24688 13954 24716 15014
rect 24766 14648 24822 14657
rect 24872 14634 24900 15914
rect 24964 15042 24992 17546
rect 25056 16289 25084 19382
rect 25148 19174 25176 20538
rect 25240 20398 25268 20839
rect 25332 20534 25360 21014
rect 25320 20528 25372 20534
rect 25320 20470 25372 20476
rect 25228 20392 25280 20398
rect 25228 20334 25280 20340
rect 25240 19990 25268 20334
rect 25318 20088 25374 20097
rect 25424 20058 25452 21082
rect 25318 20023 25374 20032
rect 25412 20052 25464 20058
rect 25228 19984 25280 19990
rect 25228 19926 25280 19932
rect 25136 19168 25188 19174
rect 25136 19110 25188 19116
rect 25136 18624 25188 18630
rect 25136 18566 25188 18572
rect 25042 16280 25098 16289
rect 25042 16215 25098 16224
rect 25044 16108 25096 16114
rect 25044 16050 25096 16056
rect 25056 15706 25084 16050
rect 25044 15700 25096 15706
rect 25044 15642 25096 15648
rect 24964 15014 25084 15042
rect 24952 14884 25004 14890
rect 24952 14826 25004 14832
rect 24822 14606 24900 14634
rect 24766 14583 24822 14592
rect 24860 14544 24912 14550
rect 24860 14486 24912 14492
rect 24872 14074 24900 14486
rect 24860 14068 24912 14074
rect 24860 14010 24912 14016
rect 23940 13524 23992 13530
rect 23940 13466 23992 13472
rect 24136 13518 24256 13546
rect 24412 13926 24716 13954
rect 23754 13424 23810 13433
rect 23938 13424 23994 13433
rect 23754 13359 23810 13368
rect 23860 13368 23938 13376
rect 23860 13359 23994 13368
rect 23768 12986 23796 13359
rect 23860 13348 23980 13359
rect 23860 13161 23888 13348
rect 24136 13308 24164 13518
rect 24412 13308 24440 13926
rect 23952 13280 24164 13308
rect 24228 13280 24440 13308
rect 23846 13152 23902 13161
rect 23846 13087 23902 13096
rect 23756 12980 23808 12986
rect 23756 12922 23808 12928
rect 23768 11830 23796 12922
rect 23848 12300 23900 12306
rect 23848 12242 23900 12248
rect 23756 11824 23808 11830
rect 23756 11766 23808 11772
rect 23756 11620 23808 11626
rect 23756 11562 23808 11568
rect 23768 11121 23796 11562
rect 23860 11354 23888 12242
rect 23848 11348 23900 11354
rect 23848 11290 23900 11296
rect 23952 11286 23980 13280
rect 24124 13184 24176 13190
rect 24124 13126 24176 13132
rect 24136 12782 24164 13126
rect 24124 12776 24176 12782
rect 24124 12718 24176 12724
rect 24032 11348 24084 11354
rect 24032 11290 24084 11296
rect 23940 11280 23992 11286
rect 23940 11222 23992 11228
rect 23754 11112 23810 11121
rect 23754 11047 23810 11056
rect 23676 10968 23888 10996
rect 23860 10656 23888 10968
rect 23952 10810 23980 11222
rect 23940 10804 23992 10810
rect 23940 10746 23992 10752
rect 23768 10628 23888 10656
rect 23662 10296 23718 10305
rect 23768 10266 23796 10628
rect 24044 10470 24072 11290
rect 24032 10464 24084 10470
rect 24032 10406 24084 10412
rect 24122 10432 24178 10441
rect 23662 10231 23718 10240
rect 23756 10260 23808 10266
rect 23676 10010 23704 10231
rect 23756 10202 23808 10208
rect 23940 10260 23992 10266
rect 23940 10202 23992 10208
rect 23754 10160 23810 10169
rect 23754 10095 23756 10104
rect 23808 10095 23810 10104
rect 23756 10066 23808 10072
rect 23848 10056 23900 10062
rect 23676 9982 23796 10010
rect 23848 9998 23900 10004
rect 23662 9752 23718 9761
rect 23662 9687 23718 9696
rect 23296 9046 23348 9052
rect 23308 8566 23336 9046
rect 23492 9030 23612 9058
rect 23296 8560 23348 8566
rect 23296 8502 23348 8508
rect 23308 8090 23336 8502
rect 23388 8288 23440 8294
rect 23388 8230 23440 8236
rect 23296 8084 23348 8090
rect 23296 8026 23348 8032
rect 23400 7954 23428 8230
rect 23388 7948 23440 7954
rect 23388 7890 23440 7896
rect 23400 7857 23428 7890
rect 23386 7848 23442 7857
rect 23386 7783 23442 7792
rect 23296 7744 23348 7750
rect 23296 7686 23348 7692
rect 23308 6882 23336 7686
rect 23400 7546 23428 7783
rect 23388 7540 23440 7546
rect 23388 7482 23440 7488
rect 23492 7313 23520 9030
rect 23570 8936 23626 8945
rect 23570 8871 23626 8880
rect 23584 7954 23612 8871
rect 23676 8634 23704 9687
rect 23664 8628 23716 8634
rect 23664 8570 23716 8576
rect 23664 8424 23716 8430
rect 23768 8401 23796 9982
rect 23664 8366 23716 8372
rect 23754 8392 23810 8401
rect 23572 7948 23624 7954
rect 23572 7890 23624 7896
rect 23478 7304 23534 7313
rect 23478 7239 23534 7248
rect 23308 6854 23520 6882
rect 23296 6792 23348 6798
rect 23296 6734 23348 6740
rect 23308 6254 23336 6734
rect 23386 6488 23442 6497
rect 23386 6423 23388 6432
rect 23440 6423 23442 6432
rect 23388 6394 23440 6400
rect 23296 6248 23348 6254
rect 23296 6190 23348 6196
rect 22940 4134 23060 4162
rect 23124 5766 23244 5794
rect 23308 5778 23336 6190
rect 23400 6186 23428 6394
rect 23388 6180 23440 6186
rect 23388 6122 23440 6128
rect 23400 5914 23428 6122
rect 23492 5914 23520 6854
rect 23388 5908 23440 5914
rect 23388 5850 23440 5856
rect 23480 5908 23532 5914
rect 23480 5850 23532 5856
rect 23572 5840 23624 5846
rect 23570 5808 23572 5817
rect 23624 5808 23626 5817
rect 23296 5772 23348 5778
rect 22650 3703 22706 3712
rect 22836 3732 22888 3738
rect 22836 3674 22888 3680
rect 21732 3470 21784 3476
rect 21272 3392 21324 3398
rect 21272 3334 21324 3340
rect 21640 3392 21692 3398
rect 21640 3334 21692 3340
rect 21178 3224 21234 3233
rect 20904 3188 20956 3194
rect 21178 3159 21180 3168
rect 20904 3130 20956 3136
rect 21232 3159 21234 3168
rect 21180 3130 21232 3136
rect 20916 2990 20944 3130
rect 20904 2984 20956 2990
rect 20904 2926 20956 2932
rect 21546 2952 21602 2961
rect 20996 2916 21048 2922
rect 21546 2887 21602 2896
rect 20996 2858 21048 2864
rect 20812 2644 20864 2650
rect 20812 2586 20864 2592
rect 20904 2576 20956 2582
rect 20904 2518 20956 2524
rect 20536 2440 20588 2446
rect 20534 2408 20536 2417
rect 20588 2408 20590 2417
rect 20534 2343 20590 2352
rect 20916 2310 20944 2518
rect 20904 2304 20956 2310
rect 20904 2246 20956 2252
rect 20916 1737 20944 2246
rect 20902 1728 20958 1737
rect 20902 1663 20958 1672
rect 21008 1193 21036 2858
rect 21180 2644 21232 2650
rect 21180 2586 21232 2592
rect 21192 2553 21220 2586
rect 21178 2544 21234 2553
rect 21178 2479 21234 2488
rect 21086 2000 21142 2009
rect 21086 1935 21142 1944
rect 21100 1737 21128 1935
rect 21086 1728 21142 1737
rect 21086 1663 21142 1672
rect 20994 1184 21050 1193
rect 20994 1119 21050 1128
rect 20916 598 21036 626
rect 14186 96 14242 105
rect 14186 31 14242 40
rect 14370 0 14426 480
rect 14922 0 14978 480
rect 15474 0 15530 480
rect 16026 0 16082 480
rect 16578 0 16634 480
rect 17130 0 17186 480
rect 17682 0 17738 480
rect 18234 0 18290 480
rect 18786 0 18842 480
rect 19338 0 19394 480
rect 19890 0 19946 480
rect 20442 0 20498 480
rect 20916 105 20944 598
rect 21008 480 21036 598
rect 21560 480 21588 2887
rect 21652 2553 21680 3334
rect 21744 3126 21772 3470
rect 22020 3466 22232 3482
rect 22008 3460 22232 3466
rect 22060 3454 22232 3460
rect 22558 3496 22614 3505
rect 22558 3431 22614 3440
rect 22008 3402 22060 3408
rect 22468 3392 22520 3398
rect 22466 3360 22468 3369
rect 22520 3360 22522 3369
rect 22466 3295 22522 3304
rect 22848 3194 22876 3674
rect 22836 3188 22888 3194
rect 22836 3130 22888 3136
rect 21732 3120 21784 3126
rect 21732 3062 21784 3068
rect 21638 2544 21694 2553
rect 21638 2479 21694 2488
rect 21744 2446 21772 3062
rect 22098 2952 22154 2961
rect 22098 2887 22154 2896
rect 21732 2440 21784 2446
rect 21732 2382 21784 2388
rect 22112 480 22140 2887
rect 22558 2816 22614 2825
rect 22558 2751 22614 2760
rect 22572 1850 22600 2751
rect 22940 2514 22968 4134
rect 23124 3738 23152 5766
rect 23296 5714 23348 5720
rect 23480 5772 23532 5778
rect 23570 5743 23626 5752
rect 23480 5714 23532 5720
rect 23202 5672 23258 5681
rect 23202 5607 23258 5616
rect 23112 3732 23164 3738
rect 23032 3692 23112 3720
rect 23032 3194 23060 3692
rect 23112 3674 23164 3680
rect 23112 3528 23164 3534
rect 23112 3470 23164 3476
rect 23020 3188 23072 3194
rect 23020 3130 23072 3136
rect 23124 3058 23152 3470
rect 23112 3052 23164 3058
rect 23112 2994 23164 3000
rect 23018 2816 23074 2825
rect 23018 2751 23074 2760
rect 23032 2650 23060 2751
rect 23020 2644 23072 2650
rect 23020 2586 23072 2592
rect 22928 2508 22980 2514
rect 22928 2450 22980 2456
rect 22572 1822 22692 1850
rect 22664 480 22692 1822
rect 23216 480 23244 5607
rect 23492 5386 23520 5714
rect 23676 5658 23704 8366
rect 23754 8327 23810 8336
rect 23860 7993 23888 9998
rect 23952 9382 23980 10202
rect 24044 9722 24072 10406
rect 24122 10367 24178 10376
rect 24032 9716 24084 9722
rect 24032 9658 24084 9664
rect 23940 9376 23992 9382
rect 23940 9318 23992 9324
rect 24136 9178 24164 10367
rect 24124 9172 24176 9178
rect 24044 9132 24124 9160
rect 23940 8832 23992 8838
rect 23940 8774 23992 8780
rect 23846 7984 23902 7993
rect 23756 7948 23808 7954
rect 23846 7919 23902 7928
rect 23756 7890 23808 7896
rect 23768 7342 23796 7890
rect 23952 7698 23980 8774
rect 24044 8090 24072 9132
rect 24124 9114 24176 9120
rect 24124 8832 24176 8838
rect 24124 8774 24176 8780
rect 24136 8673 24164 8774
rect 24122 8664 24178 8673
rect 24122 8599 24178 8608
rect 24136 8498 24164 8599
rect 24124 8492 24176 8498
rect 24124 8434 24176 8440
rect 24228 8090 24256 13280
rect 24768 13252 24820 13258
rect 24768 13194 24820 13200
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24780 12986 24808 13194
rect 24768 12980 24820 12986
rect 24768 12922 24820 12928
rect 24676 12912 24728 12918
rect 24676 12854 24728 12860
rect 24306 12608 24362 12617
rect 24306 12543 24362 12552
rect 24320 12442 24348 12543
rect 24688 12481 24716 12854
rect 24674 12472 24730 12481
rect 24308 12436 24360 12442
rect 24674 12407 24730 12416
rect 24308 12378 24360 12384
rect 24964 12374 24992 14826
rect 25056 13530 25084 15014
rect 25148 13852 25176 18566
rect 25228 17808 25280 17814
rect 25228 17750 25280 17756
rect 25240 16998 25268 17750
rect 25228 16992 25280 16998
rect 25228 16934 25280 16940
rect 25228 16720 25280 16726
rect 25226 16688 25228 16697
rect 25280 16688 25282 16697
rect 25226 16623 25282 16632
rect 25228 16244 25280 16250
rect 25228 16186 25280 16192
rect 25240 15502 25268 16186
rect 25228 15496 25280 15502
rect 25228 15438 25280 15444
rect 25228 14272 25280 14278
rect 25228 14214 25280 14220
rect 25240 13977 25268 14214
rect 25226 13968 25282 13977
rect 25226 13903 25282 13912
rect 25148 13824 25268 13852
rect 25044 13524 25096 13530
rect 25096 13484 25176 13512
rect 25044 13466 25096 13472
rect 25044 13320 25096 13326
rect 25044 13262 25096 13268
rect 25056 12889 25084 13262
rect 25148 12986 25176 13484
rect 25136 12980 25188 12986
rect 25136 12922 25188 12928
rect 25042 12880 25098 12889
rect 25042 12815 25044 12824
rect 25096 12815 25098 12824
rect 25044 12786 25096 12792
rect 25136 12776 25188 12782
rect 25136 12718 25188 12724
rect 25044 12436 25096 12442
rect 25044 12378 25096 12384
rect 24952 12368 25004 12374
rect 25056 12345 25084 12378
rect 24952 12310 25004 12316
rect 25042 12336 25098 12345
rect 24860 12300 24912 12306
rect 25042 12271 25098 12280
rect 24860 12242 24912 12248
rect 24768 12096 24820 12102
rect 24674 12064 24730 12073
rect 24289 11996 24585 12016
rect 24768 12038 24820 12044
rect 24674 11999 24730 12008
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24688 10266 24716 11999
rect 24780 10266 24808 12038
rect 24872 11694 24900 12242
rect 25148 12209 25176 12718
rect 25134 12200 25190 12209
rect 25134 12135 25190 12144
rect 25240 11914 25268 13824
rect 25148 11886 25268 11914
rect 25332 11898 25360 20023
rect 25412 19994 25464 20000
rect 25516 18426 25544 22471
rect 25686 21584 25742 21593
rect 25686 21519 25742 21528
rect 25594 21176 25650 21185
rect 25594 21111 25650 21120
rect 25504 18420 25556 18426
rect 25504 18362 25556 18368
rect 25412 16992 25464 16998
rect 25412 16934 25464 16940
rect 25504 16992 25556 16998
rect 25504 16934 25556 16940
rect 25424 16697 25452 16934
rect 25410 16688 25466 16697
rect 25410 16623 25466 16632
rect 25412 14952 25464 14958
rect 25412 14894 25464 14900
rect 25320 11892 25372 11898
rect 24860 11688 24912 11694
rect 24860 11630 24912 11636
rect 24872 11354 24900 11630
rect 24860 11348 24912 11354
rect 24860 11290 24912 11296
rect 24860 10600 24912 10606
rect 24860 10542 24912 10548
rect 24872 10305 24900 10542
rect 24858 10296 24914 10305
rect 24676 10260 24728 10266
rect 24676 10202 24728 10208
rect 24768 10260 24820 10266
rect 24858 10231 24914 10240
rect 24768 10202 24820 10208
rect 24688 10062 24716 10202
rect 24952 10124 25004 10130
rect 24952 10066 25004 10072
rect 24676 10056 24728 10062
rect 24964 10033 24992 10066
rect 24676 9998 24728 10004
rect 24950 10024 25006 10033
rect 24950 9959 25006 9968
rect 24768 9920 24820 9926
rect 24768 9862 24820 9868
rect 24952 9920 25004 9926
rect 24952 9862 25004 9868
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24780 9518 24808 9862
rect 24858 9752 24914 9761
rect 24858 9687 24914 9696
rect 24964 9704 24992 9862
rect 24872 9654 24900 9687
rect 24964 9676 25084 9704
rect 24860 9648 24912 9654
rect 24860 9590 24912 9596
rect 24768 9512 24820 9518
rect 24768 9454 24820 9460
rect 24398 9208 24454 9217
rect 24398 9143 24454 9152
rect 24412 9042 24440 9143
rect 24674 9072 24730 9081
rect 24400 9036 24452 9042
rect 24674 9007 24730 9016
rect 24400 8978 24452 8984
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24032 8084 24084 8090
rect 24032 8026 24084 8032
rect 24216 8084 24268 8090
rect 24216 8026 24268 8032
rect 24122 7984 24178 7993
rect 24122 7919 24178 7928
rect 23860 7670 23980 7698
rect 23756 7336 23808 7342
rect 23756 7278 23808 7284
rect 23756 7200 23808 7206
rect 23756 7142 23808 7148
rect 23768 6497 23796 7142
rect 23754 6488 23810 6497
rect 23754 6423 23810 6432
rect 23756 5908 23808 5914
rect 23756 5850 23808 5856
rect 23400 5370 23520 5386
rect 23388 5364 23520 5370
rect 23440 5358 23520 5364
rect 23388 5306 23440 5312
rect 23294 4992 23350 5001
rect 23294 4927 23350 4936
rect 23308 2802 23336 4927
rect 23388 4820 23440 4826
rect 23388 4762 23440 4768
rect 23400 3618 23428 4762
rect 23492 3738 23520 5358
rect 23584 5630 23704 5658
rect 23584 5302 23612 5630
rect 23662 5536 23718 5545
rect 23662 5471 23718 5480
rect 23676 5370 23704 5471
rect 23664 5364 23716 5370
rect 23664 5306 23716 5312
rect 23572 5296 23624 5302
rect 23572 5238 23624 5244
rect 23768 5234 23796 5850
rect 23860 5409 23888 7670
rect 23938 7576 23994 7585
rect 23938 7511 23940 7520
rect 23992 7511 23994 7520
rect 23940 7482 23992 7488
rect 23940 7336 23992 7342
rect 23940 7278 23992 7284
rect 23952 5828 23980 7278
rect 24136 7274 24164 7919
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24306 7304 24362 7313
rect 24124 7268 24176 7274
rect 24306 7239 24362 7248
rect 24124 7210 24176 7216
rect 23952 5800 24072 5828
rect 23938 5536 23994 5545
rect 23938 5471 23994 5480
rect 23846 5400 23902 5409
rect 23846 5335 23902 5344
rect 23848 5296 23900 5302
rect 23848 5238 23900 5244
rect 23756 5228 23808 5234
rect 23756 5170 23808 5176
rect 23664 5160 23716 5166
rect 23664 5102 23716 5108
rect 23572 4548 23624 4554
rect 23572 4490 23624 4496
rect 23480 3732 23532 3738
rect 23480 3674 23532 3680
rect 23400 3590 23520 3618
rect 23492 2922 23520 3590
rect 23480 2916 23532 2922
rect 23480 2858 23532 2864
rect 23308 2774 23520 2802
rect 23492 2417 23520 2774
rect 23478 2408 23534 2417
rect 23478 2343 23534 2352
rect 23584 2145 23612 4490
rect 23676 4026 23704 5102
rect 23768 4214 23796 5170
rect 23756 4208 23808 4214
rect 23756 4150 23808 4156
rect 23860 4026 23888 5238
rect 23952 4808 23980 5471
rect 24044 5098 24072 5800
rect 24136 5302 24164 7210
rect 24320 6712 24348 7239
rect 24228 6684 24348 6712
rect 24124 5296 24176 5302
rect 24124 5238 24176 5244
rect 24032 5092 24084 5098
rect 24084 5052 24164 5080
rect 24032 5034 24084 5040
rect 24136 4826 24164 5052
rect 24124 4820 24176 4826
rect 23952 4780 24072 4808
rect 23940 4684 23992 4690
rect 23940 4626 23992 4632
rect 23952 4321 23980 4626
rect 23938 4312 23994 4321
rect 23938 4247 23994 4256
rect 23952 4214 23980 4247
rect 23940 4208 23992 4214
rect 23940 4150 23992 4156
rect 23676 3998 23796 4026
rect 23860 3998 23980 4026
rect 23664 3936 23716 3942
rect 23662 3904 23664 3913
rect 23716 3904 23718 3913
rect 23662 3839 23718 3848
rect 23768 3194 23796 3998
rect 23756 3188 23808 3194
rect 23756 3130 23808 3136
rect 23664 3120 23716 3126
rect 23662 3088 23664 3097
rect 23716 3088 23718 3097
rect 23768 3074 23796 3130
rect 23768 3046 23888 3074
rect 23662 3023 23718 3032
rect 23860 2990 23888 3046
rect 23848 2984 23900 2990
rect 23754 2952 23810 2961
rect 23848 2926 23900 2932
rect 23754 2887 23810 2896
rect 23570 2136 23626 2145
rect 23570 2071 23626 2080
rect 23768 480 23796 2887
rect 23848 2848 23900 2854
rect 23848 2790 23900 2796
rect 23860 921 23888 2790
rect 23952 1601 23980 3998
rect 24044 3210 24072 4780
rect 24124 4762 24176 4768
rect 24124 4616 24176 4622
rect 24124 4558 24176 4564
rect 24136 4010 24164 4558
rect 24228 4146 24256 6684
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24582 6352 24638 6361
rect 24582 6287 24638 6296
rect 24596 5710 24624 6287
rect 24688 5817 24716 9007
rect 24780 6730 24808 9454
rect 24860 9036 24912 9042
rect 24860 8978 24912 8984
rect 24872 8634 24900 8978
rect 24952 8900 25004 8906
rect 24952 8842 25004 8848
rect 24964 8634 24992 8842
rect 24860 8628 24912 8634
rect 24860 8570 24912 8576
rect 24952 8628 25004 8634
rect 24952 8570 25004 8576
rect 24860 8492 24912 8498
rect 24860 8434 24912 8440
rect 24872 7818 24900 8434
rect 24952 7880 25004 7886
rect 24952 7822 25004 7828
rect 24860 7812 24912 7818
rect 24860 7754 24912 7760
rect 24872 7410 24900 7754
rect 24860 7404 24912 7410
rect 24860 7346 24912 7352
rect 24872 6934 24900 7346
rect 24964 7342 24992 7822
rect 24952 7336 25004 7342
rect 24952 7278 25004 7284
rect 25056 7018 25084 9676
rect 24964 6990 25084 7018
rect 24860 6928 24912 6934
rect 24860 6870 24912 6876
rect 24768 6724 24820 6730
rect 24768 6666 24820 6672
rect 24860 6656 24912 6662
rect 24860 6598 24912 6604
rect 24872 6254 24900 6598
rect 24860 6248 24912 6254
rect 24860 6190 24912 6196
rect 24674 5808 24730 5817
rect 24674 5743 24730 5752
rect 24768 5772 24820 5778
rect 24768 5714 24820 5720
rect 24584 5704 24636 5710
rect 24636 5652 24716 5658
rect 24584 5646 24716 5652
rect 24596 5630 24716 5646
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24688 5370 24716 5630
rect 24676 5364 24728 5370
rect 24676 5306 24728 5312
rect 24780 4978 24808 5714
rect 24860 5568 24912 5574
rect 24858 5536 24860 5545
rect 24912 5536 24914 5545
rect 24858 5471 24914 5480
rect 24860 5024 24912 5030
rect 24780 4972 24860 4978
rect 24780 4966 24912 4972
rect 24780 4950 24900 4966
rect 24676 4480 24728 4486
rect 24676 4422 24728 4428
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24688 4146 24716 4422
rect 24216 4140 24268 4146
rect 24676 4140 24728 4146
rect 24268 4100 24348 4128
rect 24216 4082 24268 4088
rect 24124 4004 24176 4010
rect 24124 3946 24176 3952
rect 24136 3466 24164 3946
rect 24216 3936 24268 3942
rect 24216 3878 24268 3884
rect 24124 3460 24176 3466
rect 24124 3402 24176 3408
rect 24228 3398 24256 3878
rect 24320 3602 24348 4100
rect 24676 4082 24728 4088
rect 24584 4072 24636 4078
rect 24584 4014 24636 4020
rect 24674 4040 24730 4049
rect 24398 3904 24454 3913
rect 24398 3839 24454 3848
rect 24412 3738 24440 3839
rect 24400 3732 24452 3738
rect 24400 3674 24452 3680
rect 24596 3641 24624 4014
rect 24674 3975 24730 3984
rect 24582 3632 24638 3641
rect 24308 3596 24360 3602
rect 24582 3567 24638 3576
rect 24308 3538 24360 3544
rect 24216 3392 24268 3398
rect 24216 3334 24268 3340
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24044 3182 24164 3210
rect 24030 3088 24086 3097
rect 24030 3023 24086 3032
rect 23938 1592 23994 1601
rect 23938 1527 23994 1536
rect 23846 912 23902 921
rect 23846 847 23902 856
rect 20902 96 20958 105
rect 20902 31 20958 40
rect 20994 0 21050 480
rect 21546 0 21602 480
rect 22098 0 22154 480
rect 22650 0 22706 480
rect 23202 0 23258 480
rect 23754 0 23810 480
rect 24044 377 24072 3023
rect 24136 2990 24164 3182
rect 24124 2984 24176 2990
rect 24124 2926 24176 2932
rect 24136 2582 24164 2926
rect 24490 2680 24546 2689
rect 24490 2615 24546 2624
rect 24504 2582 24532 2615
rect 24124 2576 24176 2582
rect 24124 2518 24176 2524
rect 24492 2576 24544 2582
rect 24492 2518 24544 2524
rect 24216 2508 24268 2514
rect 24216 2450 24268 2456
rect 24228 1057 24256 2450
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24688 1986 24716 3975
rect 24780 2650 24808 4950
rect 24860 4820 24912 4826
rect 24860 4762 24912 4768
rect 24872 4010 24900 4762
rect 24964 4078 24992 6990
rect 25044 6928 25096 6934
rect 25044 6870 25096 6876
rect 25056 6458 25084 6870
rect 25044 6452 25096 6458
rect 25044 6394 25096 6400
rect 25042 6216 25098 6225
rect 25042 6151 25044 6160
rect 25096 6151 25098 6160
rect 25044 6122 25096 6128
rect 25056 5914 25084 6122
rect 25044 5908 25096 5914
rect 25044 5850 25096 5856
rect 25056 4690 25084 5850
rect 25044 4684 25096 4690
rect 25044 4626 25096 4632
rect 25044 4480 25096 4486
rect 25044 4422 25096 4428
rect 24952 4072 25004 4078
rect 24952 4014 25004 4020
rect 24860 4004 24912 4010
rect 24860 3946 24912 3952
rect 24950 3768 25006 3777
rect 24950 3703 25006 3712
rect 24860 3528 24912 3534
rect 24860 3470 24912 3476
rect 24872 3194 24900 3470
rect 24860 3188 24912 3194
rect 24860 3130 24912 3136
rect 24872 2854 24900 3130
rect 24860 2848 24912 2854
rect 24860 2790 24912 2796
rect 24964 2666 24992 3703
rect 25056 3194 25084 4422
rect 25148 3738 25176 11886
rect 25320 11834 25372 11840
rect 25226 11792 25282 11801
rect 25226 11727 25282 11736
rect 25240 11694 25268 11727
rect 25228 11688 25280 11694
rect 25228 11630 25280 11636
rect 25226 11248 25282 11257
rect 25226 11183 25282 11192
rect 25240 8430 25268 11183
rect 25320 10260 25372 10266
rect 25320 10202 25372 10208
rect 25332 9382 25360 10202
rect 25320 9376 25372 9382
rect 25424 9353 25452 14894
rect 25516 12850 25544 16934
rect 25608 16046 25636 21111
rect 25700 16658 25728 21519
rect 25688 16652 25740 16658
rect 25688 16594 25740 16600
rect 25688 16448 25740 16454
rect 25688 16390 25740 16396
rect 25596 16040 25648 16046
rect 25596 15982 25648 15988
rect 25700 15366 25728 16390
rect 25688 15360 25740 15366
rect 25688 15302 25740 15308
rect 25700 14822 25728 15302
rect 25688 14816 25740 14822
rect 25688 14758 25740 14764
rect 25700 14074 25728 14758
rect 25688 14068 25740 14074
rect 25688 14010 25740 14016
rect 25596 13184 25648 13190
rect 25596 13126 25648 13132
rect 25504 12844 25556 12850
rect 25504 12786 25556 12792
rect 25608 12782 25636 13126
rect 25596 12776 25648 12782
rect 25596 12718 25648 12724
rect 25504 12096 25556 12102
rect 25504 12038 25556 12044
rect 25516 11558 25544 12038
rect 25504 11552 25556 11558
rect 25504 11494 25556 11500
rect 25686 11520 25742 11529
rect 25516 10470 25544 11494
rect 25686 11455 25742 11464
rect 25504 10464 25556 10470
rect 25504 10406 25556 10412
rect 25516 10266 25544 10406
rect 25504 10260 25556 10266
rect 25504 10202 25556 10208
rect 25596 10124 25648 10130
rect 25596 10066 25648 10072
rect 25608 9722 25636 10066
rect 25596 9716 25648 9722
rect 25596 9658 25648 9664
rect 25596 9580 25648 9586
rect 25596 9522 25648 9528
rect 25320 9318 25372 9324
rect 25410 9344 25466 9353
rect 25332 9178 25360 9318
rect 25410 9279 25466 9288
rect 25320 9172 25372 9178
rect 25320 9114 25372 9120
rect 25332 8945 25360 9114
rect 25318 8936 25374 8945
rect 25318 8871 25374 8880
rect 25228 8424 25280 8430
rect 25228 8366 25280 8372
rect 25412 8288 25464 8294
rect 25412 8230 25464 8236
rect 25228 7948 25280 7954
rect 25228 7890 25280 7896
rect 25240 6730 25268 7890
rect 25320 7744 25372 7750
rect 25320 7686 25372 7692
rect 25228 6724 25280 6730
rect 25228 6666 25280 6672
rect 25228 5160 25280 5166
rect 25226 5128 25228 5137
rect 25280 5128 25282 5137
rect 25226 5063 25282 5072
rect 25226 4176 25282 4185
rect 25226 4111 25282 4120
rect 25240 4078 25268 4111
rect 25228 4072 25280 4078
rect 25228 4014 25280 4020
rect 25136 3732 25188 3738
rect 25136 3674 25188 3680
rect 25044 3188 25096 3194
rect 25044 3130 25096 3136
rect 25044 2848 25096 2854
rect 25332 2836 25360 7686
rect 25424 4049 25452 8230
rect 25504 7744 25556 7750
rect 25504 7686 25556 7692
rect 25516 7342 25544 7686
rect 25504 7336 25556 7342
rect 25504 7278 25556 7284
rect 25516 5234 25544 7278
rect 25504 5228 25556 5234
rect 25504 5170 25556 5176
rect 25608 4826 25636 9522
rect 25596 4820 25648 4826
rect 25596 4762 25648 4768
rect 25410 4040 25466 4049
rect 25410 3975 25466 3984
rect 25412 3936 25464 3942
rect 25412 3878 25464 3884
rect 25424 3505 25452 3878
rect 25410 3496 25466 3505
rect 25410 3431 25466 3440
rect 25700 3398 25728 11455
rect 25792 11393 25820 24647
rect 26056 23860 26108 23866
rect 26056 23802 26108 23808
rect 25872 21344 25924 21350
rect 25872 21286 25924 21292
rect 25884 19378 25912 21286
rect 25964 20528 26016 20534
rect 25962 20496 25964 20505
rect 26016 20496 26018 20505
rect 25962 20431 26018 20440
rect 25872 19372 25924 19378
rect 25872 19314 25924 19320
rect 25964 19304 26016 19310
rect 25964 19246 26016 19252
rect 25870 19136 25926 19145
rect 25870 19071 25926 19080
rect 25884 13705 25912 19071
rect 25870 13696 25926 13705
rect 25870 13631 25926 13640
rect 25976 13433 26004 19246
rect 25962 13424 26018 13433
rect 25962 13359 26018 13368
rect 26068 12594 26096 23802
rect 26146 20768 26202 20777
rect 26146 20703 26202 20712
rect 26160 19514 26188 20703
rect 26252 20602 26280 24783
rect 27080 22409 27108 27520
rect 27632 26353 27660 27520
rect 27618 26344 27674 26353
rect 27618 26279 27674 26288
rect 27066 22400 27122 22409
rect 27066 22335 27122 22344
rect 26240 20596 26292 20602
rect 26240 20538 26292 20544
rect 26238 19816 26294 19825
rect 26238 19751 26294 19760
rect 26148 19508 26200 19514
rect 26148 19450 26200 19456
rect 26252 19310 26280 19751
rect 26332 19712 26384 19718
rect 26332 19654 26384 19660
rect 26240 19304 26292 19310
rect 26240 19246 26292 19252
rect 26148 18624 26200 18630
rect 26148 18566 26200 18572
rect 26160 17542 26188 18566
rect 26240 18080 26292 18086
rect 26238 18048 26240 18057
rect 26292 18048 26294 18057
rect 26238 17983 26294 17992
rect 26148 17536 26200 17542
rect 26148 17478 26200 17484
rect 26160 16998 26188 17478
rect 26148 16992 26200 16998
rect 26148 16934 26200 16940
rect 26160 16454 26188 16934
rect 26148 16448 26200 16454
rect 26148 16390 26200 16396
rect 26252 16182 26280 17983
rect 26344 17882 26372 19654
rect 26424 18148 26476 18154
rect 26424 18090 26476 18096
rect 26332 17876 26384 17882
rect 26332 17818 26384 17824
rect 26240 16176 26292 16182
rect 26240 16118 26292 16124
rect 26240 15904 26292 15910
rect 26240 15846 26292 15852
rect 26148 14612 26200 14618
rect 26252 14600 26280 15846
rect 26344 15706 26372 17818
rect 26332 15700 26384 15706
rect 26332 15642 26384 15648
rect 26344 15162 26372 15642
rect 26332 15156 26384 15162
rect 26332 15098 26384 15104
rect 26344 14618 26372 15098
rect 26200 14572 26280 14600
rect 26332 14612 26384 14618
rect 26148 14554 26200 14560
rect 26332 14554 26384 14560
rect 26344 14074 26372 14554
rect 26332 14068 26384 14074
rect 26332 14010 26384 14016
rect 26240 13932 26292 13938
rect 26240 13874 26292 13880
rect 26252 12986 26280 13874
rect 26344 13530 26372 14010
rect 26332 13524 26384 13530
rect 26332 13466 26384 13472
rect 26240 12980 26292 12986
rect 26240 12922 26292 12928
rect 25976 12566 26096 12594
rect 25778 11384 25834 11393
rect 25778 11319 25834 11328
rect 25976 11218 26004 12566
rect 26054 12472 26110 12481
rect 26344 12442 26372 13466
rect 26054 12407 26110 12416
rect 26332 12436 26384 12442
rect 25964 11212 26016 11218
rect 25964 11154 26016 11160
rect 25976 9586 26004 11154
rect 25964 9580 26016 9586
rect 25964 9522 26016 9528
rect 25780 9444 25832 9450
rect 25780 9386 25832 9392
rect 25792 5001 25820 9386
rect 25964 7200 26016 7206
rect 25964 7142 26016 7148
rect 25872 6724 25924 6730
rect 25872 6666 25924 6672
rect 25778 4992 25834 5001
rect 25778 4927 25834 4936
rect 25780 4684 25832 4690
rect 25780 4626 25832 4632
rect 25792 4282 25820 4626
rect 25780 4276 25832 4282
rect 25780 4218 25832 4224
rect 25884 4214 25912 6666
rect 25872 4208 25924 4214
rect 25872 4150 25924 4156
rect 25688 3392 25740 3398
rect 25688 3334 25740 3340
rect 25504 2916 25556 2922
rect 25504 2858 25556 2864
rect 25044 2790 25096 2796
rect 25240 2808 25360 2836
rect 24768 2644 24820 2650
rect 24768 2586 24820 2592
rect 24872 2638 24992 2666
rect 25056 2650 25084 2790
rect 25044 2644 25096 2650
rect 24320 1958 24716 1986
rect 24214 1048 24270 1057
rect 24214 983 24270 992
rect 24320 480 24348 1958
rect 24872 480 24900 2638
rect 25044 2586 25096 2592
rect 25056 2446 25084 2586
rect 25044 2440 25096 2446
rect 25044 2382 25096 2388
rect 25240 1578 25268 2808
rect 25516 1873 25544 2858
rect 25596 2576 25648 2582
rect 25594 2544 25596 2553
rect 25648 2544 25650 2553
rect 25594 2479 25650 2488
rect 25884 2009 25912 4150
rect 25870 2000 25926 2009
rect 25870 1935 25926 1944
rect 25502 1864 25558 1873
rect 25502 1799 25558 1808
rect 25240 1550 25452 1578
rect 25424 480 25452 1550
rect 25976 480 26004 7142
rect 26068 3194 26096 12407
rect 26332 12378 26384 12384
rect 26344 11354 26372 12378
rect 26332 11348 26384 11354
rect 26332 11290 26384 11296
rect 26436 10849 26464 18090
rect 26422 10840 26478 10849
rect 26422 10775 26478 10784
rect 26424 10260 26476 10266
rect 26424 10202 26476 10208
rect 26436 9654 26464 10202
rect 26424 9648 26476 9654
rect 26424 9590 26476 9596
rect 26436 9178 26464 9590
rect 26148 9172 26200 9178
rect 26148 9114 26200 9120
rect 26424 9172 26476 9178
rect 26424 9114 26476 9120
rect 26160 8634 26188 9114
rect 26148 8628 26200 8634
rect 26148 8570 26200 8576
rect 26160 8090 26188 8570
rect 26436 8090 26464 9114
rect 26148 8084 26200 8090
rect 26148 8026 26200 8032
rect 26424 8084 26476 8090
rect 26424 8026 26476 8032
rect 26160 7002 26188 8026
rect 26436 7546 26464 8026
rect 26424 7540 26476 7546
rect 26424 7482 26476 7488
rect 26148 6996 26200 7002
rect 26148 6938 26200 6944
rect 26160 6458 26188 6938
rect 26148 6452 26200 6458
rect 26148 6394 26200 6400
rect 26160 5914 26188 6394
rect 26148 5908 26200 5914
rect 26148 5850 26200 5856
rect 26160 5658 26188 5850
rect 26160 5630 26280 5658
rect 26252 5370 26280 5630
rect 26240 5364 26292 5370
rect 26240 5306 26292 5312
rect 26252 4826 26280 5306
rect 26240 4820 26292 4826
rect 26240 4762 26292 4768
rect 26332 4752 26384 4758
rect 26332 4694 26384 4700
rect 26240 4276 26292 4282
rect 26240 4218 26292 4224
rect 26252 3738 26280 4218
rect 26240 3732 26292 3738
rect 26240 3674 26292 3680
rect 26344 3194 26372 4694
rect 27618 3496 27674 3505
rect 27618 3431 27674 3440
rect 26056 3188 26108 3194
rect 26056 3130 26108 3136
rect 26332 3188 26384 3194
rect 26332 3130 26384 3136
rect 26068 2990 26096 3130
rect 26056 2984 26108 2990
rect 26056 2926 26108 2932
rect 26344 2650 26372 3130
rect 27066 2816 27122 2825
rect 27066 2751 27122 2760
rect 26332 2644 26384 2650
rect 26332 2586 26384 2592
rect 26514 1456 26570 1465
rect 26514 1391 26570 1400
rect 26528 480 26556 1391
rect 27080 480 27108 2751
rect 27632 480 27660 3431
rect 24030 368 24086 377
rect 24030 303 24086 312
rect 24306 0 24362 480
rect 24858 0 24914 480
rect 25410 0 25466 480
rect 25962 0 26018 480
rect 26514 0 26570 480
rect 27066 0 27122 480
rect 27618 0 27674 480
<< via2 >>
rect 1674 27648 1730 27704
rect 1490 27104 1546 27160
rect 1582 25880 1638 25936
rect 1582 24792 1638 24848
rect 846 23296 902 23352
rect 294 22752 350 22808
rect 1398 22752 1454 22808
rect 24674 27648 24730 27704
rect 1674 23196 1676 23216
rect 1676 23196 1728 23216
rect 1728 23196 1730 23216
rect 1674 23160 1730 23196
rect 1582 22480 1638 22536
rect 1398 20168 1454 20224
rect 1398 17584 1454 17640
rect 938 13096 994 13152
rect 1122 13640 1178 13696
rect 1490 16088 1546 16144
rect 2318 26560 2374 26616
rect 2042 24248 2098 24304
rect 1858 21392 1914 21448
rect 1674 20304 1730 20360
rect 2686 25336 2742 25392
rect 2226 22344 2282 22400
rect 2134 22072 2190 22128
rect 2410 22208 2466 22264
rect 2410 21140 2466 21176
rect 2410 21120 2412 21140
rect 2412 21120 2464 21140
rect 2464 21120 2466 21140
rect 2410 20984 2466 21040
rect 2318 19760 2374 19816
rect 2318 19352 2374 19408
rect 2134 18572 2136 18592
rect 2136 18572 2188 18592
rect 2188 18572 2190 18592
rect 2134 18536 2190 18572
rect 1766 16668 1768 16688
rect 1768 16668 1820 16688
rect 1820 16668 1822 16688
rect 1766 16632 1822 16668
rect 1398 14728 1454 14784
rect 1674 14592 1730 14648
rect 1950 15272 2006 15328
rect 1766 14048 1822 14104
rect 1398 11092 1400 11112
rect 1400 11092 1452 11112
rect 1452 11092 1454 11112
rect 1398 11056 1454 11092
rect 662 4528 718 4584
rect 1398 4256 1454 4312
rect 1858 13640 1914 13696
rect 2134 15136 2190 15192
rect 2042 13232 2098 13288
rect 2502 20032 2558 20088
rect 2778 23024 2834 23080
rect 3238 24112 3294 24168
rect 3514 23568 3570 23624
rect 3146 22516 3148 22536
rect 3148 22516 3200 22536
rect 3200 22516 3202 22536
rect 3146 22480 3202 22516
rect 3238 22208 3294 22264
rect 2962 21392 3018 21448
rect 3422 21528 3478 21584
rect 3514 19896 3570 19952
rect 2962 19216 3018 19272
rect 2686 15816 2742 15872
rect 2134 12688 2190 12744
rect 1950 12280 2006 12336
rect 1950 6840 2006 6896
rect 1858 4392 1914 4448
rect 1766 3732 1822 3768
rect 1766 3712 1768 3732
rect 1768 3712 1820 3732
rect 1820 3712 1822 3732
rect 1582 3168 1638 3224
rect 3422 19624 3478 19680
rect 3330 19488 3386 19544
rect 2870 15272 2926 15328
rect 2226 11464 2282 11520
rect 2594 10240 2650 10296
rect 2410 5344 2466 5400
rect 3146 15952 3202 16008
rect 2870 10920 2926 10976
rect 3882 21800 3938 21856
rect 3790 20032 3846 20088
rect 3790 19352 3846 19408
rect 4250 21528 4306 21584
rect 4066 21256 4122 21312
rect 4250 21020 4252 21040
rect 4252 21020 4304 21040
rect 4304 21020 4306 21040
rect 4250 20984 4306 21020
rect 4066 20440 4122 20496
rect 4066 19488 4122 19544
rect 4066 19352 4122 19408
rect 4066 18400 4122 18456
rect 3974 17992 4030 18048
rect 3974 17176 4030 17232
rect 3698 17040 3754 17096
rect 3514 16904 3570 16960
rect 3422 14592 3478 14648
rect 3146 13096 3202 13152
rect 3238 11600 3294 11656
rect 3054 10784 3110 10840
rect 2778 8880 2834 8936
rect 3514 13776 3570 13832
rect 3606 13504 3662 13560
rect 3422 11772 3424 11792
rect 3424 11772 3476 11792
rect 3476 11772 3478 11792
rect 3422 11736 3478 11772
rect 3238 8200 3294 8256
rect 3054 7384 3110 7440
rect 2778 6976 2834 7032
rect 3054 6024 3110 6080
rect 1858 3032 1914 3088
rect 1766 1400 1822 1456
rect 3054 3848 3110 3904
rect 2962 3712 3018 3768
rect 2870 3440 2926 3496
rect 2410 2624 2466 2680
rect 2318 2488 2374 2544
rect 1674 856 1730 912
rect 2410 2372 2466 2408
rect 2410 2352 2412 2372
rect 2412 2352 2464 2372
rect 2464 2352 2466 2372
rect 2870 1672 2926 1728
rect 2778 1264 2834 1320
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5538 24112 5594 24168
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5446 23568 5502 23624
rect 4158 17176 4214 17232
rect 4250 16768 4306 16824
rect 3790 12144 3846 12200
rect 3698 10376 3754 10432
rect 3698 8472 3754 8528
rect 4434 16768 4490 16824
rect 4342 13232 4398 13288
rect 5354 23432 5410 23488
rect 4986 22772 5042 22808
rect 4986 22752 4988 22772
rect 4988 22752 5040 22772
rect 5040 22752 5042 22772
rect 4802 21120 4858 21176
rect 4986 20848 5042 20904
rect 5078 19488 5134 19544
rect 4710 18164 4712 18184
rect 4712 18164 4764 18184
rect 4764 18164 4766 18184
rect 4710 18128 4766 18164
rect 4710 15952 4766 16008
rect 4250 12552 4306 12608
rect 4066 10648 4122 10704
rect 3882 9988 3938 10024
rect 3882 9968 3884 9988
rect 3884 9968 3936 9988
rect 3936 9968 3938 9988
rect 3974 8608 4030 8664
rect 3974 7792 4030 7848
rect 3974 7112 4030 7168
rect 3882 6296 3938 6352
rect 4526 10920 4582 10976
rect 4710 15680 4766 15736
rect 5906 23316 5962 23352
rect 5906 23296 5908 23316
rect 5908 23296 5960 23316
rect 5960 23296 5962 23316
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5538 22344 5594 22400
rect 5446 19660 5448 19680
rect 5448 19660 5500 19680
rect 5500 19660 5502 19680
rect 5446 19624 5502 19660
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5170 18672 5226 18728
rect 5262 18264 5318 18320
rect 5170 17720 5226 17776
rect 4986 16088 5042 16144
rect 4710 13948 4712 13968
rect 4712 13948 4764 13968
rect 4764 13948 4766 13968
rect 4710 13912 4766 13948
rect 5170 15816 5226 15872
rect 5078 14764 5080 14784
rect 5080 14764 5132 14784
rect 5132 14764 5134 14784
rect 5078 14728 5134 14764
rect 5262 15000 5318 15056
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5446 15544 5502 15600
rect 5446 15272 5502 15328
rect 5262 14048 5318 14104
rect 4802 11872 4858 11928
rect 4434 8356 4490 8392
rect 4434 8336 4436 8356
rect 4436 8336 4488 8356
rect 4488 8336 4490 8356
rect 5078 12552 5134 12608
rect 4894 10512 4950 10568
rect 3698 3984 3754 4040
rect 3698 1944 3754 2000
rect 4710 6160 4766 6216
rect 4618 5208 4674 5264
rect 3974 2916 4030 2952
rect 3974 2896 3976 2916
rect 3976 2896 4028 2916
rect 4028 2896 4030 2916
rect 4526 4392 4582 4448
rect 4434 2352 4490 2408
rect 4250 2216 4306 2272
rect 4986 5344 5042 5400
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5722 13640 5778 13696
rect 5538 13368 5594 13424
rect 5906 13232 5962 13288
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 6458 24384 6514 24440
rect 6182 22636 6238 22672
rect 6182 22616 6184 22636
rect 6184 22616 6236 22636
rect 6236 22616 6238 22636
rect 6366 21528 6422 21584
rect 6734 25064 6790 25120
rect 6642 23704 6698 23760
rect 7194 23840 7250 23896
rect 7654 25880 7710 25936
rect 7286 23296 7342 23352
rect 6550 22772 6606 22808
rect 6550 22752 6552 22772
rect 6552 22752 6604 22772
rect 6604 22752 6606 22772
rect 6550 20324 6606 20360
rect 6550 20304 6552 20324
rect 6552 20304 6604 20324
rect 6604 20304 6606 20324
rect 7194 23024 7250 23080
rect 7194 22616 7250 22672
rect 7378 22208 7434 22264
rect 7286 21936 7342 21992
rect 7470 21392 7526 21448
rect 7010 20476 7012 20496
rect 7012 20476 7064 20496
rect 7064 20476 7066 20496
rect 7010 20440 7066 20476
rect 6642 19488 6698 19544
rect 6550 19216 6606 19272
rect 6366 16904 6422 16960
rect 5906 12144 5962 12200
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5538 11192 5594 11248
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5722 10684 5724 10704
rect 5724 10684 5776 10704
rect 5776 10684 5778 10704
rect 5722 10648 5778 10684
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5630 9460 5632 9480
rect 5632 9460 5684 9480
rect 5684 9460 5686 9480
rect 5630 9424 5686 9460
rect 5630 8900 5686 8936
rect 5630 8880 5632 8900
rect 5632 8880 5684 8900
rect 5684 8880 5686 8900
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5538 8472 5594 8528
rect 5814 8084 5870 8120
rect 5814 8064 5816 8084
rect 5816 8064 5868 8084
rect 5868 8064 5870 8084
rect 5354 7828 5356 7848
rect 5356 7828 5408 7848
rect 5408 7828 5410 7848
rect 5354 7792 5410 7828
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5262 6432 5318 6488
rect 5262 6296 5318 6352
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 4802 3440 4858 3496
rect 5814 5636 5870 5672
rect 5814 5616 5816 5636
rect 5816 5616 5868 5636
rect 5868 5616 5870 5636
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5814 5108 5816 5128
rect 5816 5108 5868 5128
rect 5868 5108 5870 5128
rect 5814 5072 5870 5108
rect 6090 12688 6146 12744
rect 6366 13504 6422 13560
rect 6182 11872 6238 11928
rect 6182 11600 6238 11656
rect 6182 8744 6238 8800
rect 6090 6840 6146 6896
rect 5262 4256 5318 4312
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 6090 4120 6146 4176
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 6090 3168 6146 3224
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 6458 7928 6514 7984
rect 6366 7248 6422 7304
rect 6458 6704 6514 6760
rect 6458 6432 6514 6488
rect 6366 3304 6422 3360
rect 6366 3032 6422 3088
rect 7930 23024 7986 23080
rect 7562 20032 7618 20088
rect 7010 17740 7066 17776
rect 7010 17720 7012 17740
rect 7012 17720 7064 17740
rect 7064 17720 7066 17740
rect 7838 18536 7894 18592
rect 7194 17448 7250 17504
rect 6826 16360 6882 16416
rect 6826 16088 6882 16144
rect 6826 15272 6882 15328
rect 6826 15136 6882 15192
rect 7378 15952 7434 16008
rect 7286 15136 7342 15192
rect 7286 14728 7342 14784
rect 6826 14320 6882 14376
rect 6826 13640 6882 13696
rect 6642 13232 6698 13288
rect 6642 12708 6698 12744
rect 6642 12688 6644 12708
rect 6644 12688 6696 12708
rect 6696 12688 6698 12708
rect 6734 12008 6790 12064
rect 6550 2252 6552 2272
rect 6552 2252 6604 2272
rect 6604 2252 6606 2272
rect 6550 2216 6606 2252
rect 7378 13504 7434 13560
rect 7838 17856 7894 17912
rect 7654 15000 7710 15056
rect 7654 14048 7710 14104
rect 7286 11872 7342 11928
rect 6826 10412 6828 10432
rect 6828 10412 6880 10432
rect 6880 10412 6882 10432
rect 6826 10376 6882 10412
rect 6826 10240 6882 10296
rect 7194 9988 7250 10024
rect 7194 9968 7196 9988
rect 7196 9968 7248 9988
rect 7248 9968 7250 9988
rect 7102 9016 7158 9072
rect 6826 8608 6882 8664
rect 6826 2080 6882 2136
rect 7286 8336 7342 8392
rect 7286 7148 7288 7168
rect 7288 7148 7340 7168
rect 7340 7148 7342 7168
rect 7286 7112 7342 7148
rect 8482 22888 8538 22944
rect 8390 20848 8446 20904
rect 8022 19236 8078 19272
rect 8022 19216 8024 19236
rect 8024 19216 8076 19236
rect 8076 19216 8078 19236
rect 8666 24828 8668 24848
rect 8668 24828 8720 24848
rect 8720 24828 8722 24848
rect 8666 24792 8722 24828
rect 8666 21528 8722 21584
rect 8574 21392 8630 21448
rect 8022 17332 8078 17368
rect 8022 17312 8024 17332
rect 8024 17312 8076 17332
rect 8076 17312 8078 17332
rect 8390 16768 8446 16824
rect 8298 16652 8354 16688
rect 8298 16632 8300 16652
rect 8300 16632 8352 16652
rect 8352 16632 8354 16652
rect 8114 15680 8170 15736
rect 8298 15580 8300 15600
rect 8300 15580 8352 15600
rect 8352 15580 8354 15600
rect 8298 15544 8354 15580
rect 7930 13776 7986 13832
rect 7654 10004 7656 10024
rect 7656 10004 7708 10024
rect 7708 10004 7710 10024
rect 7654 9968 7710 10004
rect 7470 9696 7526 9752
rect 7378 5344 7434 5400
rect 7378 5072 7434 5128
rect 7470 4936 7526 4992
rect 7194 1944 7250 2000
rect 7470 4392 7526 4448
rect 7470 2624 7526 2680
rect 7654 8200 7710 8256
rect 7838 9696 7894 9752
rect 8482 14456 8538 14512
rect 8482 13776 8538 13832
rect 8114 12824 8170 12880
rect 8298 12724 8300 12744
rect 8300 12724 8352 12744
rect 8352 12724 8354 12744
rect 8298 12688 8354 12724
rect 8206 11736 8262 11792
rect 8206 11500 8208 11520
rect 8208 11500 8260 11520
rect 8260 11500 8262 11520
rect 8206 11464 8262 11500
rect 8298 10240 8354 10296
rect 8022 4972 8024 4992
rect 8024 4972 8076 4992
rect 8076 4972 8078 4992
rect 8022 4936 8078 4972
rect 8482 12688 8538 12744
rect 8850 20576 8906 20632
rect 8666 19352 8722 19408
rect 9954 26016 10010 26072
rect 9310 23704 9366 23760
rect 9034 21528 9090 21584
rect 9034 20884 9036 20904
rect 9036 20884 9088 20904
rect 9088 20884 9090 20904
rect 9034 20848 9090 20884
rect 9034 20304 9090 20360
rect 8758 15272 8814 15328
rect 8666 12552 8722 12608
rect 8666 8744 8722 8800
rect 8574 7248 8630 7304
rect 8390 5616 8446 5672
rect 8298 5072 8354 5128
rect 8482 4936 8538 4992
rect 8482 4528 8538 4584
rect 8666 4528 8722 4584
rect 9126 18028 9128 18048
rect 9128 18028 9180 18048
rect 9180 18028 9182 18048
rect 9126 17992 9182 18028
rect 9402 21800 9458 21856
rect 9678 24384 9734 24440
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10230 25200 10286 25256
rect 9862 23432 9918 23488
rect 9770 22480 9826 22536
rect 9310 18400 9366 18456
rect 9310 17604 9366 17640
rect 9310 17584 9312 17604
rect 9312 17584 9364 17604
rect 9364 17584 9366 17604
rect 9218 17040 9274 17096
rect 9310 16768 9366 16824
rect 9218 16224 9274 16280
rect 9126 15952 9182 16008
rect 8942 15816 8998 15872
rect 8942 14048 8998 14104
rect 8942 13932 8998 13968
rect 8942 13912 8944 13932
rect 8944 13912 8996 13932
rect 8996 13912 8998 13932
rect 9126 15036 9128 15056
rect 9128 15036 9180 15056
rect 9180 15036 9182 15056
rect 9126 15000 9182 15036
rect 9034 12552 9090 12608
rect 9218 13640 9274 13696
rect 9494 19760 9550 19816
rect 9954 21936 10010 21992
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10874 25336 10930 25392
rect 10874 25064 10930 25120
rect 10782 24248 10838 24304
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10506 22500 10562 22536
rect 10506 22480 10508 22500
rect 10508 22480 10560 22500
rect 10560 22480 10562 22500
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10598 22072 10654 22128
rect 10690 21392 10746 21448
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 9862 20168 9918 20224
rect 9494 16632 9550 16688
rect 9678 16496 9734 16552
rect 9678 16360 9734 16416
rect 9954 20032 10010 20088
rect 11150 24692 11152 24712
rect 11152 24692 11204 24712
rect 11204 24692 11206 24712
rect 11150 24656 11206 24692
rect 11242 24556 11244 24576
rect 11244 24556 11296 24576
rect 11296 24556 11298 24576
rect 11242 24520 11298 24556
rect 11242 24384 11298 24440
rect 11242 23704 11298 23760
rect 11058 23604 11060 23624
rect 11060 23604 11112 23624
rect 11112 23604 11114 23624
rect 11058 23568 11114 23604
rect 10966 23296 11022 23352
rect 11150 21936 11206 21992
rect 11058 21664 11114 21720
rect 10874 20712 10930 20768
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10414 19216 10470 19272
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 9678 14320 9734 14376
rect 9586 13096 9642 13152
rect 9034 10240 9090 10296
rect 9218 10376 9274 10432
rect 9126 9832 9182 9888
rect 8942 9460 8944 9480
rect 8944 9460 8996 9480
rect 8996 9460 8998 9480
rect 8942 9424 8998 9460
rect 8850 8372 8852 8392
rect 8852 8372 8904 8392
rect 8904 8372 8906 8392
rect 8850 8336 8906 8372
rect 8850 7792 8906 7848
rect 8942 4256 8998 4312
rect 8298 3576 8354 3632
rect 7930 3168 7986 3224
rect 7562 1536 7618 1592
rect 7746 1400 7802 1456
rect 8666 3440 8722 3496
rect 8390 2488 8446 2544
rect 9126 8200 9182 8256
rect 10782 20168 10838 20224
rect 10782 18808 10838 18864
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10138 17720 10194 17776
rect 10414 17212 10416 17232
rect 10416 17212 10468 17232
rect 10468 17212 10470 17232
rect 10414 17176 10470 17212
rect 11058 21120 11114 21176
rect 11058 20868 11114 20904
rect 11058 20848 11060 20868
rect 11060 20848 11112 20868
rect 11112 20848 11114 20868
rect 11242 21120 11298 21176
rect 11242 20032 11298 20088
rect 11058 19488 11114 19544
rect 10874 17856 10930 17912
rect 11150 18536 11206 18592
rect 11150 17992 11206 18048
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10690 16788 10746 16824
rect 10690 16768 10692 16788
rect 10692 16768 10744 16788
rect 10744 16768 10746 16788
rect 10046 14184 10102 14240
rect 9862 12316 9864 12336
rect 9864 12316 9916 12336
rect 9916 12316 9918 12336
rect 9862 12280 9918 12316
rect 9678 11872 9734 11928
rect 9678 11328 9734 11384
rect 9586 10240 9642 10296
rect 9310 8608 9366 8664
rect 9126 3884 9128 3904
rect 9128 3884 9180 3904
rect 9180 3884 9182 3904
rect 9126 3848 9182 3884
rect 9218 3068 9220 3088
rect 9220 3068 9272 3088
rect 9272 3068 9274 3088
rect 9218 3032 9274 3068
rect 9586 9832 9642 9888
rect 9678 8900 9734 8936
rect 9678 8880 9680 8900
rect 9680 8880 9732 8900
rect 9732 8880 9734 8900
rect 9770 8608 9826 8664
rect 9770 8064 9826 8120
rect 9678 5752 9734 5808
rect 9494 5092 9550 5128
rect 9770 5208 9826 5264
rect 9494 5072 9496 5092
rect 9496 5072 9548 5092
rect 9548 5072 9550 5092
rect 9678 4936 9734 4992
rect 9954 10512 10010 10568
rect 10690 15852 10692 15872
rect 10692 15852 10744 15872
rect 10744 15852 10746 15872
rect 10690 15816 10746 15852
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10046 8608 10102 8664
rect 10046 6296 10102 6352
rect 10046 5616 10102 5672
rect 9586 3712 9642 3768
rect 9862 4120 9918 4176
rect 9954 3732 10010 3768
rect 9954 3712 9956 3732
rect 9956 3712 10008 3732
rect 10008 3712 10010 3732
rect 9678 2896 9734 2952
rect 9310 2488 9366 2544
rect 9310 1672 9366 1728
rect 10322 11600 10378 11656
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10966 12960 11022 13016
rect 10230 10784 10286 10840
rect 10782 11192 10838 11248
rect 10598 11056 10654 11112
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10782 10240 10838 10296
rect 10322 9424 10378 9480
rect 10690 9324 10692 9344
rect 10692 9324 10744 9344
rect 10744 9324 10746 9344
rect 10690 9288 10746 9324
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10598 8356 10654 8392
rect 10598 8336 10600 8356
rect 10600 8336 10652 8356
rect 10652 8336 10654 8356
rect 10690 8200 10746 8256
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10690 6568 10746 6624
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10690 5752 10746 5808
rect 11518 25880 11574 25936
rect 11426 22772 11482 22808
rect 11426 22752 11428 22772
rect 11428 22752 11480 22772
rect 11480 22752 11482 22772
rect 11426 21664 11482 21720
rect 11426 21392 11482 21448
rect 11518 19488 11574 19544
rect 11518 18672 11574 18728
rect 11426 17856 11482 17912
rect 11334 16768 11390 16824
rect 12254 23976 12310 24032
rect 11702 21256 11758 21312
rect 12438 23976 12494 24032
rect 12438 23704 12494 23760
rect 12162 22616 12218 22672
rect 12162 22480 12218 22536
rect 12346 21392 12402 21448
rect 11886 19116 11888 19136
rect 11888 19116 11940 19136
rect 11940 19116 11942 19136
rect 11886 19080 11942 19116
rect 11702 18536 11758 18592
rect 11702 18264 11758 18320
rect 11426 16088 11482 16144
rect 11610 16088 11666 16144
rect 11518 14048 11574 14104
rect 11334 13776 11390 13832
rect 11426 13368 11482 13424
rect 11058 11620 11114 11656
rect 11058 11600 11060 11620
rect 11060 11600 11112 11620
rect 11112 11600 11114 11620
rect 11426 12144 11482 12200
rect 11794 14456 11850 14512
rect 11702 13232 11758 13288
rect 11702 12980 11758 13016
rect 11702 12960 11704 12980
rect 11704 12960 11756 12980
rect 11756 12960 11758 12980
rect 11702 12416 11758 12472
rect 11610 10648 11666 10704
rect 11058 7928 11114 7984
rect 10690 4936 10746 4992
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10138 3168 10194 3224
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 10138 2624 10194 2680
rect 10782 2624 10838 2680
rect 11242 5480 11298 5536
rect 11518 5908 11574 5944
rect 11518 5888 11520 5908
rect 11520 5888 11572 5908
rect 11572 5888 11574 5908
rect 11426 4936 11482 4992
rect 11334 4684 11390 4720
rect 11334 4664 11336 4684
rect 11336 4664 11388 4684
rect 11388 4664 11390 4684
rect 12162 20884 12164 20904
rect 12164 20884 12216 20904
rect 12216 20884 12218 20904
rect 12162 20848 12218 20884
rect 12438 20984 12494 21040
rect 12438 20596 12494 20632
rect 12438 20576 12440 20596
rect 12440 20576 12492 20596
rect 12492 20576 12494 20596
rect 12438 18672 12494 18728
rect 12254 17312 12310 17368
rect 12898 24656 12954 24712
rect 12714 23976 12770 24032
rect 13634 24812 13690 24848
rect 13634 24792 13636 24812
rect 13636 24792 13688 24812
rect 13688 24792 13690 24812
rect 12622 21936 12678 21992
rect 12438 17040 12494 17096
rect 12346 15816 12402 15872
rect 12530 14864 12586 14920
rect 12438 14184 12494 14240
rect 12162 13640 12218 13696
rect 11886 12180 11888 12200
rect 11888 12180 11940 12200
rect 11940 12180 11942 12200
rect 11886 12144 11942 12180
rect 11978 11736 12034 11792
rect 11794 8628 11850 8664
rect 11794 8608 11796 8628
rect 11796 8608 11848 8628
rect 11848 8608 11850 8628
rect 12530 13640 12586 13696
rect 12990 22208 13046 22264
rect 12714 21528 12770 21584
rect 12806 20848 12862 20904
rect 12806 20168 12862 20224
rect 12806 18808 12862 18864
rect 12990 20168 13046 20224
rect 12806 17584 12862 17640
rect 12806 17312 12862 17368
rect 12990 17856 13046 17912
rect 12622 13096 12678 13152
rect 12806 15308 12808 15328
rect 12808 15308 12860 15328
rect 12860 15308 12862 15328
rect 12806 15272 12862 15308
rect 12990 14864 13046 14920
rect 12898 13912 12954 13968
rect 12714 12960 12770 13016
rect 12254 10920 12310 10976
rect 11978 8608 12034 8664
rect 11886 6160 11942 6216
rect 11426 3884 11428 3904
rect 11428 3884 11480 3904
rect 11480 3884 11482 3904
rect 11426 3848 11482 3884
rect 11886 4528 11942 4584
rect 11886 4256 11942 4312
rect 11610 3984 11666 4040
rect 11058 3188 11114 3224
rect 11058 3168 11060 3188
rect 11060 3168 11112 3188
rect 11112 3168 11114 3188
rect 10966 2352 11022 2408
rect 12622 12552 12678 12608
rect 12714 10240 12770 10296
rect 12254 9152 12310 9208
rect 12714 9560 12770 9616
rect 12530 8472 12586 8528
rect 12162 7420 12164 7440
rect 12164 7420 12216 7440
rect 12216 7420 12218 7440
rect 12162 7384 12218 7420
rect 12346 7540 12402 7576
rect 12346 7520 12348 7540
rect 12348 7520 12400 7540
rect 12400 7520 12402 7540
rect 12438 7284 12440 7304
rect 12440 7284 12492 7304
rect 12492 7284 12494 7304
rect 12438 7248 12494 7284
rect 12438 5072 12494 5128
rect 12070 3576 12126 3632
rect 13542 24284 13544 24304
rect 13544 24284 13596 24304
rect 13596 24284 13598 24304
rect 13542 24248 13598 24284
rect 13450 24112 13506 24168
rect 13634 23316 13690 23352
rect 13634 23296 13636 23316
rect 13636 23296 13688 23316
rect 13688 23296 13690 23316
rect 13450 22072 13506 22128
rect 13358 19352 13414 19408
rect 13358 18420 13414 18456
rect 13358 18400 13360 18420
rect 13360 18400 13412 18420
rect 13412 18400 13414 18420
rect 13266 13912 13322 13968
rect 13358 13776 13414 13832
rect 13266 12688 13322 12744
rect 13174 8880 13230 8936
rect 13726 22208 13782 22264
rect 13634 22072 13690 22128
rect 14738 24928 14794 24984
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14094 23840 14150 23896
rect 14278 23840 14334 23896
rect 13634 20440 13690 20496
rect 14002 21800 14058 21856
rect 13910 20304 13966 20360
rect 13542 19916 13598 19952
rect 13542 19896 13544 19916
rect 13544 19896 13596 19916
rect 13596 19896 13598 19916
rect 13542 19216 13598 19272
rect 13818 18944 13874 19000
rect 13634 17604 13690 17640
rect 13634 17584 13636 17604
rect 13636 17584 13688 17604
rect 13688 17584 13690 17604
rect 13634 17312 13690 17368
rect 13634 16904 13690 16960
rect 13818 15988 13820 16008
rect 13820 15988 13872 16008
rect 13872 15988 13874 16008
rect 13818 15952 13874 15988
rect 14186 20440 14242 20496
rect 14186 19624 14242 19680
rect 14186 17448 14242 17504
rect 14186 17040 14242 17096
rect 14094 16360 14150 16416
rect 13542 14864 13598 14920
rect 13542 12552 13598 12608
rect 13450 10804 13506 10840
rect 13450 10784 13452 10804
rect 13452 10784 13504 10804
rect 13504 10784 13506 10804
rect 13358 10104 13414 10160
rect 13358 9424 13414 9480
rect 13450 7112 13506 7168
rect 13358 5752 13414 5808
rect 12806 3732 12862 3768
rect 12806 3712 12808 3732
rect 12808 3712 12860 3732
rect 12860 3712 12862 3732
rect 12622 2488 12678 2544
rect 12070 2388 12072 2408
rect 12072 2388 12124 2408
rect 12124 2388 12126 2408
rect 12070 2352 12126 2388
rect 12714 2352 12770 2408
rect 13266 3440 13322 3496
rect 13082 2216 13138 2272
rect 12990 1400 13046 1456
rect 14186 16088 14242 16144
rect 14094 14764 14096 14784
rect 14096 14764 14148 14784
rect 14148 14764 14150 14784
rect 14094 14728 14150 14764
rect 13910 13796 13966 13832
rect 13910 13776 13912 13796
rect 13912 13776 13964 13796
rect 13964 13776 13966 13796
rect 13726 12008 13782 12064
rect 13634 11736 13690 11792
rect 13910 12552 13966 12608
rect 13910 12416 13966 12472
rect 14646 24520 14702 24576
rect 14554 23704 14610 23760
rect 15106 24792 15162 24848
rect 14554 22924 14556 22944
rect 14556 22924 14608 22944
rect 14608 22924 14610 22944
rect 14554 22888 14610 22924
rect 14738 23704 14794 23760
rect 14554 22344 14610 22400
rect 14462 20440 14518 20496
rect 14370 16632 14426 16688
rect 14370 16496 14426 16552
rect 14278 14320 14334 14376
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 15106 23568 15162 23624
rect 15290 23432 15346 23488
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 15566 23296 15622 23352
rect 14094 12688 14150 12744
rect 14094 12552 14150 12608
rect 14002 11228 14004 11248
rect 14004 11228 14056 11248
rect 14056 11228 14058 11248
rect 14002 11192 14058 11228
rect 14186 11192 14242 11248
rect 13726 10376 13782 10432
rect 13726 9832 13782 9888
rect 13910 9832 13966 9888
rect 13818 9716 13874 9752
rect 13818 9696 13820 9716
rect 13820 9696 13872 9716
rect 13872 9696 13874 9716
rect 13910 8372 13912 8392
rect 13912 8372 13964 8392
rect 13964 8372 13966 8392
rect 13910 8336 13966 8372
rect 13910 7948 13966 7984
rect 13910 7928 13912 7948
rect 13912 7928 13964 7948
rect 13964 7928 13966 7948
rect 13818 5480 13874 5536
rect 13910 5208 13966 5264
rect 14738 13368 14794 13424
rect 14646 10140 14648 10160
rect 14648 10140 14700 10160
rect 14700 10140 14702 10160
rect 14646 10104 14702 10140
rect 14094 4528 14150 4584
rect 14002 3984 14058 4040
rect 14094 3848 14150 3904
rect 13450 3168 13506 3224
rect 14002 3168 14058 3224
rect 13450 3032 13506 3088
rect 13910 2896 13966 2952
rect 13450 1128 13506 1184
rect 14002 1672 14058 1728
rect 3146 312 3202 368
rect 14370 8064 14426 8120
rect 14278 7248 14334 7304
rect 14462 7404 14518 7440
rect 14462 7384 14464 7404
rect 14464 7384 14516 7404
rect 14516 7384 14518 7404
rect 14738 8744 14794 8800
rect 14738 8608 14794 8664
rect 14738 7792 14794 7848
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 15566 22616 15622 22672
rect 15566 20576 15622 20632
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 15106 19216 15162 19272
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 15290 17876 15346 17912
rect 15290 17856 15292 17876
rect 15292 17856 15344 17876
rect 15344 17856 15346 17876
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 15198 17176 15254 17232
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 15382 16088 15438 16144
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 15290 14728 15346 14784
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 15198 13776 15254 13832
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 16946 25336 17002 25392
rect 16026 24792 16082 24848
rect 15842 22480 15898 22536
rect 15750 18536 15806 18592
rect 15658 18128 15714 18184
rect 15566 13504 15622 13560
rect 16578 24792 16634 24848
rect 16394 23468 16396 23488
rect 16396 23468 16448 23488
rect 16448 23468 16450 23488
rect 16394 23432 16450 23468
rect 16394 23160 16450 23216
rect 16394 21664 16450 21720
rect 16026 17176 16082 17232
rect 15934 16224 15990 16280
rect 15290 12688 15346 12744
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 15014 9444 15070 9480
rect 15014 9424 15016 9444
rect 15016 9424 15068 9444
rect 15068 9424 15070 9444
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 15014 8492 15070 8528
rect 15014 8472 15016 8492
rect 15016 8472 15068 8492
rect 15068 8472 15070 8492
rect 14922 7928 14978 7984
rect 15382 8880 15438 8936
rect 15290 8084 15346 8120
rect 15290 8064 15292 8084
rect 15292 8064 15344 8084
rect 15344 8064 15346 8084
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14738 6160 14794 6216
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 15198 6024 15254 6080
rect 15566 11328 15622 11384
rect 15566 9968 15622 10024
rect 15658 9832 15714 9888
rect 15658 6976 15714 7032
rect 15474 6740 15476 6760
rect 15476 6740 15528 6760
rect 15528 6740 15530 6760
rect 15474 6704 15530 6740
rect 15382 6024 15438 6080
rect 14278 2372 14334 2408
rect 14278 2352 14280 2372
rect 14280 2352 14332 2372
rect 14332 2352 14334 2372
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 15658 5908 15714 5944
rect 15658 5888 15660 5908
rect 15660 5888 15712 5908
rect 15712 5888 15714 5908
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14830 3984 14886 4040
rect 14738 3884 14740 3904
rect 14740 3884 14792 3904
rect 14792 3884 14794 3904
rect 14738 3848 14794 3884
rect 14646 2624 14702 2680
rect 14462 2488 14518 2544
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 15566 5480 15622 5536
rect 15658 5208 15714 5264
rect 15658 4392 15714 4448
rect 16026 15272 16082 15328
rect 15934 13096 15990 13152
rect 15934 12280 15990 12336
rect 15934 9696 15990 9752
rect 15842 9560 15898 9616
rect 15934 9288 15990 9344
rect 15934 9016 15990 9072
rect 15842 8744 15898 8800
rect 15934 8608 15990 8664
rect 15842 8200 15898 8256
rect 16210 21256 16266 21312
rect 16762 23316 16818 23352
rect 16762 23296 16764 23316
rect 16764 23296 16816 23316
rect 16816 23296 16818 23316
rect 17314 25336 17370 25392
rect 17038 22888 17094 22944
rect 17038 22480 17094 22536
rect 16670 19080 16726 19136
rect 16946 21800 17002 21856
rect 16946 20712 17002 20768
rect 16486 17448 16542 17504
rect 16394 15408 16450 15464
rect 16302 15272 16358 15328
rect 16302 13776 16358 13832
rect 16210 12844 16266 12880
rect 16210 12824 16212 12844
rect 16212 12824 16264 12844
rect 16264 12824 16266 12844
rect 16394 11892 16450 11928
rect 16394 11872 16396 11892
rect 16396 11872 16448 11892
rect 16448 11872 16450 11892
rect 16670 17992 16726 18048
rect 16854 18300 16856 18320
rect 16856 18300 16908 18320
rect 16908 18300 16910 18320
rect 16854 18264 16910 18300
rect 16670 17312 16726 17368
rect 17038 16652 17094 16688
rect 17038 16632 17040 16652
rect 17040 16632 17092 16652
rect 17092 16632 17094 16652
rect 16854 14320 16910 14376
rect 16854 13812 16856 13832
rect 16856 13812 16908 13832
rect 16908 13812 16910 13832
rect 16854 13776 16910 13812
rect 16762 12416 16818 12472
rect 16394 10804 16450 10840
rect 16394 10784 16396 10804
rect 16396 10784 16448 10804
rect 16448 10784 16450 10804
rect 16210 10412 16212 10432
rect 16212 10412 16264 10432
rect 16264 10412 16266 10432
rect 16210 10376 16266 10412
rect 16210 9696 16266 9752
rect 16302 9288 16358 9344
rect 16302 8472 16358 8528
rect 16670 11736 16726 11792
rect 17038 13776 17094 13832
rect 16946 12144 17002 12200
rect 16486 9560 16542 9616
rect 16486 9016 16542 9072
rect 17038 11056 17094 11112
rect 16946 9968 17002 10024
rect 16026 5636 16082 5672
rect 16026 5616 16028 5636
rect 16028 5616 16080 5636
rect 16080 5616 16082 5636
rect 16026 5344 16082 5400
rect 15934 4936 15990 4992
rect 15566 2760 15622 2816
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 16394 7792 16450 7848
rect 16578 7656 16634 7712
rect 16578 6840 16634 6896
rect 16854 9832 16910 9888
rect 16854 8880 16910 8936
rect 16394 4936 16450 4992
rect 16854 6568 16910 6624
rect 16762 4664 16818 4720
rect 16670 4528 16726 4584
rect 16762 3712 16818 3768
rect 17314 24384 17370 24440
rect 18510 25064 18566 25120
rect 18418 24928 18474 24984
rect 17774 24248 17830 24304
rect 17406 23296 17462 23352
rect 17222 22092 17278 22128
rect 17222 22072 17224 22092
rect 17224 22072 17276 22092
rect 17276 22072 17278 22092
rect 17222 18808 17278 18864
rect 17222 15272 17278 15328
rect 17222 13912 17278 13968
rect 17498 21120 17554 21176
rect 17498 19896 17554 19952
rect 17406 19352 17462 19408
rect 17498 18148 17554 18184
rect 17498 18128 17500 18148
rect 17500 18128 17552 18148
rect 17552 18128 17554 18148
rect 17406 17720 17462 17776
rect 17774 22380 17776 22400
rect 17776 22380 17828 22400
rect 17828 22380 17830 22400
rect 17774 22344 17830 22380
rect 18234 22344 18290 22400
rect 18050 20984 18106 21040
rect 18050 20596 18106 20632
rect 18050 20576 18052 20596
rect 18052 20576 18104 20596
rect 18104 20576 18106 20596
rect 17774 19760 17830 19816
rect 17682 15408 17738 15464
rect 17682 14456 17738 14512
rect 17498 12980 17554 13016
rect 17498 12960 17500 12980
rect 17500 12960 17552 12980
rect 17552 12960 17554 12980
rect 17498 12688 17554 12744
rect 17222 11464 17278 11520
rect 17406 9696 17462 9752
rect 17222 7792 17278 7848
rect 17682 10920 17738 10976
rect 17682 9152 17738 9208
rect 17682 8472 17738 8528
rect 18326 19352 18382 19408
rect 18602 24928 18658 24984
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19798 24692 19800 24712
rect 19800 24692 19852 24712
rect 19852 24692 19854 24712
rect 19798 24656 19854 24692
rect 18602 24520 18658 24576
rect 18694 23704 18750 23760
rect 18878 23296 18934 23352
rect 18602 21664 18658 21720
rect 18510 21392 18566 21448
rect 18602 21256 18658 21312
rect 18510 19488 18566 19544
rect 18602 19216 18658 19272
rect 18602 18944 18658 19000
rect 18510 18400 18566 18456
rect 18050 15000 18106 15056
rect 18234 13388 18290 13424
rect 18234 13368 18236 13388
rect 18236 13368 18288 13388
rect 18288 13368 18290 13388
rect 17866 13096 17922 13152
rect 18050 13096 18106 13152
rect 17866 12824 17922 12880
rect 17498 5652 17500 5672
rect 17500 5652 17552 5672
rect 17552 5652 17554 5672
rect 17498 5616 17554 5652
rect 17314 3712 17370 3768
rect 17774 6452 17830 6488
rect 17774 6432 17776 6452
rect 17776 6432 17828 6452
rect 17828 6432 17830 6452
rect 17682 6296 17738 6352
rect 17866 6296 17922 6352
rect 18418 15952 18474 16008
rect 18326 12280 18382 12336
rect 17590 4528 17646 4584
rect 18234 9288 18290 9344
rect 18326 7964 18328 7984
rect 18328 7964 18380 7984
rect 18380 7964 18382 7984
rect 18326 7928 18382 7964
rect 18786 21936 18842 21992
rect 18694 11056 18750 11112
rect 18234 5908 18290 5944
rect 18234 5888 18236 5908
rect 18236 5888 18288 5908
rect 18288 5888 18290 5908
rect 18142 5616 18198 5672
rect 17866 4548 17922 4584
rect 17866 4528 17868 4548
rect 17868 4528 17920 4548
rect 17920 4528 17922 4548
rect 18050 3440 18106 3496
rect 18418 4664 18474 4720
rect 18326 4528 18382 4584
rect 18234 4120 18290 4176
rect 18418 3848 18474 3904
rect 18142 3032 18198 3088
rect 17774 2932 17776 2952
rect 17776 2932 17828 2952
rect 17828 2932 17830 2952
rect 17774 2896 17830 2932
rect 18326 2644 18382 2680
rect 18326 2624 18328 2644
rect 18328 2624 18380 2644
rect 18380 2624 18382 2644
rect 18234 2488 18290 2544
rect 18418 2488 18474 2544
rect 16762 2216 16818 2272
rect 16946 2252 16948 2272
rect 16948 2252 17000 2272
rect 17000 2252 17002 2272
rect 16946 2216 17002 2252
rect 16670 2080 16726 2136
rect 16762 1536 16818 1592
rect 18234 1944 18290 2000
rect 18418 1944 18474 2000
rect 17682 1808 17738 1864
rect 17590 1264 17646 1320
rect 18694 8608 18750 8664
rect 18970 22208 19026 22264
rect 18970 21664 19026 21720
rect 19062 21120 19118 21176
rect 19062 20848 19118 20904
rect 18970 20168 19026 20224
rect 18970 17196 19026 17232
rect 18970 17176 18972 17196
rect 18972 17176 19024 17196
rect 19024 17176 19026 17196
rect 19062 16360 19118 16416
rect 18970 11872 19026 11928
rect 18970 11736 19026 11792
rect 18878 11464 18934 11520
rect 18878 11056 18934 11112
rect 19246 23160 19302 23216
rect 19246 22380 19248 22400
rect 19248 22380 19300 22400
rect 19300 22380 19302 22400
rect 19246 22344 19302 22380
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 20626 26016 20682 26072
rect 21362 25200 21418 25256
rect 21270 25064 21326 25120
rect 21178 24812 21234 24848
rect 21178 24792 21180 24812
rect 21180 24792 21232 24812
rect 21232 24792 21234 24812
rect 20718 24556 20720 24576
rect 20720 24556 20772 24576
rect 20772 24556 20774 24576
rect 19982 24248 20038 24304
rect 19430 23468 19432 23488
rect 19432 23468 19484 23488
rect 19484 23468 19486 23488
rect 19430 23432 19486 23468
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19614 22888 19670 22944
rect 20166 23568 20222 23624
rect 20074 23432 20130 23488
rect 20442 23840 20498 23896
rect 20350 23296 20406 23352
rect 20166 22752 20222 22808
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19522 21392 19578 21448
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19614 20748 19616 20768
rect 19616 20748 19668 20768
rect 19668 20748 19670 20768
rect 19614 20712 19670 20748
rect 20074 21256 20130 21312
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19982 19896 20038 19952
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19430 17856 19486 17912
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19430 16768 19486 16824
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 20166 19080 20222 19136
rect 20166 18536 20222 18592
rect 20166 17312 20222 17368
rect 19982 15952 20038 16008
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19246 14048 19302 14104
rect 19154 11736 19210 11792
rect 19338 13096 19394 13152
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 20074 15272 20130 15328
rect 20166 15136 20222 15192
rect 20074 14592 20130 14648
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19522 12960 19578 13016
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19246 11600 19302 11656
rect 19246 10920 19302 10976
rect 18878 9968 18934 10024
rect 18694 5888 18750 5944
rect 18970 5752 19026 5808
rect 18694 3304 18750 3360
rect 18970 3440 19026 3496
rect 18878 3168 18934 3224
rect 20074 12860 20076 12880
rect 20076 12860 20128 12880
rect 20128 12860 20130 12880
rect 20074 12824 20130 12860
rect 20350 20440 20406 20496
rect 20350 20168 20406 20224
rect 20350 17720 20406 17776
rect 20350 17312 20406 17368
rect 20718 24520 20774 24556
rect 22466 24928 22522 24984
rect 20534 23432 20590 23488
rect 21086 24112 21142 24168
rect 20902 22108 20904 22128
rect 20904 22108 20956 22128
rect 20956 22108 20958 22128
rect 20902 22072 20958 22108
rect 20718 21548 20774 21584
rect 20718 21528 20720 21548
rect 20720 21528 20772 21548
rect 20772 21528 20774 21548
rect 20902 21392 20958 21448
rect 20718 20440 20774 20496
rect 20442 14864 20498 14920
rect 20902 20868 20958 20904
rect 20902 20848 20904 20868
rect 20904 20848 20956 20868
rect 20956 20848 20958 20868
rect 20902 19216 20958 19272
rect 20718 18400 20774 18456
rect 21822 24520 21878 24576
rect 21270 20304 21326 20360
rect 21362 19624 21418 19680
rect 21086 18128 21142 18184
rect 20994 17584 21050 17640
rect 20626 16360 20682 16416
rect 20626 15408 20682 15464
rect 20810 15272 20866 15328
rect 20902 15000 20958 15056
rect 20994 14320 21050 14376
rect 20718 13932 20774 13968
rect 20718 13912 20720 13932
rect 20720 13912 20772 13932
rect 20772 13912 20774 13932
rect 19982 11736 20038 11792
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19890 11212 19946 11248
rect 19890 11192 19892 11212
rect 19892 11192 19944 11212
rect 19944 11192 19946 11212
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19338 10240 19394 10296
rect 20258 11600 20314 11656
rect 20258 10668 20314 10704
rect 20258 10648 20260 10668
rect 20260 10648 20312 10668
rect 20312 10648 20314 10668
rect 19522 9560 19578 9616
rect 22374 24248 22430 24304
rect 22190 21684 22246 21720
rect 22190 21664 22192 21684
rect 22192 21664 22244 21684
rect 22244 21664 22246 21684
rect 22190 20984 22246 21040
rect 21914 20032 21970 20088
rect 21546 18944 21602 19000
rect 21546 18708 21548 18728
rect 21548 18708 21600 18728
rect 21600 18708 21602 18728
rect 21546 18672 21602 18708
rect 21178 16224 21234 16280
rect 20810 12416 20866 12472
rect 20718 10956 20720 10976
rect 20720 10956 20772 10976
rect 20772 10956 20774 10976
rect 20718 10920 20774 10956
rect 20902 10784 20958 10840
rect 21362 17992 21418 18048
rect 22006 19216 22062 19272
rect 21914 18944 21970 19000
rect 21362 14864 21418 14920
rect 21454 14456 21510 14512
rect 21086 12144 21142 12200
rect 21178 10784 21234 10840
rect 21270 10648 21326 10704
rect 21730 13812 21732 13832
rect 21732 13812 21784 13832
rect 21784 13812 21786 13832
rect 21730 13776 21786 13812
rect 21638 12960 21694 13016
rect 21546 10376 21602 10432
rect 21178 10104 21234 10160
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 20350 9288 20406 9344
rect 19614 8608 19670 8664
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19614 6160 19670 6216
rect 19154 6024 19210 6080
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19246 5888 19302 5944
rect 20074 5888 20130 5944
rect 19338 4936 19394 4992
rect 19246 4800 19302 4856
rect 19154 4120 19210 4176
rect 19154 3712 19210 3768
rect 19338 3984 19394 4040
rect 19062 2896 19118 2952
rect 18510 1808 18566 1864
rect 19430 2760 19486 2816
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19982 4428 19984 4448
rect 19984 4428 20036 4448
rect 20036 4428 20038 4448
rect 19982 4392 20038 4428
rect 21362 9424 21418 9480
rect 20994 9288 21050 9344
rect 20718 8372 20720 8392
rect 20720 8372 20772 8392
rect 20772 8372 20774 8392
rect 20718 8336 20774 8372
rect 20902 7928 20958 7984
rect 20350 5480 20406 5536
rect 20534 6568 20590 6624
rect 20626 5480 20682 5536
rect 21546 9424 21602 9480
rect 22006 18536 22062 18592
rect 22742 23976 22798 24032
rect 22742 22752 22798 22808
rect 22742 20596 22798 20632
rect 22742 20576 22744 20596
rect 22744 20576 22796 20596
rect 22796 20576 22798 20596
rect 22006 17856 22062 17912
rect 21914 17448 21970 17504
rect 22190 16496 22246 16552
rect 22466 17856 22522 17912
rect 21822 13096 21878 13152
rect 21546 9016 21602 9072
rect 21730 9016 21786 9072
rect 22098 14048 22154 14104
rect 21914 12416 21970 12472
rect 22006 7792 22062 7848
rect 20442 3984 20498 4040
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19890 3032 19946 3088
rect 20074 3052 20130 3088
rect 20074 3032 20076 3052
rect 20076 3032 20128 3052
rect 20128 3032 20130 3052
rect 20074 2760 20130 2816
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 19522 2216 19578 2272
rect 19798 1400 19854 1456
rect 20258 1536 20314 1592
rect 20166 1400 20222 1456
rect 20718 3848 20774 3904
rect 21454 4664 21510 4720
rect 20994 3984 21050 4040
rect 21362 3576 21418 3632
rect 22282 15136 22338 15192
rect 22282 13948 22284 13968
rect 22284 13948 22336 13968
rect 22336 13948 22338 13968
rect 22282 13912 22338 13948
rect 22282 12280 22338 12336
rect 22558 17076 22560 17096
rect 22560 17076 22612 17096
rect 22612 17076 22614 17096
rect 22558 17040 22614 17076
rect 22558 15680 22614 15736
rect 23294 23160 23350 23216
rect 23018 22924 23020 22944
rect 23020 22924 23072 22944
rect 23072 22924 23074 22944
rect 23018 22888 23074 22924
rect 23938 25336 23994 25392
rect 24582 27104 24638 27160
rect 24766 26560 24822 26616
rect 25318 25880 25374 25936
rect 24766 25744 24822 25800
rect 24766 25336 24822 25392
rect 23662 23840 23718 23896
rect 23202 21800 23258 21856
rect 23018 21392 23074 21448
rect 22834 19216 22890 19272
rect 22926 18300 22928 18320
rect 22928 18300 22980 18320
rect 22980 18300 22982 18320
rect 22926 18264 22982 18300
rect 23018 17312 23074 17368
rect 22834 16768 22890 16824
rect 23018 16496 23074 16552
rect 23018 14884 23074 14920
rect 23018 14864 23020 14884
rect 23020 14864 23072 14884
rect 23072 14864 23074 14884
rect 22926 13776 22982 13832
rect 22374 11600 22430 11656
rect 22650 11348 22706 11384
rect 22650 11328 22652 11348
rect 22652 11328 22704 11348
rect 22704 11328 22706 11348
rect 22282 9152 22338 9208
rect 22466 7384 22522 7440
rect 21730 4548 21786 4584
rect 21730 4528 21732 4548
rect 21732 4528 21784 4548
rect 21784 4528 21786 4548
rect 22374 6160 22430 6216
rect 22282 4392 22338 4448
rect 22834 10920 22890 10976
rect 23018 13640 23074 13696
rect 23846 24112 23902 24168
rect 23846 23432 23902 23488
rect 23754 22888 23810 22944
rect 23662 21664 23718 21720
rect 23846 21800 23902 21856
rect 23478 20576 23534 20632
rect 23662 21120 23718 21176
rect 23570 19352 23626 19408
rect 23294 17312 23350 17368
rect 23570 17176 23626 17232
rect 23386 15136 23442 15192
rect 23386 14456 23442 14512
rect 23386 12416 23442 12472
rect 23110 12280 23166 12336
rect 23294 12008 23350 12064
rect 23386 11056 23442 11112
rect 23110 9152 23166 9208
rect 22926 8916 22928 8936
rect 22928 8916 22980 8936
rect 22980 8916 22982 8936
rect 22926 8880 22982 8916
rect 22742 4936 22798 4992
rect 22834 4528 22890 4584
rect 22650 3712 22706 3768
rect 23294 10784 23350 10840
rect 23570 15544 23626 15600
rect 23570 12708 23626 12744
rect 23570 12688 23572 12708
rect 23572 12688 23624 12708
rect 23624 12688 23626 12708
rect 23570 12416 23626 12472
rect 23478 10512 23534 10568
rect 23478 9832 23534 9888
rect 23294 9424 23350 9480
rect 24030 19760 24086 19816
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 26238 24792 26294 24848
rect 24214 24656 24270 24712
rect 25778 24656 25834 24712
rect 24490 24268 24546 24304
rect 24490 24248 24492 24268
rect 24492 24248 24544 24268
rect 24544 24248 24546 24268
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24306 23432 24362 23488
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 25134 24132 25190 24168
rect 25134 24112 25136 24132
rect 25136 24112 25188 24132
rect 25188 24112 25190 24132
rect 25226 23704 25282 23760
rect 25410 23568 25466 23624
rect 25318 23296 25374 23352
rect 25042 22652 25044 22672
rect 25044 22652 25096 22672
rect 25096 22652 25098 22672
rect 25042 22616 25098 22652
rect 25410 23024 25466 23080
rect 25502 22480 25558 22536
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24490 20052 24546 20088
rect 24490 20032 24492 20052
rect 24492 20032 24544 20052
rect 24544 20032 24546 20052
rect 24950 20168 25006 20224
rect 24674 19624 24730 19680
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 23938 18400 23994 18456
rect 24582 18808 24638 18864
rect 24306 18672 24362 18728
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 25226 20848 25282 20904
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24214 17040 24270 17096
rect 24030 16532 24032 16552
rect 24032 16532 24084 16552
rect 24084 16532 24086 16552
rect 24030 16496 24086 16532
rect 23846 16224 23902 16280
rect 23754 16088 23810 16144
rect 23846 15852 23848 15872
rect 23848 15852 23900 15872
rect 23900 15852 23902 15872
rect 23846 15816 23902 15852
rect 24030 15272 24086 15328
rect 24122 15020 24178 15056
rect 24122 15000 24124 15020
rect 24124 15000 24176 15020
rect 24176 15000 24178 15020
rect 24122 14320 24178 14376
rect 24122 13640 24178 13696
rect 24766 17332 24822 17368
rect 24766 17312 24768 17332
rect 24768 17312 24820 17332
rect 24820 17312 24822 17332
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24306 15000 24362 15056
rect 24582 14456 24638 14512
rect 24306 14320 24362 14376
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24766 14592 24822 14648
rect 25318 20032 25374 20088
rect 25042 16224 25098 16280
rect 23754 13368 23810 13424
rect 23938 13368 23994 13424
rect 23846 13096 23902 13152
rect 23754 11056 23810 11112
rect 23662 10240 23718 10296
rect 23754 10124 23810 10160
rect 23754 10104 23756 10124
rect 23756 10104 23808 10124
rect 23808 10104 23810 10124
rect 23662 9696 23718 9752
rect 23386 7792 23442 7848
rect 23570 8880 23626 8936
rect 23478 7248 23534 7304
rect 23386 6452 23442 6488
rect 23386 6432 23388 6452
rect 23388 6432 23440 6452
rect 23440 6432 23442 6452
rect 23570 5788 23572 5808
rect 23572 5788 23624 5808
rect 23624 5788 23626 5808
rect 21178 3188 21234 3224
rect 21178 3168 21180 3188
rect 21180 3168 21232 3188
rect 21232 3168 21234 3188
rect 21546 2896 21602 2952
rect 20534 2388 20536 2408
rect 20536 2388 20588 2408
rect 20588 2388 20590 2408
rect 20534 2352 20590 2388
rect 20902 1672 20958 1728
rect 21178 2488 21234 2544
rect 21086 1944 21142 2000
rect 21086 1672 21142 1728
rect 20994 1128 21050 1184
rect 14186 40 14242 96
rect 22558 3440 22614 3496
rect 22466 3340 22468 3360
rect 22468 3340 22520 3360
rect 22520 3340 22522 3360
rect 22466 3304 22522 3340
rect 21638 2488 21694 2544
rect 22098 2896 22154 2952
rect 22558 2760 22614 2816
rect 23570 5752 23626 5788
rect 23202 5616 23258 5672
rect 23018 2760 23074 2816
rect 23754 8336 23810 8392
rect 24122 10376 24178 10432
rect 23846 7928 23902 7984
rect 24122 8608 24178 8664
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24306 12552 24362 12608
rect 24674 12416 24730 12472
rect 25226 16668 25228 16688
rect 25228 16668 25280 16688
rect 25280 16668 25282 16688
rect 25226 16632 25282 16668
rect 25226 13912 25282 13968
rect 25042 12844 25098 12880
rect 25042 12824 25044 12844
rect 25044 12824 25096 12844
rect 25096 12824 25098 12844
rect 25042 12280 25098 12336
rect 24674 12008 24730 12064
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 25134 12144 25190 12200
rect 25686 21528 25742 21584
rect 25594 21120 25650 21176
rect 25410 16632 25466 16688
rect 24858 10240 24914 10296
rect 24950 9968 25006 10024
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24858 9696 24914 9752
rect 24398 9152 24454 9208
rect 24674 9016 24730 9072
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24122 7928 24178 7984
rect 23754 6432 23810 6488
rect 23294 4936 23350 4992
rect 23662 5480 23718 5536
rect 23938 7540 23994 7576
rect 23938 7520 23940 7540
rect 23940 7520 23992 7540
rect 23992 7520 23994 7540
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24306 7248 24362 7304
rect 23938 5480 23994 5536
rect 23846 5344 23902 5400
rect 23478 2352 23534 2408
rect 23938 4256 23994 4312
rect 23662 3884 23664 3904
rect 23664 3884 23716 3904
rect 23716 3884 23718 3904
rect 23662 3848 23718 3884
rect 23662 3068 23664 3088
rect 23664 3068 23716 3088
rect 23716 3068 23718 3088
rect 23662 3032 23718 3068
rect 23754 2896 23810 2952
rect 23570 2080 23626 2136
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24582 6296 24638 6352
rect 24674 5752 24730 5808
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24858 5516 24860 5536
rect 24860 5516 24912 5536
rect 24912 5516 24914 5536
rect 24858 5480 24914 5516
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24398 3848 24454 3904
rect 24674 3984 24730 4040
rect 24582 3576 24638 3632
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24030 3032 24086 3088
rect 23938 1536 23994 1592
rect 23846 856 23902 912
rect 20902 40 20958 96
rect 24490 2624 24546 2680
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 25042 6180 25098 6216
rect 25042 6160 25044 6180
rect 25044 6160 25096 6180
rect 25096 6160 25098 6180
rect 24950 3712 25006 3768
rect 25226 11736 25282 11792
rect 25226 11192 25282 11248
rect 25686 11464 25742 11520
rect 25410 9288 25466 9344
rect 25318 8880 25374 8936
rect 25226 5108 25228 5128
rect 25228 5108 25280 5128
rect 25280 5108 25282 5128
rect 25226 5072 25282 5108
rect 25226 4120 25282 4176
rect 25410 3984 25466 4040
rect 25410 3440 25466 3496
rect 25962 20476 25964 20496
rect 25964 20476 26016 20496
rect 26016 20476 26018 20496
rect 25962 20440 26018 20476
rect 25870 19080 25926 19136
rect 25870 13640 25926 13696
rect 25962 13368 26018 13424
rect 26146 20712 26202 20768
rect 27618 26288 27674 26344
rect 27066 22344 27122 22400
rect 26238 19760 26294 19816
rect 26238 18028 26240 18048
rect 26240 18028 26292 18048
rect 26292 18028 26294 18048
rect 26238 17992 26294 18028
rect 25778 11328 25834 11384
rect 26054 12416 26110 12472
rect 25778 4936 25834 4992
rect 24214 992 24270 1048
rect 25594 2524 25596 2544
rect 25596 2524 25648 2544
rect 25648 2524 25650 2544
rect 25594 2488 25650 2524
rect 25870 1944 25926 2000
rect 25502 1808 25558 1864
rect 26422 10784 26478 10840
rect 27618 3440 27674 3496
rect 27066 2760 27122 2816
rect 26514 1400 26570 1456
rect 24030 312 24086 368
<< metal3 >>
rect 0 27706 480 27736
rect 1669 27706 1735 27709
rect 0 27704 1735 27706
rect 0 27648 1674 27704
rect 1730 27648 1735 27704
rect 0 27646 1735 27648
rect 0 27616 480 27646
rect 1669 27643 1735 27646
rect 24669 27706 24735 27709
rect 27520 27706 28000 27736
rect 24669 27704 28000 27706
rect 24669 27648 24674 27704
rect 24730 27648 28000 27704
rect 24669 27646 28000 27648
rect 24669 27643 24735 27646
rect 27520 27616 28000 27646
rect 0 27162 480 27192
rect 1485 27162 1551 27165
rect 0 27160 1551 27162
rect 0 27104 1490 27160
rect 1546 27104 1551 27160
rect 0 27102 1551 27104
rect 0 27072 480 27102
rect 1485 27099 1551 27102
rect 24577 27162 24643 27165
rect 27520 27162 28000 27192
rect 24577 27160 28000 27162
rect 24577 27104 24582 27160
rect 24638 27104 28000 27160
rect 24577 27102 28000 27104
rect 24577 27099 24643 27102
rect 27520 27072 28000 27102
rect 0 26618 480 26648
rect 2313 26618 2379 26621
rect 0 26616 2379 26618
rect 0 26560 2318 26616
rect 2374 26560 2379 26616
rect 0 26558 2379 26560
rect 0 26528 480 26558
rect 2313 26555 2379 26558
rect 24761 26618 24827 26621
rect 27520 26618 28000 26648
rect 24761 26616 28000 26618
rect 24761 26560 24766 26616
rect 24822 26560 28000 26616
rect 24761 26558 28000 26560
rect 24761 26555 24827 26558
rect 27520 26528 28000 26558
rect 8334 26284 8340 26348
rect 8404 26346 8410 26348
rect 27613 26346 27679 26349
rect 8404 26344 27679 26346
rect 8404 26288 27618 26344
rect 27674 26288 27679 26344
rect 8404 26286 27679 26288
rect 8404 26284 8410 26286
rect 27613 26283 27679 26286
rect 9949 26074 10015 26077
rect 20621 26074 20687 26077
rect 9949 26072 20687 26074
rect 9949 26016 9954 26072
rect 10010 26016 20626 26072
rect 20682 26016 20687 26072
rect 9949 26014 20687 26016
rect 9949 26011 10015 26014
rect 20621 26011 20687 26014
rect 0 25938 480 25968
rect 1577 25938 1643 25941
rect 0 25936 1643 25938
rect 0 25880 1582 25936
rect 1638 25880 1643 25936
rect 0 25878 1643 25880
rect 0 25848 480 25878
rect 1577 25875 1643 25878
rect 7649 25938 7715 25941
rect 8334 25938 8340 25940
rect 7649 25936 8340 25938
rect 7649 25880 7654 25936
rect 7710 25880 8340 25936
rect 7649 25878 8340 25880
rect 7649 25875 7715 25878
rect 8334 25876 8340 25878
rect 8404 25876 8410 25940
rect 11513 25938 11579 25941
rect 25313 25938 25379 25941
rect 27520 25938 28000 25968
rect 11513 25936 25379 25938
rect 11513 25880 11518 25936
rect 11574 25880 25318 25936
rect 25374 25880 25379 25936
rect 11513 25878 25379 25880
rect 11513 25875 11579 25878
rect 25313 25875 25379 25878
rect 25454 25878 28000 25938
rect 24761 25802 24827 25805
rect 25454 25802 25514 25878
rect 27520 25848 28000 25878
rect 24761 25800 25514 25802
rect 24761 25744 24766 25800
rect 24822 25744 25514 25800
rect 24761 25742 25514 25744
rect 24761 25739 24827 25742
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 0 25394 480 25424
rect 2681 25394 2747 25397
rect 0 25392 2747 25394
rect 0 25336 2686 25392
rect 2742 25336 2747 25392
rect 0 25334 2747 25336
rect 0 25304 480 25334
rect 2681 25331 2747 25334
rect 10869 25394 10935 25397
rect 16941 25394 17007 25397
rect 10869 25392 17007 25394
rect 10869 25336 10874 25392
rect 10930 25336 16946 25392
rect 17002 25336 17007 25392
rect 10869 25334 17007 25336
rect 10869 25331 10935 25334
rect 16941 25331 17007 25334
rect 17309 25394 17375 25397
rect 23933 25394 23999 25397
rect 17309 25392 23999 25394
rect 17309 25336 17314 25392
rect 17370 25336 23938 25392
rect 23994 25336 23999 25392
rect 17309 25334 23999 25336
rect 17309 25331 17375 25334
rect 23933 25331 23999 25334
rect 24761 25394 24827 25397
rect 27520 25394 28000 25424
rect 24761 25392 28000 25394
rect 24761 25336 24766 25392
rect 24822 25336 28000 25392
rect 24761 25334 28000 25336
rect 24761 25331 24827 25334
rect 27520 25304 28000 25334
rect 10225 25258 10291 25261
rect 21357 25258 21423 25261
rect 10225 25256 21423 25258
rect 10225 25200 10230 25256
rect 10286 25200 21362 25256
rect 21418 25200 21423 25256
rect 10225 25198 21423 25200
rect 10225 25195 10291 25198
rect 21357 25195 21423 25198
rect 6729 25122 6795 25125
rect 10869 25122 10935 25125
rect 6729 25120 10935 25122
rect 6729 25064 6734 25120
rect 6790 25064 10874 25120
rect 10930 25064 10935 25120
rect 6729 25062 10935 25064
rect 6729 25059 6795 25062
rect 10869 25059 10935 25062
rect 18505 25122 18571 25125
rect 21265 25122 21331 25125
rect 18505 25120 21331 25122
rect 18505 25064 18510 25120
rect 18566 25064 21270 25120
rect 21326 25064 21331 25120
rect 18505 25062 21331 25064
rect 18505 25059 18571 25062
rect 21265 25059 21331 25062
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 14733 24986 14799 24989
rect 18413 24986 18479 24989
rect 14733 24984 14842 24986
rect 14733 24928 14738 24984
rect 14794 24928 14842 24984
rect 14733 24923 14842 24928
rect 0 24850 480 24880
rect 1577 24850 1643 24853
rect 0 24848 1643 24850
rect 0 24792 1582 24848
rect 1638 24792 1643 24848
rect 0 24790 1643 24792
rect 0 24760 480 24790
rect 1577 24787 1643 24790
rect 8661 24850 8727 24853
rect 13629 24850 13695 24853
rect 8661 24848 13695 24850
rect 8661 24792 8666 24848
rect 8722 24792 13634 24848
rect 13690 24792 13695 24848
rect 8661 24790 13695 24792
rect 14782 24850 14842 24923
rect 15334 24984 18479 24986
rect 15334 24928 18418 24984
rect 18474 24928 18479 24984
rect 15334 24926 18479 24928
rect 15101 24850 15167 24853
rect 15334 24850 15394 24926
rect 18413 24923 18479 24926
rect 18597 24986 18663 24989
rect 22461 24986 22527 24989
rect 18597 24984 22527 24986
rect 18597 24928 18602 24984
rect 18658 24928 22466 24984
rect 22522 24928 22527 24984
rect 18597 24926 22527 24928
rect 18597 24923 18663 24926
rect 22461 24923 22527 24926
rect 14782 24848 15394 24850
rect 14782 24792 15106 24848
rect 15162 24792 15394 24848
rect 14782 24790 15394 24792
rect 8661 24787 8727 24790
rect 13629 24787 13695 24790
rect 15101 24787 15167 24790
rect 15878 24788 15884 24852
rect 15948 24850 15954 24852
rect 16021 24850 16087 24853
rect 15948 24848 16087 24850
rect 15948 24792 16026 24848
rect 16082 24792 16087 24848
rect 15948 24790 16087 24792
rect 15948 24788 15954 24790
rect 16021 24787 16087 24790
rect 16573 24850 16639 24853
rect 21173 24850 21239 24853
rect 16573 24848 21239 24850
rect 16573 24792 16578 24848
rect 16634 24792 21178 24848
rect 21234 24792 21239 24848
rect 16573 24790 21239 24792
rect 16573 24787 16639 24790
rect 21173 24787 21239 24790
rect 26233 24850 26299 24853
rect 27520 24850 28000 24880
rect 26233 24848 28000 24850
rect 26233 24792 26238 24848
rect 26294 24792 28000 24848
rect 26233 24790 28000 24792
rect 26233 24787 26299 24790
rect 27520 24760 28000 24790
rect 11145 24716 11211 24717
rect 11094 24652 11100 24716
rect 11164 24714 11211 24716
rect 12893 24714 12959 24717
rect 19793 24714 19859 24717
rect 11164 24712 11256 24714
rect 11206 24656 11256 24712
rect 11164 24654 11256 24656
rect 12893 24712 19859 24714
rect 12893 24656 12898 24712
rect 12954 24656 19798 24712
rect 19854 24656 19859 24712
rect 12893 24654 19859 24656
rect 11164 24652 11211 24654
rect 11145 24651 11211 24652
rect 12893 24651 12959 24654
rect 19793 24651 19859 24654
rect 24209 24714 24275 24717
rect 25773 24714 25839 24717
rect 24209 24712 25839 24714
rect 24209 24656 24214 24712
rect 24270 24656 25778 24712
rect 25834 24656 25839 24712
rect 24209 24654 25839 24656
rect 24209 24651 24275 24654
rect 25773 24651 25839 24654
rect 11237 24580 11303 24581
rect 11237 24578 11284 24580
rect 11192 24576 11284 24578
rect 11192 24520 11242 24576
rect 11192 24518 11284 24520
rect 11237 24516 11284 24518
rect 11348 24516 11354 24580
rect 14641 24578 14707 24581
rect 18597 24578 18663 24581
rect 14641 24576 18663 24578
rect 14641 24520 14646 24576
rect 14702 24520 18602 24576
rect 18658 24520 18663 24576
rect 14641 24518 18663 24520
rect 11237 24515 11303 24516
rect 14641 24515 14707 24518
rect 18597 24515 18663 24518
rect 20478 24516 20484 24580
rect 20548 24578 20554 24580
rect 20713 24578 20779 24581
rect 20548 24576 20779 24578
rect 20548 24520 20718 24576
rect 20774 24520 20779 24576
rect 20548 24518 20779 24520
rect 20548 24516 20554 24518
rect 20713 24515 20779 24518
rect 21817 24578 21883 24581
rect 21950 24578 21956 24580
rect 21817 24576 21956 24578
rect 21817 24520 21822 24576
rect 21878 24520 21956 24576
rect 21817 24518 21956 24520
rect 21817 24515 21883 24518
rect 21950 24516 21956 24518
rect 22020 24516 22026 24580
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 6453 24442 6519 24445
rect 9673 24442 9739 24445
rect 6453 24440 9739 24442
rect 6453 24384 6458 24440
rect 6514 24384 9678 24440
rect 9734 24384 9739 24440
rect 6453 24382 9739 24384
rect 6453 24379 6519 24382
rect 9673 24379 9739 24382
rect 11237 24442 11303 24445
rect 17309 24442 17375 24445
rect 11237 24440 17375 24442
rect 11237 24384 11242 24440
rect 11298 24384 17314 24440
rect 17370 24384 17375 24440
rect 11237 24382 17375 24384
rect 11237 24379 11303 24382
rect 17309 24379 17375 24382
rect 2037 24306 2103 24309
rect 10777 24306 10843 24309
rect 13537 24306 13603 24309
rect 2037 24304 7666 24306
rect 2037 24248 2042 24304
rect 2098 24248 7666 24304
rect 2037 24246 7666 24248
rect 2037 24243 2103 24246
rect 0 24170 480 24200
rect 3233 24170 3299 24173
rect 0 24168 3299 24170
rect 0 24112 3238 24168
rect 3294 24112 3299 24168
rect 0 24110 3299 24112
rect 0 24080 480 24110
rect 3233 24107 3299 24110
rect 5533 24170 5599 24173
rect 7606 24170 7666 24246
rect 10777 24304 13603 24306
rect 10777 24248 10782 24304
rect 10838 24248 13542 24304
rect 13598 24248 13603 24304
rect 10777 24246 13603 24248
rect 10777 24243 10843 24246
rect 13537 24243 13603 24246
rect 17769 24306 17835 24309
rect 19977 24306 20043 24309
rect 17769 24304 20043 24306
rect 17769 24248 17774 24304
rect 17830 24248 19982 24304
rect 20038 24248 20043 24304
rect 17769 24246 20043 24248
rect 17769 24243 17835 24246
rect 19977 24243 20043 24246
rect 22369 24306 22435 24309
rect 24485 24306 24551 24309
rect 22369 24304 24551 24306
rect 22369 24248 22374 24304
rect 22430 24248 24490 24304
rect 24546 24248 24551 24304
rect 22369 24246 24551 24248
rect 22369 24243 22435 24246
rect 24485 24243 24551 24246
rect 12566 24170 12572 24172
rect 5533 24168 7482 24170
rect 5533 24112 5538 24168
rect 5594 24112 7482 24168
rect 5533 24110 7482 24112
rect 7606 24110 12572 24170
rect 5533 24107 5599 24110
rect 7422 24034 7482 24110
rect 12566 24108 12572 24110
rect 12636 24170 12642 24172
rect 13445 24170 13511 24173
rect 21081 24170 21147 24173
rect 23841 24172 23907 24173
rect 12636 24168 13511 24170
rect 12636 24112 13450 24168
rect 13506 24112 13511 24168
rect 12636 24110 13511 24112
rect 12636 24108 12642 24110
rect 13445 24107 13511 24110
rect 14782 24168 21147 24170
rect 14782 24112 21086 24168
rect 21142 24112 21147 24168
rect 14782 24110 21147 24112
rect 12014 24034 12020 24036
rect 7422 23974 12020 24034
rect 12014 23972 12020 23974
rect 12084 23972 12090 24036
rect 12249 24034 12315 24037
rect 12433 24034 12499 24037
rect 12249 24032 12499 24034
rect 12249 23976 12254 24032
rect 12310 23976 12438 24032
rect 12494 23976 12499 24032
rect 12249 23974 12499 23976
rect 12249 23971 12315 23974
rect 12433 23971 12499 23974
rect 12709 24034 12775 24037
rect 14782 24034 14842 24110
rect 21081 24107 21147 24110
rect 23790 24108 23796 24172
rect 23860 24170 23907 24172
rect 25129 24170 25195 24173
rect 27520 24170 28000 24200
rect 23860 24168 23952 24170
rect 23902 24112 23952 24168
rect 23860 24110 23952 24112
rect 25129 24168 28000 24170
rect 25129 24112 25134 24168
rect 25190 24112 28000 24168
rect 25129 24110 28000 24112
rect 23860 24108 23907 24110
rect 23841 24107 23907 24108
rect 25129 24107 25195 24110
rect 27520 24080 28000 24110
rect 12709 24032 14842 24034
rect 12709 23976 12714 24032
rect 12770 23976 14842 24032
rect 12709 23974 14842 23976
rect 12709 23971 12775 23974
rect 15510 23972 15516 24036
rect 15580 24034 15586 24036
rect 22737 24034 22803 24037
rect 15580 24032 22803 24034
rect 15580 23976 22742 24032
rect 22798 23976 22803 24032
rect 15580 23974 22803 23976
rect 15580 23972 15586 23974
rect 22737 23971 22803 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 7189 23898 7255 23901
rect 14089 23898 14155 23901
rect 7189 23896 14155 23898
rect 7189 23840 7194 23896
rect 7250 23840 14094 23896
rect 14150 23840 14155 23896
rect 7189 23838 14155 23840
rect 7189 23835 7255 23838
rect 14089 23835 14155 23838
rect 14273 23898 14339 23901
rect 14774 23898 14780 23900
rect 14273 23896 14780 23898
rect 14273 23840 14278 23896
rect 14334 23840 14780 23896
rect 14273 23838 14780 23840
rect 14273 23835 14339 23838
rect 14774 23836 14780 23838
rect 14844 23836 14850 23900
rect 20437 23898 20503 23901
rect 23657 23898 23723 23901
rect 20437 23896 23723 23898
rect 20437 23840 20442 23896
rect 20498 23840 23662 23896
rect 23718 23840 23723 23896
rect 20437 23838 23723 23840
rect 20437 23835 20503 23838
rect 23657 23835 23723 23838
rect 6637 23762 6703 23765
rect 9305 23762 9371 23765
rect 11237 23762 11303 23765
rect 6637 23760 9371 23762
rect 6637 23704 6642 23760
rect 6698 23704 9310 23760
rect 9366 23704 9371 23760
rect 6637 23702 9371 23704
rect 6637 23699 6703 23702
rect 9305 23699 9371 23702
rect 10550 23760 11303 23762
rect 10550 23704 11242 23760
rect 11298 23704 11303 23760
rect 10550 23702 11303 23704
rect 0 23626 480 23656
rect 3509 23626 3575 23629
rect 0 23624 3575 23626
rect 0 23568 3514 23624
rect 3570 23568 3575 23624
rect 0 23566 3575 23568
rect 0 23536 480 23566
rect 3509 23563 3575 23566
rect 5441 23626 5507 23629
rect 10550 23626 10610 23702
rect 11237 23699 11303 23702
rect 12433 23762 12499 23765
rect 14549 23762 14615 23765
rect 12433 23760 14615 23762
rect 12433 23704 12438 23760
rect 12494 23704 14554 23760
rect 14610 23704 14615 23760
rect 12433 23702 14615 23704
rect 12433 23699 12499 23702
rect 14549 23699 14615 23702
rect 14733 23762 14799 23765
rect 16798 23762 16804 23764
rect 14733 23760 16804 23762
rect 14733 23704 14738 23760
rect 14794 23704 16804 23760
rect 14733 23702 16804 23704
rect 14733 23699 14799 23702
rect 16798 23700 16804 23702
rect 16868 23700 16874 23764
rect 18689 23762 18755 23765
rect 25221 23762 25287 23765
rect 18689 23760 25287 23762
rect 18689 23704 18694 23760
rect 18750 23704 25226 23760
rect 25282 23704 25287 23760
rect 18689 23702 25287 23704
rect 18689 23699 18755 23702
rect 25221 23699 25287 23702
rect 5441 23624 10610 23626
rect 5441 23568 5446 23624
rect 5502 23568 10610 23624
rect 5441 23566 10610 23568
rect 11053 23626 11119 23629
rect 13854 23626 13860 23628
rect 11053 23624 13860 23626
rect 11053 23568 11058 23624
rect 11114 23568 13860 23624
rect 11053 23566 13860 23568
rect 5441 23563 5507 23566
rect 11053 23563 11119 23566
rect 13854 23564 13860 23566
rect 13924 23564 13930 23628
rect 15101 23626 15167 23629
rect 16246 23626 16252 23628
rect 15101 23624 16252 23626
rect 15101 23568 15106 23624
rect 15162 23568 16252 23624
rect 15101 23566 16252 23568
rect 15101 23563 15167 23566
rect 16246 23564 16252 23566
rect 16316 23564 16322 23628
rect 20161 23626 20227 23629
rect 24710 23626 24716 23628
rect 20161 23624 24716 23626
rect 20161 23568 20166 23624
rect 20222 23568 24716 23624
rect 20161 23566 24716 23568
rect 20161 23563 20227 23566
rect 24710 23564 24716 23566
rect 24780 23564 24786 23628
rect 25405 23626 25471 23629
rect 27520 23626 28000 23656
rect 25405 23624 28000 23626
rect 25405 23568 25410 23624
rect 25466 23568 28000 23624
rect 25405 23566 28000 23568
rect 25405 23563 25471 23566
rect 27520 23536 28000 23566
rect 5349 23490 5415 23493
rect 9857 23490 9923 23493
rect 5349 23488 9923 23490
rect 5349 23432 5354 23488
rect 5410 23432 9862 23488
rect 9918 23432 9923 23488
rect 5349 23430 9923 23432
rect 5349 23427 5415 23430
rect 9857 23427 9923 23430
rect 15285 23492 15351 23493
rect 15285 23488 15332 23492
rect 15396 23490 15402 23492
rect 16389 23490 16455 23493
rect 19425 23492 19491 23493
rect 15285 23432 15290 23488
rect 15285 23428 15332 23432
rect 15396 23430 15442 23490
rect 16389 23488 19074 23490
rect 16389 23432 16394 23488
rect 16450 23432 19074 23488
rect 16389 23430 19074 23432
rect 15396 23428 15402 23430
rect 15285 23427 15351 23428
rect 16389 23427 16455 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 841 23354 907 23357
rect 5901 23354 5967 23357
rect 841 23352 5967 23354
rect 841 23296 846 23352
rect 902 23296 5906 23352
rect 5962 23296 5967 23352
rect 841 23294 5967 23296
rect 841 23291 907 23294
rect 5901 23291 5967 23294
rect 6126 23292 6132 23356
rect 6196 23354 6202 23356
rect 7281 23354 7347 23357
rect 6196 23352 7347 23354
rect 6196 23296 7286 23352
rect 7342 23296 7347 23352
rect 6196 23294 7347 23296
rect 6196 23292 6202 23294
rect 7281 23291 7347 23294
rect 10961 23354 11027 23357
rect 11462 23354 11468 23356
rect 10961 23352 11468 23354
rect 10961 23296 10966 23352
rect 11022 23296 11468 23352
rect 10961 23294 11468 23296
rect 10961 23291 11027 23294
rect 11462 23292 11468 23294
rect 11532 23292 11538 23356
rect 13629 23354 13695 23357
rect 15561 23354 15627 23357
rect 16757 23354 16823 23357
rect 13629 23352 16823 23354
rect 13629 23296 13634 23352
rect 13690 23296 15566 23352
rect 15622 23296 16762 23352
rect 16818 23296 16823 23352
rect 13629 23294 16823 23296
rect 13629 23291 13695 23294
rect 15561 23291 15627 23294
rect 16757 23291 16823 23294
rect 17401 23354 17467 23357
rect 18873 23354 18939 23357
rect 17401 23352 18939 23354
rect 17401 23296 17406 23352
rect 17462 23296 18878 23352
rect 18934 23296 18939 23352
rect 17401 23294 18939 23296
rect 17401 23291 17467 23294
rect 18873 23291 18939 23294
rect 1669 23218 1735 23221
rect 16389 23218 16455 23221
rect 1669 23216 16455 23218
rect 1669 23160 1674 23216
rect 1730 23160 16394 23216
rect 16450 23160 16455 23216
rect 1669 23158 16455 23160
rect 1669 23155 1735 23158
rect 16389 23155 16455 23158
rect 0 23082 480 23112
rect 2773 23082 2839 23085
rect 0 23080 2839 23082
rect 0 23024 2778 23080
rect 2834 23024 2839 23080
rect 0 23022 2839 23024
rect 0 22992 480 23022
rect 2773 23019 2839 23022
rect 7189 23082 7255 23085
rect 7925 23082 7991 23085
rect 19014 23082 19074 23430
rect 19374 23428 19380 23492
rect 19444 23490 19491 23492
rect 20069 23492 20135 23493
rect 20069 23490 20116 23492
rect 19444 23488 19536 23490
rect 19486 23432 19536 23488
rect 19444 23430 19536 23432
rect 20024 23488 20116 23490
rect 20024 23432 20074 23488
rect 20024 23430 20116 23432
rect 19444 23428 19491 23430
rect 19425 23427 19491 23428
rect 20069 23428 20116 23430
rect 20180 23428 20186 23492
rect 20529 23490 20595 23493
rect 23841 23490 23907 23493
rect 20529 23488 23907 23490
rect 20529 23432 20534 23488
rect 20590 23432 23846 23488
rect 23902 23432 23907 23488
rect 20529 23430 23907 23432
rect 20069 23427 20135 23428
rect 20529 23427 20595 23430
rect 23841 23427 23907 23430
rect 24301 23490 24367 23493
rect 24894 23490 24900 23492
rect 24301 23488 24900 23490
rect 24301 23432 24306 23488
rect 24362 23432 24900 23488
rect 24301 23430 24900 23432
rect 24301 23427 24367 23430
rect 24894 23428 24900 23430
rect 24964 23428 24970 23492
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 20345 23354 20411 23357
rect 25313 23354 25379 23357
rect 20345 23352 25379 23354
rect 20345 23296 20350 23352
rect 20406 23296 25318 23352
rect 25374 23296 25379 23352
rect 20345 23294 25379 23296
rect 20345 23291 20411 23294
rect 25313 23291 25379 23294
rect 19241 23218 19307 23221
rect 23289 23218 23355 23221
rect 19241 23216 23355 23218
rect 19241 23160 19246 23216
rect 19302 23160 23294 23216
rect 23350 23160 23355 23216
rect 19241 23158 23355 23160
rect 19241 23155 19307 23158
rect 23289 23155 23355 23158
rect 23422 23082 23428 23084
rect 7189 23080 7991 23082
rect 7189 23024 7194 23080
rect 7250 23024 7930 23080
rect 7986 23024 7991 23080
rect 7189 23022 7991 23024
rect 7189 23019 7255 23022
rect 7925 23019 7991 23022
rect 14782 23022 16866 23082
rect 19014 23022 23428 23082
rect 8477 22946 8543 22949
rect 14549 22946 14615 22949
rect 8477 22944 14615 22946
rect 8477 22888 8482 22944
rect 8538 22888 14554 22944
rect 14610 22888 14615 22944
rect 8477 22886 14615 22888
rect 8477 22883 8543 22886
rect 14549 22883 14615 22886
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 289 22810 355 22813
rect 1393 22810 1459 22813
rect 4981 22810 5047 22813
rect 289 22808 1226 22810
rect 289 22752 294 22808
rect 350 22752 1226 22808
rect 289 22750 1226 22752
rect 289 22747 355 22750
rect 1166 22674 1226 22750
rect 1393 22808 5047 22810
rect 1393 22752 1398 22808
rect 1454 22752 4986 22808
rect 5042 22752 5047 22808
rect 1393 22750 5047 22752
rect 1393 22747 1459 22750
rect 4981 22747 5047 22750
rect 6545 22810 6611 22813
rect 11421 22810 11487 22813
rect 14782 22810 14842 23022
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 6545 22808 11487 22810
rect 6545 22752 6550 22808
rect 6606 22752 11426 22808
rect 11482 22752 11487 22808
rect 6545 22750 11487 22752
rect 6545 22747 6611 22750
rect 11421 22747 11487 22750
rect 11654 22750 14842 22810
rect 16806 22810 16866 23022
rect 23422 23020 23428 23022
rect 23492 23020 23498 23084
rect 25405 23082 25471 23085
rect 27520 23082 28000 23112
rect 25405 23080 28000 23082
rect 25405 23024 25410 23080
rect 25466 23024 28000 23080
rect 25405 23022 28000 23024
rect 25405 23019 25471 23022
rect 27520 22992 28000 23022
rect 17033 22946 17099 22949
rect 19609 22946 19675 22949
rect 17033 22944 19675 22946
rect 17033 22888 17038 22944
rect 17094 22888 19614 22944
rect 19670 22888 19675 22944
rect 17033 22886 19675 22888
rect 17033 22883 17099 22886
rect 19609 22883 19675 22886
rect 23013 22946 23079 22949
rect 23606 22946 23612 22948
rect 23013 22944 23612 22946
rect 23013 22888 23018 22944
rect 23074 22888 23612 22944
rect 23013 22886 23612 22888
rect 23013 22883 23079 22886
rect 23606 22884 23612 22886
rect 23676 22946 23682 22948
rect 23749 22946 23815 22949
rect 23676 22944 23815 22946
rect 23676 22888 23754 22944
rect 23810 22888 23815 22944
rect 23676 22886 23815 22888
rect 23676 22884 23682 22886
rect 23749 22883 23815 22886
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 20161 22810 20227 22813
rect 16806 22808 20227 22810
rect 16806 22752 20166 22808
rect 20222 22752 20227 22808
rect 16806 22750 20227 22752
rect 6177 22674 6243 22677
rect 1166 22672 6243 22674
rect 1166 22616 6182 22672
rect 6238 22616 6243 22672
rect 1166 22614 6243 22616
rect 6177 22611 6243 22614
rect 7189 22674 7255 22677
rect 11654 22674 11714 22750
rect 20161 22747 20227 22750
rect 22737 22810 22803 22813
rect 23054 22810 23060 22812
rect 22737 22808 23060 22810
rect 22737 22752 22742 22808
rect 22798 22752 23060 22808
rect 22737 22750 23060 22752
rect 22737 22747 22803 22750
rect 23054 22748 23060 22750
rect 23124 22748 23130 22812
rect 7189 22672 11714 22674
rect 7189 22616 7194 22672
rect 7250 22616 11714 22672
rect 7189 22614 11714 22616
rect 12157 22674 12223 22677
rect 15561 22674 15627 22677
rect 12157 22672 15627 22674
rect 12157 22616 12162 22672
rect 12218 22616 15566 22672
rect 15622 22616 15627 22672
rect 12157 22614 15627 22616
rect 7189 22611 7255 22614
rect 12157 22611 12223 22614
rect 15561 22611 15627 22614
rect 19190 22612 19196 22676
rect 19260 22674 19266 22676
rect 25037 22674 25103 22677
rect 19260 22672 25103 22674
rect 19260 22616 25042 22672
rect 25098 22616 25103 22672
rect 19260 22614 25103 22616
rect 19260 22612 19266 22614
rect 25037 22611 25103 22614
rect 0 22538 480 22568
rect 1577 22538 1643 22541
rect 0 22536 1643 22538
rect 0 22480 1582 22536
rect 1638 22480 1643 22536
rect 0 22478 1643 22480
rect 0 22448 480 22478
rect 1577 22475 1643 22478
rect 3141 22538 3207 22541
rect 9765 22538 9831 22541
rect 10501 22538 10567 22541
rect 3141 22536 9831 22538
rect 3141 22480 3146 22536
rect 3202 22480 9770 22536
rect 9826 22480 9831 22536
rect 3141 22478 9831 22480
rect 3141 22475 3207 22478
rect 9765 22475 9831 22478
rect 9952 22536 10567 22538
rect 9952 22480 10506 22536
rect 10562 22480 10567 22536
rect 9952 22478 10567 22480
rect 2221 22402 2287 22405
rect 5533 22402 5599 22405
rect 9952 22402 10012 22478
rect 10501 22475 10567 22478
rect 12157 22538 12223 22541
rect 15837 22538 15903 22541
rect 12157 22536 15903 22538
rect 12157 22480 12162 22536
rect 12218 22480 15842 22536
rect 15898 22480 15903 22536
rect 12157 22478 15903 22480
rect 12157 22475 12223 22478
rect 15837 22475 15903 22478
rect 17033 22538 17099 22541
rect 25497 22538 25563 22541
rect 27520 22538 28000 22568
rect 17033 22536 23122 22538
rect 17033 22480 17038 22536
rect 17094 22480 23122 22536
rect 17033 22478 23122 22480
rect 17033 22475 17099 22478
rect 2221 22400 5599 22402
rect 2221 22344 2226 22400
rect 2282 22344 5538 22400
rect 5594 22344 5599 22400
rect 2221 22342 5599 22344
rect 2221 22339 2287 22342
rect 5533 22339 5599 22342
rect 7238 22342 10012 22402
rect 14549 22402 14615 22405
rect 17769 22402 17835 22405
rect 14549 22400 17835 22402
rect 14549 22344 14554 22400
rect 14610 22344 17774 22400
rect 17830 22344 17835 22400
rect 14549 22342 17835 22344
rect 2405 22268 2471 22269
rect 2405 22266 2452 22268
rect 2360 22264 2452 22266
rect 2360 22208 2410 22264
rect 2360 22206 2452 22208
rect 2405 22204 2452 22206
rect 2516 22204 2522 22268
rect 3233 22266 3299 22269
rect 7238 22266 7298 22342
rect 14549 22339 14615 22342
rect 17769 22339 17835 22342
rect 18229 22402 18295 22405
rect 19241 22402 19307 22405
rect 18229 22400 19307 22402
rect 18229 22344 18234 22400
rect 18290 22344 19246 22400
rect 19302 22344 19307 22400
rect 18229 22342 19307 22344
rect 23062 22402 23122 22478
rect 25497 22536 28000 22538
rect 25497 22480 25502 22536
rect 25558 22480 28000 22536
rect 25497 22478 28000 22480
rect 25497 22475 25563 22478
rect 27520 22448 28000 22478
rect 27061 22402 27127 22405
rect 23062 22400 27127 22402
rect 23062 22344 27066 22400
rect 27122 22344 27127 22400
rect 23062 22342 27127 22344
rect 18229 22339 18295 22342
rect 19241 22339 19307 22342
rect 27061 22339 27127 22342
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 3233 22264 7298 22266
rect 3233 22208 3238 22264
rect 3294 22208 7298 22264
rect 3233 22206 7298 22208
rect 7373 22266 7439 22269
rect 9622 22266 9628 22268
rect 7373 22264 9628 22266
rect 7373 22208 7378 22264
rect 7434 22208 9628 22264
rect 7373 22206 9628 22208
rect 2405 22203 2471 22204
rect 3233 22203 3299 22206
rect 7373 22203 7439 22206
rect 9622 22204 9628 22206
rect 9692 22204 9698 22268
rect 12985 22266 13051 22269
rect 13721 22268 13787 22269
rect 13670 22266 13676 22268
rect 10734 22264 13051 22266
rect 10734 22208 12990 22264
rect 13046 22208 13051 22264
rect 10734 22206 13051 22208
rect 13630 22206 13676 22266
rect 13740 22264 13787 22268
rect 13782 22208 13787 22264
rect 2129 22130 2195 22133
rect 10593 22130 10659 22133
rect 10734 22130 10794 22206
rect 12985 22203 13051 22206
rect 13670 22204 13676 22206
rect 13740 22204 13787 22208
rect 14774 22204 14780 22268
rect 14844 22266 14850 22268
rect 18965 22266 19031 22269
rect 14844 22264 19031 22266
rect 14844 22208 18970 22264
rect 19026 22208 19031 22264
rect 14844 22206 19031 22208
rect 14844 22204 14850 22206
rect 13721 22203 13787 22204
rect 18965 22203 19031 22206
rect 2129 22128 10426 22130
rect 2129 22072 2134 22128
rect 2190 22072 10426 22128
rect 2129 22070 10426 22072
rect 2129 22067 2195 22070
rect 7281 21994 7347 21997
rect 9949 21994 10015 21997
rect 7281 21992 10015 21994
rect 7281 21936 7286 21992
rect 7342 21936 9954 21992
rect 10010 21936 10015 21992
rect 7281 21934 10015 21936
rect 10366 21994 10426 22070
rect 10593 22128 10794 22130
rect 10593 22072 10598 22128
rect 10654 22072 10794 22128
rect 10593 22070 10794 22072
rect 10593 22067 10659 22070
rect 12014 22068 12020 22132
rect 12084 22130 12090 22132
rect 13445 22130 13511 22133
rect 12084 22128 13511 22130
rect 12084 22072 13450 22128
rect 13506 22072 13511 22128
rect 12084 22070 13511 22072
rect 12084 22068 12090 22070
rect 13445 22067 13511 22070
rect 13629 22128 13695 22133
rect 13629 22072 13634 22128
rect 13690 22072 13695 22128
rect 13629 22067 13695 22072
rect 17217 22130 17283 22133
rect 20897 22130 20963 22133
rect 17217 22128 20963 22130
rect 17217 22072 17222 22128
rect 17278 22072 20902 22128
rect 20958 22072 20963 22128
rect 17217 22070 20963 22072
rect 17217 22067 17283 22070
rect 20897 22067 20963 22070
rect 11145 21994 11211 21997
rect 12617 21996 12683 21997
rect 10366 21992 11211 21994
rect 10366 21936 11150 21992
rect 11206 21936 11211 21992
rect 10366 21934 11211 21936
rect 7281 21931 7347 21934
rect 9949 21931 10015 21934
rect 11145 21931 11211 21934
rect 12566 21932 12572 21996
rect 12636 21994 12683 21996
rect 12636 21992 12728 21994
rect 12678 21936 12728 21992
rect 12636 21934 12728 21936
rect 12636 21932 12683 21934
rect 12617 21931 12683 21932
rect 0 21858 480 21888
rect 3877 21858 3943 21861
rect 0 21856 3943 21858
rect 0 21800 3882 21856
rect 3938 21800 3943 21856
rect 0 21798 3943 21800
rect 0 21768 480 21798
rect 3877 21795 3943 21798
rect 9397 21858 9463 21861
rect 13302 21858 13308 21860
rect 9397 21856 13308 21858
rect 9397 21800 9402 21856
rect 9458 21800 13308 21856
rect 9397 21798 13308 21800
rect 9397 21795 9463 21798
rect 13302 21796 13308 21798
rect 13372 21796 13378 21860
rect 13632 21858 13692 22067
rect 18781 21994 18847 21997
rect 19190 21994 19196 21996
rect 18781 21992 19196 21994
rect 18781 21936 18786 21992
rect 18842 21936 19196 21992
rect 18781 21934 19196 21936
rect 18781 21931 18847 21934
rect 19190 21932 19196 21934
rect 19260 21932 19266 21996
rect 13997 21858 14063 21861
rect 13632 21856 14063 21858
rect 13632 21800 14002 21856
rect 14058 21800 14063 21856
rect 13632 21798 14063 21800
rect 13997 21795 14063 21798
rect 16941 21858 17007 21861
rect 20478 21858 20484 21860
rect 16941 21856 20484 21858
rect 16941 21800 16946 21856
rect 17002 21800 20484 21856
rect 16941 21798 20484 21800
rect 16941 21795 17007 21798
rect 20478 21796 20484 21798
rect 20548 21796 20554 21860
rect 23197 21858 23263 21861
rect 23841 21858 23907 21861
rect 27520 21858 28000 21888
rect 23197 21856 23907 21858
rect 23197 21800 23202 21856
rect 23258 21800 23846 21856
rect 23902 21800 23907 21856
rect 23197 21798 23907 21800
rect 23197 21795 23263 21798
rect 23841 21795 23907 21798
rect 25822 21798 28000 21858
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 11053 21722 11119 21725
rect 6134 21720 11119 21722
rect 6134 21664 11058 21720
rect 11114 21664 11119 21720
rect 6134 21662 11119 21664
rect 3417 21586 3483 21589
rect 4245 21586 4311 21589
rect 6134 21586 6194 21662
rect 11053 21659 11119 21662
rect 11421 21722 11487 21725
rect 16389 21722 16455 21725
rect 18597 21722 18663 21725
rect 11421 21720 14842 21722
rect 11421 21664 11426 21720
rect 11482 21664 14842 21720
rect 11421 21662 14842 21664
rect 11421 21659 11487 21662
rect 3417 21584 6194 21586
rect 3417 21528 3422 21584
rect 3478 21528 4250 21584
rect 4306 21528 6194 21584
rect 3417 21526 6194 21528
rect 6361 21586 6427 21589
rect 8661 21586 8727 21589
rect 6361 21584 8727 21586
rect 6361 21528 6366 21584
rect 6422 21528 8666 21584
rect 8722 21528 8727 21584
rect 6361 21526 8727 21528
rect 3417 21523 3483 21526
rect 4245 21523 4311 21526
rect 6361 21523 6427 21526
rect 8661 21523 8727 21526
rect 9029 21586 9095 21589
rect 12709 21586 12775 21589
rect 9029 21584 12775 21586
rect 9029 21528 9034 21584
rect 9090 21528 12714 21584
rect 12770 21528 12775 21584
rect 9029 21526 12775 21528
rect 14782 21586 14842 21662
rect 16389 21720 18663 21722
rect 16389 21664 16394 21720
rect 16450 21664 18602 21720
rect 18658 21664 18663 21720
rect 16389 21662 18663 21664
rect 16389 21659 16455 21662
rect 18597 21659 18663 21662
rect 18965 21722 19031 21725
rect 22185 21722 22251 21725
rect 18965 21720 22251 21722
rect 18965 21664 18970 21720
rect 19026 21664 22190 21720
rect 22246 21664 22251 21720
rect 18965 21662 22251 21664
rect 18965 21659 19031 21662
rect 22185 21659 22251 21662
rect 23657 21722 23723 21725
rect 23657 21720 24042 21722
rect 23657 21664 23662 21720
rect 23718 21664 24042 21720
rect 23657 21662 24042 21664
rect 23657 21659 23723 21662
rect 20713 21586 20779 21589
rect 14782 21584 20779 21586
rect 14782 21528 20718 21584
rect 20774 21528 20779 21584
rect 14782 21526 20779 21528
rect 23982 21586 24042 21662
rect 25681 21586 25747 21589
rect 23982 21584 25747 21586
rect 23982 21528 25686 21584
rect 25742 21528 25747 21584
rect 23982 21526 25747 21528
rect 9029 21523 9095 21526
rect 12709 21523 12775 21526
rect 20713 21523 20779 21526
rect 25681 21523 25747 21526
rect 1853 21450 1919 21453
rect 2957 21450 3023 21453
rect 7465 21450 7531 21453
rect 1853 21448 7531 21450
rect 1853 21392 1858 21448
rect 1914 21392 2962 21448
rect 3018 21392 7470 21448
rect 7526 21392 7531 21448
rect 1853 21390 7531 21392
rect 1853 21387 1919 21390
rect 2957 21387 3023 21390
rect 7465 21387 7531 21390
rect 8569 21450 8635 21453
rect 10685 21450 10751 21453
rect 11421 21450 11487 21453
rect 8569 21448 11487 21450
rect 8569 21392 8574 21448
rect 8630 21392 10690 21448
rect 10746 21392 11426 21448
rect 11482 21392 11487 21448
rect 8569 21390 11487 21392
rect 8569 21387 8635 21390
rect 10685 21387 10751 21390
rect 11421 21387 11487 21390
rect 12341 21450 12407 21453
rect 18505 21450 18571 21453
rect 12341 21448 18571 21450
rect 12341 21392 12346 21448
rect 12402 21392 18510 21448
rect 18566 21392 18571 21448
rect 12341 21390 18571 21392
rect 12341 21387 12407 21390
rect 18505 21387 18571 21390
rect 19374 21388 19380 21452
rect 19444 21450 19450 21452
rect 19517 21450 19583 21453
rect 20897 21452 20963 21453
rect 20846 21450 20852 21452
rect 19444 21448 19583 21450
rect 19444 21392 19522 21448
rect 19578 21392 19583 21448
rect 19444 21390 19583 21392
rect 20806 21390 20852 21450
rect 20916 21448 20963 21452
rect 20958 21392 20963 21448
rect 19444 21388 19450 21390
rect 19517 21387 19583 21390
rect 20846 21388 20852 21390
rect 20916 21388 20963 21392
rect 20897 21387 20963 21388
rect 23013 21450 23079 21453
rect 25822 21450 25882 21798
rect 27520 21768 28000 21798
rect 23013 21448 25882 21450
rect 23013 21392 23018 21448
rect 23074 21392 25882 21448
rect 23013 21390 25882 21392
rect 23013 21387 23079 21390
rect 0 21314 480 21344
rect 4061 21314 4127 21317
rect 0 21312 4127 21314
rect 0 21256 4066 21312
rect 4122 21256 4127 21312
rect 0 21254 4127 21256
rect 0 21224 480 21254
rect 4061 21251 4127 21254
rect 11697 21314 11763 21317
rect 16205 21314 16271 21317
rect 18597 21314 18663 21317
rect 11697 21312 18663 21314
rect 11697 21256 11702 21312
rect 11758 21256 16210 21312
rect 16266 21256 18602 21312
rect 18658 21256 18663 21312
rect 11697 21254 18663 21256
rect 11697 21251 11763 21254
rect 16205 21251 16271 21254
rect 18597 21251 18663 21254
rect 20069 21314 20135 21317
rect 27520 21314 28000 21344
rect 20069 21312 28000 21314
rect 20069 21256 20074 21312
rect 20130 21256 28000 21312
rect 20069 21254 28000 21256
rect 20069 21251 20135 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 27520 21224 28000 21254
rect 19610 21183 19930 21184
rect 2405 21178 2471 21181
rect 4797 21178 4863 21181
rect 2405 21176 4863 21178
rect 2405 21120 2410 21176
rect 2466 21120 4802 21176
rect 4858 21120 4863 21176
rect 2405 21118 4863 21120
rect 2405 21115 2471 21118
rect 4797 21115 4863 21118
rect 11053 21178 11119 21181
rect 11237 21178 11303 21181
rect 11053 21176 11303 21178
rect 11053 21120 11058 21176
rect 11114 21120 11242 21176
rect 11298 21120 11303 21176
rect 11053 21118 11303 21120
rect 11053 21115 11119 21118
rect 11237 21115 11303 21118
rect 17166 21116 17172 21180
rect 17236 21178 17242 21180
rect 17493 21178 17559 21181
rect 19057 21178 19123 21181
rect 17236 21176 19123 21178
rect 17236 21120 17498 21176
rect 17554 21120 19062 21176
rect 19118 21120 19123 21176
rect 17236 21118 19123 21120
rect 17236 21116 17242 21118
rect 17493 21115 17559 21118
rect 19057 21115 19123 21118
rect 23657 21178 23723 21181
rect 25589 21178 25655 21181
rect 23657 21176 25655 21178
rect 23657 21120 23662 21176
rect 23718 21120 25594 21176
rect 25650 21120 25655 21176
rect 23657 21118 25655 21120
rect 23657 21115 23723 21118
rect 25589 21115 25655 21118
rect 2405 21042 2471 21045
rect 4245 21042 4311 21045
rect 12433 21042 12499 21045
rect 18045 21042 18111 21045
rect 22185 21042 22251 21045
rect 2405 21040 3066 21042
rect 2405 20984 2410 21040
rect 2466 20984 3066 21040
rect 2405 20982 3066 20984
rect 2405 20979 2471 20982
rect 3006 20906 3066 20982
rect 4245 21040 12499 21042
rect 4245 20984 4250 21040
rect 4306 20984 12438 21040
rect 12494 20984 12499 21040
rect 4245 20982 12499 20984
rect 4245 20979 4311 20982
rect 12433 20979 12499 20982
rect 14414 20982 17786 21042
rect 4981 20906 5047 20909
rect 8385 20906 8451 20909
rect 3006 20904 5047 20906
rect 3006 20848 4986 20904
rect 5042 20848 5047 20904
rect 3006 20846 5047 20848
rect 4981 20843 5047 20846
rect 5398 20904 8451 20906
rect 5398 20848 8390 20904
rect 8446 20848 8451 20904
rect 5398 20846 8451 20848
rect 0 20770 480 20800
rect 5398 20770 5458 20846
rect 8385 20843 8451 20846
rect 9029 20906 9095 20909
rect 11053 20906 11119 20909
rect 9029 20904 11119 20906
rect 9029 20848 9034 20904
rect 9090 20848 11058 20904
rect 11114 20848 11119 20904
rect 9029 20846 11119 20848
rect 9029 20843 9095 20846
rect 11053 20843 11119 20846
rect 12157 20906 12223 20909
rect 12801 20906 12867 20909
rect 14414 20906 14474 20982
rect 12157 20904 14474 20906
rect 12157 20848 12162 20904
rect 12218 20848 12806 20904
rect 12862 20848 14474 20904
rect 12157 20846 14474 20848
rect 17726 20906 17786 20982
rect 18045 21040 22251 21042
rect 18045 20984 18050 21040
rect 18106 20984 22190 21040
rect 22246 20984 22251 21040
rect 18045 20982 22251 20984
rect 18045 20979 18111 20982
rect 22185 20979 22251 20982
rect 19057 20906 19123 20909
rect 17726 20904 19123 20906
rect 17726 20848 19062 20904
rect 19118 20848 19123 20904
rect 17726 20846 19123 20848
rect 12157 20843 12223 20846
rect 12801 20843 12867 20846
rect 19057 20843 19123 20846
rect 20897 20906 20963 20909
rect 25221 20906 25287 20909
rect 20897 20904 25287 20906
rect 20897 20848 20902 20904
rect 20958 20848 25226 20904
rect 25282 20848 25287 20904
rect 20897 20846 25287 20848
rect 20897 20843 20963 20846
rect 25221 20843 25287 20846
rect 0 20710 5458 20770
rect 10869 20770 10935 20773
rect 12198 20770 12204 20772
rect 10869 20768 12204 20770
rect 10869 20712 10874 20768
rect 10930 20712 12204 20768
rect 10869 20710 12204 20712
rect 0 20680 480 20710
rect 10869 20707 10935 20710
rect 12198 20708 12204 20710
rect 12268 20708 12274 20772
rect 16941 20770 17007 20773
rect 19609 20770 19675 20773
rect 16941 20768 19675 20770
rect 16941 20712 16946 20768
rect 17002 20712 19614 20768
rect 19670 20712 19675 20768
rect 16941 20710 19675 20712
rect 16941 20707 17007 20710
rect 19609 20707 19675 20710
rect 26141 20770 26207 20773
rect 27520 20770 28000 20800
rect 26141 20768 28000 20770
rect 26141 20712 26146 20768
rect 26202 20712 28000 20768
rect 26141 20710 28000 20712
rect 26141 20707 26207 20710
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 27520 20680 28000 20710
rect 24277 20639 24597 20640
rect 8845 20634 8911 20637
rect 12433 20634 12499 20637
rect 8845 20632 12499 20634
rect 8845 20576 8850 20632
rect 8906 20576 12438 20632
rect 12494 20576 12499 20632
rect 8845 20574 12499 20576
rect 8845 20571 8911 20574
rect 12433 20571 12499 20574
rect 15561 20634 15627 20637
rect 18045 20634 18111 20637
rect 15561 20632 18111 20634
rect 15561 20576 15566 20632
rect 15622 20576 18050 20632
rect 18106 20576 18111 20632
rect 15561 20574 18111 20576
rect 15561 20571 15627 20574
rect 18045 20571 18111 20574
rect 22737 20634 22803 20637
rect 23473 20634 23539 20637
rect 22737 20632 23539 20634
rect 22737 20576 22742 20632
rect 22798 20576 23478 20632
rect 23534 20576 23539 20632
rect 22737 20574 23539 20576
rect 22737 20571 22803 20574
rect 23473 20571 23539 20574
rect 4061 20498 4127 20501
rect 7005 20498 7071 20501
rect 4061 20496 7071 20498
rect 4061 20440 4066 20496
rect 4122 20440 7010 20496
rect 7066 20440 7071 20496
rect 4061 20438 7071 20440
rect 4061 20435 4127 20438
rect 7005 20435 7071 20438
rect 13629 20498 13695 20501
rect 14181 20498 14247 20501
rect 13629 20496 14247 20498
rect 13629 20440 13634 20496
rect 13690 20440 14186 20496
rect 14242 20440 14247 20496
rect 13629 20438 14247 20440
rect 13629 20435 13695 20438
rect 14181 20435 14247 20438
rect 14457 20498 14523 20501
rect 20345 20498 20411 20501
rect 14457 20496 20411 20498
rect 14457 20440 14462 20496
rect 14518 20440 20350 20496
rect 20406 20440 20411 20496
rect 14457 20438 20411 20440
rect 14457 20435 14523 20438
rect 20345 20435 20411 20438
rect 20713 20498 20779 20501
rect 25957 20498 26023 20501
rect 20713 20496 26023 20498
rect 20713 20440 20718 20496
rect 20774 20440 25962 20496
rect 26018 20440 26023 20496
rect 20713 20438 26023 20440
rect 20713 20435 20779 20438
rect 25957 20435 26023 20438
rect 1669 20362 1735 20365
rect 6545 20362 6611 20365
rect 1669 20360 6611 20362
rect 1669 20304 1674 20360
rect 1730 20304 6550 20360
rect 6606 20304 6611 20360
rect 1669 20302 6611 20304
rect 1669 20299 1735 20302
rect 6545 20299 6611 20302
rect 9029 20362 9095 20365
rect 13905 20362 13971 20365
rect 21265 20362 21331 20365
rect 9029 20360 13971 20362
rect 9029 20304 9034 20360
rect 9090 20304 13910 20360
rect 13966 20304 13971 20360
rect 9029 20302 13971 20304
rect 9029 20299 9095 20302
rect 13905 20299 13971 20302
rect 19382 20360 21331 20362
rect 19382 20304 21270 20360
rect 21326 20304 21331 20360
rect 19382 20302 21331 20304
rect 1393 20226 1459 20229
rect 9857 20226 9923 20229
rect 1393 20224 9923 20226
rect 1393 20168 1398 20224
rect 1454 20168 9862 20224
rect 9918 20168 9923 20224
rect 1393 20166 9923 20168
rect 1393 20163 1459 20166
rect 9857 20163 9923 20166
rect 10777 20226 10843 20229
rect 12801 20226 12867 20229
rect 10777 20224 12867 20226
rect 10777 20168 10782 20224
rect 10838 20168 12806 20224
rect 12862 20168 12867 20224
rect 10777 20166 12867 20168
rect 10777 20163 10843 20166
rect 12801 20163 12867 20166
rect 12985 20226 13051 20229
rect 18965 20226 19031 20229
rect 12985 20224 19031 20226
rect 12985 20168 12990 20224
rect 13046 20168 18970 20224
rect 19026 20168 19031 20224
rect 12985 20166 19031 20168
rect 12985 20163 13051 20166
rect 18965 20163 19031 20166
rect 10277 20160 10597 20161
rect 0 20090 480 20120
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 2497 20090 2563 20093
rect 0 20088 2563 20090
rect 0 20032 2502 20088
rect 2558 20032 2563 20088
rect 0 20030 2563 20032
rect 0 20000 480 20030
rect 2497 20027 2563 20030
rect 3785 20090 3851 20093
rect 7557 20090 7623 20093
rect 9949 20092 10015 20093
rect 9949 20090 9996 20092
rect 3785 20088 7623 20090
rect 3785 20032 3790 20088
rect 3846 20032 7562 20088
rect 7618 20032 7623 20088
rect 3785 20030 7623 20032
rect 9904 20088 9996 20090
rect 9904 20032 9954 20088
rect 9904 20030 9996 20032
rect 3785 20027 3851 20030
rect 7557 20027 7623 20030
rect 9949 20028 9996 20030
rect 10060 20028 10066 20092
rect 11237 20090 11303 20093
rect 19382 20090 19442 20302
rect 21265 20299 21331 20302
rect 20345 20226 20411 20229
rect 24945 20226 25011 20229
rect 20345 20224 25011 20226
rect 20345 20168 20350 20224
rect 20406 20168 24950 20224
rect 25006 20168 25011 20224
rect 20345 20166 25011 20168
rect 20345 20163 20411 20166
rect 24945 20163 25011 20166
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 11237 20088 19442 20090
rect 11237 20032 11242 20088
rect 11298 20032 19442 20088
rect 11237 20030 19442 20032
rect 21909 20090 21975 20093
rect 24485 20090 24551 20093
rect 21909 20088 24551 20090
rect 21909 20032 21914 20088
rect 21970 20032 24490 20088
rect 24546 20032 24551 20088
rect 21909 20030 24551 20032
rect 9949 20027 10015 20028
rect 11237 20027 11303 20030
rect 21909 20027 21975 20030
rect 24485 20027 24551 20030
rect 25313 20090 25379 20093
rect 27520 20090 28000 20120
rect 25313 20088 28000 20090
rect 25313 20032 25318 20088
rect 25374 20032 28000 20088
rect 25313 20030 28000 20032
rect 25313 20027 25379 20030
rect 27520 20000 28000 20030
rect 3509 19954 3575 19957
rect 13537 19954 13603 19957
rect 3509 19952 13603 19954
rect 3509 19896 3514 19952
rect 3570 19896 13542 19952
rect 13598 19896 13603 19952
rect 3509 19894 13603 19896
rect 3509 19891 3575 19894
rect 13537 19891 13603 19894
rect 17493 19954 17559 19957
rect 19977 19954 20043 19957
rect 17493 19952 20043 19954
rect 17493 19896 17498 19952
rect 17554 19896 19982 19952
rect 20038 19896 20043 19952
rect 17493 19894 20043 19896
rect 17493 19891 17559 19894
rect 19977 19891 20043 19894
rect 2313 19818 2379 19821
rect 9489 19818 9555 19821
rect 17769 19818 17835 19821
rect 2313 19816 7666 19818
rect 2313 19760 2318 19816
rect 2374 19760 7666 19816
rect 2313 19758 7666 19760
rect 2313 19755 2379 19758
rect 3417 19682 3483 19685
rect 5441 19682 5507 19685
rect 3417 19680 5507 19682
rect 3417 19624 3422 19680
rect 3478 19624 5446 19680
rect 5502 19624 5507 19680
rect 3417 19622 5507 19624
rect 7606 19682 7666 19758
rect 9489 19816 17835 19818
rect 9489 19760 9494 19816
rect 9550 19760 17774 19816
rect 17830 19760 17835 19816
rect 9489 19758 17835 19760
rect 9489 19755 9555 19758
rect 17769 19755 17835 19758
rect 24025 19818 24091 19821
rect 26233 19818 26299 19821
rect 24025 19816 26299 19818
rect 24025 19760 24030 19816
rect 24086 19760 26238 19816
rect 26294 19760 26299 19816
rect 24025 19758 26299 19760
rect 24025 19755 24091 19758
rect 26233 19755 26299 19758
rect 14181 19682 14247 19685
rect 21357 19682 21423 19685
rect 7606 19680 14247 19682
rect 7606 19624 14186 19680
rect 14242 19624 14247 19680
rect 7606 19622 14247 19624
rect 3417 19619 3483 19622
rect 5441 19619 5507 19622
rect 14181 19619 14247 19622
rect 15334 19680 21423 19682
rect 15334 19624 21362 19680
rect 21418 19624 21423 19680
rect 15334 19622 21423 19624
rect 5610 19616 5930 19617
rect 0 19546 480 19576
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 3325 19546 3391 19549
rect 0 19544 3391 19546
rect 0 19488 3330 19544
rect 3386 19488 3391 19544
rect 0 19486 3391 19488
rect 0 19456 480 19486
rect 3325 19483 3391 19486
rect 4061 19546 4127 19549
rect 5073 19546 5139 19549
rect 4061 19544 5139 19546
rect 4061 19488 4066 19544
rect 4122 19488 5078 19544
rect 5134 19488 5139 19544
rect 4061 19486 5139 19488
rect 4061 19483 4127 19486
rect 5073 19483 5139 19486
rect 6637 19546 6703 19549
rect 11053 19546 11119 19549
rect 11513 19546 11579 19549
rect 6637 19544 11579 19546
rect 6637 19488 6642 19544
rect 6698 19488 11058 19544
rect 11114 19488 11518 19544
rect 11574 19488 11579 19544
rect 6637 19486 11579 19488
rect 6637 19483 6703 19486
rect 11053 19483 11119 19486
rect 11513 19483 11579 19486
rect 2313 19410 2379 19413
rect 3785 19410 3851 19413
rect 2313 19408 3851 19410
rect 2313 19352 2318 19408
rect 2374 19352 3790 19408
rect 3846 19352 3851 19408
rect 2313 19350 3851 19352
rect 2313 19347 2379 19350
rect 3785 19347 3851 19350
rect 4061 19410 4127 19413
rect 8661 19410 8727 19413
rect 13353 19410 13419 19413
rect 15334 19410 15394 19622
rect 21357 19619 21423 19622
rect 24669 19682 24735 19685
rect 24894 19682 24900 19684
rect 24669 19680 24900 19682
rect 24669 19624 24674 19680
rect 24730 19624 24900 19680
rect 24669 19622 24900 19624
rect 24669 19619 24735 19622
rect 24894 19620 24900 19622
rect 24964 19620 24970 19684
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 18270 19484 18276 19548
rect 18340 19546 18346 19548
rect 18505 19546 18571 19549
rect 18340 19544 18571 19546
rect 18340 19488 18510 19544
rect 18566 19488 18571 19544
rect 18340 19486 18571 19488
rect 18340 19484 18346 19486
rect 18505 19483 18571 19486
rect 25078 19484 25084 19548
rect 25148 19546 25154 19548
rect 27520 19546 28000 19576
rect 25148 19486 28000 19546
rect 25148 19484 25154 19486
rect 27520 19456 28000 19486
rect 4061 19408 8727 19410
rect 4061 19352 4066 19408
rect 4122 19352 8666 19408
rect 8722 19352 8727 19408
rect 4061 19350 8727 19352
rect 4061 19347 4127 19350
rect 8661 19347 8727 19350
rect 9998 19350 11530 19410
rect 2957 19274 3023 19277
rect 6545 19274 6611 19277
rect 2957 19272 6611 19274
rect 2957 19216 2962 19272
rect 3018 19216 6550 19272
rect 6606 19216 6611 19272
rect 2957 19214 6611 19216
rect 2957 19211 3023 19214
rect 6545 19211 6611 19214
rect 8017 19274 8083 19277
rect 9998 19274 10058 19350
rect 8017 19272 9736 19274
rect 8017 19216 8022 19272
rect 8078 19240 9736 19272
rect 9860 19240 10058 19274
rect 8078 19216 10058 19240
rect 8017 19214 10058 19216
rect 10409 19274 10475 19277
rect 10910 19274 10916 19276
rect 10409 19272 10916 19274
rect 10409 19216 10414 19272
rect 10470 19216 10916 19272
rect 10409 19214 10916 19216
rect 8017 19211 8083 19214
rect 9676 19180 9920 19214
rect 10409 19211 10475 19214
rect 10910 19212 10916 19214
rect 10980 19212 10986 19276
rect 11470 19274 11530 19350
rect 13353 19408 15394 19410
rect 13353 19352 13358 19408
rect 13414 19352 15394 19408
rect 13353 19350 15394 19352
rect 17401 19410 17467 19413
rect 18321 19410 18387 19413
rect 23565 19410 23631 19413
rect 17401 19408 23631 19410
rect 17401 19352 17406 19408
rect 17462 19352 18326 19408
rect 18382 19352 23570 19408
rect 23626 19352 23631 19408
rect 17401 19350 23631 19352
rect 13353 19347 13419 19350
rect 17401 19347 17467 19350
rect 18321 19347 18387 19350
rect 23565 19347 23631 19350
rect 13537 19274 13603 19277
rect 11470 19272 13603 19274
rect 11470 19216 13542 19272
rect 13598 19216 13603 19272
rect 11470 19214 13603 19216
rect 13537 19211 13603 19214
rect 15101 19274 15167 19277
rect 18597 19274 18663 19277
rect 20897 19274 20963 19277
rect 15101 19272 20963 19274
rect 15101 19216 15106 19272
rect 15162 19216 18602 19272
rect 18658 19216 20902 19272
rect 20958 19216 20963 19272
rect 15101 19214 20963 19216
rect 15101 19211 15167 19214
rect 18597 19211 18663 19214
rect 20897 19211 20963 19214
rect 22001 19274 22067 19277
rect 22829 19274 22895 19277
rect 22001 19272 22895 19274
rect 22001 19216 22006 19272
rect 22062 19216 22834 19272
rect 22890 19216 22895 19272
rect 22001 19214 22895 19216
rect 22001 19211 22067 19214
rect 22829 19211 22895 19214
rect 11881 19140 11947 19141
rect 11830 19076 11836 19140
rect 11900 19138 11947 19140
rect 11900 19136 11992 19138
rect 11942 19080 11992 19136
rect 11900 19078 11992 19080
rect 11900 19076 11947 19078
rect 12934 19076 12940 19140
rect 13004 19138 13010 19140
rect 16665 19138 16731 19141
rect 13004 19136 16731 19138
rect 13004 19080 16670 19136
rect 16726 19080 16731 19136
rect 13004 19078 16731 19080
rect 13004 19076 13010 19078
rect 11881 19075 11947 19076
rect 16665 19075 16731 19078
rect 20161 19138 20227 19141
rect 25865 19138 25931 19141
rect 20161 19136 25931 19138
rect 20161 19080 20166 19136
rect 20222 19080 25870 19136
rect 25926 19080 25931 19136
rect 20161 19078 25931 19080
rect 20161 19075 20227 19078
rect 25865 19075 25931 19078
rect 10277 19072 10597 19073
rect 0 19002 480 19032
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 13813 19002 13879 19005
rect 18597 19002 18663 19005
rect 0 18942 4906 19002
rect 0 18912 480 18942
rect 4846 18866 4906 18942
rect 13813 19000 18663 19002
rect 13813 18944 13818 19000
rect 13874 18944 18602 19000
rect 18658 18944 18663 19000
rect 13813 18942 18663 18944
rect 13813 18939 13879 18942
rect 18597 18939 18663 18942
rect 21541 19002 21607 19005
rect 21909 19002 21975 19005
rect 27520 19002 28000 19032
rect 21541 19000 21975 19002
rect 21541 18944 21546 19000
rect 21602 18944 21914 19000
rect 21970 18944 21975 19000
rect 21541 18942 21975 18944
rect 21541 18939 21607 18942
rect 21909 18939 21975 18942
rect 23476 18942 28000 19002
rect 10777 18866 10843 18869
rect 4846 18864 10843 18866
rect 4846 18808 10782 18864
rect 10838 18808 10843 18864
rect 4846 18806 10843 18808
rect 10777 18803 10843 18806
rect 12801 18866 12867 18869
rect 16430 18866 16436 18868
rect 12801 18864 16436 18866
rect 12801 18808 12806 18864
rect 12862 18808 16436 18864
rect 12801 18806 16436 18808
rect 12801 18803 12867 18806
rect 16430 18804 16436 18806
rect 16500 18804 16506 18868
rect 17217 18866 17283 18869
rect 23476 18866 23536 18942
rect 27520 18912 28000 18942
rect 17217 18864 23536 18866
rect 17217 18808 17222 18864
rect 17278 18808 23536 18864
rect 17217 18806 23536 18808
rect 17217 18803 17283 18806
rect 23974 18804 23980 18868
rect 24044 18866 24050 18868
rect 24577 18866 24643 18869
rect 24044 18864 24643 18866
rect 24044 18808 24582 18864
rect 24638 18808 24643 18864
rect 24044 18806 24643 18808
rect 24044 18804 24050 18806
rect 24577 18803 24643 18806
rect 5165 18730 5231 18733
rect 11513 18730 11579 18733
rect 5165 18728 11579 18730
rect 5165 18672 5170 18728
rect 5226 18672 11518 18728
rect 11574 18672 11579 18728
rect 5165 18670 11579 18672
rect 5165 18667 5231 18670
rect 11513 18667 11579 18670
rect 12433 18730 12499 18733
rect 21541 18730 21607 18733
rect 12433 18728 21607 18730
rect 12433 18672 12438 18728
rect 12494 18672 21546 18728
rect 21602 18672 21607 18728
rect 12433 18670 21607 18672
rect 12433 18667 12499 18670
rect 21541 18667 21607 18670
rect 22870 18668 22876 18732
rect 22940 18730 22946 18732
rect 24301 18730 24367 18733
rect 22940 18728 24367 18730
rect 22940 18672 24306 18728
rect 24362 18672 24367 18728
rect 22940 18670 24367 18672
rect 22940 18668 22946 18670
rect 24301 18667 24367 18670
rect 2129 18594 2195 18597
rect 2630 18594 2636 18596
rect 2129 18592 2636 18594
rect 2129 18536 2134 18592
rect 2190 18536 2636 18592
rect 2129 18534 2636 18536
rect 2129 18531 2195 18534
rect 2630 18532 2636 18534
rect 2700 18532 2706 18596
rect 7833 18594 7899 18597
rect 11145 18594 11211 18597
rect 11697 18596 11763 18597
rect 11646 18594 11652 18596
rect 7833 18592 11211 18594
rect 7833 18536 7838 18592
rect 7894 18536 11150 18592
rect 11206 18536 11211 18592
rect 7833 18534 11211 18536
rect 11606 18534 11652 18594
rect 11716 18592 11763 18596
rect 11758 18536 11763 18592
rect 7833 18531 7899 18534
rect 11145 18531 11211 18534
rect 11646 18532 11652 18534
rect 11716 18532 11763 18536
rect 11697 18531 11763 18532
rect 15745 18594 15811 18597
rect 20161 18594 20227 18597
rect 22001 18594 22067 18597
rect 15745 18592 20227 18594
rect 15745 18536 15750 18592
rect 15806 18536 20166 18592
rect 20222 18536 20227 18592
rect 15745 18534 20227 18536
rect 15745 18531 15811 18534
rect 20161 18531 20227 18534
rect 20302 18592 22067 18594
rect 20302 18536 22006 18592
rect 22062 18536 22067 18592
rect 20302 18534 22067 18536
rect 5610 18528 5930 18529
rect 0 18458 480 18488
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 4061 18458 4127 18461
rect 0 18456 4127 18458
rect 0 18400 4066 18456
rect 4122 18400 4127 18456
rect 0 18398 4127 18400
rect 0 18368 480 18398
rect 4061 18395 4127 18398
rect 9305 18458 9371 18461
rect 13353 18458 13419 18461
rect 9305 18456 13419 18458
rect 9305 18400 9310 18456
rect 9366 18400 13358 18456
rect 13414 18400 13419 18456
rect 9305 18398 13419 18400
rect 9305 18395 9371 18398
rect 13353 18395 13419 18398
rect 18505 18458 18571 18461
rect 20302 18458 20362 18534
rect 22001 18531 22067 18534
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 18505 18456 20362 18458
rect 18505 18400 18510 18456
rect 18566 18400 20362 18456
rect 18505 18398 20362 18400
rect 20713 18458 20779 18461
rect 23933 18458 23999 18461
rect 27520 18458 28000 18488
rect 20713 18456 23999 18458
rect 20713 18400 20718 18456
rect 20774 18400 23938 18456
rect 23994 18400 23999 18456
rect 20713 18398 23999 18400
rect 18505 18395 18571 18398
rect 20713 18395 20779 18398
rect 23933 18395 23999 18398
rect 24902 18398 28000 18458
rect 5257 18322 5323 18325
rect 11697 18322 11763 18325
rect 5257 18320 11763 18322
rect 5257 18264 5262 18320
rect 5318 18264 11702 18320
rect 11758 18264 11763 18320
rect 5257 18262 11763 18264
rect 5257 18259 5323 18262
rect 11697 18259 11763 18262
rect 16849 18322 16915 18325
rect 22921 18322 22987 18325
rect 16849 18320 22987 18322
rect 16849 18264 16854 18320
rect 16910 18264 22926 18320
rect 22982 18264 22987 18320
rect 16849 18262 22987 18264
rect 16849 18259 16915 18262
rect 22921 18259 22987 18262
rect 4705 18186 4771 18189
rect 15653 18186 15719 18189
rect 4705 18184 15719 18186
rect 4705 18128 4710 18184
rect 4766 18128 15658 18184
rect 15714 18128 15719 18184
rect 4705 18126 15719 18128
rect 4705 18123 4771 18126
rect 15653 18123 15719 18126
rect 17493 18186 17559 18189
rect 20846 18186 20852 18188
rect 17493 18184 20852 18186
rect 17493 18128 17498 18184
rect 17554 18128 20852 18184
rect 17493 18126 20852 18128
rect 17493 18123 17559 18126
rect 20846 18124 20852 18126
rect 20916 18124 20922 18188
rect 21081 18186 21147 18189
rect 24902 18186 24962 18398
rect 27520 18368 28000 18398
rect 21081 18184 24962 18186
rect 21081 18128 21086 18184
rect 21142 18128 24962 18184
rect 21081 18126 24962 18128
rect 21081 18123 21147 18126
rect 3969 18050 4035 18053
rect 9121 18050 9187 18053
rect 3969 18048 9187 18050
rect 3969 17992 3974 18048
rect 4030 17992 9126 18048
rect 9182 17992 9187 18048
rect 3969 17990 9187 17992
rect 3969 17987 4035 17990
rect 9121 17987 9187 17990
rect 11145 18050 11211 18053
rect 16665 18050 16731 18053
rect 11145 18048 16731 18050
rect 11145 17992 11150 18048
rect 11206 17992 16670 18048
rect 16726 17992 16731 18048
rect 11145 17990 16731 17992
rect 11145 17987 11211 17990
rect 16665 17987 16731 17990
rect 21357 18050 21423 18053
rect 26233 18050 26299 18053
rect 21357 18048 23858 18050
rect 21357 17992 21362 18048
rect 21418 17992 23858 18048
rect 21357 17990 23858 17992
rect 21357 17987 21423 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 7833 17914 7899 17917
rect 4984 17912 7899 17914
rect 4984 17856 7838 17912
rect 7894 17856 7899 17912
rect 4984 17854 7899 17856
rect 0 17778 480 17808
rect 4984 17778 5044 17854
rect 7833 17851 7899 17854
rect 10869 17914 10935 17917
rect 11421 17914 11487 17917
rect 10869 17912 11487 17914
rect 10869 17856 10874 17912
rect 10930 17856 11426 17912
rect 11482 17856 11487 17912
rect 10869 17854 11487 17856
rect 10869 17851 10935 17854
rect 11421 17851 11487 17854
rect 12985 17914 13051 17917
rect 13118 17914 13124 17916
rect 12985 17912 13124 17914
rect 12985 17856 12990 17912
rect 13046 17856 13124 17912
rect 12985 17854 13124 17856
rect 12985 17851 13051 17854
rect 13118 17852 13124 17854
rect 13188 17852 13194 17916
rect 15285 17914 15351 17917
rect 19425 17914 19491 17917
rect 15285 17912 19491 17914
rect 15285 17856 15290 17912
rect 15346 17856 19430 17912
rect 19486 17856 19491 17912
rect 15285 17854 19491 17856
rect 15285 17851 15351 17854
rect 19425 17851 19491 17854
rect 20478 17852 20484 17916
rect 20548 17914 20554 17916
rect 22001 17914 22067 17917
rect 20548 17912 22067 17914
rect 20548 17856 22006 17912
rect 22062 17856 22067 17912
rect 20548 17854 22067 17856
rect 20548 17852 20554 17854
rect 22001 17851 22067 17854
rect 22461 17916 22527 17917
rect 22461 17912 22508 17916
rect 22572 17914 22578 17916
rect 23798 17914 23858 17990
rect 24304 18048 26299 18050
rect 24304 17992 26238 18048
rect 26294 17992 26299 18048
rect 24304 17990 26299 17992
rect 24304 17914 24364 17990
rect 26233 17987 26299 17990
rect 22461 17856 22466 17912
rect 22461 17852 22508 17856
rect 22572 17854 22618 17914
rect 23798 17854 24364 17914
rect 22572 17852 22578 17854
rect 22461 17851 22527 17852
rect 5165 17780 5231 17781
rect 5165 17778 5212 17780
rect 0 17718 5044 17778
rect 5120 17776 5212 17778
rect 5120 17720 5170 17776
rect 5120 17718 5212 17720
rect 0 17688 480 17718
rect 5165 17716 5212 17718
rect 5276 17716 5282 17780
rect 7005 17778 7071 17781
rect 10133 17778 10199 17781
rect 10726 17778 10732 17780
rect 7005 17776 9506 17778
rect 7005 17720 7010 17776
rect 7066 17720 9506 17776
rect 7005 17718 9506 17720
rect 5165 17715 5231 17716
rect 7005 17715 7071 17718
rect 1393 17642 1459 17645
rect 9305 17642 9371 17645
rect 1393 17640 9371 17642
rect 1393 17584 1398 17640
rect 1454 17584 9310 17640
rect 9366 17584 9371 17640
rect 1393 17582 9371 17584
rect 9446 17642 9506 17718
rect 10133 17776 10732 17778
rect 10133 17720 10138 17776
rect 10194 17720 10732 17776
rect 10133 17718 10732 17720
rect 10133 17715 10199 17718
rect 10726 17716 10732 17718
rect 10796 17716 10802 17780
rect 17401 17778 17467 17781
rect 20345 17778 20411 17781
rect 17401 17776 20411 17778
rect 17401 17720 17406 17776
rect 17462 17720 20350 17776
rect 20406 17720 20411 17776
rect 17401 17718 20411 17720
rect 17401 17715 17467 17718
rect 20345 17715 20411 17718
rect 20662 17716 20668 17780
rect 20732 17778 20738 17780
rect 27520 17778 28000 17808
rect 20732 17718 28000 17778
rect 20732 17716 20738 17718
rect 27520 17688 28000 17718
rect 12801 17642 12867 17645
rect 9446 17640 12867 17642
rect 9446 17584 12806 17640
rect 12862 17584 12867 17640
rect 9446 17582 12867 17584
rect 1393 17579 1459 17582
rect 9305 17579 9371 17582
rect 12801 17579 12867 17582
rect 13629 17642 13695 17645
rect 20989 17642 21055 17645
rect 13629 17640 21055 17642
rect 13629 17584 13634 17640
rect 13690 17584 20994 17640
rect 21050 17584 21055 17640
rect 13629 17582 21055 17584
rect 13629 17579 13695 17582
rect 20989 17579 21055 17582
rect 7189 17506 7255 17509
rect 7782 17506 7788 17508
rect 7189 17504 7788 17506
rect 7189 17448 7194 17504
rect 7250 17448 7788 17504
rect 7189 17446 7788 17448
rect 7189 17443 7255 17446
rect 7782 17444 7788 17446
rect 7852 17506 7858 17508
rect 14181 17506 14247 17509
rect 7852 17504 14247 17506
rect 7852 17448 14186 17504
rect 14242 17448 14247 17504
rect 7852 17446 14247 17448
rect 7852 17444 7858 17446
rect 14181 17443 14247 17446
rect 16481 17506 16547 17509
rect 21909 17506 21975 17509
rect 16481 17504 21975 17506
rect 16481 17448 16486 17504
rect 16542 17448 21914 17504
rect 21970 17448 21975 17504
rect 16481 17446 21975 17448
rect 16481 17443 16547 17446
rect 21909 17443 21975 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 8017 17370 8083 17373
rect 12249 17370 12315 17373
rect 8017 17368 12315 17370
rect 8017 17312 8022 17368
rect 8078 17312 12254 17368
rect 12310 17312 12315 17368
rect 8017 17310 12315 17312
rect 8017 17307 8083 17310
rect 12249 17307 12315 17310
rect 12801 17370 12867 17373
rect 13629 17372 13695 17373
rect 13629 17370 13676 17372
rect 12801 17368 13676 17370
rect 13740 17370 13746 17372
rect 16665 17370 16731 17373
rect 20161 17370 20227 17373
rect 12801 17312 12806 17368
rect 12862 17312 13634 17368
rect 12801 17310 13676 17312
rect 12801 17307 12867 17310
rect 13629 17308 13676 17310
rect 13740 17310 13822 17370
rect 16665 17368 20227 17370
rect 16665 17312 16670 17368
rect 16726 17312 20166 17368
rect 20222 17312 20227 17368
rect 16665 17310 20227 17312
rect 13740 17308 13746 17310
rect 13629 17307 13695 17308
rect 16665 17307 16731 17310
rect 20161 17307 20227 17310
rect 20345 17370 20411 17373
rect 23013 17370 23079 17373
rect 23289 17372 23355 17373
rect 20345 17368 23079 17370
rect 20345 17312 20350 17368
rect 20406 17312 23018 17368
rect 23074 17312 23079 17368
rect 20345 17310 23079 17312
rect 20345 17307 20411 17310
rect 23013 17307 23079 17310
rect 23238 17308 23244 17372
rect 23308 17370 23355 17372
rect 24761 17370 24827 17373
rect 25078 17370 25084 17372
rect 23308 17368 23400 17370
rect 23350 17312 23400 17368
rect 23308 17310 23400 17312
rect 24761 17368 25084 17370
rect 24761 17312 24766 17368
rect 24822 17312 25084 17368
rect 24761 17310 25084 17312
rect 23308 17308 23355 17310
rect 23289 17307 23355 17308
rect 24761 17307 24827 17310
rect 25078 17308 25084 17310
rect 25148 17308 25154 17372
rect 0 17234 480 17264
rect 3969 17234 4035 17237
rect 0 17232 4035 17234
rect 0 17176 3974 17232
rect 4030 17176 4035 17232
rect 0 17174 4035 17176
rect 0 17144 480 17174
rect 3969 17171 4035 17174
rect 4153 17234 4219 17237
rect 10409 17234 10475 17237
rect 15193 17234 15259 17237
rect 4153 17232 9506 17234
rect 4153 17176 4158 17232
rect 4214 17176 9506 17232
rect 4153 17174 9506 17176
rect 4153 17171 4219 17174
rect 3693 17098 3759 17101
rect 9213 17098 9279 17101
rect 3693 17096 9279 17098
rect 3693 17040 3698 17096
rect 3754 17040 9218 17096
rect 9274 17040 9279 17096
rect 3693 17038 9279 17040
rect 9446 17098 9506 17174
rect 10409 17232 15259 17234
rect 10409 17176 10414 17232
rect 10470 17176 15198 17232
rect 15254 17176 15259 17232
rect 10409 17174 15259 17176
rect 10409 17171 10475 17174
rect 15193 17171 15259 17174
rect 16021 17234 16087 17237
rect 18965 17234 19031 17237
rect 16021 17232 23306 17234
rect 16021 17176 16026 17232
rect 16082 17176 18970 17232
rect 19026 17176 23306 17232
rect 16021 17174 23306 17176
rect 16021 17171 16087 17174
rect 18965 17171 19031 17174
rect 12433 17098 12499 17101
rect 9446 17096 12499 17098
rect 9446 17040 12438 17096
rect 12494 17040 12499 17096
rect 9446 17038 12499 17040
rect 3693 17035 3759 17038
rect 9213 17035 9279 17038
rect 12433 17035 12499 17038
rect 14181 17098 14247 17101
rect 22553 17098 22619 17101
rect 14181 17096 22619 17098
rect 14181 17040 14186 17096
rect 14242 17040 22558 17096
rect 22614 17040 22619 17096
rect 14181 17038 22619 17040
rect 23246 17098 23306 17174
rect 23422 17172 23428 17236
rect 23492 17234 23498 17236
rect 23565 17234 23631 17237
rect 27520 17234 28000 17264
rect 23492 17232 23631 17234
rect 23492 17176 23570 17232
rect 23626 17176 23631 17232
rect 23492 17174 23631 17176
rect 23492 17172 23498 17174
rect 23565 17171 23631 17174
rect 24350 17174 28000 17234
rect 24209 17098 24275 17101
rect 23246 17096 24275 17098
rect 23246 17040 24214 17096
rect 24270 17040 24275 17096
rect 23246 17038 24275 17040
rect 14181 17035 14247 17038
rect 22553 17035 22619 17038
rect 24209 17035 24275 17038
rect 3509 16962 3575 16965
rect 6361 16962 6427 16965
rect 3509 16960 6427 16962
rect 3509 16904 3514 16960
rect 3570 16904 6366 16960
rect 6422 16904 6427 16960
rect 3509 16902 6427 16904
rect 3509 16899 3575 16902
rect 6361 16899 6427 16902
rect 13629 16962 13695 16965
rect 16614 16962 16620 16964
rect 13629 16960 16620 16962
rect 13629 16904 13634 16960
rect 13690 16904 16620 16960
rect 13629 16902 16620 16904
rect 13629 16899 13695 16902
rect 16614 16900 16620 16902
rect 16684 16900 16690 16964
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 4245 16826 4311 16829
rect 1350 16824 4311 16826
rect 1350 16768 4250 16824
rect 4306 16768 4311 16824
rect 1350 16766 4311 16768
rect 0 16690 480 16720
rect 1350 16690 1410 16766
rect 4245 16763 4311 16766
rect 4429 16826 4495 16829
rect 8385 16826 8451 16829
rect 9305 16826 9371 16829
rect 4429 16824 9371 16826
rect 4429 16768 4434 16824
rect 4490 16768 8390 16824
rect 8446 16768 9310 16824
rect 9366 16768 9371 16824
rect 4429 16766 9371 16768
rect 4429 16763 4495 16766
rect 8385 16763 8451 16766
rect 9305 16763 9371 16766
rect 10685 16826 10751 16829
rect 11329 16826 11395 16829
rect 19425 16826 19491 16829
rect 10685 16824 19491 16826
rect 10685 16768 10690 16824
rect 10746 16768 11334 16824
rect 11390 16768 19430 16824
rect 19486 16768 19491 16824
rect 10685 16766 19491 16768
rect 10685 16763 10751 16766
rect 11329 16763 11395 16766
rect 19425 16763 19491 16766
rect 22829 16826 22895 16829
rect 24350 16826 24410 17174
rect 27520 17144 28000 17174
rect 22829 16824 24410 16826
rect 22829 16768 22834 16824
rect 22890 16768 24410 16824
rect 22829 16766 24410 16768
rect 22829 16763 22895 16766
rect 0 16630 1410 16690
rect 1761 16690 1827 16693
rect 8293 16690 8359 16693
rect 1761 16688 8359 16690
rect 1761 16632 1766 16688
rect 1822 16632 8298 16688
rect 8354 16632 8359 16688
rect 1761 16630 8359 16632
rect 0 16600 480 16630
rect 1761 16627 1827 16630
rect 8293 16627 8359 16630
rect 8886 16628 8892 16692
rect 8956 16690 8962 16692
rect 9489 16690 9555 16693
rect 8956 16688 9555 16690
rect 8956 16632 9494 16688
rect 9550 16632 9555 16688
rect 8956 16630 9555 16632
rect 8956 16628 8962 16630
rect 9489 16627 9555 16630
rect 13486 16628 13492 16692
rect 13556 16690 13562 16692
rect 14365 16690 14431 16693
rect 13556 16688 14431 16690
rect 13556 16632 14370 16688
rect 14426 16632 14431 16688
rect 13556 16630 14431 16632
rect 13556 16628 13562 16630
rect 14365 16627 14431 16630
rect 17033 16690 17099 16693
rect 25221 16690 25287 16693
rect 17033 16688 25287 16690
rect 17033 16632 17038 16688
rect 17094 16632 25226 16688
rect 25282 16632 25287 16688
rect 17033 16630 25287 16632
rect 17033 16627 17099 16630
rect 25221 16627 25287 16630
rect 25405 16690 25471 16693
rect 27520 16690 28000 16720
rect 25405 16688 28000 16690
rect 25405 16632 25410 16688
rect 25466 16632 28000 16688
rect 25405 16630 28000 16632
rect 25405 16627 25471 16630
rect 27520 16600 28000 16630
rect 8518 16492 8524 16556
rect 8588 16554 8594 16556
rect 9673 16554 9739 16557
rect 8588 16552 9739 16554
rect 8588 16496 9678 16552
rect 9734 16496 9739 16552
rect 8588 16494 9739 16496
rect 8588 16492 8594 16494
rect 9673 16491 9739 16494
rect 14365 16554 14431 16557
rect 22185 16554 22251 16557
rect 14365 16552 22251 16554
rect 14365 16496 14370 16552
rect 14426 16496 22190 16552
rect 22246 16496 22251 16552
rect 14365 16494 22251 16496
rect 14365 16491 14431 16494
rect 22185 16491 22251 16494
rect 23013 16554 23079 16557
rect 24025 16554 24091 16557
rect 23013 16552 24091 16554
rect 23013 16496 23018 16552
rect 23074 16496 24030 16552
rect 24086 16496 24091 16552
rect 23013 16494 24091 16496
rect 23013 16491 23079 16494
rect 24025 16491 24091 16494
rect 6821 16418 6887 16421
rect 9673 16418 9739 16421
rect 6821 16416 9739 16418
rect 6821 16360 6826 16416
rect 6882 16360 9678 16416
rect 9734 16360 9739 16416
rect 6821 16358 9739 16360
rect 6821 16355 6887 16358
rect 9673 16355 9739 16358
rect 9990 16356 9996 16420
rect 10060 16418 10066 16420
rect 14089 16418 14155 16421
rect 10060 16416 14155 16418
rect 10060 16360 14094 16416
rect 14150 16360 14155 16416
rect 10060 16358 14155 16360
rect 10060 16356 10066 16358
rect 14089 16355 14155 16358
rect 19057 16418 19123 16421
rect 20621 16418 20687 16421
rect 19057 16416 20687 16418
rect 19057 16360 19062 16416
rect 19118 16360 20626 16416
rect 20682 16360 20687 16416
rect 19057 16358 20687 16360
rect 19057 16355 19123 16358
rect 20621 16355 20687 16358
rect 20854 16358 24042 16418
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 9213 16282 9279 16285
rect 12750 16282 12756 16284
rect 6686 16222 9138 16282
rect 1485 16148 1551 16149
rect 1485 16146 1532 16148
rect 1440 16144 1532 16146
rect 1440 16088 1490 16144
rect 1440 16086 1532 16088
rect 1485 16084 1532 16086
rect 1596 16084 1602 16148
rect 4981 16146 5047 16149
rect 6686 16146 6746 16222
rect 4981 16144 6746 16146
rect 4981 16088 4986 16144
rect 5042 16088 6746 16144
rect 4981 16086 6746 16088
rect 6821 16146 6887 16149
rect 9078 16146 9138 16222
rect 9213 16280 12756 16282
rect 9213 16224 9218 16280
rect 9274 16224 12756 16280
rect 9213 16222 12756 16224
rect 9213 16219 9279 16222
rect 12750 16220 12756 16222
rect 12820 16282 12826 16284
rect 14774 16282 14780 16284
rect 12820 16222 14780 16282
rect 12820 16220 12826 16222
rect 14774 16220 14780 16222
rect 14844 16220 14850 16284
rect 15929 16282 15995 16285
rect 20854 16282 20914 16358
rect 15929 16280 20914 16282
rect 15929 16224 15934 16280
rect 15990 16224 20914 16280
rect 15929 16222 20914 16224
rect 21173 16282 21239 16285
rect 23841 16282 23907 16285
rect 21173 16280 23907 16282
rect 21173 16224 21178 16280
rect 21234 16224 23846 16280
rect 23902 16224 23907 16280
rect 21173 16222 23907 16224
rect 15929 16219 15995 16222
rect 21173 16219 21239 16222
rect 23841 16219 23907 16222
rect 11421 16146 11487 16149
rect 6821 16144 7666 16146
rect 6821 16088 6826 16144
rect 6882 16088 7666 16144
rect 6821 16086 7666 16088
rect 9078 16144 11487 16146
rect 9078 16088 11426 16144
rect 11482 16088 11487 16144
rect 9078 16086 11487 16088
rect 1485 16083 1551 16084
rect 4981 16083 5047 16086
rect 6821 16083 6887 16086
rect 0 16010 480 16040
rect 3141 16010 3207 16013
rect 4705 16010 4771 16013
rect 7373 16010 7439 16013
rect 0 16008 3207 16010
rect 0 15952 3146 16008
rect 3202 15952 3207 16008
rect 0 15950 3207 15952
rect 0 15920 480 15950
rect 3141 15947 3207 15950
rect 4662 16008 7439 16010
rect 4662 15952 4710 16008
rect 4766 15952 7378 16008
rect 7434 15952 7439 16008
rect 4662 15950 7439 15952
rect 7606 16010 7666 16086
rect 11421 16083 11487 16086
rect 11605 16146 11671 16149
rect 14181 16146 14247 16149
rect 15377 16146 15443 16149
rect 23749 16146 23815 16149
rect 11605 16144 14106 16146
rect 11605 16088 11610 16144
rect 11666 16088 14106 16144
rect 11605 16086 14106 16088
rect 11605 16083 11671 16086
rect 9121 16010 9187 16013
rect 13813 16010 13879 16013
rect 7606 16008 13879 16010
rect 7606 15952 9126 16008
rect 9182 15952 13818 16008
rect 13874 15952 13879 16008
rect 7606 15950 13879 15952
rect 4662 15947 4771 15950
rect 7373 15947 7439 15950
rect 9121 15947 9187 15950
rect 13813 15947 13879 15950
rect 2681 15874 2747 15877
rect 4662 15874 4722 15947
rect 2681 15872 4722 15874
rect 2681 15816 2686 15872
rect 2742 15816 4722 15872
rect 2681 15814 4722 15816
rect 5165 15874 5231 15877
rect 8937 15874 9003 15877
rect 5165 15872 9003 15874
rect 5165 15816 5170 15872
rect 5226 15816 8942 15872
rect 8998 15816 9003 15872
rect 5165 15814 9003 15816
rect 2681 15811 2747 15814
rect 5165 15811 5231 15814
rect 8937 15811 9003 15814
rect 10685 15874 10751 15877
rect 12341 15874 12407 15877
rect 10685 15872 12407 15874
rect 10685 15816 10690 15872
rect 10746 15816 12346 15872
rect 12402 15816 12407 15872
rect 10685 15814 12407 15816
rect 14046 15874 14106 16086
rect 14181 16144 23815 16146
rect 14181 16088 14186 16144
rect 14242 16088 15382 16144
rect 15438 16088 23754 16144
rect 23810 16088 23815 16144
rect 14181 16086 23815 16088
rect 14181 16083 14247 16086
rect 15377 16083 15443 16086
rect 23749 16083 23815 16086
rect 17902 15948 17908 16012
rect 17972 16010 17978 16012
rect 18413 16010 18479 16013
rect 17972 16008 18479 16010
rect 17972 15952 18418 16008
rect 18474 15952 18479 16008
rect 17972 15950 18479 15952
rect 17972 15948 17978 15950
rect 18413 15947 18479 15950
rect 19977 16010 20043 16013
rect 20662 16010 20668 16012
rect 19977 16008 20668 16010
rect 19977 15952 19982 16008
rect 20038 15952 20668 16008
rect 19977 15950 20668 15952
rect 19977 15947 20043 15950
rect 20662 15948 20668 15950
rect 20732 15948 20738 16012
rect 23982 16010 24042 16358
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 24894 16220 24900 16284
rect 24964 16282 24970 16284
rect 25037 16282 25103 16285
rect 24964 16280 25103 16282
rect 24964 16224 25042 16280
rect 25098 16224 25103 16280
rect 24964 16222 25103 16224
rect 24964 16220 24970 16222
rect 25037 16219 25103 16222
rect 27520 16010 28000 16040
rect 23982 15950 28000 16010
rect 27520 15920 28000 15950
rect 23841 15874 23907 15877
rect 23974 15874 23980 15876
rect 14046 15814 17050 15874
rect 10685 15811 10751 15814
rect 12341 15811 12407 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 4705 15738 4771 15741
rect 8109 15738 8175 15741
rect 4705 15736 8175 15738
rect 4705 15680 4710 15736
rect 4766 15680 8114 15736
rect 8170 15680 8175 15736
rect 4705 15678 8175 15680
rect 4705 15675 4771 15678
rect 8109 15675 8175 15678
rect 5441 15602 5507 15605
rect 8293 15602 8359 15605
rect 9446 15604 9874 15636
rect 5441 15600 8359 15602
rect 5441 15544 5446 15600
rect 5502 15544 8298 15600
rect 8354 15544 8359 15600
rect 5441 15542 8359 15544
rect 5441 15539 5507 15542
rect 8293 15539 8359 15542
rect 9438 15540 9444 15604
rect 9508 15602 9874 15604
rect 12934 15602 12940 15604
rect 9508 15576 12940 15602
rect 9508 15540 9514 15576
rect 9814 15542 12940 15576
rect 12934 15540 12940 15542
rect 13004 15540 13010 15604
rect 16990 15602 17050 15814
rect 23841 15872 23980 15874
rect 23841 15816 23846 15872
rect 23902 15816 23980 15872
rect 23841 15814 23980 15816
rect 23841 15811 23907 15814
rect 23974 15812 23980 15814
rect 24044 15812 24050 15876
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 22553 15738 22619 15741
rect 23238 15738 23244 15740
rect 22553 15736 23244 15738
rect 22553 15680 22558 15736
rect 22614 15680 23244 15736
rect 22553 15678 23244 15680
rect 22553 15675 22619 15678
rect 23238 15676 23244 15678
rect 23308 15676 23314 15740
rect 23422 15676 23428 15740
rect 23492 15738 23498 15740
rect 23790 15738 23796 15740
rect 23492 15678 23796 15738
rect 23492 15676 23498 15678
rect 23790 15676 23796 15678
rect 23860 15676 23866 15740
rect 23565 15602 23631 15605
rect 16990 15600 23631 15602
rect 16990 15544 23570 15600
rect 23626 15544 23631 15600
rect 16990 15542 23631 15544
rect 23565 15539 23631 15542
rect 0 15466 480 15496
rect 16389 15466 16455 15469
rect 0 15464 16455 15466
rect 0 15408 16394 15464
rect 16450 15408 16455 15464
rect 0 15406 16455 15408
rect 0 15376 480 15406
rect 16389 15403 16455 15406
rect 17677 15466 17743 15469
rect 20621 15466 20687 15469
rect 17677 15464 20687 15466
rect 17677 15408 17682 15464
rect 17738 15408 20626 15464
rect 20682 15408 20687 15464
rect 17677 15406 20687 15408
rect 17677 15403 17743 15406
rect 20621 15403 20687 15406
rect 23974 15404 23980 15468
rect 24044 15466 24050 15468
rect 27520 15466 28000 15496
rect 24044 15406 28000 15466
rect 24044 15404 24050 15406
rect 27520 15376 28000 15406
rect 1945 15330 2011 15333
rect 2865 15330 2931 15333
rect 5441 15330 5507 15333
rect 6821 15332 6887 15333
rect 6821 15330 6868 15332
rect 1945 15328 2931 15330
rect 1945 15272 1950 15328
rect 2006 15272 2870 15328
rect 2926 15272 2931 15328
rect 1945 15270 2931 15272
rect 1945 15267 2011 15270
rect 2865 15267 2931 15270
rect 3006 15328 5507 15330
rect 3006 15272 5446 15328
rect 5502 15272 5507 15328
rect 3006 15270 5507 15272
rect 6776 15328 6868 15330
rect 6776 15272 6826 15328
rect 6776 15270 6868 15272
rect 2129 15194 2195 15197
rect 3006 15194 3066 15270
rect 5441 15267 5507 15270
rect 6821 15268 6868 15270
rect 6932 15268 6938 15332
rect 8753 15330 8819 15333
rect 12801 15330 12867 15333
rect 8753 15328 12867 15330
rect 8753 15272 8758 15328
rect 8814 15272 12806 15328
rect 12862 15272 12867 15328
rect 8753 15270 12867 15272
rect 6821 15267 6887 15268
rect 8753 15267 8819 15270
rect 12801 15267 12867 15270
rect 16021 15330 16087 15333
rect 16297 15332 16363 15333
rect 16246 15330 16252 15332
rect 16021 15328 16252 15330
rect 16316 15330 16363 15332
rect 17217 15330 17283 15333
rect 20069 15330 20135 15333
rect 16316 15328 16408 15330
rect 16021 15272 16026 15328
rect 16082 15272 16252 15328
rect 16358 15272 16408 15328
rect 16021 15270 16252 15272
rect 16021 15267 16087 15270
rect 16246 15268 16252 15270
rect 16316 15270 16408 15272
rect 17217 15328 20135 15330
rect 17217 15272 17222 15328
rect 17278 15272 20074 15328
rect 20130 15272 20135 15328
rect 17217 15270 20135 15272
rect 16316 15268 16363 15270
rect 16297 15267 16363 15268
rect 17217 15267 17283 15270
rect 20069 15267 20135 15270
rect 20805 15330 20871 15333
rect 24025 15330 24091 15333
rect 20805 15328 24091 15330
rect 20805 15272 20810 15328
rect 20866 15272 24030 15328
rect 24086 15272 24091 15328
rect 20805 15270 24091 15272
rect 20805 15267 20871 15270
rect 24025 15267 24091 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 2129 15192 3066 15194
rect 2129 15136 2134 15192
rect 2190 15136 3066 15192
rect 2129 15134 3066 15136
rect 6821 15194 6887 15197
rect 7281 15194 7347 15197
rect 6821 15192 7347 15194
rect 6821 15136 6826 15192
rect 6882 15136 7286 15192
rect 7342 15136 7347 15192
rect 6821 15134 7347 15136
rect 2129 15131 2195 15134
rect 6821 15131 6887 15134
rect 7281 15131 7347 15134
rect 20161 15194 20227 15197
rect 22277 15194 22343 15197
rect 23381 15194 23447 15197
rect 20161 15192 23447 15194
rect 20161 15136 20166 15192
rect 20222 15136 22282 15192
rect 22338 15136 23386 15192
rect 23442 15136 23447 15192
rect 20161 15134 23447 15136
rect 20161 15131 20227 15134
rect 22277 15131 22343 15134
rect 23381 15131 23447 15134
rect 5257 15058 5323 15061
rect 7649 15058 7715 15061
rect 9121 15058 9187 15061
rect 5257 15056 9187 15058
rect 5257 15000 5262 15056
rect 5318 15000 7654 15056
rect 7710 15000 9126 15056
rect 9182 15000 9187 15056
rect 5257 14998 9187 15000
rect 5257 14995 5323 14998
rect 7649 14995 7715 14998
rect 9121 14995 9187 14998
rect 14590 14996 14596 15060
rect 14660 15058 14666 15060
rect 18045 15058 18111 15061
rect 20897 15058 20963 15061
rect 24117 15058 24183 15061
rect 14660 15056 20730 15058
rect 14660 15000 18050 15056
rect 18106 15000 20730 15056
rect 14660 14998 20730 15000
rect 14660 14996 14666 14998
rect 18045 14995 18111 14998
rect 0 14922 480 14952
rect 8702 14922 8708 14924
rect 0 14862 8708 14922
rect 0 14832 480 14862
rect 8702 14860 8708 14862
rect 8772 14860 8778 14924
rect 9308 14922 9690 14956
rect 12525 14922 12591 14925
rect 9308 14920 12591 14922
rect 9308 14896 12530 14920
rect 1393 14786 1459 14789
rect 5073 14786 5139 14789
rect 1393 14784 5139 14786
rect 1393 14728 1398 14784
rect 1454 14728 5078 14784
rect 5134 14728 5139 14784
rect 1393 14726 5139 14728
rect 1393 14723 1459 14726
rect 5073 14723 5139 14726
rect 7281 14786 7347 14789
rect 9308 14786 9368 14896
rect 9630 14864 12530 14896
rect 12586 14864 12591 14920
rect 9630 14862 12591 14864
rect 12525 14859 12591 14862
rect 12985 14922 13051 14925
rect 13537 14922 13603 14925
rect 20437 14922 20503 14925
rect 12985 14920 20503 14922
rect 12985 14864 12990 14920
rect 13046 14864 13542 14920
rect 13598 14864 20442 14920
rect 20498 14864 20503 14920
rect 12985 14862 20503 14864
rect 12985 14859 13051 14862
rect 13537 14859 13603 14862
rect 20437 14859 20503 14862
rect 9990 14786 9996 14788
rect 7281 14784 9368 14786
rect 7281 14728 7286 14784
rect 7342 14728 9368 14784
rect 7281 14726 9368 14728
rect 9492 14726 9996 14786
rect 7281 14723 7347 14726
rect 1669 14650 1735 14653
rect 1894 14650 1900 14652
rect 1669 14648 1900 14650
rect 1669 14592 1674 14648
rect 1730 14592 1900 14648
rect 1669 14590 1900 14592
rect 1669 14587 1735 14590
rect 1894 14588 1900 14590
rect 1964 14588 1970 14652
rect 3417 14650 3483 14653
rect 8518 14650 8524 14652
rect 3417 14648 8524 14650
rect 3417 14592 3422 14648
rect 3478 14592 8524 14648
rect 3417 14590 8524 14592
rect 3417 14587 3483 14590
rect 8518 14588 8524 14590
rect 8588 14588 8594 14652
rect 8702 14588 8708 14652
rect 8772 14650 8778 14652
rect 9492 14650 9552 14726
rect 9990 14724 9996 14726
rect 10060 14724 10066 14788
rect 14089 14786 14155 14789
rect 14222 14786 14228 14788
rect 11976 14784 14228 14786
rect 11976 14728 14094 14784
rect 14150 14728 14228 14784
rect 11976 14726 14228 14728
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 8772 14590 9552 14650
rect 8772 14588 8778 14590
rect 8477 14514 8543 14517
rect 11789 14514 11855 14517
rect 8477 14512 11855 14514
rect 8477 14456 8482 14512
rect 8538 14456 11794 14512
rect 11850 14456 11855 14512
rect 8477 14454 11855 14456
rect 8477 14451 8543 14454
rect 11789 14451 11855 14454
rect 0 14378 480 14408
rect 6821 14378 6887 14381
rect 9673 14378 9739 14381
rect 0 14318 6746 14378
rect 0 14288 480 14318
rect 6686 14242 6746 14318
rect 6821 14376 9739 14378
rect 6821 14320 6826 14376
rect 6882 14320 9678 14376
rect 9734 14320 9739 14376
rect 6821 14318 9739 14320
rect 6821 14315 6887 14318
rect 9673 14315 9739 14318
rect 9806 14316 9812 14380
rect 9876 14378 9882 14380
rect 11976 14378 12036 14726
rect 14089 14723 14155 14726
rect 14222 14724 14228 14726
rect 14292 14724 14298 14788
rect 14774 14724 14780 14788
rect 14844 14786 14850 14788
rect 15285 14786 15351 14789
rect 14844 14784 15351 14786
rect 14844 14728 15290 14784
rect 15346 14728 15351 14784
rect 14844 14726 15351 14728
rect 20670 14786 20730 14998
rect 20897 15056 24183 15058
rect 20897 15000 20902 15056
rect 20958 15000 24122 15056
rect 24178 15000 24183 15056
rect 20897 14998 24183 15000
rect 20897 14995 20963 14998
rect 24117 14995 24183 14998
rect 24301 15058 24367 15061
rect 24301 15056 24962 15058
rect 24301 15000 24306 15056
rect 24362 15000 24962 15056
rect 24301 14998 24962 15000
rect 24301 14995 24367 14998
rect 21357 14922 21423 14925
rect 23013 14922 23079 14925
rect 21357 14920 23079 14922
rect 21357 14864 21362 14920
rect 21418 14864 23018 14920
rect 23074 14864 23079 14920
rect 21357 14862 23079 14864
rect 21357 14859 21423 14862
rect 23013 14859 23079 14862
rect 23974 14860 23980 14924
rect 24044 14922 24050 14924
rect 24710 14922 24716 14924
rect 24044 14862 24716 14922
rect 24044 14860 24050 14862
rect 24710 14860 24716 14862
rect 24780 14860 24786 14924
rect 24902 14922 24962 14998
rect 27520 14922 28000 14952
rect 24902 14862 28000 14922
rect 27520 14832 28000 14862
rect 20670 14726 24962 14786
rect 14844 14724 14850 14726
rect 15285 14723 15351 14726
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 20069 14650 20135 14653
rect 24761 14650 24827 14653
rect 20069 14648 24827 14650
rect 20069 14592 20074 14648
rect 20130 14592 24766 14648
rect 24822 14592 24827 14648
rect 20069 14590 24827 14592
rect 20069 14587 20135 14590
rect 24761 14587 24827 14590
rect 17677 14514 17743 14517
rect 21449 14514 21515 14517
rect 17677 14512 21515 14514
rect 17677 14456 17682 14512
rect 17738 14456 21454 14512
rect 21510 14456 21515 14512
rect 17677 14454 21515 14456
rect 17677 14451 17743 14454
rect 21449 14451 21515 14454
rect 23381 14514 23447 14517
rect 24577 14514 24643 14517
rect 23381 14512 24643 14514
rect 23381 14456 23386 14512
rect 23442 14456 24582 14512
rect 24638 14456 24643 14512
rect 23381 14454 24643 14456
rect 23381 14451 23447 14454
rect 24577 14451 24643 14454
rect 9876 14318 12036 14378
rect 14273 14378 14339 14381
rect 14406 14378 14412 14380
rect 14273 14376 14412 14378
rect 14273 14320 14278 14376
rect 14334 14320 14412 14376
rect 14273 14318 14412 14320
rect 9876 14316 9882 14318
rect 14273 14315 14339 14318
rect 14406 14316 14412 14318
rect 14476 14316 14482 14380
rect 16849 14378 16915 14381
rect 20989 14378 21055 14381
rect 16849 14376 21055 14378
rect 16849 14320 16854 14376
rect 16910 14320 20994 14376
rect 21050 14320 21055 14376
rect 16849 14318 21055 14320
rect 16849 14315 16915 14318
rect 20989 14315 21055 14318
rect 24117 14378 24183 14381
rect 24301 14378 24367 14381
rect 24117 14376 24367 14378
rect 24117 14320 24122 14376
rect 24178 14320 24306 14376
rect 24362 14320 24367 14376
rect 24117 14318 24367 14320
rect 24902 14378 24962 14726
rect 27520 14378 28000 14408
rect 24902 14318 28000 14378
rect 24117 14315 24183 14318
rect 24301 14315 24367 14318
rect 27520 14288 28000 14318
rect 10041 14242 10107 14245
rect 12433 14242 12499 14245
rect 6686 14182 9138 14242
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 1761 14106 1827 14109
rect 5257 14106 5323 14109
rect 7649 14106 7715 14109
rect 8937 14106 9003 14109
rect 1761 14104 5323 14106
rect 1761 14048 1766 14104
rect 1822 14048 5262 14104
rect 5318 14048 5323 14104
rect 1761 14046 5323 14048
rect 1761 14043 1827 14046
rect 5257 14043 5323 14046
rect 7606 14104 9003 14106
rect 7606 14048 7654 14104
rect 7710 14048 8942 14104
rect 8998 14048 9003 14104
rect 7606 14046 9003 14048
rect 9078 14106 9138 14182
rect 10041 14240 12499 14242
rect 10041 14184 10046 14240
rect 10102 14184 12438 14240
rect 12494 14184 12499 14240
rect 10041 14182 12499 14184
rect 10041 14179 10107 14182
rect 12433 14179 12499 14182
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 11513 14106 11579 14109
rect 11646 14106 11652 14108
rect 9078 14104 11652 14106
rect 9078 14048 11518 14104
rect 11574 14048 11652 14104
rect 9078 14046 11652 14048
rect 7606 14043 7715 14046
rect 8937 14043 9003 14046
rect 11513 14043 11579 14046
rect 11646 14044 11652 14046
rect 11716 14044 11722 14108
rect 19241 14106 19307 14109
rect 22093 14106 22159 14109
rect 19241 14104 22159 14106
rect 19241 14048 19246 14104
rect 19302 14048 22098 14104
rect 22154 14048 22159 14104
rect 19241 14046 22159 14048
rect 19241 14043 19307 14046
rect 22093 14043 22159 14046
rect 4705 13970 4771 13973
rect 7606 13970 7666 14043
rect 4705 13968 7666 13970
rect 4705 13912 4710 13968
rect 4766 13912 7666 13968
rect 4705 13910 7666 13912
rect 8937 13970 9003 13973
rect 12893 13970 12959 13973
rect 8937 13968 12959 13970
rect 8937 13912 8942 13968
rect 8998 13912 12898 13968
rect 12954 13912 12959 13968
rect 8937 13910 12959 13912
rect 4705 13907 4771 13910
rect 8937 13907 9003 13910
rect 12893 13907 12959 13910
rect 13261 13970 13327 13973
rect 17217 13970 17283 13973
rect 20713 13972 20779 13973
rect 13261 13968 17283 13970
rect 13261 13912 13266 13968
rect 13322 13912 17222 13968
rect 17278 13912 17283 13968
rect 13261 13910 17283 13912
rect 13261 13907 13327 13910
rect 17217 13907 17283 13910
rect 20662 13908 20668 13972
rect 20732 13970 20779 13972
rect 22277 13970 22343 13973
rect 25221 13970 25287 13973
rect 20732 13968 20824 13970
rect 20774 13912 20824 13968
rect 20732 13910 20824 13912
rect 22277 13968 25287 13970
rect 22277 13912 22282 13968
rect 22338 13912 25226 13968
rect 25282 13912 25287 13968
rect 22277 13910 25287 13912
rect 20732 13908 20779 13910
rect 20713 13907 20779 13908
rect 22277 13907 22343 13910
rect 25221 13907 25287 13910
rect 3509 13834 3575 13837
rect 7925 13834 7991 13837
rect 3509 13832 7991 13834
rect 3509 13776 3514 13832
rect 3570 13776 7930 13832
rect 7986 13776 7991 13832
rect 3509 13774 7991 13776
rect 3509 13771 3575 13774
rect 7925 13771 7991 13774
rect 8477 13834 8543 13837
rect 9438 13834 9444 13836
rect 8477 13832 9444 13834
rect 8477 13776 8482 13832
rect 8538 13776 9444 13832
rect 8477 13774 9444 13776
rect 8477 13771 8543 13774
rect 9438 13772 9444 13774
rect 9508 13772 9514 13836
rect 11329 13834 11395 13837
rect 13353 13834 13419 13837
rect 11329 13832 13419 13834
rect 11329 13776 11334 13832
rect 11390 13776 13358 13832
rect 13414 13776 13419 13832
rect 11329 13774 13419 13776
rect 11329 13771 11395 13774
rect 13353 13771 13419 13774
rect 13905 13834 13971 13837
rect 15193 13834 15259 13837
rect 13905 13832 15259 13834
rect 13905 13776 13910 13832
rect 13966 13776 15198 13832
rect 15254 13776 15259 13832
rect 13905 13774 15259 13776
rect 13905 13771 13971 13774
rect 15193 13771 15259 13774
rect 16297 13834 16363 13837
rect 16849 13834 16915 13837
rect 16297 13832 16915 13834
rect 16297 13776 16302 13832
rect 16358 13776 16854 13832
rect 16910 13776 16915 13832
rect 16297 13774 16915 13776
rect 16297 13771 16363 13774
rect 16849 13771 16915 13774
rect 17033 13834 17099 13837
rect 17350 13834 17356 13836
rect 17033 13832 17356 13834
rect 17033 13776 17038 13832
rect 17094 13776 17356 13832
rect 17033 13774 17356 13776
rect 17033 13771 17099 13774
rect 17350 13772 17356 13774
rect 17420 13772 17426 13836
rect 21725 13834 21791 13837
rect 22921 13834 22987 13837
rect 19382 13774 20178 13834
rect 0 13698 480 13728
rect 1117 13698 1183 13701
rect 0 13696 1183 13698
rect 0 13640 1122 13696
rect 1178 13640 1183 13696
rect 0 13638 1183 13640
rect 0 13608 480 13638
rect 1117 13635 1183 13638
rect 1853 13698 1919 13701
rect 5717 13698 5783 13701
rect 1853 13696 5783 13698
rect 1853 13640 1858 13696
rect 1914 13640 5722 13696
rect 5778 13640 5783 13696
rect 1853 13638 5783 13640
rect 1853 13635 1919 13638
rect 5717 13635 5783 13638
rect 6821 13698 6887 13701
rect 9213 13698 9279 13701
rect 6821 13696 9279 13698
rect 6821 13640 6826 13696
rect 6882 13640 9218 13696
rect 9274 13640 9279 13696
rect 6821 13638 9279 13640
rect 6821 13635 6887 13638
rect 9213 13635 9279 13638
rect 12157 13698 12223 13701
rect 12525 13698 12591 13701
rect 19382 13698 19442 13774
rect 12157 13696 19442 13698
rect 12157 13640 12162 13696
rect 12218 13640 12530 13696
rect 12586 13640 19442 13696
rect 12157 13638 19442 13640
rect 20118 13698 20178 13774
rect 21725 13832 22987 13834
rect 21725 13776 21730 13832
rect 21786 13776 22926 13832
rect 22982 13776 22987 13832
rect 21725 13774 22987 13776
rect 21725 13771 21791 13774
rect 22921 13771 22987 13774
rect 23013 13698 23079 13701
rect 24117 13698 24183 13701
rect 20118 13696 24183 13698
rect 20118 13640 23018 13696
rect 23074 13640 24122 13696
rect 24178 13640 24183 13696
rect 20118 13638 24183 13640
rect 12157 13635 12223 13638
rect 12525 13635 12591 13638
rect 23013 13635 23079 13638
rect 24117 13635 24183 13638
rect 25865 13698 25931 13701
rect 27520 13698 28000 13728
rect 25865 13696 28000 13698
rect 25865 13640 25870 13696
rect 25926 13640 28000 13696
rect 25865 13638 28000 13640
rect 25865 13635 25931 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 27520 13608 28000 13638
rect 19610 13567 19930 13568
rect 3601 13562 3667 13565
rect 6361 13562 6427 13565
rect 7373 13564 7439 13565
rect 7373 13562 7420 13564
rect 3601 13560 6427 13562
rect 3601 13504 3606 13560
rect 3662 13504 6366 13560
rect 6422 13504 6427 13560
rect 3601 13502 6427 13504
rect 7328 13560 7420 13562
rect 7328 13504 7378 13560
rect 7328 13502 7420 13504
rect 3601 13499 3667 13502
rect 6361 13499 6427 13502
rect 7373 13500 7420 13502
rect 7484 13500 7490 13564
rect 9254 13500 9260 13564
rect 9324 13562 9330 13564
rect 9990 13562 9996 13564
rect 9324 13502 9996 13562
rect 9324 13500 9330 13502
rect 9990 13500 9996 13502
rect 10060 13500 10066 13564
rect 15561 13562 15627 13565
rect 15561 13560 18522 13562
rect 15561 13504 15566 13560
rect 15622 13504 18522 13560
rect 15561 13502 18522 13504
rect 7373 13499 7439 13500
rect 15561 13499 15627 13502
rect 5533 13426 5599 13429
rect 11421 13426 11487 13429
rect 14590 13426 14596 13428
rect 5533 13424 11487 13426
rect 5533 13368 5538 13424
rect 5594 13368 11426 13424
rect 11482 13368 11487 13424
rect 5533 13366 11487 13368
rect 5533 13363 5599 13366
rect 11421 13363 11487 13366
rect 11700 13366 14596 13426
rect 11700 13293 11760 13366
rect 14590 13364 14596 13366
rect 14660 13364 14666 13428
rect 14733 13426 14799 13429
rect 18229 13426 18295 13429
rect 14733 13424 18295 13426
rect 14733 13368 14738 13424
rect 14794 13368 18234 13424
rect 18290 13368 18295 13424
rect 14733 13366 18295 13368
rect 18462 13426 18522 13502
rect 21030 13500 21036 13564
rect 21100 13562 21106 13564
rect 24710 13562 24716 13564
rect 21100 13502 24716 13562
rect 21100 13500 21106 13502
rect 24710 13500 24716 13502
rect 24780 13500 24786 13564
rect 23749 13426 23815 13429
rect 18462 13424 23815 13426
rect 18462 13368 23754 13424
rect 23810 13368 23815 13424
rect 18462 13366 23815 13368
rect 14733 13363 14799 13366
rect 18229 13363 18295 13366
rect 23749 13363 23815 13366
rect 23933 13426 23999 13429
rect 25957 13426 26023 13429
rect 23933 13424 26023 13426
rect 23933 13368 23938 13424
rect 23994 13368 25962 13424
rect 26018 13368 26023 13424
rect 23933 13366 26023 13368
rect 23933 13363 23999 13366
rect 25957 13363 26023 13366
rect 1894 13228 1900 13292
rect 1964 13290 1970 13292
rect 2037 13290 2103 13293
rect 1964 13288 2103 13290
rect 1964 13232 2042 13288
rect 2098 13232 2103 13288
rect 1964 13230 2103 13232
rect 1964 13228 1970 13230
rect 2037 13227 2103 13230
rect 3734 13228 3740 13292
rect 3804 13290 3810 13292
rect 4337 13290 4403 13293
rect 5901 13290 5967 13293
rect 3804 13288 5967 13290
rect 3804 13232 4342 13288
rect 4398 13232 5906 13288
rect 5962 13232 5967 13288
rect 3804 13230 5967 13232
rect 3804 13228 3810 13230
rect 4337 13227 4403 13230
rect 5901 13227 5967 13230
rect 6637 13290 6703 13293
rect 11697 13290 11763 13293
rect 6637 13288 11763 13290
rect 6637 13232 6642 13288
rect 6698 13232 11702 13288
rect 11758 13232 11763 13288
rect 6637 13230 11763 13232
rect 6637 13227 6703 13230
rect 11697 13227 11763 13230
rect 12390 13230 24962 13290
rect 0 13154 480 13184
rect 933 13154 999 13157
rect 3141 13154 3207 13157
rect 0 13152 3207 13154
rect 0 13096 938 13152
rect 994 13096 3146 13152
rect 3202 13096 3207 13152
rect 0 13094 3207 13096
rect 0 13064 480 13094
rect 933 13091 999 13094
rect 3141 13091 3207 13094
rect 9581 13154 9647 13157
rect 12390 13154 12450 13230
rect 12617 13156 12683 13157
rect 12566 13154 12572 13156
rect 9581 13152 12450 13154
rect 9581 13096 9586 13152
rect 9642 13096 12450 13152
rect 9581 13094 12450 13096
rect 12526 13094 12572 13154
rect 12636 13152 12683 13156
rect 12678 13096 12683 13152
rect 9581 13091 9647 13094
rect 12566 13092 12572 13094
rect 12636 13092 12683 13096
rect 12617 13091 12683 13092
rect 15929 13154 15995 13157
rect 17861 13154 17927 13157
rect 15929 13152 17927 13154
rect 15929 13096 15934 13152
rect 15990 13096 17866 13152
rect 17922 13096 17927 13152
rect 15929 13094 17927 13096
rect 15929 13091 15995 13094
rect 17861 13091 17927 13094
rect 18045 13154 18111 13157
rect 19333 13154 19399 13157
rect 18045 13152 19399 13154
rect 18045 13096 18050 13152
rect 18106 13096 19338 13152
rect 19394 13096 19399 13152
rect 18045 13094 19399 13096
rect 18045 13091 18111 13094
rect 19333 13091 19399 13094
rect 20662 13092 20668 13156
rect 20732 13154 20738 13156
rect 21817 13154 21883 13157
rect 23841 13154 23907 13157
rect 20732 13152 23907 13154
rect 20732 13096 21822 13152
rect 21878 13096 23846 13152
rect 23902 13096 23907 13152
rect 20732 13094 23907 13096
rect 24902 13154 24962 13230
rect 27520 13154 28000 13184
rect 24902 13094 28000 13154
rect 20732 13092 20738 13094
rect 21817 13091 21883 13094
rect 23841 13091 23907 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 27520 13064 28000 13094
rect 24277 13023 24597 13024
rect 10961 13020 11027 13021
rect 1526 12956 1532 13020
rect 1596 13018 1602 13020
rect 10910 13018 10916 13020
rect 1596 12958 4906 13018
rect 10834 12958 10916 13018
rect 10980 13018 11027 13020
rect 11697 13018 11763 13021
rect 10980 13016 11763 13018
rect 11022 12960 11702 13016
rect 11758 12960 11763 13016
rect 1596 12956 1602 12958
rect 1894 12684 1900 12748
rect 1964 12746 1970 12748
rect 2129 12746 2195 12749
rect 1964 12744 2195 12746
rect 1964 12688 2134 12744
rect 2190 12688 2195 12744
rect 1964 12686 2195 12688
rect 4846 12746 4906 12958
rect 10910 12956 10916 12958
rect 10980 12958 11763 12960
rect 10980 12956 11027 12958
rect 10961 12955 11027 12956
rect 11697 12955 11763 12958
rect 12709 13018 12775 13021
rect 13302 13018 13308 13020
rect 12709 13016 13308 13018
rect 12709 12960 12714 13016
rect 12770 12960 13308 13016
rect 12709 12958 13308 12960
rect 12709 12955 12775 12958
rect 13302 12956 13308 12958
rect 13372 12956 13378 13020
rect 17493 13018 17559 13021
rect 19517 13018 19583 13021
rect 21633 13018 21699 13021
rect 17493 13016 21699 13018
rect 17493 12960 17498 13016
rect 17554 12960 19522 13016
rect 19578 12960 21638 13016
rect 21694 12960 21699 13016
rect 17493 12958 21699 12960
rect 17493 12955 17559 12958
rect 19517 12955 19583 12958
rect 21633 12955 21699 12958
rect 8109 12882 8175 12885
rect 16205 12882 16271 12885
rect 8109 12880 16271 12882
rect 8109 12824 8114 12880
rect 8170 12824 16210 12880
rect 16266 12824 16271 12880
rect 8109 12822 16271 12824
rect 8109 12819 8175 12822
rect 16205 12819 16271 12822
rect 17861 12882 17927 12885
rect 20069 12882 20135 12885
rect 17861 12880 20135 12882
rect 17861 12824 17866 12880
rect 17922 12824 20074 12880
rect 20130 12824 20135 12880
rect 17861 12822 20135 12824
rect 17861 12819 17927 12822
rect 20069 12819 20135 12822
rect 20294 12820 20300 12884
rect 20364 12882 20370 12884
rect 25037 12882 25103 12885
rect 20364 12880 25103 12882
rect 20364 12824 25042 12880
rect 25098 12824 25103 12880
rect 20364 12822 25103 12824
rect 20364 12820 20370 12822
rect 25037 12819 25103 12822
rect 6085 12746 6151 12749
rect 4846 12744 6151 12746
rect 4846 12688 6090 12744
rect 6146 12688 6151 12744
rect 4846 12686 6151 12688
rect 1964 12684 1970 12686
rect 2129 12683 2195 12686
rect 6085 12683 6151 12686
rect 6637 12746 6703 12749
rect 8293 12746 8359 12749
rect 6637 12744 8359 12746
rect 6637 12688 6642 12744
rect 6698 12688 8298 12744
rect 8354 12688 8359 12744
rect 6637 12686 8359 12688
rect 6637 12683 6703 12686
rect 8293 12683 8359 12686
rect 8477 12746 8543 12749
rect 13261 12746 13327 12749
rect 8477 12744 13327 12746
rect 8477 12688 8482 12744
rect 8538 12688 13266 12744
rect 13322 12688 13327 12744
rect 8477 12686 13327 12688
rect 8477 12683 8543 12686
rect 13261 12683 13327 12686
rect 14089 12746 14155 12749
rect 15285 12746 15351 12749
rect 15878 12746 15884 12748
rect 14089 12744 14290 12746
rect 14089 12688 14094 12744
rect 14150 12688 14290 12744
rect 14089 12686 14290 12688
rect 14089 12683 14155 12686
rect 0 12610 480 12640
rect 3366 12610 3372 12612
rect 0 12550 3372 12610
rect 0 12520 480 12550
rect 3366 12548 3372 12550
rect 3436 12548 3442 12612
rect 4245 12610 4311 12613
rect 5073 12610 5139 12613
rect 8661 12610 8727 12613
rect 4245 12608 4538 12610
rect 4245 12552 4250 12608
rect 4306 12552 4538 12608
rect 4245 12550 4538 12552
rect 4245 12547 4311 12550
rect 4478 12474 4538 12550
rect 5073 12608 8727 12610
rect 5073 12552 5078 12608
rect 5134 12552 8666 12608
rect 8722 12552 8727 12608
rect 5073 12550 8727 12552
rect 5073 12547 5139 12550
rect 8661 12547 8727 12550
rect 9029 12610 9095 12613
rect 9254 12610 9260 12612
rect 9029 12608 9260 12610
rect 9029 12552 9034 12608
rect 9090 12552 9260 12608
rect 9029 12550 9260 12552
rect 9029 12547 9095 12550
rect 9254 12548 9260 12550
rect 9324 12548 9330 12612
rect 12617 12610 12683 12613
rect 12750 12610 12756 12612
rect 12617 12608 12756 12610
rect 12617 12552 12622 12608
rect 12678 12552 12756 12608
rect 12617 12550 12756 12552
rect 12617 12547 12683 12550
rect 12750 12548 12756 12550
rect 12820 12548 12826 12612
rect 13537 12608 13603 12613
rect 13537 12552 13542 12608
rect 13598 12552 13603 12608
rect 13537 12547 13603 12552
rect 13905 12610 13971 12613
rect 14089 12610 14155 12613
rect 13905 12608 14155 12610
rect 13905 12552 13910 12608
rect 13966 12552 14094 12608
rect 14150 12552 14155 12608
rect 13905 12550 14155 12552
rect 13905 12547 13971 12550
rect 14089 12547 14155 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 9806 12474 9812 12476
rect 4478 12414 9812 12474
rect 9806 12412 9812 12414
rect 9876 12412 9882 12476
rect 11697 12474 11763 12477
rect 13540 12474 13600 12547
rect 11697 12472 13600 12474
rect 11697 12416 11702 12472
rect 11758 12416 13600 12472
rect 11697 12414 13600 12416
rect 13905 12474 13971 12477
rect 14230 12474 14290 12686
rect 15285 12744 15884 12746
rect 15285 12688 15290 12744
rect 15346 12688 15884 12744
rect 15285 12686 15884 12688
rect 15285 12683 15351 12686
rect 15878 12684 15884 12686
rect 15948 12684 15954 12748
rect 17493 12746 17559 12749
rect 23565 12746 23631 12749
rect 17493 12744 23631 12746
rect 17493 12688 17498 12744
rect 17554 12688 23570 12744
rect 23626 12688 23631 12744
rect 17493 12686 23631 12688
rect 17493 12683 17559 12686
rect 23565 12683 23631 12686
rect 15326 12548 15332 12612
rect 15396 12610 15402 12612
rect 15878 12610 15884 12612
rect 15396 12550 15884 12610
rect 15396 12548 15402 12550
rect 15878 12548 15884 12550
rect 15948 12548 15954 12612
rect 24301 12610 24367 12613
rect 27520 12610 28000 12640
rect 24301 12608 28000 12610
rect 24301 12552 24306 12608
rect 24362 12552 28000 12608
rect 24301 12550 28000 12552
rect 24301 12547 24367 12550
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 27520 12520 28000 12550
rect 19610 12479 19930 12480
rect 13905 12472 14290 12474
rect 13905 12416 13910 12472
rect 13966 12416 14290 12472
rect 13905 12414 14290 12416
rect 11697 12411 11763 12414
rect 13905 12411 13971 12414
rect 16430 12412 16436 12476
rect 16500 12474 16506 12476
rect 16757 12474 16823 12477
rect 20805 12474 20871 12477
rect 16500 12472 16823 12474
rect 16500 12416 16762 12472
rect 16818 12416 16823 12472
rect 16500 12414 16823 12416
rect 16500 12412 16506 12414
rect 16757 12411 16823 12414
rect 20118 12472 20871 12474
rect 20118 12416 20810 12472
rect 20866 12416 20871 12472
rect 20118 12414 20871 12416
rect 1945 12340 2011 12341
rect 1894 12276 1900 12340
rect 1964 12338 2011 12340
rect 1964 12336 2056 12338
rect 2006 12280 2056 12336
rect 1964 12278 2056 12280
rect 1964 12276 2011 12278
rect 9622 12276 9628 12340
rect 9692 12338 9698 12340
rect 9857 12338 9923 12341
rect 9692 12336 9923 12338
rect 9692 12280 9862 12336
rect 9918 12280 9923 12336
rect 9692 12278 9923 12280
rect 9692 12276 9698 12278
rect 1945 12275 2011 12276
rect 9857 12275 9923 12278
rect 15929 12338 15995 12341
rect 18321 12338 18387 12341
rect 20118 12338 20178 12414
rect 20805 12411 20871 12414
rect 21030 12412 21036 12476
rect 21100 12474 21106 12476
rect 21909 12474 21975 12477
rect 23381 12474 23447 12477
rect 23565 12474 23631 12477
rect 21100 12472 22340 12474
rect 21100 12416 21914 12472
rect 21970 12416 22340 12472
rect 21100 12414 22340 12416
rect 21100 12412 21106 12414
rect 21909 12411 21975 12414
rect 22280 12341 22340 12414
rect 23381 12472 23631 12474
rect 23381 12416 23386 12472
rect 23442 12416 23570 12472
rect 23626 12416 23631 12472
rect 23381 12414 23631 12416
rect 23381 12411 23447 12414
rect 23565 12411 23631 12414
rect 24669 12474 24735 12477
rect 26049 12474 26115 12477
rect 24669 12472 26115 12474
rect 24669 12416 24674 12472
rect 24730 12416 26054 12472
rect 26110 12416 26115 12472
rect 24669 12414 26115 12416
rect 24669 12411 24735 12414
rect 26049 12411 26115 12414
rect 15929 12336 20178 12338
rect 15929 12280 15934 12336
rect 15990 12280 18326 12336
rect 18382 12280 20178 12336
rect 15929 12278 20178 12280
rect 22277 12336 22343 12341
rect 22277 12280 22282 12336
rect 22338 12280 22343 12336
rect 15929 12275 15995 12278
rect 18321 12275 18387 12278
rect 22277 12275 22343 12280
rect 23105 12338 23171 12341
rect 25037 12338 25103 12341
rect 23105 12336 25103 12338
rect 23105 12280 23110 12336
rect 23166 12280 25042 12336
rect 25098 12280 25103 12336
rect 23105 12278 25103 12280
rect 23105 12275 23171 12278
rect 25037 12275 25103 12278
rect 3785 12204 3851 12205
rect 3734 12140 3740 12204
rect 3804 12202 3851 12204
rect 5901 12202 5967 12205
rect 6494 12202 6500 12204
rect 3804 12200 3896 12202
rect 3846 12144 3896 12200
rect 3804 12142 3896 12144
rect 5901 12200 6500 12202
rect 5901 12144 5906 12200
rect 5962 12144 6500 12200
rect 5901 12142 6500 12144
rect 3804 12140 3851 12142
rect 3785 12139 3851 12140
rect 5901 12139 5967 12142
rect 6494 12140 6500 12142
rect 6564 12140 6570 12204
rect 11421 12202 11487 12205
rect 9584 12200 11487 12202
rect 9584 12144 11426 12200
rect 11482 12144 11487 12200
rect 9584 12142 11487 12144
rect 9584 12100 9644 12142
rect 11421 12139 11487 12142
rect 11881 12202 11947 12205
rect 13486 12202 13492 12204
rect 11881 12200 13492 12202
rect 11881 12144 11886 12200
rect 11942 12144 13492 12200
rect 11881 12142 13492 12144
rect 11881 12139 11947 12142
rect 13486 12140 13492 12142
rect 13556 12140 13562 12204
rect 16941 12202 17007 12205
rect 14782 12200 17007 12202
rect 14782 12144 16946 12200
rect 17002 12144 17007 12200
rect 14782 12142 17007 12144
rect 6729 12066 6795 12069
rect 6862 12066 6868 12068
rect 6729 12064 6868 12066
rect 6729 12008 6734 12064
rect 6790 12008 6868 12064
rect 6729 12006 6868 12008
rect 6729 12003 6795 12006
rect 6862 12004 6868 12006
rect 6932 12004 6938 12068
rect 9492 12066 9644 12100
rect 7054 12040 9644 12066
rect 13721 12066 13787 12069
rect 14782 12066 14842 12142
rect 16941 12139 17007 12142
rect 21081 12202 21147 12205
rect 25129 12202 25195 12205
rect 21081 12200 25195 12202
rect 21081 12144 21086 12200
rect 21142 12144 25134 12200
rect 25190 12144 25195 12200
rect 21081 12142 25195 12144
rect 21081 12139 21147 12142
rect 25129 12139 25195 12142
rect 23289 12066 23355 12069
rect 13721 12064 14842 12066
rect 7054 12006 9552 12040
rect 13721 12008 13726 12064
rect 13782 12008 14842 12064
rect 13721 12006 14842 12008
rect 15334 12064 23355 12066
rect 15334 12008 23294 12064
rect 23350 12008 23355 12064
rect 15334 12006 23355 12008
rect 5610 12000 5930 12001
rect 0 11930 480 11960
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 4797 11930 4863 11933
rect 0 11928 4863 11930
rect 0 11872 4802 11928
rect 4858 11872 4863 11928
rect 0 11870 4863 11872
rect 0 11840 480 11870
rect 4797 11867 4863 11870
rect 6177 11930 6243 11933
rect 7054 11930 7114 12006
rect 13721 12003 13787 12006
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 6177 11928 7114 11930
rect 6177 11872 6182 11928
rect 6238 11872 7114 11928
rect 6177 11870 7114 11872
rect 7281 11930 7347 11933
rect 9673 11930 9739 11933
rect 7281 11928 13876 11930
rect 7281 11872 7286 11928
rect 7342 11872 9678 11928
rect 9734 11872 13876 11928
rect 7281 11870 13876 11872
rect 6177 11867 6243 11870
rect 7281 11867 7347 11870
rect 9673 11867 9739 11870
rect 3417 11794 3483 11797
rect 7782 11794 7788 11796
rect 3417 11792 7788 11794
rect 3417 11736 3422 11792
rect 3478 11736 7788 11792
rect 3417 11734 7788 11736
rect 3417 11731 3483 11734
rect 7782 11732 7788 11734
rect 7852 11732 7858 11796
rect 8201 11794 8267 11797
rect 11973 11794 12039 11797
rect 8201 11792 12039 11794
rect 8201 11736 8206 11792
rect 8262 11736 11978 11792
rect 12034 11736 12039 11792
rect 8201 11734 12039 11736
rect 8201 11731 8267 11734
rect 11973 11731 12039 11734
rect 13118 11732 13124 11796
rect 13188 11794 13194 11796
rect 13629 11794 13695 11797
rect 13188 11792 13695 11794
rect 13188 11736 13634 11792
rect 13690 11736 13695 11792
rect 13188 11734 13695 11736
rect 13816 11794 13876 11870
rect 15334 11794 15394 12006
rect 23289 12003 23355 12006
rect 24669 12066 24735 12069
rect 24894 12066 24900 12068
rect 24669 12064 24900 12066
rect 24669 12008 24674 12064
rect 24730 12008 24900 12064
rect 24669 12006 24900 12008
rect 24669 12003 24735 12006
rect 24894 12004 24900 12006
rect 24964 12004 24970 12068
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 16389 11930 16455 11933
rect 18965 11930 19031 11933
rect 27520 11930 28000 11960
rect 16389 11928 19031 11930
rect 16389 11872 16394 11928
rect 16450 11872 18970 11928
rect 19026 11872 19031 11928
rect 16389 11870 19031 11872
rect 16389 11867 16455 11870
rect 18965 11867 19031 11870
rect 24902 11870 28000 11930
rect 13816 11734 15394 11794
rect 16665 11794 16731 11797
rect 18965 11794 19031 11797
rect 19149 11794 19215 11797
rect 16665 11792 19215 11794
rect 16665 11736 16670 11792
rect 16726 11736 18970 11792
rect 19026 11736 19154 11792
rect 19210 11736 19215 11792
rect 16665 11734 19215 11736
rect 13188 11732 13194 11734
rect 13629 11731 13695 11734
rect 16665 11731 16731 11734
rect 18965 11731 19031 11734
rect 19149 11731 19215 11734
rect 19977 11794 20043 11797
rect 24902 11794 24962 11870
rect 27520 11840 28000 11870
rect 19977 11792 24962 11794
rect 19977 11736 19982 11792
rect 20038 11736 24962 11792
rect 19977 11734 24962 11736
rect 25221 11794 25287 11797
rect 25814 11794 25820 11796
rect 25221 11792 25820 11794
rect 25221 11736 25226 11792
rect 25282 11736 25820 11792
rect 25221 11734 25820 11736
rect 19977 11731 20043 11734
rect 25221 11731 25287 11734
rect 25814 11732 25820 11734
rect 25884 11732 25890 11796
rect 3233 11658 3299 11661
rect 5206 11658 5212 11660
rect 3233 11656 5212 11658
rect 3233 11600 3238 11656
rect 3294 11600 5212 11656
rect 3233 11598 5212 11600
rect 3233 11595 3299 11598
rect 5206 11596 5212 11598
rect 5276 11658 5282 11660
rect 6177 11658 6243 11661
rect 5276 11656 6243 11658
rect 5276 11600 6182 11656
rect 6238 11600 6243 11656
rect 5276 11598 6243 11600
rect 5276 11596 5282 11598
rect 6177 11595 6243 11598
rect 6862 11596 6868 11660
rect 6932 11658 6938 11660
rect 10317 11658 10383 11661
rect 11053 11658 11119 11661
rect 19241 11658 19307 11661
rect 20253 11658 20319 11661
rect 22369 11658 22435 11661
rect 6932 11656 19307 11658
rect 6932 11600 10322 11656
rect 10378 11600 11058 11656
rect 11114 11600 19246 11656
rect 19302 11600 19307 11656
rect 6932 11598 19307 11600
rect 6932 11596 6938 11598
rect 10317 11595 10383 11598
rect 11053 11595 11119 11598
rect 19241 11595 19307 11598
rect 19382 11598 20178 11658
rect 2221 11522 2287 11525
rect 8201 11522 8267 11525
rect 2221 11520 8267 11522
rect 2221 11464 2226 11520
rect 2282 11464 8206 11520
rect 8262 11464 8267 11520
rect 2221 11462 8267 11464
rect 2221 11459 2287 11462
rect 8201 11459 8267 11462
rect 17217 11522 17283 11525
rect 18873 11522 18939 11525
rect 19382 11522 19442 11598
rect 17217 11520 19442 11522
rect 17217 11464 17222 11520
rect 17278 11464 18878 11520
rect 18934 11464 19442 11520
rect 17217 11462 19442 11464
rect 17217 11459 17283 11462
rect 18873 11459 18939 11462
rect 10277 11456 10597 11457
rect 0 11386 480 11416
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 9673 11386 9739 11389
rect 0 11384 9739 11386
rect 0 11328 9678 11384
rect 9734 11328 9739 11384
rect 0 11326 9739 11328
rect 0 11296 480 11326
rect 9673 11323 9739 11326
rect 13486 11324 13492 11388
rect 13556 11386 13562 11388
rect 15561 11386 15627 11389
rect 13556 11384 15627 11386
rect 13556 11328 15566 11384
rect 15622 11328 15627 11384
rect 13556 11326 15627 11328
rect 13556 11324 13562 11326
rect 15561 11323 15627 11326
rect 5533 11250 5599 11253
rect 6494 11250 6500 11252
rect 5533 11248 6500 11250
rect 5533 11192 5538 11248
rect 5594 11192 6500 11248
rect 5533 11190 6500 11192
rect 5533 11187 5599 11190
rect 6494 11188 6500 11190
rect 6564 11188 6570 11252
rect 10777 11250 10843 11253
rect 13997 11250 14063 11253
rect 10777 11248 14063 11250
rect 10777 11192 10782 11248
rect 10838 11192 14002 11248
rect 14058 11192 14063 11248
rect 10777 11190 14063 11192
rect 10777 11187 10843 11190
rect 13997 11187 14063 11190
rect 14181 11250 14247 11253
rect 19885 11250 19951 11253
rect 14181 11248 19951 11250
rect 14181 11192 14186 11248
rect 14242 11192 19890 11248
rect 19946 11192 19951 11248
rect 14181 11190 19951 11192
rect 20118 11250 20178 11598
rect 20253 11656 22435 11658
rect 20253 11600 20258 11656
rect 20314 11600 22374 11656
rect 22430 11600 22435 11656
rect 20253 11598 22435 11600
rect 20253 11595 20319 11598
rect 22369 11595 22435 11598
rect 24710 11460 24716 11524
rect 24780 11522 24786 11524
rect 25681 11522 25747 11525
rect 24780 11520 26066 11522
rect 24780 11464 25686 11520
rect 25742 11464 26066 11520
rect 24780 11462 26066 11464
rect 24780 11460 24786 11462
rect 25681 11459 25747 11462
rect 22645 11386 22711 11389
rect 25773 11386 25839 11389
rect 22645 11384 25839 11386
rect 22645 11328 22650 11384
rect 22706 11328 25778 11384
rect 25834 11328 25839 11384
rect 22645 11326 25839 11328
rect 26006 11386 26066 11462
rect 27520 11386 28000 11416
rect 26006 11326 28000 11386
rect 22645 11323 22711 11326
rect 25773 11323 25839 11326
rect 27520 11296 28000 11326
rect 25221 11250 25287 11253
rect 20118 11248 25287 11250
rect 20118 11192 25226 11248
rect 25282 11192 25287 11248
rect 20118 11190 25287 11192
rect 14181 11187 14247 11190
rect 19885 11187 19951 11190
rect 25221 11187 25287 11190
rect 1393 11114 1459 11117
rect 10593 11114 10659 11117
rect 1393 11112 10659 11114
rect 1393 11056 1398 11112
rect 1454 11056 10598 11112
rect 10654 11056 10659 11112
rect 1393 11054 10659 11056
rect 1393 11051 1459 11054
rect 10593 11051 10659 11054
rect 17033 11114 17099 11117
rect 18689 11114 18755 11117
rect 17033 11112 18755 11114
rect 17033 11056 17038 11112
rect 17094 11056 18694 11112
rect 18750 11056 18755 11112
rect 17033 11054 18755 11056
rect 17033 11051 17099 11054
rect 18689 11051 18755 11054
rect 18873 11114 18939 11117
rect 23381 11114 23447 11117
rect 18873 11112 23447 11114
rect 18873 11056 18878 11112
rect 18934 11056 23386 11112
rect 23442 11056 23447 11112
rect 18873 11054 23447 11056
rect 18873 11051 18939 11054
rect 23381 11051 23447 11054
rect 23606 11052 23612 11116
rect 23676 11114 23682 11116
rect 23749 11114 23815 11117
rect 23676 11112 23815 11114
rect 23676 11056 23754 11112
rect 23810 11056 23815 11112
rect 23676 11054 23815 11056
rect 23676 11052 23682 11054
rect 23749 11051 23815 11054
rect 2865 10978 2931 10981
rect 4521 10978 4587 10981
rect 2865 10976 4587 10978
rect 2865 10920 2870 10976
rect 2926 10920 4526 10976
rect 4582 10920 4587 10976
rect 2865 10918 4587 10920
rect 2865 10915 2931 10918
rect 4521 10915 4587 10918
rect 9254 10916 9260 10980
rect 9324 10978 9330 10980
rect 12249 10978 12315 10981
rect 9324 10976 12315 10978
rect 9324 10920 12254 10976
rect 12310 10920 12315 10976
rect 9324 10918 12315 10920
rect 9324 10916 9330 10918
rect 12249 10915 12315 10918
rect 16430 10916 16436 10980
rect 16500 10978 16506 10980
rect 17677 10978 17743 10981
rect 16500 10976 17743 10978
rect 16500 10920 17682 10976
rect 17738 10920 17743 10976
rect 16500 10918 17743 10920
rect 16500 10916 16506 10918
rect 17677 10915 17743 10918
rect 19241 10978 19307 10981
rect 20713 10978 20779 10981
rect 19241 10976 20779 10978
rect 19241 10920 19246 10976
rect 19302 10920 20718 10976
rect 20774 10920 20779 10976
rect 19241 10918 20779 10920
rect 19241 10915 19307 10918
rect 20713 10915 20779 10918
rect 22502 10916 22508 10980
rect 22572 10978 22578 10980
rect 22829 10978 22895 10981
rect 22572 10976 22895 10978
rect 22572 10920 22834 10976
rect 22890 10920 22895 10976
rect 22572 10918 22895 10920
rect 22572 10916 22578 10918
rect 22829 10915 22895 10918
rect 5610 10912 5930 10913
rect 0 10842 480 10872
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 3049 10842 3115 10845
rect 0 10840 3115 10842
rect 0 10784 3054 10840
rect 3110 10784 3115 10840
rect 0 10782 3115 10784
rect 0 10752 480 10782
rect 3049 10779 3115 10782
rect 10225 10842 10291 10845
rect 13445 10842 13511 10845
rect 10225 10840 13511 10842
rect 10225 10784 10230 10840
rect 10286 10784 13450 10840
rect 13506 10784 13511 10840
rect 10225 10782 13511 10784
rect 10225 10779 10291 10782
rect 13445 10779 13511 10782
rect 16389 10842 16455 10845
rect 20897 10842 20963 10845
rect 16389 10840 20963 10842
rect 16389 10784 16394 10840
rect 16450 10784 20902 10840
rect 20958 10784 20963 10840
rect 16389 10782 20963 10784
rect 16389 10779 16455 10782
rect 20897 10779 20963 10782
rect 21173 10842 21239 10845
rect 23289 10842 23355 10845
rect 21173 10840 23355 10842
rect 21173 10784 21178 10840
rect 21234 10784 23294 10840
rect 23350 10784 23355 10840
rect 21173 10782 23355 10784
rect 21173 10779 21239 10782
rect 23289 10779 23355 10782
rect 24894 10780 24900 10844
rect 24964 10842 24970 10844
rect 26417 10842 26483 10845
rect 27520 10842 28000 10872
rect 24964 10840 28000 10842
rect 24964 10784 26422 10840
rect 26478 10784 28000 10840
rect 24964 10782 28000 10784
rect 24964 10780 24970 10782
rect 26417 10779 26483 10782
rect 27520 10752 28000 10782
rect 4061 10706 4127 10709
rect 5717 10706 5783 10709
rect 4061 10704 5783 10706
rect 4061 10648 4066 10704
rect 4122 10648 5722 10704
rect 5778 10648 5783 10704
rect 4061 10646 5783 10648
rect 4061 10643 4127 10646
rect 5717 10643 5783 10646
rect 11605 10706 11671 10709
rect 12566 10706 12572 10708
rect 11605 10704 12572 10706
rect 11605 10648 11610 10704
rect 11666 10648 12572 10704
rect 11605 10646 12572 10648
rect 11605 10643 11671 10646
rect 12566 10644 12572 10646
rect 12636 10706 12642 10708
rect 13486 10706 13492 10708
rect 12636 10646 13492 10706
rect 12636 10644 12642 10646
rect 13486 10644 13492 10646
rect 13556 10644 13562 10708
rect 20253 10706 20319 10709
rect 21265 10706 21331 10709
rect 20253 10704 21331 10706
rect 20253 10648 20258 10704
rect 20314 10648 21270 10704
rect 21326 10648 21331 10704
rect 20253 10646 21331 10648
rect 20253 10643 20319 10646
rect 21265 10643 21331 10646
rect 4889 10570 4955 10573
rect 9949 10570 10015 10573
rect 4889 10568 10015 10570
rect 4889 10512 4894 10568
rect 4950 10512 9954 10568
rect 10010 10512 10015 10568
rect 4889 10510 10015 10512
rect 4889 10507 4955 10510
rect 9949 10507 10015 10510
rect 23473 10570 23539 10573
rect 23473 10568 24778 10570
rect 23473 10512 23478 10568
rect 23534 10512 24778 10568
rect 23473 10510 24778 10512
rect 23473 10507 23539 10510
rect 3693 10434 3759 10437
rect 6678 10434 6684 10436
rect 3693 10432 6684 10434
rect 3693 10376 3698 10432
rect 3754 10376 6684 10432
rect 3693 10374 6684 10376
rect 3693 10371 3759 10374
rect 6678 10372 6684 10374
rect 6748 10372 6754 10436
rect 6821 10434 6887 10437
rect 9213 10434 9279 10437
rect 6821 10432 9279 10434
rect 6821 10376 6826 10432
rect 6882 10376 9218 10432
rect 9274 10376 9279 10432
rect 6821 10374 9279 10376
rect 6821 10371 6887 10374
rect 9213 10371 9279 10374
rect 13721 10434 13787 10437
rect 16205 10434 16271 10437
rect 13721 10432 16271 10434
rect 13721 10376 13726 10432
rect 13782 10376 16210 10432
rect 16266 10376 16271 10432
rect 13721 10374 16271 10376
rect 13721 10371 13787 10374
rect 16205 10371 16271 10374
rect 21541 10434 21607 10437
rect 24117 10434 24183 10437
rect 21541 10432 24183 10434
rect 21541 10376 21546 10432
rect 21602 10376 24122 10432
rect 24178 10376 24183 10432
rect 21541 10374 24183 10376
rect 21541 10371 21607 10374
rect 24117 10371 24183 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 2589 10298 2655 10301
rect 6821 10298 6887 10301
rect 2589 10296 6887 10298
rect 2589 10240 2594 10296
rect 2650 10240 6826 10296
rect 6882 10240 6887 10296
rect 2589 10238 6887 10240
rect 2589 10235 2655 10238
rect 6821 10235 6887 10238
rect 8293 10298 8359 10301
rect 9029 10298 9095 10301
rect 9581 10298 9647 10301
rect 10777 10300 10843 10301
rect 8293 10296 9647 10298
rect 8293 10240 8298 10296
rect 8354 10240 9034 10296
rect 9090 10240 9586 10296
rect 9642 10240 9647 10296
rect 8293 10238 9647 10240
rect 8293 10235 8359 10238
rect 9029 10235 9095 10238
rect 9581 10235 9647 10238
rect 10726 10236 10732 10300
rect 10796 10298 10843 10300
rect 12709 10298 12775 10301
rect 19333 10298 19399 10301
rect 10796 10296 10888 10298
rect 10838 10240 10888 10296
rect 10796 10238 10888 10240
rect 12709 10296 19399 10298
rect 12709 10240 12714 10296
rect 12770 10240 19338 10296
rect 19394 10240 19399 10296
rect 12709 10238 19399 10240
rect 10796 10236 10843 10238
rect 10777 10235 10843 10236
rect 12709 10235 12775 10238
rect 19333 10235 19399 10238
rect 22686 10236 22692 10300
rect 22756 10298 22762 10300
rect 23657 10298 23723 10301
rect 24718 10300 24778 10510
rect 24853 10300 24919 10301
rect 22756 10296 23723 10298
rect 22756 10240 23662 10296
rect 23718 10240 23723 10296
rect 22756 10238 23723 10240
rect 22756 10236 22762 10238
rect 23657 10235 23723 10238
rect 24710 10236 24716 10300
rect 24780 10236 24786 10300
rect 24853 10296 24900 10300
rect 24964 10298 24970 10300
rect 24853 10240 24858 10296
rect 24853 10236 24900 10240
rect 24964 10238 25010 10298
rect 24964 10236 24970 10238
rect 24853 10235 24919 10236
rect 0 10162 480 10192
rect 13353 10162 13419 10165
rect 0 10160 13419 10162
rect 0 10104 13358 10160
rect 13414 10104 13419 10160
rect 0 10102 13419 10104
rect 0 10072 480 10102
rect 13353 10099 13419 10102
rect 14641 10162 14707 10165
rect 21173 10162 21239 10165
rect 14641 10160 21239 10162
rect 14641 10104 14646 10160
rect 14702 10104 21178 10160
rect 21234 10104 21239 10160
rect 14641 10102 21239 10104
rect 14641 10099 14707 10102
rect 21173 10099 21239 10102
rect 23749 10162 23815 10165
rect 27520 10162 28000 10192
rect 23749 10160 28000 10162
rect 23749 10104 23754 10160
rect 23810 10104 28000 10160
rect 23749 10102 28000 10104
rect 23749 10099 23815 10102
rect 27520 10072 28000 10102
rect 3877 10026 3943 10029
rect 7189 10026 7255 10029
rect 3877 10024 7255 10026
rect 3877 9968 3882 10024
rect 3938 9968 7194 10024
rect 7250 9968 7255 10024
rect 3877 9966 7255 9968
rect 3877 9963 3943 9966
rect 7189 9963 7255 9966
rect 7649 10026 7715 10029
rect 15561 10026 15627 10029
rect 16941 10026 17007 10029
rect 7649 10024 15627 10026
rect 7649 9968 7654 10024
rect 7710 9968 15566 10024
rect 15622 9968 15627 10024
rect 7649 9966 15627 9968
rect 7649 9963 7715 9966
rect 15561 9963 15627 9966
rect 16254 10024 17007 10026
rect 16254 9968 16946 10024
rect 17002 9968 17007 10024
rect 16254 9966 17007 9968
rect 8886 9828 8892 9892
rect 8956 9890 8962 9892
rect 9121 9890 9187 9893
rect 8956 9888 9187 9890
rect 8956 9832 9126 9888
rect 9182 9832 9187 9888
rect 8956 9830 9187 9832
rect 8956 9828 8962 9830
rect 9121 9827 9187 9830
rect 9581 9890 9647 9893
rect 13721 9890 13787 9893
rect 9581 9888 13787 9890
rect 9581 9832 9586 9888
rect 9642 9832 13726 9888
rect 13782 9832 13787 9888
rect 9581 9830 13787 9832
rect 9581 9827 9647 9830
rect 13721 9827 13787 9830
rect 13905 9890 13971 9893
rect 14774 9890 14780 9892
rect 13905 9888 14780 9890
rect 13905 9832 13910 9888
rect 13966 9832 14780 9888
rect 13905 9830 14780 9832
rect 13905 9827 13971 9830
rect 14774 9828 14780 9830
rect 14844 9828 14850 9892
rect 15653 9890 15719 9893
rect 16254 9892 16314 9966
rect 16941 9963 17007 9966
rect 18873 10026 18939 10029
rect 24945 10026 25011 10029
rect 18873 10024 25011 10026
rect 18873 9968 18878 10024
rect 18934 9968 24950 10024
rect 25006 9968 25011 10024
rect 18873 9966 25011 9968
rect 18873 9963 18939 9966
rect 24945 9963 25011 9966
rect 16246 9890 16252 9892
rect 15653 9888 16252 9890
rect 15653 9832 15658 9888
rect 15714 9832 16252 9888
rect 15653 9830 16252 9832
rect 15653 9827 15719 9830
rect 16246 9828 16252 9830
rect 16316 9828 16322 9892
rect 16849 9890 16915 9893
rect 22870 9890 22876 9892
rect 16849 9888 22876 9890
rect 16849 9832 16854 9888
rect 16910 9832 22876 9888
rect 16849 9830 22876 9832
rect 16849 9827 16915 9830
rect 22870 9828 22876 9830
rect 22940 9828 22946 9892
rect 23473 9890 23539 9893
rect 23246 9888 23539 9890
rect 23246 9832 23478 9888
rect 23534 9832 23539 9888
rect 23246 9830 23539 9832
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 7465 9754 7531 9757
rect 7833 9754 7899 9757
rect 13813 9754 13879 9757
rect 7465 9752 13879 9754
rect 7465 9696 7470 9752
rect 7526 9696 7838 9752
rect 7894 9696 13818 9752
rect 13874 9696 13879 9752
rect 7465 9694 13879 9696
rect 7465 9691 7531 9694
rect 7833 9691 7899 9694
rect 13813 9691 13879 9694
rect 15929 9754 15995 9757
rect 16205 9754 16271 9757
rect 17401 9754 17467 9757
rect 23246 9754 23306 9830
rect 23473 9827 23539 9830
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 15929 9752 16130 9754
rect 15929 9696 15934 9752
rect 15990 9696 16130 9752
rect 15929 9694 16130 9696
rect 15929 9691 15995 9694
rect 0 9618 480 9648
rect 12709 9618 12775 9621
rect 15837 9618 15903 9621
rect 0 9558 7666 9618
rect 0 9528 480 9558
rect 5625 9482 5691 9485
rect 6126 9482 6132 9484
rect 5625 9480 6132 9482
rect 5625 9424 5630 9480
rect 5686 9424 6132 9480
rect 5625 9422 6132 9424
rect 5625 9419 5691 9422
rect 6126 9420 6132 9422
rect 6196 9420 6202 9484
rect 0 9074 480 9104
rect 7097 9074 7163 9077
rect 0 9072 7163 9074
rect 0 9016 7102 9072
rect 7158 9016 7163 9072
rect 0 9014 7163 9016
rect 7606 9074 7666 9558
rect 12709 9616 15903 9618
rect 12709 9560 12714 9616
rect 12770 9560 15842 9616
rect 15898 9560 15903 9616
rect 12709 9558 15903 9560
rect 16070 9618 16130 9694
rect 16205 9752 23306 9754
rect 16205 9696 16210 9752
rect 16266 9696 17406 9752
rect 17462 9696 23306 9752
rect 16205 9694 23306 9696
rect 16205 9691 16271 9694
rect 17401 9691 17467 9694
rect 23422 9692 23428 9756
rect 23492 9754 23498 9756
rect 23657 9754 23723 9757
rect 24853 9756 24919 9757
rect 24853 9754 24900 9756
rect 23492 9752 23723 9754
rect 23492 9696 23662 9752
rect 23718 9696 23723 9752
rect 23492 9694 23723 9696
rect 24808 9752 24900 9754
rect 24808 9696 24858 9752
rect 24808 9694 24900 9696
rect 23492 9692 23498 9694
rect 23657 9691 23723 9694
rect 24853 9692 24900 9694
rect 24964 9692 24970 9756
rect 24853 9691 24919 9692
rect 16481 9618 16547 9621
rect 16070 9616 16547 9618
rect 16070 9560 16486 9616
rect 16542 9560 16547 9616
rect 16070 9558 16547 9560
rect 12709 9555 12775 9558
rect 15837 9555 15903 9558
rect 16481 9555 16547 9558
rect 16614 9556 16620 9620
rect 16684 9618 16690 9620
rect 19517 9618 19583 9621
rect 27520 9618 28000 9648
rect 16684 9616 19583 9618
rect 16684 9560 19522 9616
rect 19578 9560 19583 9616
rect 16684 9558 19583 9560
rect 16684 9556 16690 9558
rect 19517 9555 19583 9558
rect 22142 9558 28000 9618
rect 8937 9482 9003 9485
rect 10317 9482 10383 9485
rect 13353 9482 13419 9485
rect 8937 9480 13419 9482
rect 8937 9424 8942 9480
rect 8998 9424 10322 9480
rect 10378 9424 13358 9480
rect 13414 9424 13419 9480
rect 8937 9422 13419 9424
rect 8937 9419 9003 9422
rect 10317 9419 10383 9422
rect 13353 9419 13419 9422
rect 14774 9420 14780 9484
rect 14844 9482 14850 9484
rect 15009 9482 15075 9485
rect 21357 9482 21423 9485
rect 14844 9480 15075 9482
rect 14844 9424 15014 9480
rect 15070 9424 15075 9480
rect 14844 9422 15075 9424
rect 14844 9420 14850 9422
rect 15009 9419 15075 9422
rect 18232 9480 21423 9482
rect 18232 9424 21362 9480
rect 21418 9424 21423 9480
rect 18232 9422 21423 9424
rect 18232 9349 18292 9422
rect 21357 9419 21423 9422
rect 21541 9482 21607 9485
rect 22142 9482 22202 9558
rect 27520 9528 28000 9558
rect 21541 9480 22202 9482
rect 21541 9424 21546 9480
rect 21602 9424 22202 9480
rect 21541 9422 22202 9424
rect 21541 9419 21607 9422
rect 23054 9420 23060 9484
rect 23124 9482 23130 9484
rect 23289 9482 23355 9485
rect 23124 9480 23355 9482
rect 23124 9424 23294 9480
rect 23350 9424 23355 9480
rect 23124 9422 23355 9424
rect 23124 9420 23130 9422
rect 23289 9419 23355 9422
rect 10685 9346 10751 9349
rect 15929 9346 15995 9349
rect 10685 9344 15995 9346
rect 10685 9288 10690 9344
rect 10746 9288 15934 9344
rect 15990 9288 15995 9344
rect 10685 9286 15995 9288
rect 10685 9283 10751 9286
rect 15929 9283 15995 9286
rect 16297 9346 16363 9349
rect 18229 9346 18295 9349
rect 20345 9348 20411 9349
rect 16297 9344 18295 9346
rect 16297 9288 16302 9344
rect 16358 9288 18234 9344
rect 18290 9288 18295 9344
rect 16297 9286 18295 9288
rect 16297 9283 16363 9286
rect 18229 9283 18295 9286
rect 20294 9284 20300 9348
rect 20364 9346 20411 9348
rect 20989 9346 21055 9349
rect 25405 9346 25471 9349
rect 20364 9344 20456 9346
rect 20406 9288 20456 9344
rect 20364 9286 20456 9288
rect 20989 9344 25471 9346
rect 20989 9288 20994 9344
rect 21050 9288 25410 9344
rect 25466 9288 25471 9344
rect 20989 9286 25471 9288
rect 20364 9284 20411 9286
rect 20345 9283 20411 9284
rect 20989 9283 21055 9286
rect 25405 9283 25471 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 12249 9210 12315 9213
rect 17677 9210 17743 9213
rect 12249 9208 17743 9210
rect 12249 9152 12254 9208
rect 12310 9152 17682 9208
rect 17738 9152 17743 9208
rect 12249 9150 17743 9152
rect 12249 9147 12315 9150
rect 17677 9147 17743 9150
rect 22277 9210 22343 9213
rect 23105 9210 23171 9213
rect 24393 9210 24459 9213
rect 22277 9208 24459 9210
rect 22277 9152 22282 9208
rect 22338 9152 23110 9208
rect 23166 9152 24398 9208
rect 24454 9152 24459 9208
rect 22277 9150 24459 9152
rect 22277 9147 22343 9150
rect 23105 9147 23171 9150
rect 24393 9147 24459 9150
rect 15929 9074 15995 9077
rect 16481 9074 16547 9077
rect 21541 9074 21607 9077
rect 7606 9072 15995 9074
rect 7606 9016 15934 9072
rect 15990 9016 15995 9072
rect 7606 9014 15995 9016
rect 0 8984 480 9014
rect 7097 9011 7163 9014
rect 15929 9011 15995 9014
rect 16070 9072 21607 9074
rect 16070 9016 16486 9072
rect 16542 9016 21546 9072
rect 21602 9016 21607 9072
rect 16070 9014 21607 9016
rect 2773 8938 2839 8941
rect 5625 8938 5691 8941
rect 9673 8938 9739 8941
rect 2773 8936 9739 8938
rect 2773 8880 2778 8936
rect 2834 8880 5630 8936
rect 5686 8880 9678 8936
rect 9734 8880 9739 8936
rect 2773 8878 9739 8880
rect 2773 8875 2839 8878
rect 5625 8875 5691 8878
rect 9673 8875 9739 8878
rect 13169 8938 13235 8941
rect 15377 8938 15443 8941
rect 13169 8936 15443 8938
rect 13169 8880 13174 8936
rect 13230 8880 15382 8936
rect 15438 8880 15443 8936
rect 13169 8878 15443 8880
rect 13169 8875 13235 8878
rect 15377 8875 15443 8878
rect 15694 8876 15700 8940
rect 15764 8938 15770 8940
rect 16070 8938 16130 9014
rect 16481 9011 16547 9014
rect 21541 9011 21607 9014
rect 21725 9074 21791 9077
rect 24669 9074 24735 9077
rect 27520 9074 28000 9104
rect 21725 9072 23628 9074
rect 21725 9016 21730 9072
rect 21786 9016 23628 9072
rect 21725 9014 23628 9016
rect 21725 9011 21791 9014
rect 23568 8941 23628 9014
rect 24669 9072 28000 9074
rect 24669 9016 24674 9072
rect 24730 9016 28000 9072
rect 24669 9014 28000 9016
rect 24669 9011 24735 9014
rect 27520 8984 28000 9014
rect 15764 8878 16130 8938
rect 16849 8938 16915 8941
rect 22921 8938 22987 8941
rect 16849 8936 22987 8938
rect 16849 8880 16854 8936
rect 16910 8880 22926 8936
rect 22982 8880 22987 8936
rect 16849 8878 22987 8880
rect 15764 8876 15770 8878
rect 16849 8875 16915 8878
rect 22921 8875 22987 8878
rect 23565 8936 23631 8941
rect 25313 8938 25379 8941
rect 23565 8880 23570 8936
rect 23626 8880 23631 8936
rect 23565 8875 23631 8880
rect 23798 8936 25379 8938
rect 23798 8880 25318 8936
rect 25374 8880 25379 8936
rect 23798 8878 25379 8880
rect 6177 8802 6243 8805
rect 8661 8802 8727 8805
rect 6177 8800 8727 8802
rect 6177 8744 6182 8800
rect 6238 8744 8666 8800
rect 8722 8744 8727 8800
rect 6177 8742 8727 8744
rect 6177 8739 6243 8742
rect 8661 8739 8727 8742
rect 14406 8740 14412 8804
rect 14476 8802 14482 8804
rect 14733 8802 14799 8805
rect 14476 8800 14799 8802
rect 14476 8744 14738 8800
rect 14794 8744 14799 8800
rect 14476 8742 14799 8744
rect 14476 8740 14482 8742
rect 14733 8739 14799 8742
rect 15837 8802 15903 8805
rect 16982 8802 16988 8804
rect 15837 8800 16988 8802
rect 15837 8744 15842 8800
rect 15898 8744 16988 8800
rect 15837 8742 16988 8744
rect 15837 8739 15903 8742
rect 16982 8740 16988 8742
rect 17052 8740 17058 8804
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 2814 8604 2820 8668
rect 2884 8666 2890 8668
rect 3969 8666 4035 8669
rect 2884 8664 4035 8666
rect 2884 8608 3974 8664
rect 4030 8608 4035 8664
rect 2884 8606 4035 8608
rect 2884 8604 2890 8606
rect 3969 8603 4035 8606
rect 6821 8666 6887 8669
rect 9305 8666 9371 8669
rect 9765 8666 9831 8669
rect 6821 8664 9831 8666
rect 6821 8608 6826 8664
rect 6882 8608 9310 8664
rect 9366 8608 9770 8664
rect 9826 8608 9831 8664
rect 6821 8606 9831 8608
rect 6821 8603 6887 8606
rect 9305 8603 9371 8606
rect 9765 8603 9831 8606
rect 10041 8666 10107 8669
rect 11789 8666 11855 8669
rect 10041 8664 11855 8666
rect 10041 8608 10046 8664
rect 10102 8608 11794 8664
rect 11850 8608 11855 8664
rect 10041 8606 11855 8608
rect 10041 8603 10107 8606
rect 11789 8603 11855 8606
rect 11973 8666 12039 8669
rect 14733 8666 14799 8669
rect 11973 8664 14799 8666
rect 11973 8608 11978 8664
rect 12034 8608 14738 8664
rect 14794 8608 14799 8664
rect 11973 8606 14799 8608
rect 11973 8603 12039 8606
rect 14733 8603 14799 8606
rect 15929 8666 15995 8669
rect 18689 8666 18755 8669
rect 15929 8664 18755 8666
rect 15929 8608 15934 8664
rect 15990 8608 18694 8664
rect 18750 8608 18755 8664
rect 15929 8606 18755 8608
rect 15929 8603 15995 8606
rect 18689 8603 18755 8606
rect 19609 8666 19675 8669
rect 23798 8666 23858 8878
rect 25313 8875 25379 8878
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 19609 8664 23858 8666
rect 19609 8608 19614 8664
rect 19670 8608 23858 8664
rect 19609 8606 23858 8608
rect 19609 8603 19675 8606
rect 23974 8604 23980 8668
rect 24044 8666 24050 8668
rect 24117 8666 24183 8669
rect 24044 8664 24183 8666
rect 24044 8608 24122 8664
rect 24178 8608 24183 8664
rect 24044 8606 24183 8608
rect 24044 8604 24050 8606
rect 24117 8603 24183 8606
rect 0 8530 480 8560
rect 3693 8530 3759 8533
rect 0 8528 3759 8530
rect 0 8472 3698 8528
rect 3754 8472 3759 8528
rect 0 8470 3759 8472
rect 0 8440 480 8470
rect 3693 8467 3759 8470
rect 5533 8530 5599 8533
rect 12525 8530 12591 8533
rect 15009 8530 15075 8533
rect 16297 8530 16363 8533
rect 5533 8528 14842 8530
rect 5533 8472 5538 8528
rect 5594 8472 12530 8528
rect 12586 8472 14842 8528
rect 5533 8470 14842 8472
rect 5533 8467 5599 8470
rect 12525 8467 12591 8470
rect 4429 8394 4495 8397
rect 7281 8394 7347 8397
rect 8845 8396 8911 8397
rect 8845 8394 8892 8396
rect 4429 8392 7347 8394
rect 4429 8336 4434 8392
rect 4490 8336 7286 8392
rect 7342 8336 7347 8392
rect 4429 8334 7347 8336
rect 8800 8392 8892 8394
rect 8800 8336 8850 8392
rect 8800 8334 8892 8336
rect 4429 8331 4495 8334
rect 7281 8331 7347 8334
rect 8845 8332 8892 8334
rect 8956 8332 8962 8396
rect 10593 8394 10659 8397
rect 9124 8392 10659 8394
rect 9124 8336 10598 8392
rect 10654 8336 10659 8392
rect 9124 8334 10659 8336
rect 8845 8331 8911 8332
rect 9124 8261 9184 8334
rect 10593 8331 10659 8334
rect 13905 8394 13971 8397
rect 14590 8394 14596 8396
rect 13905 8392 14596 8394
rect 13905 8336 13910 8392
rect 13966 8336 14596 8392
rect 13905 8334 14596 8336
rect 13905 8331 13971 8334
rect 14590 8332 14596 8334
rect 14660 8332 14666 8396
rect 14782 8394 14842 8470
rect 15009 8528 16363 8530
rect 15009 8472 15014 8528
rect 15070 8472 16302 8528
rect 16358 8472 16363 8528
rect 15009 8470 16363 8472
rect 15009 8467 15075 8470
rect 16297 8467 16363 8470
rect 17677 8530 17743 8533
rect 27520 8530 28000 8560
rect 17677 8528 28000 8530
rect 17677 8472 17682 8528
rect 17738 8472 28000 8528
rect 17677 8470 28000 8472
rect 17677 8467 17743 8470
rect 27520 8440 28000 8470
rect 20713 8394 20779 8397
rect 14782 8392 20779 8394
rect 14782 8336 20718 8392
rect 20774 8336 20779 8392
rect 14782 8334 20779 8336
rect 20713 8331 20779 8334
rect 23749 8394 23815 8397
rect 23974 8394 23980 8396
rect 23749 8392 23980 8394
rect 23749 8336 23754 8392
rect 23810 8336 23980 8392
rect 23749 8334 23980 8336
rect 23749 8331 23815 8334
rect 23974 8332 23980 8334
rect 24044 8332 24050 8396
rect 2446 8196 2452 8260
rect 2516 8258 2522 8260
rect 3233 8258 3299 8261
rect 2516 8256 3299 8258
rect 2516 8200 3238 8256
rect 3294 8200 3299 8256
rect 2516 8198 3299 8200
rect 2516 8196 2522 8198
rect 3233 8195 3299 8198
rect 7649 8258 7715 8261
rect 7782 8258 7788 8260
rect 7649 8256 7788 8258
rect 7649 8200 7654 8256
rect 7710 8200 7788 8256
rect 7649 8198 7788 8200
rect 7649 8195 7715 8198
rect 7782 8196 7788 8198
rect 7852 8196 7858 8260
rect 9121 8256 9187 8261
rect 9121 8200 9126 8256
rect 9182 8200 9187 8256
rect 9121 8195 9187 8200
rect 10685 8258 10751 8261
rect 15837 8258 15903 8261
rect 10685 8256 15903 8258
rect 10685 8200 10690 8256
rect 10746 8200 15842 8256
rect 15898 8200 15903 8256
rect 10685 8198 15903 8200
rect 10685 8195 10751 8198
rect 15837 8195 15903 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 5809 8122 5875 8125
rect 9765 8122 9831 8125
rect 14365 8122 14431 8125
rect 5809 8120 9831 8122
rect 5809 8064 5814 8120
rect 5870 8064 9770 8120
rect 9826 8064 9831 8120
rect 5809 8062 9831 8064
rect 5809 8059 5875 8062
rect 9765 8059 9831 8062
rect 10734 8120 14431 8122
rect 10734 8064 14370 8120
rect 14426 8064 14431 8120
rect 10734 8062 14431 8064
rect 6453 7986 6519 7989
rect 10734 7986 10794 8062
rect 14365 8059 14431 8062
rect 15285 8122 15351 8125
rect 15510 8122 15516 8124
rect 15285 8120 15516 8122
rect 15285 8064 15290 8120
rect 15346 8064 15516 8120
rect 15285 8062 15516 8064
rect 15285 8059 15351 8062
rect 15510 8060 15516 8062
rect 15580 8060 15586 8124
rect 6453 7984 10794 7986
rect 6453 7928 6458 7984
rect 6514 7928 10794 7984
rect 6453 7926 10794 7928
rect 11053 7986 11119 7989
rect 13905 7986 13971 7989
rect 11053 7984 13971 7986
rect 11053 7928 11058 7984
rect 11114 7928 13910 7984
rect 13966 7928 13971 7984
rect 11053 7926 13971 7928
rect 6453 7923 6519 7926
rect 11053 7923 11119 7926
rect 13905 7923 13971 7926
rect 14774 7924 14780 7988
rect 14844 7986 14850 7988
rect 14917 7986 14983 7989
rect 14844 7984 14983 7986
rect 14844 7928 14922 7984
rect 14978 7928 14983 7984
rect 14844 7926 14983 7928
rect 14844 7924 14850 7926
rect 14917 7923 14983 7926
rect 18321 7986 18387 7989
rect 20897 7986 20963 7989
rect 18321 7984 20963 7986
rect 18321 7928 18326 7984
rect 18382 7928 20902 7984
rect 20958 7928 20963 7984
rect 18321 7926 20963 7928
rect 18321 7923 18387 7926
rect 20897 7923 20963 7926
rect 23841 7986 23907 7989
rect 24117 7986 24183 7989
rect 23841 7984 24183 7986
rect 23841 7928 23846 7984
rect 23902 7928 24122 7984
rect 24178 7928 24183 7984
rect 23841 7926 24183 7928
rect 23841 7923 23907 7926
rect 24117 7923 24183 7926
rect 0 7850 480 7880
rect 3969 7850 4035 7853
rect 0 7848 4035 7850
rect 0 7792 3974 7848
rect 4030 7792 4035 7848
rect 0 7790 4035 7792
rect 0 7760 480 7790
rect 3969 7787 4035 7790
rect 5349 7850 5415 7853
rect 8845 7850 8911 7853
rect 5349 7848 8911 7850
rect 5349 7792 5354 7848
rect 5410 7792 8850 7848
rect 8906 7792 8911 7848
rect 5349 7790 8911 7792
rect 5349 7787 5415 7790
rect 8845 7787 8911 7790
rect 14733 7850 14799 7853
rect 16389 7850 16455 7853
rect 17217 7850 17283 7853
rect 22001 7850 22067 7853
rect 14733 7848 15394 7850
rect 14733 7792 14738 7848
rect 14794 7792 15394 7848
rect 14733 7790 15394 7792
rect 14733 7787 14799 7790
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 11830 7516 11836 7580
rect 11900 7578 11906 7580
rect 12341 7578 12407 7581
rect 15334 7578 15394 7790
rect 16389 7848 22067 7850
rect 16389 7792 16394 7848
rect 16450 7792 17222 7848
rect 17278 7792 22006 7848
rect 22062 7792 22067 7848
rect 16389 7790 22067 7792
rect 16389 7787 16455 7790
rect 17217 7787 17283 7790
rect 22001 7787 22067 7790
rect 23238 7788 23244 7852
rect 23308 7850 23314 7852
rect 23381 7850 23447 7853
rect 27520 7850 28000 7880
rect 23308 7848 23447 7850
rect 23308 7792 23386 7848
rect 23442 7792 23447 7848
rect 23308 7790 23447 7792
rect 23308 7788 23314 7790
rect 23381 7787 23447 7790
rect 24120 7790 28000 7850
rect 16573 7714 16639 7717
rect 24120 7714 24180 7790
rect 27520 7760 28000 7790
rect 16573 7712 24180 7714
rect 16573 7656 16578 7712
rect 16634 7656 24180 7712
rect 16573 7654 24180 7656
rect 16573 7651 16639 7654
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 11900 7576 14152 7578
rect 11900 7520 12346 7576
rect 12402 7520 14152 7576
rect 11900 7518 14152 7520
rect 15334 7518 23674 7578
rect 11900 7516 11906 7518
rect 12341 7515 12407 7518
rect 3049 7442 3115 7445
rect 12157 7442 12223 7445
rect 3049 7440 12223 7442
rect 3049 7384 3054 7440
rect 3110 7384 12162 7440
rect 12218 7384 12223 7440
rect 3049 7382 12223 7384
rect 3049 7379 3115 7382
rect 12157 7379 12223 7382
rect 0 7306 480 7336
rect 3918 7306 3924 7308
rect 0 7246 3924 7306
rect 0 7216 480 7246
rect 3918 7244 3924 7246
rect 3988 7244 3994 7308
rect 6361 7306 6427 7309
rect 7782 7306 7788 7308
rect 6361 7304 7788 7306
rect 6361 7248 6366 7304
rect 6422 7248 7788 7304
rect 6361 7246 7788 7248
rect 6361 7243 6427 7246
rect 7782 7244 7788 7246
rect 7852 7244 7858 7308
rect 8569 7306 8635 7309
rect 12433 7306 12499 7309
rect 8569 7304 12499 7306
rect 8569 7248 8574 7304
rect 8630 7248 12438 7304
rect 12494 7248 12499 7304
rect 8569 7246 12499 7248
rect 8569 7243 8635 7246
rect 12433 7243 12499 7246
rect 3969 7170 4035 7173
rect 7281 7170 7347 7173
rect 3969 7168 7347 7170
rect 3969 7112 3974 7168
rect 4030 7112 7286 7168
rect 7342 7112 7347 7168
rect 3969 7110 7347 7112
rect 3969 7107 4035 7110
rect 7281 7107 7347 7110
rect 13302 7108 13308 7172
rect 13372 7170 13378 7172
rect 13445 7170 13511 7173
rect 14092 7170 14152 7518
rect 14457 7442 14523 7445
rect 22461 7442 22527 7445
rect 14457 7440 22527 7442
rect 14457 7384 14462 7440
rect 14518 7384 22466 7440
rect 22522 7384 22527 7440
rect 14457 7382 22527 7384
rect 14457 7379 14523 7382
rect 22461 7379 22527 7382
rect 14273 7306 14339 7309
rect 23473 7306 23539 7309
rect 14273 7304 23539 7306
rect 14273 7248 14278 7304
rect 14334 7248 23478 7304
rect 23534 7248 23539 7304
rect 14273 7246 23539 7248
rect 23614 7306 23674 7518
rect 23790 7516 23796 7580
rect 23860 7578 23866 7580
rect 23933 7578 23999 7581
rect 23860 7576 23999 7578
rect 23860 7520 23938 7576
rect 23994 7520 23999 7576
rect 23860 7518 23999 7520
rect 23860 7516 23866 7518
rect 23933 7515 23999 7518
rect 24301 7306 24367 7309
rect 27520 7306 28000 7336
rect 23614 7304 28000 7306
rect 23614 7248 24306 7304
rect 24362 7248 28000 7304
rect 23614 7246 28000 7248
rect 14273 7243 14339 7246
rect 23473 7243 23539 7246
rect 24301 7243 24367 7246
rect 27520 7216 28000 7246
rect 13372 7168 13968 7170
rect 13372 7112 13450 7168
rect 13506 7112 13968 7168
rect 13372 7110 13968 7112
rect 14092 7110 18154 7170
rect 13372 7108 13378 7110
rect 13445 7107 13511 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 2773 7034 2839 7037
rect 13908 7034 13968 7110
rect 15653 7034 15719 7037
rect 2773 7032 10196 7034
rect 2773 6976 2778 7032
rect 2834 6976 10196 7032
rect 2773 6974 10196 6976
rect 13908 7032 15719 7034
rect 13908 6976 15658 7032
rect 15714 6976 15719 7032
rect 13908 6974 15719 6976
rect 2773 6971 2839 6974
rect 1945 6898 2011 6901
rect 6085 6898 6151 6901
rect 1945 6896 6151 6898
rect 1945 6840 1950 6896
rect 2006 6840 6090 6896
rect 6146 6840 6151 6896
rect 1945 6838 6151 6840
rect 10136 6898 10196 6974
rect 15653 6971 15719 6974
rect 11830 6898 11836 6900
rect 10136 6838 11836 6898
rect 1945 6835 2011 6838
rect 6085 6835 6151 6838
rect 11830 6836 11836 6838
rect 11900 6836 11906 6900
rect 16573 6898 16639 6901
rect 13678 6896 16639 6898
rect 13678 6840 16578 6896
rect 16634 6840 16639 6896
rect 13678 6838 16639 6840
rect 0 6762 480 6792
rect 3918 6762 3924 6764
rect 0 6702 3924 6762
rect 0 6672 480 6702
rect 3918 6700 3924 6702
rect 3988 6700 3994 6764
rect 6453 6762 6519 6765
rect 13678 6762 13738 6838
rect 16573 6835 16639 6838
rect 15469 6762 15535 6765
rect 6453 6760 13738 6762
rect 6453 6704 6458 6760
rect 6514 6704 13738 6760
rect 6453 6702 13738 6704
rect 13816 6760 15535 6762
rect 13816 6704 15474 6760
rect 15530 6704 15535 6760
rect 13816 6702 15535 6704
rect 18094 6762 18154 7110
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 19374 6836 19380 6900
rect 19444 6898 19450 6900
rect 20294 6898 20300 6900
rect 19444 6838 20300 6898
rect 19444 6836 19450 6838
rect 20294 6836 20300 6838
rect 20364 6836 20370 6900
rect 27520 6762 28000 6792
rect 18094 6702 28000 6762
rect 6453 6699 6519 6702
rect 10685 6626 10751 6629
rect 13816 6626 13876 6702
rect 15469 6699 15535 6702
rect 27520 6672 28000 6702
rect 10685 6624 13876 6626
rect 10685 6568 10690 6624
rect 10746 6568 13876 6624
rect 10685 6566 13876 6568
rect 16849 6626 16915 6629
rect 20529 6626 20595 6629
rect 16849 6624 20595 6626
rect 16849 6568 16854 6624
rect 16910 6568 20534 6624
rect 20590 6568 20595 6624
rect 16849 6566 20595 6568
rect 10685 6563 10751 6566
rect 16849 6563 16915 6566
rect 20529 6563 20595 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 5257 6490 5323 6493
rect 5390 6490 5396 6492
rect 5257 6488 5396 6490
rect 5257 6432 5262 6488
rect 5318 6432 5396 6488
rect 5257 6430 5396 6432
rect 5257 6427 5323 6430
rect 5390 6428 5396 6430
rect 5460 6428 5466 6492
rect 6453 6490 6519 6493
rect 17769 6492 17835 6493
rect 6453 6488 13692 6490
rect 6453 6432 6458 6488
rect 6514 6432 13692 6488
rect 6453 6430 13692 6432
rect 6453 6427 6519 6430
rect 3877 6354 3943 6357
rect 5257 6354 5323 6357
rect 10041 6354 10107 6357
rect 3877 6352 10107 6354
rect 3877 6296 3882 6352
rect 3938 6296 5262 6352
rect 5318 6296 10046 6352
rect 10102 6296 10107 6352
rect 3877 6294 10107 6296
rect 13632 6354 13692 6430
rect 17718 6428 17724 6492
rect 17788 6490 17835 6492
rect 17788 6488 17880 6490
rect 17830 6432 17880 6488
rect 17788 6430 17880 6432
rect 17788 6428 17835 6430
rect 20110 6428 20116 6492
rect 20180 6490 20186 6492
rect 23381 6490 23447 6493
rect 23749 6492 23815 6493
rect 23749 6490 23796 6492
rect 20180 6488 23447 6490
rect 20180 6432 23386 6488
rect 23442 6432 23447 6488
rect 20180 6430 23447 6432
rect 23704 6488 23796 6490
rect 23704 6432 23754 6488
rect 23704 6430 23796 6432
rect 20180 6428 20186 6430
rect 17769 6427 17835 6428
rect 23381 6427 23447 6430
rect 23749 6428 23796 6430
rect 23860 6428 23866 6492
rect 23749 6427 23815 6428
rect 17677 6354 17743 6357
rect 13632 6352 17743 6354
rect 13632 6296 17682 6352
rect 17738 6296 17743 6352
rect 13632 6294 17743 6296
rect 3877 6291 3943 6294
rect 5257 6291 5323 6294
rect 10041 6291 10107 6294
rect 17677 6291 17743 6294
rect 17861 6354 17927 6357
rect 24577 6354 24643 6357
rect 17861 6352 24643 6354
rect 17861 6296 17866 6352
rect 17922 6296 24582 6352
rect 24638 6296 24643 6352
rect 17861 6294 24643 6296
rect 17861 6291 17927 6294
rect 24577 6291 24643 6294
rect 4705 6218 4771 6221
rect 11881 6218 11947 6221
rect 4705 6216 11947 6218
rect 4705 6160 4710 6216
rect 4766 6160 11886 6216
rect 11942 6160 11947 6216
rect 4705 6158 11947 6160
rect 4705 6155 4771 6158
rect 11881 6155 11947 6158
rect 14733 6218 14799 6221
rect 19609 6218 19675 6221
rect 14733 6216 19675 6218
rect 14733 6160 14738 6216
rect 14794 6160 19614 6216
rect 19670 6160 19675 6216
rect 14733 6158 19675 6160
rect 14733 6155 14799 6158
rect 19609 6155 19675 6158
rect 22369 6218 22435 6221
rect 25037 6218 25103 6221
rect 22369 6216 25103 6218
rect 22369 6160 22374 6216
rect 22430 6160 25042 6216
rect 25098 6160 25103 6216
rect 22369 6158 25103 6160
rect 22369 6155 22435 6158
rect 25037 6155 25103 6158
rect 0 6082 480 6112
rect 3049 6082 3115 6085
rect 0 6080 3115 6082
rect 0 6024 3054 6080
rect 3110 6024 3115 6080
rect 0 6022 3115 6024
rect 0 5992 480 6022
rect 3049 6019 3115 6022
rect 14774 6020 14780 6084
rect 14844 6082 14850 6084
rect 15193 6082 15259 6085
rect 14844 6080 15259 6082
rect 14844 6024 15198 6080
rect 15254 6024 15259 6080
rect 14844 6022 15259 6024
rect 14844 6020 14850 6022
rect 15193 6019 15259 6022
rect 15377 6082 15443 6085
rect 19149 6082 19215 6085
rect 15377 6080 19215 6082
rect 15377 6024 15382 6080
rect 15438 6024 19154 6080
rect 19210 6024 19215 6080
rect 15377 6022 19215 6024
rect 15377 6019 15443 6022
rect 19149 6019 19215 6022
rect 20294 6020 20300 6084
rect 20364 6082 20370 6084
rect 27520 6082 28000 6112
rect 20364 6022 28000 6082
rect 20364 6020 20370 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 27520 5992 28000 6022
rect 19610 5951 19930 5952
rect 11513 5948 11579 5949
rect 11462 5884 11468 5948
rect 11532 5946 11579 5948
rect 11532 5944 11624 5946
rect 11574 5888 11624 5944
rect 11532 5886 11624 5888
rect 11532 5884 11579 5886
rect 11830 5884 11836 5948
rect 11900 5946 11906 5948
rect 15653 5946 15719 5949
rect 18229 5946 18295 5949
rect 11900 5944 15719 5946
rect 11900 5888 15658 5944
rect 15714 5888 15719 5944
rect 11900 5886 15719 5888
rect 11900 5884 11906 5886
rect 11513 5883 11579 5884
rect 15653 5883 15719 5886
rect 16254 5944 18295 5946
rect 16254 5888 18234 5944
rect 18290 5888 18295 5944
rect 16254 5886 18295 5888
rect 9673 5810 9739 5813
rect 10685 5810 10751 5813
rect 9673 5808 10751 5810
rect 9673 5752 9678 5808
rect 9734 5752 10690 5808
rect 10746 5752 10751 5808
rect 9673 5750 10751 5752
rect 9673 5747 9739 5750
rect 10685 5747 10751 5750
rect 13353 5810 13419 5813
rect 16254 5810 16314 5886
rect 18229 5883 18295 5886
rect 18689 5946 18755 5949
rect 19241 5948 19307 5949
rect 19190 5946 19196 5948
rect 18689 5944 19196 5946
rect 19260 5946 19307 5948
rect 20069 5946 20135 5949
rect 19260 5944 19352 5946
rect 18689 5888 18694 5944
rect 18750 5888 19196 5944
rect 19302 5888 19352 5944
rect 18689 5886 19196 5888
rect 18689 5883 18755 5886
rect 19190 5884 19196 5886
rect 19260 5886 19352 5888
rect 20069 5944 23858 5946
rect 20069 5888 20074 5944
rect 20130 5888 23858 5944
rect 20069 5886 23858 5888
rect 19260 5884 19307 5886
rect 19241 5883 19307 5884
rect 20069 5883 20135 5886
rect 13353 5808 16314 5810
rect 13353 5752 13358 5808
rect 13414 5752 16314 5808
rect 13353 5750 16314 5752
rect 18965 5810 19031 5813
rect 23565 5810 23631 5813
rect 18965 5808 23631 5810
rect 18965 5752 18970 5808
rect 19026 5752 23570 5808
rect 23626 5752 23631 5808
rect 18965 5750 23631 5752
rect 13353 5747 13419 5750
rect 18965 5747 19031 5750
rect 23565 5747 23631 5750
rect 5809 5674 5875 5677
rect 8385 5674 8451 5677
rect 10041 5674 10107 5677
rect 5809 5672 10107 5674
rect 5809 5616 5814 5672
rect 5870 5616 8390 5672
rect 8446 5616 10046 5672
rect 10102 5616 10107 5672
rect 5809 5614 10107 5616
rect 5809 5611 5875 5614
rect 8385 5611 8451 5614
rect 10041 5611 10107 5614
rect 16021 5674 16087 5677
rect 17493 5676 17559 5677
rect 16021 5672 17418 5674
rect 16021 5616 16026 5672
rect 16082 5616 17418 5672
rect 16021 5614 17418 5616
rect 16021 5611 16087 5614
rect 0 5538 480 5568
rect 2998 5538 3004 5540
rect 0 5478 3004 5538
rect 0 5448 480 5478
rect 2998 5476 3004 5478
rect 3068 5476 3074 5540
rect 11237 5538 11303 5541
rect 6088 5536 11303 5538
rect 6088 5480 11242 5536
rect 11298 5480 11303 5536
rect 6088 5478 11303 5480
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 2405 5402 2471 5405
rect 4981 5402 5047 5405
rect 2405 5400 5047 5402
rect 2405 5344 2410 5400
rect 2466 5344 4986 5400
rect 5042 5344 5047 5400
rect 2405 5342 5047 5344
rect 2405 5339 2471 5342
rect 4981 5339 5047 5342
rect 4613 5266 4679 5269
rect 6088 5266 6148 5478
rect 11237 5475 11303 5478
rect 11462 5476 11468 5540
rect 11532 5538 11538 5540
rect 13813 5538 13879 5541
rect 11532 5536 13879 5538
rect 11532 5480 13818 5536
rect 13874 5480 13879 5536
rect 11532 5478 13879 5480
rect 11532 5476 11538 5478
rect 7373 5402 7439 5405
rect 7598 5402 7604 5404
rect 7373 5400 7604 5402
rect 7373 5344 7378 5400
rect 7434 5344 7604 5400
rect 7373 5342 7604 5344
rect 7373 5339 7439 5342
rect 7598 5340 7604 5342
rect 7668 5340 7674 5404
rect 11094 5340 11100 5404
rect 11164 5402 11170 5404
rect 11470 5402 11530 5476
rect 13813 5475 13879 5478
rect 15561 5538 15627 5541
rect 16246 5538 16252 5540
rect 15561 5536 16252 5538
rect 15561 5480 15566 5536
rect 15622 5480 16252 5536
rect 15561 5478 16252 5480
rect 15561 5475 15627 5478
rect 16246 5476 16252 5478
rect 16316 5476 16322 5540
rect 17358 5538 17418 5614
rect 17493 5672 17540 5676
rect 17604 5674 17610 5676
rect 18137 5674 18203 5677
rect 23197 5674 23263 5677
rect 17493 5616 17498 5672
rect 17493 5612 17540 5616
rect 17604 5614 17650 5674
rect 18137 5672 23263 5674
rect 18137 5616 18142 5672
rect 18198 5616 23202 5672
rect 23258 5616 23263 5672
rect 18137 5614 23263 5616
rect 17604 5612 17610 5614
rect 17493 5611 17559 5612
rect 18137 5611 18203 5614
rect 23197 5611 23263 5614
rect 20345 5538 20411 5541
rect 17358 5536 20411 5538
rect 17358 5480 20350 5536
rect 20406 5480 20411 5536
rect 17358 5478 20411 5480
rect 20345 5475 20411 5478
rect 20621 5538 20687 5541
rect 23657 5538 23723 5541
rect 20621 5536 23723 5538
rect 20621 5480 20626 5536
rect 20682 5480 23662 5536
rect 23718 5480 23723 5536
rect 20621 5478 23723 5480
rect 23798 5538 23858 5886
rect 24669 5810 24735 5813
rect 24894 5810 24900 5812
rect 24669 5808 24900 5810
rect 24669 5752 24674 5808
rect 24730 5752 24900 5808
rect 24669 5750 24900 5752
rect 24669 5747 24735 5750
rect 24894 5748 24900 5750
rect 24964 5748 24970 5812
rect 23933 5538 23999 5541
rect 23798 5536 23999 5538
rect 23798 5480 23938 5536
rect 23994 5480 23999 5536
rect 23798 5478 23999 5480
rect 20621 5475 20687 5478
rect 23657 5475 23723 5478
rect 23933 5475 23999 5478
rect 24853 5538 24919 5541
rect 27520 5538 28000 5568
rect 24853 5536 28000 5538
rect 24853 5480 24858 5536
rect 24914 5480 28000 5536
rect 24853 5478 28000 5480
rect 24853 5475 24919 5478
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 27520 5448 28000 5478
rect 24277 5407 24597 5408
rect 11164 5342 11530 5402
rect 16021 5402 16087 5405
rect 23841 5402 23907 5405
rect 16021 5400 23907 5402
rect 16021 5344 16026 5400
rect 16082 5344 23846 5400
rect 23902 5344 23907 5400
rect 16021 5342 23907 5344
rect 11164 5340 11170 5342
rect 16021 5339 16087 5342
rect 23841 5339 23907 5342
rect 4613 5264 6148 5266
rect 4613 5208 4618 5264
rect 4674 5208 6148 5264
rect 4613 5206 6148 5208
rect 9765 5266 9831 5269
rect 13905 5266 13971 5269
rect 15653 5268 15719 5269
rect 15653 5266 15700 5268
rect 9765 5264 13971 5266
rect 9765 5208 9770 5264
rect 9826 5208 13910 5264
rect 13966 5208 13971 5264
rect 9765 5206 13971 5208
rect 15608 5264 15700 5266
rect 15608 5208 15658 5264
rect 15608 5206 15700 5208
rect 4613 5203 4679 5206
rect 9765 5203 9831 5206
rect 13905 5203 13971 5206
rect 15653 5204 15700 5206
rect 15764 5204 15770 5268
rect 17350 5204 17356 5268
rect 17420 5266 17426 5268
rect 21766 5266 21772 5268
rect 17420 5206 21772 5266
rect 17420 5204 17426 5206
rect 21766 5204 21772 5206
rect 21836 5204 21842 5268
rect 15653 5203 15719 5204
rect 5809 5130 5875 5133
rect 7373 5130 7439 5133
rect 8293 5130 8359 5133
rect 9489 5132 9555 5133
rect 5809 5128 8359 5130
rect 5809 5072 5814 5128
rect 5870 5072 7378 5128
rect 7434 5072 8298 5128
rect 8354 5072 8359 5128
rect 5809 5070 8359 5072
rect 5809 5067 5875 5070
rect 7373 5067 7439 5070
rect 8293 5067 8359 5070
rect 9438 5068 9444 5132
rect 9508 5130 9555 5132
rect 12433 5130 12499 5133
rect 25221 5130 25287 5133
rect 9508 5128 9600 5130
rect 9550 5072 9600 5128
rect 9508 5070 9600 5072
rect 12433 5128 25287 5130
rect 12433 5072 12438 5128
rect 12494 5072 25226 5128
rect 25282 5072 25287 5128
rect 12433 5070 25287 5072
rect 9508 5068 9555 5070
rect 9489 5067 9555 5068
rect 12433 5067 12499 5070
rect 25221 5067 25287 5070
rect 0 4994 480 5024
rect 7465 4994 7531 4997
rect 0 4992 7531 4994
rect 0 4936 7470 4992
rect 7526 4936 7531 4992
rect 0 4934 7531 4936
rect 0 4904 480 4934
rect 7465 4931 7531 4934
rect 8017 4994 8083 4997
rect 8477 4994 8543 4997
rect 9673 4994 9739 4997
rect 8017 4992 9739 4994
rect 8017 4936 8022 4992
rect 8078 4936 8482 4992
rect 8538 4936 9678 4992
rect 9734 4936 9739 4992
rect 8017 4934 9739 4936
rect 8017 4931 8083 4934
rect 8477 4931 8543 4934
rect 9673 4931 9739 4934
rect 10685 4994 10751 4997
rect 11421 4994 11487 4997
rect 15929 4994 15995 4997
rect 10685 4992 15995 4994
rect 10685 4936 10690 4992
rect 10746 4936 11426 4992
rect 11482 4936 15934 4992
rect 15990 4936 15995 4992
rect 10685 4934 15995 4936
rect 10685 4931 10751 4934
rect 11421 4931 11487 4934
rect 15929 4931 15995 4934
rect 16389 4994 16455 4997
rect 19333 4994 19399 4997
rect 16389 4992 19399 4994
rect 16389 4936 16394 4992
rect 16450 4936 19338 4992
rect 19394 4936 19399 4992
rect 16389 4934 19399 4936
rect 16389 4931 16455 4934
rect 19333 4931 19399 4934
rect 22737 4994 22803 4997
rect 23289 4994 23355 4997
rect 22737 4992 23355 4994
rect 22737 4936 22742 4992
rect 22798 4936 23294 4992
rect 23350 4936 23355 4992
rect 22737 4934 23355 4936
rect 22737 4931 22803 4934
rect 23289 4931 23355 4934
rect 25773 4994 25839 4997
rect 27520 4994 28000 5024
rect 25773 4992 28000 4994
rect 25773 4936 25778 4992
rect 25834 4936 28000 4992
rect 25773 4934 28000 4936
rect 25773 4931 25839 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 27520 4904 28000 4934
rect 19610 4863 19930 4864
rect 16982 4796 16988 4860
rect 17052 4858 17058 4860
rect 19241 4858 19307 4861
rect 17052 4856 19307 4858
rect 17052 4800 19246 4856
rect 19302 4800 19307 4856
rect 17052 4798 19307 4800
rect 17052 4796 17058 4798
rect 19241 4795 19307 4798
rect 11329 4722 11395 4725
rect 16757 4722 16823 4725
rect 11329 4720 16823 4722
rect 11329 4664 11334 4720
rect 11390 4664 16762 4720
rect 16818 4664 16823 4720
rect 11329 4662 16823 4664
rect 11329 4659 11395 4662
rect 16757 4659 16823 4662
rect 18413 4722 18479 4725
rect 21449 4722 21515 4725
rect 18413 4720 21515 4722
rect 18413 4664 18418 4720
rect 18474 4664 21454 4720
rect 21510 4664 21515 4720
rect 18413 4662 21515 4664
rect 18413 4659 18479 4662
rect 21449 4659 21515 4662
rect 657 4586 723 4589
rect 8477 4586 8543 4589
rect 657 4584 8543 4586
rect 657 4528 662 4584
rect 718 4528 8482 4584
rect 8538 4528 8543 4584
rect 657 4526 8543 4528
rect 657 4523 723 4526
rect 8477 4523 8543 4526
rect 8661 4586 8727 4589
rect 11881 4586 11947 4589
rect 8661 4584 11947 4586
rect 8661 4528 8666 4584
rect 8722 4528 11886 4584
rect 11942 4528 11947 4584
rect 8661 4526 11947 4528
rect 8661 4523 8727 4526
rect 11881 4523 11947 4526
rect 14089 4586 14155 4589
rect 16665 4586 16731 4589
rect 17585 4586 17651 4589
rect 17861 4586 17927 4589
rect 14089 4584 15578 4586
rect 14089 4528 14094 4584
rect 14150 4528 15578 4584
rect 14089 4526 15578 4528
rect 14089 4523 14155 4526
rect 0 4450 480 4480
rect 1853 4450 1919 4453
rect 0 4448 1919 4450
rect 0 4392 1858 4448
rect 1914 4392 1919 4448
rect 0 4390 1919 4392
rect 0 4360 480 4390
rect 1853 4387 1919 4390
rect 4521 4450 4587 4453
rect 4654 4450 4660 4452
rect 4521 4448 4660 4450
rect 4521 4392 4526 4448
rect 4582 4392 4660 4448
rect 4521 4390 4660 4392
rect 4521 4387 4587 4390
rect 4654 4388 4660 4390
rect 4724 4388 4730 4452
rect 7465 4450 7531 4453
rect 11462 4450 11468 4452
rect 7465 4448 11468 4450
rect 7465 4392 7470 4448
rect 7526 4392 11468 4448
rect 7465 4390 11468 4392
rect 7465 4387 7531 4390
rect 11462 4388 11468 4390
rect 11532 4388 11538 4452
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 1393 4314 1459 4317
rect 5257 4314 5323 4317
rect 1393 4312 5323 4314
rect 1393 4256 1398 4312
rect 1454 4256 5262 4312
rect 5318 4256 5323 4312
rect 1393 4254 5323 4256
rect 1393 4251 1459 4254
rect 5257 4251 5323 4254
rect 8937 4314 9003 4317
rect 11881 4314 11947 4317
rect 15518 4314 15578 4526
rect 16665 4584 17927 4586
rect 16665 4528 16670 4584
rect 16726 4528 17590 4584
rect 17646 4528 17866 4584
rect 17922 4528 17927 4584
rect 16665 4526 17927 4528
rect 16665 4523 16731 4526
rect 17585 4523 17651 4526
rect 17861 4523 17927 4526
rect 18321 4586 18387 4589
rect 21725 4586 21791 4589
rect 18321 4584 21791 4586
rect 18321 4528 18326 4584
rect 18382 4528 21730 4584
rect 21786 4528 21791 4584
rect 18321 4526 21791 4528
rect 18321 4523 18387 4526
rect 21725 4523 21791 4526
rect 22686 4524 22692 4588
rect 22756 4586 22762 4588
rect 22829 4586 22895 4589
rect 22756 4584 22895 4586
rect 22756 4528 22834 4584
rect 22890 4528 22895 4584
rect 22756 4526 22895 4528
rect 22756 4524 22762 4526
rect 22829 4523 22895 4526
rect 23016 4526 24732 4586
rect 15653 4450 15719 4453
rect 19977 4450 20043 4453
rect 15653 4448 20043 4450
rect 15653 4392 15658 4448
rect 15714 4392 19982 4448
rect 20038 4392 20043 4448
rect 15653 4390 20043 4392
rect 15653 4387 15719 4390
rect 19977 4387 20043 4390
rect 22277 4450 22343 4453
rect 23016 4450 23076 4526
rect 22277 4448 23076 4450
rect 22277 4392 22282 4448
rect 22338 4392 23076 4448
rect 22277 4390 23076 4392
rect 24672 4450 24732 4526
rect 27520 4450 28000 4480
rect 24672 4390 28000 4450
rect 22277 4387 22343 4390
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 27520 4360 28000 4390
rect 24277 4319 24597 4320
rect 23933 4314 23999 4317
rect 8937 4312 14658 4314
rect 8937 4256 8942 4312
rect 8998 4256 11886 4312
rect 11942 4256 14658 4312
rect 8937 4254 14658 4256
rect 15518 4312 23999 4314
rect 15518 4256 23938 4312
rect 23994 4256 23999 4312
rect 15518 4254 23999 4256
rect 8937 4251 9003 4254
rect 11881 4251 11947 4254
rect 6085 4178 6151 4181
rect 9857 4178 9923 4181
rect 6085 4176 9923 4178
rect 6085 4120 6090 4176
rect 6146 4120 9862 4176
rect 9918 4120 9923 4176
rect 6085 4118 9923 4120
rect 14598 4178 14658 4254
rect 23933 4251 23999 4254
rect 18229 4178 18295 4181
rect 14598 4176 18295 4178
rect 14598 4120 18234 4176
rect 18290 4120 18295 4176
rect 14598 4118 18295 4120
rect 6085 4115 6151 4118
rect 9857 4115 9923 4118
rect 18229 4115 18295 4118
rect 19149 4178 19215 4181
rect 25221 4178 25287 4181
rect 19149 4176 19626 4178
rect 19149 4120 19154 4176
rect 19210 4120 19626 4176
rect 19149 4118 19626 4120
rect 19149 4115 19215 4118
rect 3693 4042 3759 4045
rect 11605 4042 11671 4045
rect 3693 4040 11671 4042
rect 3693 3984 3698 4040
rect 3754 3984 11610 4040
rect 11666 3984 11671 4040
rect 3693 3982 11671 3984
rect 3693 3979 3759 3982
rect 11605 3979 11671 3982
rect 13854 3980 13860 4044
rect 13924 4042 13930 4044
rect 13997 4042 14063 4045
rect 13924 4040 14063 4042
rect 13924 3984 14002 4040
rect 14058 3984 14063 4040
rect 13924 3982 14063 3984
rect 13924 3980 13930 3982
rect 13997 3979 14063 3982
rect 14825 4042 14891 4045
rect 19333 4042 19399 4045
rect 14825 4040 19399 4042
rect 14825 3984 14830 4040
rect 14886 3984 19338 4040
rect 19394 3984 19399 4040
rect 14825 3982 19399 3984
rect 19566 4042 19626 4118
rect 22004 4176 25287 4178
rect 22004 4120 25226 4176
rect 25282 4120 25287 4176
rect 22004 4118 25287 4120
rect 20437 4042 20503 4045
rect 19566 4040 20503 4042
rect 19566 3984 20442 4040
rect 20498 3984 20503 4040
rect 19566 3982 20503 3984
rect 14825 3979 14891 3982
rect 19333 3979 19399 3982
rect 20437 3979 20503 3982
rect 20989 4042 21055 4045
rect 22004 4042 22064 4118
rect 25221 4115 25287 4118
rect 20989 4040 22064 4042
rect 20989 3984 20994 4040
rect 21050 3984 22064 4040
rect 20989 3982 22064 3984
rect 20989 3979 21055 3982
rect 23054 3980 23060 4044
rect 23124 4042 23130 4044
rect 24669 4042 24735 4045
rect 25405 4042 25471 4045
rect 23124 3982 24594 4042
rect 23124 3980 23130 3982
rect 3049 3906 3115 3909
rect 9121 3906 9187 3909
rect 3049 3904 9187 3906
rect 3049 3848 3054 3904
rect 3110 3848 9126 3904
rect 9182 3848 9187 3904
rect 3049 3846 9187 3848
rect 3049 3843 3115 3846
rect 9121 3843 9187 3846
rect 11421 3906 11487 3909
rect 13670 3906 13676 3908
rect 11421 3904 13676 3906
rect 11421 3848 11426 3904
rect 11482 3848 13676 3904
rect 11421 3846 13676 3848
rect 11421 3843 11487 3846
rect 13670 3844 13676 3846
rect 13740 3844 13746 3908
rect 14089 3906 14155 3909
rect 14406 3906 14412 3908
rect 14089 3904 14412 3906
rect 14089 3848 14094 3904
rect 14150 3848 14412 3904
rect 14089 3846 14412 3848
rect 14089 3843 14155 3846
rect 14406 3844 14412 3846
rect 14476 3844 14482 3908
rect 14733 3906 14799 3909
rect 18413 3906 18479 3909
rect 14733 3904 18479 3906
rect 14733 3848 14738 3904
rect 14794 3848 18418 3904
rect 18474 3848 18479 3904
rect 14733 3846 18479 3848
rect 14733 3843 14799 3846
rect 18413 3843 18479 3846
rect 20713 3906 20779 3909
rect 23657 3906 23723 3909
rect 20713 3904 23723 3906
rect 20713 3848 20718 3904
rect 20774 3848 23662 3904
rect 23718 3848 23723 3904
rect 20713 3846 23723 3848
rect 20713 3843 20779 3846
rect 23657 3843 23723 3846
rect 23974 3844 23980 3908
rect 24044 3906 24050 3908
rect 24393 3906 24459 3909
rect 24044 3904 24459 3906
rect 24044 3848 24398 3904
rect 24454 3848 24459 3904
rect 24044 3846 24459 3848
rect 24534 3906 24594 3982
rect 24669 4040 25471 4042
rect 24669 3984 24674 4040
rect 24730 3984 25410 4040
rect 25466 3984 25471 4040
rect 24669 3982 25471 3984
rect 24669 3979 24735 3982
rect 25405 3979 25471 3982
rect 24534 3846 25146 3906
rect 24044 3844 24050 3846
rect 24393 3843 24459 3846
rect 10277 3840 10597 3841
rect 0 3770 480 3800
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 1761 3770 1827 3773
rect 0 3768 1827 3770
rect 0 3712 1766 3768
rect 1822 3712 1827 3768
rect 0 3710 1827 3712
rect 0 3680 480 3710
rect 1761 3707 1827 3710
rect 2957 3770 3023 3773
rect 9581 3770 9647 3773
rect 9949 3770 10015 3773
rect 2957 3768 10015 3770
rect 2957 3712 2962 3768
rect 3018 3712 9586 3768
rect 9642 3712 9954 3768
rect 10010 3712 10015 3768
rect 2957 3710 10015 3712
rect 2957 3707 3023 3710
rect 9581 3707 9647 3710
rect 9949 3707 10015 3710
rect 12198 3708 12204 3772
rect 12268 3770 12274 3772
rect 12801 3770 12867 3773
rect 16757 3772 16823 3773
rect 16757 3770 16804 3772
rect 12268 3768 12867 3770
rect 12268 3712 12806 3768
rect 12862 3712 12867 3768
rect 12268 3710 12867 3712
rect 16712 3768 16804 3770
rect 16712 3712 16762 3768
rect 16712 3710 16804 3712
rect 12268 3708 12274 3710
rect 12801 3707 12867 3710
rect 16757 3708 16804 3710
rect 16868 3708 16874 3772
rect 17309 3770 17375 3773
rect 19149 3770 19215 3773
rect 17309 3768 19215 3770
rect 17309 3712 17314 3768
rect 17370 3712 19154 3768
rect 19210 3712 19215 3768
rect 17309 3710 19215 3712
rect 16757 3707 16823 3708
rect 17309 3707 17375 3710
rect 19149 3707 19215 3710
rect 22645 3770 22711 3773
rect 24945 3770 25011 3773
rect 22645 3768 25011 3770
rect 22645 3712 22650 3768
rect 22706 3712 24950 3768
rect 25006 3712 25011 3768
rect 22645 3710 25011 3712
rect 25086 3770 25146 3846
rect 27520 3770 28000 3800
rect 25086 3710 28000 3770
rect 22645 3707 22711 3710
rect 24945 3707 25011 3710
rect 27520 3680 28000 3710
rect 8293 3634 8359 3637
rect 12065 3634 12131 3637
rect 21357 3634 21423 3637
rect 24577 3634 24643 3637
rect 8293 3632 21423 3634
rect 8293 3576 8298 3632
rect 8354 3576 12070 3632
rect 12126 3576 21362 3632
rect 21418 3576 21423 3632
rect 8293 3574 21423 3576
rect 8293 3571 8359 3574
rect 12065 3571 12131 3574
rect 21357 3571 21423 3574
rect 21590 3632 24643 3634
rect 21590 3576 24582 3632
rect 24638 3576 24643 3632
rect 21590 3574 24643 3576
rect 2865 3498 2931 3501
rect 4797 3498 4863 3501
rect 8661 3498 8727 3501
rect 2865 3496 8727 3498
rect 2865 3440 2870 3496
rect 2926 3440 4802 3496
rect 4858 3440 8666 3496
rect 8722 3440 8727 3496
rect 2865 3438 8727 3440
rect 2865 3435 2931 3438
rect 4797 3435 4863 3438
rect 8661 3435 8727 3438
rect 13261 3498 13327 3501
rect 18045 3498 18111 3501
rect 13261 3496 18111 3498
rect 13261 3440 13266 3496
rect 13322 3440 18050 3496
rect 18106 3440 18111 3496
rect 13261 3438 18111 3440
rect 13261 3435 13327 3438
rect 18045 3435 18111 3438
rect 18965 3498 19031 3501
rect 21590 3498 21650 3574
rect 24577 3571 24643 3574
rect 18965 3496 21650 3498
rect 18965 3440 18970 3496
rect 19026 3440 21650 3496
rect 18965 3438 21650 3440
rect 22553 3498 22619 3501
rect 25405 3498 25471 3501
rect 27613 3498 27679 3501
rect 22553 3496 24732 3498
rect 22553 3440 22558 3496
rect 22614 3440 24732 3496
rect 22553 3438 24732 3440
rect 18965 3435 19031 3438
rect 22553 3435 22619 3438
rect 6361 3362 6427 3365
rect 18689 3362 18755 3365
rect 22461 3362 22527 3365
rect 6361 3360 11300 3362
rect 6361 3304 6366 3360
rect 6422 3304 11300 3360
rect 6361 3302 11300 3304
rect 6361 3299 6427 3302
rect 5610 3296 5930 3297
rect 0 3226 480 3256
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 1577 3226 1643 3229
rect 0 3224 1643 3226
rect 0 3168 1582 3224
rect 1638 3168 1643 3224
rect 0 3166 1643 3168
rect 0 3136 480 3166
rect 1577 3163 1643 3166
rect 6085 3226 6151 3229
rect 7925 3226 7991 3229
rect 6085 3224 7991 3226
rect 6085 3168 6090 3224
rect 6146 3168 7930 3224
rect 7986 3168 7991 3224
rect 6085 3166 7991 3168
rect 6085 3163 6151 3166
rect 7925 3163 7991 3166
rect 10133 3226 10199 3229
rect 11053 3226 11119 3229
rect 10133 3224 11119 3226
rect 10133 3168 10138 3224
rect 10194 3168 11058 3224
rect 11114 3168 11119 3224
rect 10133 3166 11119 3168
rect 11240 3226 11300 3302
rect 18689 3360 22527 3362
rect 18689 3304 18694 3360
rect 18750 3304 22466 3360
rect 22522 3304 22527 3360
rect 18689 3302 22527 3304
rect 18689 3299 18755 3302
rect 22461 3299 22527 3302
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 13445 3226 13511 3229
rect 13997 3226 14063 3229
rect 11240 3224 14063 3226
rect 11240 3168 13450 3224
rect 13506 3168 14002 3224
rect 14058 3168 14063 3224
rect 11240 3166 14063 3168
rect 10133 3163 10199 3166
rect 11053 3163 11119 3166
rect 13445 3163 13511 3166
rect 13997 3163 14063 3166
rect 18873 3226 18939 3229
rect 21173 3226 21239 3229
rect 18873 3224 21239 3226
rect 18873 3168 18878 3224
rect 18934 3168 21178 3224
rect 21234 3168 21239 3224
rect 18873 3166 21239 3168
rect 24672 3226 24732 3438
rect 25405 3496 27679 3498
rect 25405 3440 25410 3496
rect 25466 3440 27618 3496
rect 27674 3440 27679 3496
rect 25405 3438 27679 3440
rect 25405 3435 25471 3438
rect 27613 3435 27679 3438
rect 27520 3226 28000 3256
rect 24672 3166 28000 3226
rect 18873 3163 18939 3166
rect 21173 3163 21239 3166
rect 27520 3136 28000 3166
rect 1853 3090 1919 3093
rect 6361 3090 6427 3093
rect 1853 3088 6427 3090
rect 1853 3032 1858 3088
rect 1914 3032 6366 3088
rect 6422 3032 6427 3088
rect 1853 3030 6427 3032
rect 1853 3027 1919 3030
rect 6361 3027 6427 3030
rect 9213 3090 9279 3093
rect 11278 3090 11284 3092
rect 9213 3088 11284 3090
rect 9213 3032 9218 3088
rect 9274 3032 11284 3088
rect 9213 3030 11284 3032
rect 9213 3027 9279 3030
rect 11278 3028 11284 3030
rect 11348 3090 11354 3092
rect 13445 3090 13511 3093
rect 11348 3088 13511 3090
rect 11348 3032 13450 3088
rect 13506 3032 13511 3088
rect 11348 3030 13511 3032
rect 11348 3028 11354 3030
rect 13445 3027 13511 3030
rect 18137 3090 18203 3093
rect 19885 3090 19951 3093
rect 18137 3088 19951 3090
rect 18137 3032 18142 3088
rect 18198 3032 19890 3088
rect 19946 3032 19951 3088
rect 18137 3030 19951 3032
rect 18137 3027 18203 3030
rect 19885 3027 19951 3030
rect 20069 3090 20135 3093
rect 23657 3090 23723 3093
rect 20069 3088 23723 3090
rect 20069 3032 20074 3088
rect 20130 3032 23662 3088
rect 23718 3032 23723 3088
rect 20069 3030 23723 3032
rect 20069 3027 20135 3030
rect 23657 3027 23723 3030
rect 23790 3028 23796 3092
rect 23860 3090 23866 3092
rect 24025 3090 24091 3093
rect 23860 3088 24091 3090
rect 23860 3032 24030 3088
rect 24086 3032 24091 3088
rect 23860 3030 24091 3032
rect 23860 3028 23866 3030
rect 24025 3027 24091 3030
rect 3969 2954 4035 2957
rect 9673 2954 9739 2957
rect 13905 2954 13971 2957
rect 17769 2954 17835 2957
rect 3969 2952 9739 2954
rect 3969 2896 3974 2952
rect 4030 2896 9678 2952
rect 9734 2896 9739 2952
rect 3969 2894 9739 2896
rect 3969 2891 4035 2894
rect 9673 2891 9739 2894
rect 13862 2952 17835 2954
rect 13862 2896 13910 2952
rect 13966 2896 17774 2952
rect 17830 2896 17835 2952
rect 13862 2894 17835 2896
rect 13862 2891 13971 2894
rect 17769 2891 17835 2894
rect 19057 2954 19123 2957
rect 21541 2954 21607 2957
rect 19057 2952 21607 2954
rect 19057 2896 19062 2952
rect 19118 2896 21546 2952
rect 21602 2896 21607 2952
rect 19057 2894 21607 2896
rect 19057 2891 19123 2894
rect 21541 2891 21607 2894
rect 21766 2892 21772 2956
rect 21836 2954 21842 2956
rect 22093 2954 22159 2957
rect 21836 2952 22159 2954
rect 21836 2896 22098 2952
rect 22154 2896 22159 2952
rect 21836 2894 22159 2896
rect 21836 2892 21842 2894
rect 22093 2891 22159 2894
rect 23422 2892 23428 2956
rect 23492 2954 23498 2956
rect 23749 2954 23815 2957
rect 23492 2952 23815 2954
rect 23492 2896 23754 2952
rect 23810 2896 23815 2952
rect 23492 2894 23815 2896
rect 23492 2892 23498 2894
rect 23749 2891 23815 2894
rect 10277 2752 10597 2753
rect 0 2682 480 2712
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 2405 2682 2471 2685
rect 0 2680 2471 2682
rect 0 2624 2410 2680
rect 2466 2624 2471 2680
rect 0 2622 2471 2624
rect 0 2592 480 2622
rect 2405 2619 2471 2622
rect 7465 2682 7531 2685
rect 10133 2682 10199 2685
rect 7465 2680 10199 2682
rect 7465 2624 7470 2680
rect 7526 2624 10138 2680
rect 10194 2624 10199 2680
rect 7465 2622 10199 2624
rect 7465 2619 7531 2622
rect 10133 2619 10199 2622
rect 10777 2682 10843 2685
rect 13862 2682 13922 2891
rect 15561 2818 15627 2821
rect 19425 2818 19491 2821
rect 15561 2816 19491 2818
rect 15561 2760 15566 2816
rect 15622 2760 19430 2816
rect 19486 2760 19491 2816
rect 15561 2758 19491 2760
rect 15561 2755 15627 2758
rect 19425 2755 19491 2758
rect 20069 2818 20135 2821
rect 22553 2818 22619 2821
rect 20069 2816 22619 2818
rect 20069 2760 20074 2816
rect 20130 2760 22558 2816
rect 22614 2760 22619 2816
rect 20069 2758 22619 2760
rect 20069 2755 20135 2758
rect 22553 2755 22619 2758
rect 23013 2818 23079 2821
rect 27061 2818 27127 2821
rect 23013 2816 27127 2818
rect 23013 2760 23018 2816
rect 23074 2760 27066 2816
rect 27122 2760 27127 2816
rect 23013 2758 27127 2760
rect 23013 2755 23079 2758
rect 27061 2755 27127 2758
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 10777 2680 13922 2682
rect 10777 2624 10782 2680
rect 10838 2624 13922 2680
rect 10777 2622 13922 2624
rect 14641 2682 14707 2685
rect 18321 2682 18387 2685
rect 14641 2680 18387 2682
rect 14641 2624 14646 2680
rect 14702 2624 18326 2680
rect 18382 2624 18387 2680
rect 14641 2622 18387 2624
rect 10777 2619 10843 2622
rect 14641 2619 14707 2622
rect 18321 2619 18387 2622
rect 24485 2682 24551 2685
rect 24710 2682 24716 2684
rect 24485 2680 24716 2682
rect 24485 2624 24490 2680
rect 24546 2624 24716 2680
rect 24485 2622 24716 2624
rect 24485 2619 24551 2622
rect 24710 2620 24716 2622
rect 24780 2620 24786 2684
rect 27520 2682 28000 2712
rect 26926 2622 28000 2682
rect 2313 2546 2379 2549
rect 8385 2546 8451 2549
rect 2313 2544 8451 2546
rect 2313 2488 2318 2544
rect 2374 2488 8390 2544
rect 8446 2488 8451 2544
rect 2313 2486 8451 2488
rect 2313 2483 2379 2486
rect 8385 2483 8451 2486
rect 9305 2546 9371 2549
rect 12617 2546 12683 2549
rect 9305 2544 12683 2546
rect 9305 2488 9310 2544
rect 9366 2488 12622 2544
rect 12678 2488 12683 2544
rect 9305 2486 12683 2488
rect 9305 2483 9371 2486
rect 12617 2483 12683 2486
rect 14457 2546 14523 2549
rect 14457 2544 15532 2546
rect 14457 2488 14462 2544
rect 14518 2488 15532 2544
rect 14457 2486 15532 2488
rect 14457 2483 14523 2486
rect 2405 2410 2471 2413
rect 4429 2410 4495 2413
rect 10961 2410 11027 2413
rect 2405 2408 4495 2410
rect 2405 2352 2410 2408
rect 2466 2352 4434 2408
rect 4490 2352 4495 2408
rect 2405 2350 4495 2352
rect 2405 2347 2471 2350
rect 4429 2347 4495 2350
rect 4662 2408 11027 2410
rect 4662 2352 10966 2408
rect 11022 2352 11027 2408
rect 4662 2350 11027 2352
rect 4245 2274 4311 2277
rect 4662 2274 4722 2350
rect 10961 2347 11027 2350
rect 12065 2410 12131 2413
rect 12709 2410 12775 2413
rect 14273 2410 14339 2413
rect 15472 2410 15532 2486
rect 16614 2484 16620 2548
rect 16684 2546 16690 2548
rect 18229 2546 18295 2549
rect 16684 2544 18295 2546
rect 16684 2488 18234 2544
rect 18290 2488 18295 2544
rect 16684 2486 18295 2488
rect 16684 2484 16690 2486
rect 18229 2483 18295 2486
rect 18413 2546 18479 2549
rect 21173 2546 21239 2549
rect 18413 2544 21239 2546
rect 18413 2488 18418 2544
rect 18474 2488 21178 2544
rect 21234 2488 21239 2544
rect 18413 2486 21239 2488
rect 18413 2483 18479 2486
rect 21173 2483 21239 2486
rect 21633 2546 21699 2549
rect 25589 2546 25655 2549
rect 21633 2544 25655 2546
rect 21633 2488 21638 2544
rect 21694 2488 25594 2544
rect 25650 2488 25655 2544
rect 21633 2486 25655 2488
rect 21633 2483 21699 2486
rect 25589 2483 25655 2486
rect 20529 2410 20595 2413
rect 12065 2408 15394 2410
rect 12065 2352 12070 2408
rect 12126 2352 12714 2408
rect 12770 2352 14278 2408
rect 14334 2352 15394 2408
rect 12065 2350 15394 2352
rect 15472 2408 20595 2410
rect 15472 2352 20534 2408
rect 20590 2352 20595 2408
rect 15472 2350 20595 2352
rect 12065 2347 12131 2350
rect 12709 2347 12775 2350
rect 14273 2347 14339 2350
rect 4245 2272 4722 2274
rect 4245 2216 4250 2272
rect 4306 2216 4722 2272
rect 4245 2214 4722 2216
rect 6545 2274 6611 2277
rect 13077 2274 13143 2277
rect 6545 2272 13143 2274
rect 6545 2216 6550 2272
rect 6606 2216 13082 2272
rect 13138 2216 13143 2272
rect 6545 2214 13143 2216
rect 15334 2274 15394 2350
rect 20529 2347 20595 2350
rect 23473 2410 23539 2413
rect 26926 2410 26986 2622
rect 27520 2592 28000 2622
rect 23473 2408 26986 2410
rect 23473 2352 23478 2408
rect 23534 2352 26986 2408
rect 23473 2350 26986 2352
rect 23473 2347 23539 2350
rect 16757 2274 16823 2277
rect 15334 2272 16823 2274
rect 15334 2216 16762 2272
rect 16818 2216 16823 2272
rect 15334 2214 16823 2216
rect 4245 2211 4311 2214
rect 6545 2211 6611 2214
rect 13077 2211 13143 2214
rect 16757 2211 16823 2214
rect 16941 2274 17007 2277
rect 19517 2274 19583 2277
rect 16941 2272 19583 2274
rect 16941 2216 16946 2272
rect 17002 2216 19522 2272
rect 19578 2216 19583 2272
rect 16941 2214 19583 2216
rect 16941 2211 17007 2214
rect 19517 2211 19583 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 6821 2138 6887 2141
rect 16665 2138 16731 2141
rect 23565 2138 23631 2141
rect 6821 2136 9874 2138
rect 6821 2080 6826 2136
rect 6882 2080 9874 2136
rect 6821 2078 9874 2080
rect 6821 2075 6887 2078
rect 0 2002 480 2032
rect 3693 2002 3759 2005
rect 0 2000 3759 2002
rect 0 1944 3698 2000
rect 3754 1944 3759 2000
rect 0 1942 3759 1944
rect 0 1912 480 1942
rect 3693 1939 3759 1942
rect 7189 2002 7255 2005
rect 9814 2002 9874 2078
rect 16665 2136 23631 2138
rect 16665 2080 16670 2136
rect 16726 2080 23570 2136
rect 23626 2080 23631 2136
rect 16665 2078 23631 2080
rect 16665 2075 16731 2078
rect 23565 2075 23631 2078
rect 18229 2002 18295 2005
rect 7189 2000 9690 2002
rect 7189 1944 7194 2000
rect 7250 1944 9690 2000
rect 7189 1942 9690 1944
rect 9814 2000 18295 2002
rect 9814 1944 18234 2000
rect 18290 1944 18295 2000
rect 9814 1942 18295 1944
rect 7189 1939 7255 1942
rect 9630 1866 9690 1942
rect 18229 1939 18295 1942
rect 18413 2002 18479 2005
rect 21081 2002 21147 2005
rect 18413 2000 21147 2002
rect 18413 1944 18418 2000
rect 18474 1944 21086 2000
rect 21142 1944 21147 2000
rect 18413 1942 21147 1944
rect 18413 1939 18479 1942
rect 21081 1939 21147 1942
rect 25865 2002 25931 2005
rect 27520 2002 28000 2032
rect 25865 2000 28000 2002
rect 25865 1944 25870 2000
rect 25926 1944 28000 2000
rect 25865 1942 28000 1944
rect 25865 1939 25931 1942
rect 27520 1912 28000 1942
rect 17677 1866 17743 1869
rect 9630 1864 17743 1866
rect 9630 1808 17682 1864
rect 17738 1808 17743 1864
rect 9630 1806 17743 1808
rect 17677 1803 17743 1806
rect 18505 1866 18571 1869
rect 25497 1866 25563 1869
rect 18505 1864 25563 1866
rect 18505 1808 18510 1864
rect 18566 1808 25502 1864
rect 25558 1808 25563 1864
rect 18505 1806 25563 1808
rect 18505 1803 18571 1806
rect 25497 1803 25563 1806
rect 2865 1730 2931 1733
rect 9305 1730 9371 1733
rect 2865 1728 9371 1730
rect 2865 1672 2870 1728
rect 2926 1672 9310 1728
rect 9366 1672 9371 1728
rect 2865 1670 9371 1672
rect 2865 1667 2931 1670
rect 9305 1667 9371 1670
rect 13997 1730 14063 1733
rect 20897 1730 20963 1733
rect 13997 1728 20963 1730
rect 13997 1672 14002 1728
rect 14058 1672 20902 1728
rect 20958 1672 20963 1728
rect 13997 1670 20963 1672
rect 13997 1667 14063 1670
rect 20897 1667 20963 1670
rect 21081 1730 21147 1733
rect 24710 1730 24716 1732
rect 21081 1728 24716 1730
rect 21081 1672 21086 1728
rect 21142 1672 24716 1728
rect 21081 1670 24716 1672
rect 21081 1667 21147 1670
rect 24710 1668 24716 1670
rect 24780 1668 24786 1732
rect 7557 1594 7623 1597
rect 16614 1594 16620 1596
rect 7557 1592 16620 1594
rect 7557 1536 7562 1592
rect 7618 1536 16620 1592
rect 7557 1534 16620 1536
rect 7557 1531 7623 1534
rect 16614 1532 16620 1534
rect 16684 1532 16690 1596
rect 16757 1594 16823 1597
rect 20253 1594 20319 1597
rect 16757 1592 20319 1594
rect 16757 1536 16762 1592
rect 16818 1536 20258 1592
rect 20314 1536 20319 1592
rect 16757 1534 20319 1536
rect 16757 1531 16823 1534
rect 20253 1531 20319 1534
rect 23933 1594 23999 1597
rect 23933 1592 26986 1594
rect 23933 1536 23938 1592
rect 23994 1536 26986 1592
rect 23933 1534 26986 1536
rect 23933 1531 23999 1534
rect 0 1458 480 1488
rect 1761 1458 1827 1461
rect 0 1456 1827 1458
rect 0 1400 1766 1456
rect 1822 1400 1827 1456
rect 0 1398 1827 1400
rect 0 1368 480 1398
rect 1761 1395 1827 1398
rect 7598 1396 7604 1460
rect 7668 1458 7674 1460
rect 7741 1458 7807 1461
rect 7668 1456 7807 1458
rect 7668 1400 7746 1456
rect 7802 1400 7807 1456
rect 7668 1398 7807 1400
rect 7668 1396 7674 1398
rect 7741 1395 7807 1398
rect 12985 1458 13051 1461
rect 19793 1458 19859 1461
rect 12985 1456 19859 1458
rect 12985 1400 12990 1456
rect 13046 1400 19798 1456
rect 19854 1400 19859 1456
rect 12985 1398 19859 1400
rect 12985 1395 13051 1398
rect 19793 1395 19859 1398
rect 20161 1458 20227 1461
rect 26509 1458 26575 1461
rect 20161 1456 26575 1458
rect 20161 1400 20166 1456
rect 20222 1400 26514 1456
rect 26570 1400 26575 1456
rect 20161 1398 26575 1400
rect 26926 1458 26986 1534
rect 27520 1458 28000 1488
rect 26926 1398 28000 1458
rect 20161 1395 20227 1398
rect 26509 1395 26575 1398
rect 27520 1368 28000 1398
rect 2773 1322 2839 1325
rect 17585 1322 17651 1325
rect 2773 1320 17651 1322
rect 2773 1264 2778 1320
rect 2834 1264 17590 1320
rect 17646 1264 17651 1320
rect 2773 1262 17651 1264
rect 2773 1259 2839 1262
rect 17585 1259 17651 1262
rect 13445 1186 13511 1189
rect 20989 1186 21055 1189
rect 13445 1184 21055 1186
rect 13445 1128 13450 1184
rect 13506 1128 20994 1184
rect 21050 1128 21055 1184
rect 13445 1126 21055 1128
rect 13445 1123 13511 1126
rect 20989 1123 21055 1126
rect 15878 988 15884 1052
rect 15948 1050 15954 1052
rect 24209 1050 24275 1053
rect 15948 1048 24275 1050
rect 15948 992 24214 1048
rect 24270 992 24275 1048
rect 15948 990 24275 992
rect 15948 988 15954 990
rect 24209 987 24275 990
rect 0 914 480 944
rect 1669 914 1735 917
rect 0 912 1735 914
rect 0 856 1674 912
rect 1730 856 1735 912
rect 0 854 1735 856
rect 0 824 480 854
rect 1669 851 1735 854
rect 23841 914 23907 917
rect 27520 914 28000 944
rect 23841 912 28000 914
rect 23841 856 23846 912
rect 23902 856 28000 912
rect 23841 854 28000 856
rect 23841 851 23907 854
rect 27520 824 28000 854
rect 0 370 480 400
rect 3141 370 3207 373
rect 0 368 3207 370
rect 0 312 3146 368
rect 3202 312 3207 368
rect 0 310 3207 312
rect 0 280 480 310
rect 3141 307 3207 310
rect 24025 370 24091 373
rect 27520 370 28000 400
rect 24025 368 28000 370
rect 24025 312 24030 368
rect 24086 312 28000 368
rect 24025 310 28000 312
rect 24025 307 24091 310
rect 27520 280 28000 310
rect 14181 98 14247 101
rect 20897 98 20963 101
rect 14181 96 20963 98
rect 14181 40 14186 96
rect 14242 40 20902 96
rect 20958 40 20963 96
rect 14181 38 20963 40
rect 14181 35 14247 38
rect 20897 35 20963 38
<< via3 >>
rect 8340 26284 8404 26348
rect 8340 25876 8404 25940
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 15884 24788 15948 24852
rect 11100 24712 11164 24716
rect 11100 24656 11150 24712
rect 11150 24656 11164 24712
rect 11100 24652 11164 24656
rect 11284 24576 11348 24580
rect 11284 24520 11298 24576
rect 11298 24520 11348 24576
rect 11284 24516 11348 24520
rect 20484 24516 20548 24580
rect 21956 24516 22020 24580
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 12572 24108 12636 24172
rect 12020 23972 12084 24036
rect 23796 24168 23860 24172
rect 23796 24112 23846 24168
rect 23846 24112 23860 24168
rect 23796 24108 23860 24112
rect 15516 23972 15580 24036
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 14780 23836 14844 23900
rect 16804 23700 16868 23764
rect 13860 23564 13924 23628
rect 16252 23564 16316 23628
rect 24716 23564 24780 23628
rect 15332 23488 15396 23492
rect 15332 23432 15346 23488
rect 15346 23432 15396 23488
rect 15332 23428 15396 23432
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 6132 23292 6196 23356
rect 11468 23292 11532 23356
rect 19380 23488 19444 23492
rect 19380 23432 19430 23488
rect 19430 23432 19444 23488
rect 19380 23428 19444 23432
rect 20116 23488 20180 23492
rect 20116 23432 20130 23488
rect 20130 23432 20180 23488
rect 20116 23428 20180 23432
rect 24900 23428 24964 23492
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 23428 23020 23492 23084
rect 23612 22884 23676 22948
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 23060 22748 23124 22812
rect 19196 22612 19260 22676
rect 2452 22264 2516 22268
rect 2452 22208 2466 22264
rect 2466 22208 2516 22264
rect 2452 22204 2516 22208
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 9628 22204 9692 22268
rect 13676 22264 13740 22268
rect 13676 22208 13726 22264
rect 13726 22208 13740 22264
rect 13676 22204 13740 22208
rect 14780 22204 14844 22268
rect 12020 22068 12084 22132
rect 12572 21992 12636 21996
rect 12572 21936 12622 21992
rect 12622 21936 12636 21992
rect 12572 21932 12636 21936
rect 13308 21796 13372 21860
rect 19196 21932 19260 21996
rect 20484 21796 20548 21860
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 19380 21388 19444 21452
rect 20852 21448 20916 21452
rect 20852 21392 20902 21448
rect 20902 21392 20916 21448
rect 20852 21388 20916 21392
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 17172 21116 17236 21180
rect 12204 20708 12268 20772
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 9996 20088 10060 20092
rect 9996 20032 10010 20088
rect 10010 20032 10060 20088
rect 9996 20028 10060 20032
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24900 19620 24964 19684
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 18276 19484 18340 19548
rect 25084 19484 25148 19548
rect 10916 19212 10980 19276
rect 11836 19136 11900 19140
rect 11836 19080 11886 19136
rect 11886 19080 11900 19136
rect 11836 19076 11900 19080
rect 12940 19076 13004 19140
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 16436 18804 16500 18868
rect 23980 18804 24044 18868
rect 22876 18668 22940 18732
rect 2636 18532 2700 18596
rect 11652 18592 11716 18596
rect 11652 18536 11702 18592
rect 11702 18536 11716 18592
rect 11652 18532 11716 18536
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 20852 18124 20916 18188
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 13124 17852 13188 17916
rect 20484 17852 20548 17916
rect 22508 17912 22572 17916
rect 22508 17856 22522 17912
rect 22522 17856 22572 17912
rect 22508 17852 22572 17856
rect 5212 17776 5276 17780
rect 5212 17720 5226 17776
rect 5226 17720 5276 17776
rect 5212 17716 5276 17720
rect 10732 17716 10796 17780
rect 20668 17716 20732 17780
rect 7788 17444 7852 17508
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 13676 17368 13740 17372
rect 13676 17312 13690 17368
rect 13690 17312 13740 17368
rect 13676 17308 13740 17312
rect 23244 17368 23308 17372
rect 23244 17312 23294 17368
rect 23294 17312 23308 17368
rect 23244 17308 23308 17312
rect 25084 17308 25148 17372
rect 23428 17172 23492 17236
rect 16620 16900 16684 16964
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 8892 16628 8956 16692
rect 13492 16628 13556 16692
rect 8524 16492 8588 16556
rect 9996 16356 10060 16420
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 1532 16144 1596 16148
rect 1532 16088 1546 16144
rect 1546 16088 1596 16144
rect 1532 16084 1596 16088
rect 12756 16220 12820 16284
rect 14780 16220 14844 16284
rect 17908 15948 17972 16012
rect 20668 15948 20732 16012
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 24900 16220 24964 16284
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 9444 15540 9508 15604
rect 12940 15540 13004 15604
rect 23980 15812 24044 15876
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 23244 15676 23308 15740
rect 23428 15676 23492 15740
rect 23796 15676 23860 15740
rect 23980 15404 24044 15468
rect 6868 15328 6932 15332
rect 6868 15272 6882 15328
rect 6882 15272 6932 15328
rect 6868 15268 6932 15272
rect 16252 15328 16316 15332
rect 16252 15272 16302 15328
rect 16302 15272 16316 15328
rect 16252 15268 16316 15272
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 14596 14996 14660 15060
rect 8708 14860 8772 14924
rect 1900 14588 1964 14652
rect 8524 14588 8588 14652
rect 8708 14588 8772 14652
rect 9996 14724 10060 14788
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 9812 14316 9876 14380
rect 14228 14724 14292 14788
rect 14780 14724 14844 14788
rect 23980 14860 24044 14924
rect 24716 14860 24780 14924
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 14412 14316 14476 14380
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 11652 14044 11716 14108
rect 20668 13968 20732 13972
rect 20668 13912 20718 13968
rect 20718 13912 20732 13968
rect 20668 13908 20732 13912
rect 9444 13772 9508 13836
rect 17356 13772 17420 13836
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 7420 13560 7484 13564
rect 7420 13504 7434 13560
rect 7434 13504 7484 13560
rect 7420 13500 7484 13504
rect 9260 13500 9324 13564
rect 9996 13500 10060 13564
rect 14596 13364 14660 13428
rect 21036 13500 21100 13564
rect 24716 13500 24780 13564
rect 1900 13228 1964 13292
rect 3740 13228 3804 13292
rect 12572 13152 12636 13156
rect 12572 13096 12622 13152
rect 12622 13096 12636 13152
rect 12572 13092 12636 13096
rect 20668 13092 20732 13156
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 1532 12956 1596 13020
rect 10916 13016 10980 13020
rect 10916 12960 10966 13016
rect 10966 12960 10980 13016
rect 1900 12684 1964 12748
rect 10916 12956 10980 12960
rect 13308 12956 13372 13020
rect 20300 12820 20364 12884
rect 3372 12548 3436 12612
rect 9260 12548 9324 12612
rect 12756 12548 12820 12612
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 9812 12412 9876 12476
rect 15884 12684 15948 12748
rect 15332 12548 15396 12612
rect 15884 12548 15948 12612
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 16436 12412 16500 12476
rect 1900 12336 1964 12340
rect 1900 12280 1950 12336
rect 1950 12280 1964 12336
rect 1900 12276 1964 12280
rect 9628 12276 9692 12340
rect 21036 12412 21100 12476
rect 3740 12200 3804 12204
rect 3740 12144 3790 12200
rect 3790 12144 3804 12200
rect 3740 12140 3804 12144
rect 6500 12140 6564 12204
rect 13492 12140 13556 12204
rect 6868 12004 6932 12068
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 7788 11732 7852 11796
rect 13124 11732 13188 11796
rect 24900 12004 24964 12068
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 25820 11732 25884 11796
rect 5212 11596 5276 11660
rect 6868 11596 6932 11660
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 13492 11324 13556 11388
rect 6500 11188 6564 11252
rect 24716 11460 24780 11524
rect 23612 11052 23676 11116
rect 9260 10916 9324 10980
rect 16436 10916 16500 10980
rect 22508 10916 22572 10980
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 24900 10780 24964 10844
rect 12572 10644 12636 10708
rect 13492 10644 13556 10708
rect 6684 10372 6748 10436
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 10732 10296 10796 10300
rect 10732 10240 10782 10296
rect 10782 10240 10796 10296
rect 10732 10236 10796 10240
rect 22692 10236 22756 10300
rect 24716 10236 24780 10300
rect 24900 10296 24964 10300
rect 24900 10240 24914 10296
rect 24914 10240 24964 10296
rect 24900 10236 24964 10240
rect 8892 9828 8956 9892
rect 14780 9828 14844 9892
rect 16252 9828 16316 9892
rect 22876 9828 22940 9892
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 6132 9420 6196 9484
rect 23428 9692 23492 9756
rect 24900 9752 24964 9756
rect 24900 9696 24914 9752
rect 24914 9696 24964 9752
rect 24900 9692 24964 9696
rect 16620 9556 16684 9620
rect 14780 9420 14844 9484
rect 23060 9420 23124 9484
rect 20300 9344 20364 9348
rect 20300 9288 20350 9344
rect 20350 9288 20364 9344
rect 20300 9284 20364 9288
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 15700 8876 15764 8940
rect 14412 8740 14476 8804
rect 16988 8740 17052 8804
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 2820 8604 2884 8668
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 23980 8604 24044 8668
rect 8892 8392 8956 8396
rect 8892 8336 8906 8392
rect 8906 8336 8956 8392
rect 8892 8332 8956 8336
rect 14596 8332 14660 8396
rect 23980 8332 24044 8396
rect 2452 8196 2516 8260
rect 7788 8196 7852 8260
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 15516 8060 15580 8124
rect 14780 7924 14844 7988
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 11836 7516 11900 7580
rect 23244 7788 23308 7852
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 3924 7244 3988 7308
rect 7788 7244 7852 7308
rect 13308 7108 13372 7172
rect 23796 7516 23860 7580
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 11836 6836 11900 6900
rect 3924 6700 3988 6764
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 19380 6836 19444 6900
rect 20300 6836 20364 6900
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 5396 6428 5460 6492
rect 17724 6488 17788 6492
rect 17724 6432 17774 6488
rect 17774 6432 17788 6488
rect 17724 6428 17788 6432
rect 20116 6428 20180 6492
rect 23796 6488 23860 6492
rect 23796 6432 23810 6488
rect 23810 6432 23860 6488
rect 23796 6428 23860 6432
rect 14780 6020 14844 6084
rect 20300 6020 20364 6084
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 11468 5944 11532 5948
rect 11468 5888 11518 5944
rect 11518 5888 11532 5944
rect 11468 5884 11532 5888
rect 11836 5884 11900 5948
rect 19196 5944 19260 5948
rect 19196 5888 19246 5944
rect 19246 5888 19260 5944
rect 19196 5884 19260 5888
rect 3004 5476 3068 5540
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 11468 5476 11532 5540
rect 7604 5340 7668 5404
rect 11100 5340 11164 5404
rect 16252 5476 16316 5540
rect 17540 5672 17604 5676
rect 17540 5616 17554 5672
rect 17554 5616 17604 5672
rect 17540 5612 17604 5616
rect 24900 5748 24964 5812
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 15700 5264 15764 5268
rect 15700 5208 15714 5264
rect 15714 5208 15764 5264
rect 15700 5204 15764 5208
rect 17356 5204 17420 5268
rect 21772 5204 21836 5268
rect 9444 5128 9508 5132
rect 9444 5072 9494 5128
rect 9494 5072 9508 5128
rect 9444 5068 9508 5072
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 16988 4796 17052 4860
rect 4660 4388 4724 4452
rect 11468 4388 11532 4452
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 22692 4524 22756 4588
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 13860 3980 13924 4044
rect 23060 3980 23124 4044
rect 13676 3844 13740 3908
rect 14412 3844 14476 3908
rect 23980 3844 24044 3908
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 12204 3708 12268 3772
rect 16804 3768 16868 3772
rect 16804 3712 16818 3768
rect 16818 3712 16868 3768
rect 16804 3708 16868 3712
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 11284 3028 11348 3092
rect 23796 3028 23860 3092
rect 21772 2892 21836 2956
rect 23428 2892 23492 2956
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 24716 2620 24780 2684
rect 16620 2484 16684 2548
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
rect 24716 1668 24780 1732
rect 16620 1532 16684 1596
rect 7604 1396 7668 1460
rect 15884 988 15948 1052
<< metal4 >>
rect 8339 26348 8405 26349
rect 8339 26284 8340 26348
rect 8404 26284 8405 26348
rect 8339 26283 8405 26284
rect 8342 25941 8402 26283
rect 8339 25940 8405 25941
rect 8339 25876 8340 25940
rect 8404 25876 8405 25940
rect 8339 25875 8405 25876
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 11099 24716 11165 24717
rect 11099 24652 11100 24716
rect 11164 24652 11165 24716
rect 11099 24651 11165 24652
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 6131 23356 6197 23357
rect 6131 23292 6132 23356
rect 6196 23292 6197 23356
rect 6131 23291 6197 23292
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 2451 22268 2517 22269
rect 2451 22204 2452 22268
rect 2516 22204 2517 22268
rect 2451 22203 2517 22204
rect 1531 16148 1597 16149
rect 1531 16084 1532 16148
rect 1596 16084 1597 16148
rect 1531 16083 1597 16084
rect 1534 13021 1594 16083
rect 1899 14652 1965 14653
rect 1899 14588 1900 14652
rect 1964 14588 1965 14652
rect 1899 14587 1965 14588
rect 1902 13293 1962 14587
rect 1899 13292 1965 13293
rect 1899 13228 1900 13292
rect 1964 13228 1965 13292
rect 1899 13227 1965 13228
rect 1531 13020 1597 13021
rect 1531 12956 1532 13020
rect 1596 12956 1597 13020
rect 1531 12955 1597 12956
rect 1899 12748 1965 12749
rect 1899 12684 1900 12748
rect 1964 12684 1965 12748
rect 1899 12683 1965 12684
rect 1902 12341 1962 12683
rect 1899 12340 1965 12341
rect 1899 12276 1900 12340
rect 1964 12276 1965 12340
rect 1899 12275 1965 12276
rect 2454 8261 2514 22203
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 2635 18596 2701 18597
rect 2635 18532 2636 18596
rect 2700 18532 2701 18596
rect 2635 18531 2701 18532
rect 2638 10570 2698 18531
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5211 17780 5277 17781
rect 5211 17716 5212 17780
rect 5276 17716 5277 17780
rect 5211 17715 5277 17716
rect 3739 13292 3805 13293
rect 3739 13228 3740 13292
rect 3804 13228 3805 13292
rect 3739 13227 3805 13228
rect 3374 12613 3434 13142
rect 3371 12612 3437 12613
rect 3371 12548 3372 12612
rect 3436 12548 3437 12612
rect 3371 12547 3437 12548
rect 3742 12205 3802 13227
rect 3739 12204 3805 12205
rect 3739 12140 3740 12204
rect 3804 12140 3805 12204
rect 3739 12139 3805 12140
rect 5214 11661 5274 17715
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5211 11660 5277 11661
rect 5211 11596 5212 11660
rect 5276 11596 5277 11660
rect 5211 11595 5277 11596
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 2638 10510 2882 10570
rect 2822 8669 2882 10510
rect 5610 9824 5931 10848
rect 6134 9978 6194 23291
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 9627 22268 9693 22269
rect 9627 22204 9628 22268
rect 9692 22204 9693 22268
rect 9627 22203 9693 22204
rect 9630 20178 9690 22203
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 9995 20092 10061 20093
rect 9995 20028 9996 20092
rect 10060 20028 10061 20092
rect 9995 20027 10061 20028
rect 7787 17508 7853 17509
rect 7787 17444 7788 17508
rect 7852 17444 7853 17508
rect 7787 17443 7853 17444
rect 6867 15332 6933 15333
rect 6867 15268 6868 15332
rect 6932 15268 6933 15332
rect 6867 15267 6933 15268
rect 6870 14058 6930 15267
rect 6499 12204 6565 12205
rect 6499 12140 6500 12204
rect 6564 12140 6565 12204
rect 6499 12139 6565 12140
rect 6502 12018 6562 12139
rect 6870 12069 6930 13822
rect 7422 13565 7482 15862
rect 7419 13564 7485 13565
rect 7419 13500 7420 13564
rect 7484 13500 7485 13564
rect 7419 13499 7485 13500
rect 6867 12068 6933 12069
rect 6867 12004 6868 12068
rect 6932 12004 6933 12068
rect 6867 12003 6933 12004
rect 7790 11797 7850 17443
rect 8891 16692 8957 16693
rect 8891 16628 8892 16692
rect 8956 16628 8957 16692
rect 8891 16627 8957 16628
rect 8523 16556 8589 16557
rect 8523 16492 8524 16556
rect 8588 16492 8589 16556
rect 8523 16491 8589 16492
rect 8526 14653 8586 16491
rect 8707 14924 8773 14925
rect 8707 14860 8708 14924
rect 8772 14860 8773 14924
rect 8707 14859 8773 14860
rect 8710 14653 8770 14859
rect 8523 14652 8589 14653
rect 8523 14588 8524 14652
rect 8588 14588 8589 14652
rect 8523 14587 8589 14588
rect 8707 14652 8773 14653
rect 8707 14588 8708 14652
rect 8772 14588 8773 14652
rect 8707 14587 8773 14588
rect 7787 11796 7853 11797
rect 6502 11253 6562 11782
rect 7787 11732 7788 11796
rect 7852 11732 7853 11796
rect 7787 11731 7853 11732
rect 6867 11660 6933 11661
rect 6867 11596 6868 11660
rect 6932 11596 6933 11660
rect 6867 11595 6933 11596
rect 6499 11252 6565 11253
rect 6499 11188 6500 11252
rect 6564 11188 6565 11252
rect 6499 11187 6565 11188
rect 6870 10570 6930 11595
rect 6686 10510 6930 10570
rect 6686 10437 6746 10510
rect 6683 10436 6749 10437
rect 6683 10372 6684 10436
rect 6748 10372 6749 10436
rect 6683 10371 6749 10372
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 8894 9893 8954 16627
rect 9443 15604 9509 15605
rect 9443 15540 9444 15604
rect 9508 15540 9509 15604
rect 9443 15539 9509 15540
rect 9446 13837 9506 15539
rect 9443 13836 9509 13837
rect 9443 13772 9444 13836
rect 9508 13772 9509 13836
rect 9443 13771 9509 13772
rect 9259 13564 9325 13565
rect 9259 13500 9260 13564
rect 9324 13500 9325 13564
rect 9259 13499 9325 13500
rect 9262 13378 9322 13499
rect 9259 12612 9325 12613
rect 9259 12548 9260 12612
rect 9324 12548 9325 12612
rect 9259 12547 9325 12548
rect 9262 10981 9322 12547
rect 9630 12341 9690 17222
rect 9998 16690 10058 20027
rect 9814 16630 10058 16690
rect 10277 19072 10597 20096
rect 10915 19276 10981 19277
rect 10915 19212 10916 19276
rect 10980 19212 10981 19276
rect 10915 19211 10981 19212
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10731 17780 10797 17781
rect 10731 17716 10732 17780
rect 10796 17716 10797 17780
rect 10731 17715 10797 17716
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 9814 14650 9874 16630
rect 9995 16420 10061 16421
rect 9995 16356 9996 16420
rect 10060 16356 10061 16420
rect 9995 16355 10061 16356
rect 9998 14789 10058 16355
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 9995 14788 10061 14789
rect 9995 14724 9996 14788
rect 10060 14724 10061 14788
rect 9995 14723 10061 14724
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 9814 14590 10058 14650
rect 9811 14380 9877 14381
rect 9811 14316 9812 14380
rect 9876 14316 9877 14380
rect 9811 14315 9877 14316
rect 9814 12477 9874 14315
rect 9998 13565 10058 14590
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 9995 13564 10061 13565
rect 9995 13500 9996 13564
rect 10060 13500 10061 13564
rect 9995 13499 10061 13500
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 9811 12476 9877 12477
rect 9811 12412 9812 12476
rect 9876 12412 9877 12476
rect 9811 12411 9877 12412
rect 9627 12340 9693 12341
rect 9627 12276 9628 12340
rect 9692 12276 9693 12340
rect 9627 12275 9693 12276
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 9259 10980 9325 10981
rect 9259 10916 9260 10980
rect 9324 10916 9325 10980
rect 9259 10915 9325 10916
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 8891 9892 8957 9893
rect 8891 9828 8892 9892
rect 8956 9828 8957 9892
rect 8891 9827 8957 9828
rect 6134 9485 6194 9742
rect 6131 9484 6197 9485
rect 6131 9420 6132 9484
rect 6196 9420 6197 9484
rect 6131 9419 6197 9420
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 2819 8668 2885 8669
rect 2819 8604 2820 8668
rect 2884 8604 2885 8668
rect 2819 8603 2885 8604
rect 2451 8260 2517 8261
rect 2451 8196 2452 8260
rect 2516 8196 2517 8260
rect 2451 8195 2517 8196
rect 5610 7648 5931 8672
rect 10277 9280 10597 10304
rect 10734 10301 10794 17715
rect 10918 13021 10978 19211
rect 10915 13020 10981 13021
rect 10915 12956 10916 13020
rect 10980 12956 10981 13020
rect 10915 12955 10981 12956
rect 10731 10300 10797 10301
rect 10731 10236 10732 10300
rect 10796 10236 10797 10300
rect 10731 10235 10797 10236
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 8891 8332 8892 8382
rect 8956 8332 8957 8382
rect 8891 8331 8957 8332
rect 7787 8260 7853 8261
rect 7787 8196 7788 8260
rect 7852 8196 7853 8260
rect 7787 8195 7853 8196
rect 7790 7938 7850 8195
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 3923 7308 3989 7309
rect 3923 7258 3924 7308
rect 3988 7258 3989 7308
rect 3923 6764 3989 6765
rect 3923 6700 3924 6764
rect 3988 6700 3989 6764
rect 3923 6699 3989 6700
rect 3926 5898 3986 6699
rect 5610 6560 5931 7584
rect 7790 7309 7850 7702
rect 7787 7308 7853 7309
rect 7787 7244 7788 7308
rect 7852 7244 7853 7308
rect 7787 7243 7853 7244
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 3003 5540 3069 5541
rect 3003 5476 3004 5540
rect 3068 5476 3069 5540
rect 3003 5475 3069 5476
rect 3006 2498 3066 5475
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 7603 5404 7669 5405
rect 7603 5340 7604 5404
rect 7668 5340 7669 5404
rect 7603 5339 7669 5340
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 7606 1461 7666 5339
rect 10277 4928 10597 5952
rect 11102 5405 11162 24651
rect 11283 24580 11349 24581
rect 11283 24516 11284 24580
rect 11348 24516 11349 24580
rect 11283 24515 11349 24516
rect 11099 5404 11165 5405
rect 11099 5340 11100 5404
rect 11164 5340 11165 5404
rect 11099 5339 11165 5340
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 11286 3093 11346 24515
rect 12571 24172 12637 24173
rect 12571 24108 12572 24172
rect 12636 24108 12637 24172
rect 12571 24107 12637 24108
rect 12019 24036 12085 24037
rect 12019 23972 12020 24036
rect 12084 23972 12085 24036
rect 12019 23971 12085 23972
rect 12022 23578 12082 23971
rect 11467 23356 11533 23357
rect 11467 23292 11468 23356
rect 11532 23292 11533 23356
rect 11467 23291 11533 23292
rect 11470 5949 11530 23291
rect 12022 22133 12082 23342
rect 12019 22132 12085 22133
rect 12019 22068 12020 22132
rect 12084 22068 12085 22132
rect 12019 22067 12085 22068
rect 12574 21997 12634 24107
rect 14944 23968 15264 24992
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 15883 24852 15949 24853
rect 15883 24788 15884 24852
rect 15948 24788 15949 24852
rect 15883 24787 15949 24788
rect 15515 24036 15581 24037
rect 15515 23972 15516 24036
rect 15580 23972 15581 24036
rect 15515 23971 15581 23972
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14779 23900 14845 23901
rect 14779 23836 14780 23900
rect 14844 23836 14845 23900
rect 14779 23835 14845 23836
rect 13859 23628 13925 23629
rect 13859 23564 13860 23628
rect 13924 23564 13925 23628
rect 13859 23563 13925 23564
rect 13675 22268 13741 22269
rect 13675 22204 13676 22268
rect 13740 22204 13741 22268
rect 13675 22203 13741 22204
rect 12571 21996 12637 21997
rect 12571 21932 12572 21996
rect 12636 21932 12637 21996
rect 12571 21931 12637 21932
rect 13307 21860 13373 21861
rect 13307 21796 13308 21860
rect 13372 21796 13373 21860
rect 13307 21795 13373 21796
rect 13310 21538 13370 21795
rect 12203 20772 12269 20773
rect 12203 20708 12204 20772
rect 12268 20708 12269 20772
rect 12203 20707 12269 20708
rect 11835 19140 11901 19141
rect 11835 19076 11836 19140
rect 11900 19076 11901 19140
rect 11835 19075 11901 19076
rect 11651 18596 11717 18597
rect 11651 18532 11652 18596
rect 11716 18532 11717 18596
rect 11651 18531 11717 18532
rect 11654 14109 11714 18531
rect 11651 14108 11717 14109
rect 11651 14044 11652 14108
rect 11716 14044 11717 14108
rect 11651 14043 11717 14044
rect 11838 7581 11898 19075
rect 11835 7580 11901 7581
rect 11835 7516 11836 7580
rect 11900 7516 11901 7580
rect 11835 7515 11901 7516
rect 11835 6900 11901 6901
rect 11835 6836 11836 6900
rect 11900 6836 11901 6900
rect 11835 6835 11901 6836
rect 11838 5949 11898 6835
rect 11467 5948 11533 5949
rect 11467 5884 11468 5948
rect 11532 5884 11533 5948
rect 11467 5883 11533 5884
rect 11835 5948 11901 5949
rect 11835 5884 11836 5948
rect 11900 5884 11901 5948
rect 11835 5883 11901 5884
rect 11467 5540 11533 5541
rect 11467 5476 11468 5540
rect 11532 5476 11533 5540
rect 11467 5475 11533 5476
rect 11470 4453 11530 5475
rect 11467 4452 11533 4453
rect 11467 4388 11468 4452
rect 11532 4388 11533 4452
rect 11467 4387 11533 4388
rect 12206 3773 12266 20707
rect 12939 19140 13005 19141
rect 12939 19076 12940 19140
rect 13004 19076 13005 19140
rect 12939 19075 13005 19076
rect 12755 16284 12821 16285
rect 12755 16220 12756 16284
rect 12820 16220 12821 16284
rect 12755 16219 12821 16220
rect 12571 13156 12637 13157
rect 12571 13092 12572 13156
rect 12636 13092 12637 13156
rect 12571 13091 12637 13092
rect 12574 10709 12634 13091
rect 12758 12613 12818 16219
rect 12942 15605 13002 19075
rect 13123 17916 13189 17917
rect 13123 17852 13124 17916
rect 13188 17852 13189 17916
rect 13123 17851 13189 17852
rect 12939 15604 13005 15605
rect 12939 15540 12940 15604
rect 13004 15540 13005 15604
rect 12939 15539 13005 15540
rect 12755 12612 12821 12613
rect 12755 12548 12756 12612
rect 12820 12548 12821 12612
rect 12755 12547 12821 12548
rect 13126 11797 13186 17851
rect 13310 13021 13370 21302
rect 13678 17373 13738 22203
rect 13675 17372 13741 17373
rect 13675 17308 13676 17372
rect 13740 17308 13741 17372
rect 13675 17307 13741 17308
rect 13491 16692 13557 16693
rect 13491 16628 13492 16692
rect 13556 16628 13557 16692
rect 13491 16627 13557 16628
rect 13307 13020 13373 13021
rect 13307 12956 13308 13020
rect 13372 12956 13373 13020
rect 13307 12955 13373 12956
rect 13494 12698 13554 16627
rect 13494 12205 13554 12462
rect 13491 12204 13557 12205
rect 13491 12140 13492 12204
rect 13556 12140 13557 12204
rect 13491 12139 13557 12140
rect 13123 11796 13189 11797
rect 13123 11732 13124 11796
rect 13188 11732 13189 11796
rect 13123 11731 13189 11732
rect 13494 11389 13554 11782
rect 13491 11388 13557 11389
rect 13491 11324 13492 11388
rect 13556 11324 13557 11388
rect 13491 11323 13557 11324
rect 12571 10708 12637 10709
rect 12571 10644 12572 10708
rect 12636 10644 12637 10708
rect 13491 10708 13557 10709
rect 13491 10658 13492 10708
rect 13556 10658 13557 10708
rect 12571 10643 12637 10644
rect 13862 4045 13922 23563
rect 14782 22269 14842 23835
rect 14944 22880 15264 23904
rect 15331 23492 15397 23493
rect 15331 23428 15332 23492
rect 15396 23428 15397 23492
rect 15331 23427 15397 23428
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14779 22268 14845 22269
rect 14779 22204 14780 22268
rect 14844 22204 14845 22268
rect 14779 22203 14845 22204
rect 14782 16285 14842 22203
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14779 16284 14845 16285
rect 14779 16220 14780 16284
rect 14844 16220 14845 16284
rect 14779 16219 14845 16220
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14595 15060 14661 15061
rect 14595 14996 14596 15060
rect 14660 14996 14661 15060
rect 14595 14995 14661 14996
rect 14227 14788 14293 14789
rect 14227 14738 14228 14788
rect 14292 14738 14293 14788
rect 14411 14380 14477 14381
rect 14411 14316 14412 14380
rect 14476 14316 14477 14380
rect 14411 14315 14477 14316
rect 14414 8805 14474 14315
rect 14598 13429 14658 14995
rect 14779 14788 14845 14789
rect 14779 14724 14780 14788
rect 14844 14724 14845 14788
rect 14779 14723 14845 14724
rect 14595 13428 14661 13429
rect 14595 13364 14596 13428
rect 14660 13364 14661 13428
rect 14595 13363 14661 13364
rect 14782 9893 14842 14723
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 15334 12613 15394 23427
rect 15331 12612 15397 12613
rect 15331 12548 15332 12612
rect 15396 12548 15397 12612
rect 15331 12547 15397 12548
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14779 9892 14845 9893
rect 14779 9828 14780 9892
rect 14844 9828 14845 9892
rect 14779 9827 14845 9828
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14779 9484 14845 9485
rect 14779 9420 14780 9484
rect 14844 9420 14845 9484
rect 14779 9419 14845 9420
rect 14411 8804 14477 8805
rect 14411 8740 14412 8804
rect 14476 8740 14477 8804
rect 14411 8739 14477 8740
rect 13859 4044 13925 4045
rect 13859 3980 13860 4044
rect 13924 3980 13925 4044
rect 13859 3979 13925 3980
rect 14414 3909 14474 8739
rect 14595 8396 14661 8397
rect 14595 8332 14596 8396
rect 14660 8394 14661 8396
rect 14782 8394 14842 9419
rect 14660 8334 14842 8394
rect 14660 8332 14661 8334
rect 14595 8331 14661 8332
rect 14782 7989 14842 8334
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14779 7988 14845 7989
rect 14779 7924 14780 7988
rect 14844 7924 14845 7988
rect 14779 7923 14845 7924
rect 14782 6085 14842 7923
rect 14944 7648 15264 8672
rect 15518 8125 15578 23971
rect 15886 12749 15946 24787
rect 19610 24512 19930 25536
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 20483 24580 20549 24581
rect 20483 24516 20484 24580
rect 20548 24516 20549 24580
rect 20483 24515 20549 24516
rect 21955 24580 22021 24581
rect 21955 24516 21956 24580
rect 22020 24516 22021 24580
rect 21955 24515 22021 24516
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 16803 23764 16869 23765
rect 16803 23700 16804 23764
rect 16868 23700 16869 23764
rect 16803 23699 16869 23700
rect 16251 23628 16317 23629
rect 16251 23564 16252 23628
rect 16316 23564 16317 23628
rect 16251 23563 16317 23564
rect 16254 20858 16314 23563
rect 16438 18869 16498 19262
rect 16435 18868 16501 18869
rect 16435 18804 16436 18868
rect 16500 18804 16501 18868
rect 16435 18803 16501 18804
rect 16619 16964 16685 16965
rect 16619 16900 16620 16964
rect 16684 16900 16685 16964
rect 16619 16899 16685 16900
rect 15883 12748 15949 12749
rect 15883 12684 15884 12748
rect 15948 12684 15949 12748
rect 15883 12683 15949 12684
rect 15883 12612 15949 12613
rect 15883 12548 15884 12612
rect 15948 12548 15949 12612
rect 15883 12547 15949 12548
rect 15699 8940 15765 8941
rect 15699 8876 15700 8940
rect 15764 8876 15765 8940
rect 15699 8875 15765 8876
rect 15515 8124 15581 8125
rect 15515 8060 15516 8124
rect 15580 8060 15581 8124
rect 15515 8059 15581 8060
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14779 6084 14845 6085
rect 14779 6020 14780 6084
rect 14844 6020 14845 6084
rect 14779 6019 14845 6020
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 15702 5269 15762 8875
rect 15699 5268 15765 5269
rect 15699 5204 15700 5268
rect 15764 5204 15765 5268
rect 15699 5203 15765 5204
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 13675 3908 13741 3909
rect 13675 3844 13676 3908
rect 13740 3844 13741 3908
rect 13675 3843 13741 3844
rect 14411 3908 14477 3909
rect 14411 3844 14412 3908
rect 14476 3844 14477 3908
rect 14411 3843 14477 3844
rect 12203 3772 12269 3773
rect 12203 3708 12204 3772
rect 12268 3708 12269 3772
rect 12203 3707 12269 3708
rect 13678 3178 13738 3843
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 11283 3092 11349 3093
rect 11283 3028 11284 3092
rect 11348 3028 11349 3092
rect 11283 3027 11349 3028
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 7603 1460 7669 1461
rect 7603 1396 7604 1460
rect 7668 1396 7669 1460
rect 7603 1395 7669 1396
rect 15886 1053 15946 12547
rect 16435 12476 16501 12477
rect 16435 12412 16436 12476
rect 16500 12412 16501 12476
rect 16435 12411 16501 12412
rect 16438 10981 16498 12411
rect 16435 10980 16501 10981
rect 16435 10916 16436 10980
rect 16500 10916 16501 10980
rect 16435 10915 16501 10916
rect 16622 9621 16682 16899
rect 16619 9620 16685 9621
rect 16619 9556 16620 9620
rect 16684 9556 16685 9620
rect 16619 9555 16685 9556
rect 16254 5541 16314 7022
rect 16251 5540 16317 5541
rect 16251 5476 16252 5540
rect 16316 5476 16317 5540
rect 16251 5475 16317 5476
rect 16806 3773 16866 23699
rect 19610 23424 19930 24448
rect 20115 23492 20181 23493
rect 20115 23428 20116 23492
rect 20180 23428 20181 23492
rect 20115 23427 20181 23428
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19195 22676 19261 22677
rect 19195 22612 19196 22676
rect 19260 22612 19261 22676
rect 19195 22611 19261 22612
rect 19198 21997 19258 22611
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19195 21996 19261 21997
rect 19195 21932 19196 21996
rect 19260 21932 19261 21996
rect 19195 21931 19261 21932
rect 19379 21452 19445 21453
rect 19379 21388 19380 21452
rect 19444 21388 19445 21452
rect 19379 21387 19445 21388
rect 17171 21180 17237 21181
rect 17171 21116 17172 21180
rect 17236 21116 17237 21180
rect 17171 21115 17237 21116
rect 16987 8804 17053 8805
rect 16987 8740 16988 8804
rect 17052 8740 17053 8804
rect 16987 8739 17053 8740
rect 16990 4861 17050 8739
rect 16987 4860 17053 4861
rect 16987 4796 16988 4860
rect 17052 4796 17053 4860
rect 16987 4795 17053 4796
rect 16803 3772 16869 3773
rect 16803 3708 16804 3772
rect 16868 3708 16869 3772
rect 16803 3707 16869 3708
rect 16619 2548 16685 2549
rect 16619 2484 16620 2548
rect 16684 2484 16685 2548
rect 17174 2498 17234 21115
rect 18278 19549 18338 19942
rect 18275 19548 18341 19549
rect 18275 19484 18276 19548
rect 18340 19484 18341 19548
rect 18275 19483 18341 19484
rect 19382 14738 19442 21387
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 17355 13836 17421 13837
rect 17355 13772 17356 13836
rect 17420 13772 17421 13836
rect 17355 13771 17421 13772
rect 17358 5269 17418 13771
rect 17726 8618 17786 11782
rect 19382 6901 19442 14502
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19379 6900 19445 6901
rect 19379 6836 19380 6900
rect 19444 6836 19445 6900
rect 19379 6835 19445 6836
rect 19610 6016 19930 7040
rect 20118 6493 20178 23427
rect 20486 21861 20546 24515
rect 20483 21860 20549 21861
rect 20483 21796 20484 21860
rect 20548 21796 20549 21860
rect 20483 21795 20549 21796
rect 20486 17917 20546 21795
rect 20851 18188 20917 18189
rect 20851 18124 20852 18188
rect 20916 18124 20917 18188
rect 20851 18123 20917 18124
rect 20854 18050 20914 18123
rect 20854 17990 21098 18050
rect 20483 17916 20549 17917
rect 20483 17852 20484 17916
rect 20548 17852 20549 17916
rect 20483 17851 20549 17852
rect 20667 17780 20733 17781
rect 20667 17716 20668 17780
rect 20732 17716 20733 17780
rect 20667 17715 20733 17716
rect 20670 16013 20730 17715
rect 20667 16012 20733 16013
rect 20667 15948 20668 16012
rect 20732 15948 20733 16012
rect 20667 15947 20733 15948
rect 21038 13565 21098 17990
rect 21035 13564 21101 13565
rect 21035 13500 21036 13564
rect 21100 13500 21101 13564
rect 21035 13499 21101 13500
rect 20667 13092 20668 13142
rect 20732 13092 20733 13142
rect 20667 13091 20733 13092
rect 20299 12884 20365 12885
rect 20299 12820 20300 12884
rect 20364 12820 20365 12884
rect 20299 12819 20365 12820
rect 20302 9349 20362 12819
rect 21035 12412 21036 12462
rect 21100 12412 21101 12462
rect 21035 12411 21101 12412
rect 21958 12018 22018 24515
rect 23795 24172 23861 24173
rect 23795 24108 23796 24172
rect 23860 24108 23861 24172
rect 23795 24107 23861 24108
rect 23427 23084 23493 23085
rect 23427 23020 23428 23084
rect 23492 23020 23493 23084
rect 23427 23019 23493 23020
rect 23059 22812 23125 22813
rect 23059 22748 23060 22812
rect 23124 22748 23125 22812
rect 23059 22747 23125 22748
rect 22507 17916 22573 17917
rect 22507 17852 22508 17916
rect 22572 17852 22573 17916
rect 22507 17851 22573 17852
rect 22510 10981 22570 17851
rect 22507 10980 22573 10981
rect 22507 10916 22508 10980
rect 22572 10916 22573 10980
rect 22507 10915 22573 10916
rect 22694 10301 22754 20622
rect 22875 18732 22941 18733
rect 22875 18668 22876 18732
rect 22940 18668 22941 18732
rect 22875 18667 22941 18668
rect 22691 10300 22757 10301
rect 22691 10236 22692 10300
rect 22756 10236 22757 10300
rect 22691 10235 22757 10236
rect 22878 9893 22938 18667
rect 22875 9892 22941 9893
rect 22875 9828 22876 9892
rect 22940 9828 22941 9892
rect 22875 9827 22941 9828
rect 20299 9348 20365 9349
rect 20299 9284 20300 9348
rect 20364 9284 20365 9348
rect 20299 9283 20365 9284
rect 22878 7170 22938 9827
rect 23062 9485 23122 22747
rect 23243 17372 23309 17373
rect 23243 17308 23244 17372
rect 23308 17308 23309 17372
rect 23243 17307 23309 17308
rect 23246 15741 23306 17307
rect 23430 17237 23490 23019
rect 23611 22948 23677 22949
rect 23611 22884 23612 22948
rect 23676 22884 23677 22948
rect 23611 22883 23677 22884
rect 23427 17236 23493 17237
rect 23427 17172 23428 17236
rect 23492 17172 23493 17236
rect 23427 17171 23493 17172
rect 23243 15740 23309 15741
rect 23243 15676 23244 15740
rect 23308 15676 23309 15740
rect 23243 15675 23309 15676
rect 23427 15740 23493 15741
rect 23427 15676 23428 15740
rect 23492 15676 23493 15740
rect 23427 15675 23493 15676
rect 23430 9757 23490 15675
rect 23614 14650 23674 22883
rect 23798 15741 23858 24107
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24715 23628 24781 23629
rect 24715 23564 24716 23628
rect 24780 23564 24781 23628
rect 24715 23563 24781 23564
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 23979 18868 24045 18869
rect 23979 18804 23980 18868
rect 24044 18804 24045 18868
rect 23979 18803 24045 18804
rect 23982 15877 24042 18803
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 23979 15876 24045 15877
rect 23979 15812 23980 15876
rect 24044 15812 24045 15876
rect 23979 15811 24045 15812
rect 23795 15740 23861 15741
rect 23795 15676 23796 15740
rect 23860 15676 23861 15740
rect 23795 15675 23861 15676
rect 23979 15468 24045 15469
rect 23979 15418 23980 15468
rect 24044 15418 24045 15468
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 23979 14924 24045 14925
rect 23979 14860 23980 14924
rect 24044 14860 24045 14924
rect 23979 14859 24045 14860
rect 23614 14590 23858 14650
rect 23611 11116 23677 11117
rect 23611 11052 23612 11116
rect 23676 11052 23677 11116
rect 23611 11051 23677 11052
rect 23427 9756 23493 9757
rect 23427 9692 23428 9756
rect 23492 9692 23493 9756
rect 23427 9691 23493 9692
rect 23059 9484 23125 9485
rect 23059 9420 23060 9484
rect 23124 9420 23125 9484
rect 23059 9419 23125 9420
rect 23614 7258 23674 11051
rect 23798 7581 23858 14590
rect 23982 8669 24042 14859
rect 24277 14176 24597 15200
rect 24718 14925 24778 23563
rect 24899 23492 24965 23493
rect 24899 23428 24900 23492
rect 24964 23428 24965 23492
rect 24899 23427 24965 23428
rect 24902 19685 24962 23427
rect 24899 19684 24965 19685
rect 24899 19620 24900 19684
rect 24964 19620 24965 19684
rect 24899 19619 24965 19620
rect 25083 19548 25149 19549
rect 25083 19498 25084 19548
rect 25148 19498 25149 19548
rect 24899 16284 24965 16285
rect 24899 16220 24900 16284
rect 24964 16220 24965 16284
rect 24899 16219 24965 16220
rect 24715 14924 24781 14925
rect 24715 14860 24716 14924
rect 24780 14860 24781 14924
rect 24715 14859 24781 14860
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24715 13564 24781 13565
rect 24715 13500 24716 13564
rect 24780 13500 24781 13564
rect 24715 13499 24781 13500
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24718 11525 24778 13499
rect 24902 12069 24962 16219
rect 24899 12068 24965 12069
rect 24899 12004 24900 12068
rect 24964 12004 24965 12068
rect 24899 12003 24965 12004
rect 25819 11732 25820 11782
rect 25884 11732 25885 11782
rect 25819 11731 25885 11732
rect 24715 11524 24781 11525
rect 24715 11460 24716 11524
rect 24780 11460 24781 11524
rect 24715 11459 24781 11460
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24899 10844 24965 10845
rect 24899 10780 24900 10844
rect 24964 10780 24965 10844
rect 24899 10779 24965 10780
rect 24902 10658 24962 10779
rect 24715 10300 24781 10301
rect 24715 10236 24716 10300
rect 24780 10236 24781 10300
rect 24715 10235 24781 10236
rect 24899 10300 24965 10301
rect 24899 10236 24900 10300
rect 24964 10236 24965 10300
rect 24899 10235 24965 10236
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 23979 8668 24045 8669
rect 23979 8604 23980 8668
rect 24044 8604 24045 8668
rect 23979 8603 24045 8604
rect 23979 8396 24045 8397
rect 23979 8332 23980 8396
rect 24044 8332 24045 8396
rect 23979 8331 24045 8332
rect 23795 7580 23861 7581
rect 23795 7516 23796 7580
rect 23860 7516 23861 7580
rect 23795 7515 23861 7516
rect 22878 7110 23122 7170
rect 20299 6900 20365 6901
rect 20299 6836 20300 6900
rect 20364 6836 20365 6900
rect 20299 6835 20365 6836
rect 20115 6492 20181 6493
rect 20115 6428 20116 6492
rect 20180 6428 20181 6492
rect 20115 6427 20181 6428
rect 20302 6085 20362 6835
rect 20299 6084 20365 6085
rect 20299 6020 20300 6084
rect 20364 6020 20365 6084
rect 20299 6019 20365 6020
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19195 5948 19261 5949
rect 19195 5898 19196 5948
rect 19260 5898 19261 5948
rect 17539 5676 17605 5677
rect 17539 5612 17540 5676
rect 17604 5612 17605 5676
rect 17539 5611 17605 5612
rect 17355 5268 17421 5269
rect 17355 5204 17356 5268
rect 17420 5204 17421 5268
rect 17355 5203 17421 5204
rect 17542 4538 17602 5611
rect 19610 4928 19930 5952
rect 21771 5268 21837 5269
rect 21771 5204 21772 5268
rect 21836 5204 21837 5268
rect 21771 5203 21837 5204
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 21774 2957 21834 5203
rect 22694 4589 22754 4982
rect 22691 4588 22757 4589
rect 22691 4524 22692 4588
rect 22756 4524 22757 4588
rect 22691 4523 22757 4524
rect 23062 4045 23122 7110
rect 23795 6492 23861 6493
rect 23795 6428 23796 6492
rect 23860 6428 23861 6492
rect 23795 6427 23861 6428
rect 23059 4044 23125 4045
rect 23059 3980 23060 4044
rect 23124 3980 23125 4044
rect 23059 3979 23125 3980
rect 21771 2956 21837 2957
rect 21771 2892 21772 2956
rect 21836 2892 21837 2956
rect 23798 3093 23858 6427
rect 23982 3909 24042 8331
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 23979 3908 24045 3909
rect 23979 3844 23980 3908
rect 24044 3844 24045 3908
rect 23979 3843 24045 3844
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 23795 3092 23861 3093
rect 23795 3028 23796 3092
rect 23860 3028 23861 3092
rect 23795 3027 23861 3028
rect 21771 2891 21837 2892
rect 23427 2892 23428 2942
rect 23492 2892 23493 2942
rect 23427 2891 23493 2892
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 16619 2483 16685 2484
rect 16622 1597 16682 2483
rect 19610 2128 19930 2688
rect 24277 2208 24597 3232
rect 24718 2685 24778 10235
rect 24902 9757 24962 10235
rect 24899 9756 24965 9757
rect 24899 9692 24900 9756
rect 24964 9692 24965 9756
rect 24899 9691 24965 9692
rect 24899 5812 24965 5813
rect 24899 5748 24900 5812
rect 24964 5748 24965 5812
rect 24899 5747 24965 5748
rect 24715 2684 24781 2685
rect 24715 2620 24716 2684
rect 24780 2620 24781 2684
rect 24715 2619 24781 2620
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
rect 24715 1732 24781 1733
rect 24715 1668 24716 1732
rect 24780 1730 24781 1732
rect 24902 1730 24962 5747
rect 24780 1670 24962 1730
rect 24780 1668 24781 1670
rect 24715 1667 24781 1668
rect 16619 1596 16685 1597
rect 16619 1532 16620 1596
rect 16684 1532 16685 1596
rect 16619 1531 16685 1532
rect 15883 1052 15949 1053
rect 15883 988 15884 1052
rect 15948 988 15949 1052
rect 15883 987 15949 988
<< via4 >>
rect 3286 13142 3522 13378
rect 9542 19942 9778 20178
rect 7334 15862 7570 16098
rect 6782 13822 7018 14058
rect 6414 11782 6650 12018
rect 9542 17222 9778 17458
rect 6046 9742 6282 9978
rect 9174 13142 9410 13378
rect 8806 8396 9042 8618
rect 8806 8382 8892 8396
rect 8892 8382 8956 8396
rect 8956 8382 9042 8396
rect 7702 7702 7938 7938
rect 3838 7244 3924 7258
rect 3924 7244 3988 7258
rect 3988 7244 4074 7258
rect 3838 7022 4074 7244
rect 5310 6492 5546 6578
rect 5310 6428 5396 6492
rect 5396 6428 5460 6492
rect 5460 6428 5546 6492
rect 5310 6342 5546 6428
rect 3838 5662 4074 5898
rect 4574 4452 4810 4538
rect 4574 4388 4660 4452
rect 4660 4388 4724 4452
rect 4724 4388 4810 4452
rect 4574 4302 4810 4388
rect 2918 2262 3154 2498
rect 9358 5132 9594 5218
rect 9358 5068 9444 5132
rect 9444 5068 9508 5132
rect 9508 5068 9594 5132
rect 9358 4982 9594 5068
rect 11934 23342 12170 23578
rect 13222 21302 13458 21538
rect 13406 12462 13642 12698
rect 13406 11782 13642 12018
rect 13406 10644 13492 10658
rect 13492 10644 13556 10658
rect 13556 10644 13642 10658
rect 13406 10422 13642 10644
rect 13222 7172 13458 7258
rect 13222 7108 13308 7172
rect 13308 7108 13372 7172
rect 13372 7108 13458 7172
rect 13222 7022 13458 7108
rect 14142 14724 14228 14738
rect 14228 14724 14292 14738
rect 14292 14724 14378 14738
rect 14142 14502 14378 14724
rect 16166 20622 16402 20858
rect 16350 19262 16586 19498
rect 16166 15332 16402 15418
rect 16166 15268 16252 15332
rect 16252 15268 16316 15332
rect 16316 15268 16402 15332
rect 16166 15182 16402 15268
rect 13590 2942 13826 3178
rect 16166 9892 16402 9978
rect 16166 9828 16252 9892
rect 16252 9828 16316 9892
rect 16316 9828 16402 9892
rect 16166 9742 16402 9828
rect 16166 7022 16402 7258
rect 19294 23492 19530 23578
rect 19294 23428 19380 23492
rect 19380 23428 19444 23492
rect 19444 23428 19530 23492
rect 19294 23342 19530 23428
rect 18190 19942 18426 20178
rect 17822 16012 18058 16098
rect 17822 15948 17908 16012
rect 17908 15948 17972 16012
rect 17972 15948 18058 16012
rect 17822 15862 18058 15948
rect 19294 14502 19530 14738
rect 17638 11782 17874 12018
rect 17638 8382 17874 8618
rect 17638 6492 17874 6578
rect 17638 6428 17724 6492
rect 17724 6428 17788 6492
rect 17788 6428 17874 6492
rect 17638 6342 17874 6428
rect 20766 21452 21002 21538
rect 20766 21388 20852 21452
rect 20852 21388 20916 21452
rect 20916 21388 21002 21452
rect 20766 21302 21002 21388
rect 20582 13972 20818 14058
rect 20582 13908 20668 13972
rect 20668 13908 20732 13972
rect 20732 13908 20818 13972
rect 20582 13822 20818 13908
rect 20582 13156 20818 13378
rect 20582 13142 20668 13156
rect 20668 13142 20732 13156
rect 20732 13142 20818 13156
rect 20950 12476 21186 12698
rect 20950 12462 21036 12476
rect 21036 12462 21100 12476
rect 21100 12462 21186 12476
rect 22606 20622 22842 20858
rect 21870 11782 22106 12018
rect 23894 15404 23980 15418
rect 23980 15404 24044 15418
rect 24044 15404 24130 15418
rect 23894 15182 24130 15404
rect 23158 7852 23394 7938
rect 23158 7788 23244 7852
rect 23244 7788 23308 7852
rect 23308 7788 23394 7852
rect 23158 7702 23394 7788
rect 24998 19484 25084 19498
rect 25084 19484 25148 19498
rect 25148 19484 25234 19498
rect 24998 19262 25234 19484
rect 24998 17372 25234 17458
rect 24998 17308 25084 17372
rect 25084 17308 25148 17372
rect 25148 17308 25234 17372
rect 24998 17222 25234 17308
rect 25734 11796 25970 12018
rect 25734 11782 25820 11796
rect 25820 11782 25884 11796
rect 25884 11782 25970 11796
rect 24814 10422 25050 10658
rect 19110 5884 19196 5898
rect 19196 5884 19260 5898
rect 19260 5884 19346 5898
rect 19110 5662 19346 5884
rect 17454 4302 17690 4538
rect 22606 4982 22842 5218
rect 23526 7022 23762 7258
rect 23342 2956 23578 3178
rect 23342 2942 23428 2956
rect 23428 2942 23492 2956
rect 23492 2942 23578 2956
rect 17086 2262 17322 2498
<< metal5 >>
rect 11892 23578 19572 23620
rect 11892 23342 11934 23578
rect 12170 23342 19294 23578
rect 19530 23342 19572 23578
rect 11892 23300 19572 23342
rect 13180 21538 21044 21580
rect 13180 21302 13222 21538
rect 13458 21302 20766 21538
rect 21002 21302 21044 21538
rect 13180 21260 21044 21302
rect 16124 20858 22884 20900
rect 16124 20622 16166 20858
rect 16402 20622 22606 20858
rect 22842 20622 22884 20858
rect 16124 20580 22884 20622
rect 9500 20178 18468 20220
rect 9500 19942 9542 20178
rect 9778 19942 18190 20178
rect 18426 19942 18468 20178
rect 9500 19900 18468 19942
rect 16308 19498 25276 19540
rect 16308 19262 16350 19498
rect 16586 19262 24998 19498
rect 25234 19262 25276 19498
rect 16308 19220 25276 19262
rect 9500 17458 25276 17500
rect 9500 17222 9542 17458
rect 9778 17222 24998 17458
rect 25234 17222 25276 17458
rect 9500 17180 25276 17222
rect 7292 16098 18100 16140
rect 7292 15862 7334 16098
rect 7570 15862 17822 16098
rect 18058 15862 18100 16098
rect 7292 15820 18100 15862
rect 16124 15418 24172 15460
rect 16124 15182 16166 15418
rect 16402 15182 23894 15418
rect 24130 15182 24172 15418
rect 16124 15140 24172 15182
rect 14100 14738 19572 14780
rect 14100 14502 14142 14738
rect 14378 14502 19294 14738
rect 19530 14502 19572 14738
rect 14100 14460 19572 14502
rect 6740 14058 20860 14100
rect 6740 13822 6782 14058
rect 7018 13822 20582 14058
rect 20818 13822 20860 14058
rect 6740 13780 20860 13822
rect 3244 13378 20860 13420
rect 3244 13142 3286 13378
rect 3522 13142 9174 13378
rect 9410 13142 20582 13378
rect 20818 13142 20860 13378
rect 3244 13100 20860 13142
rect 13364 12698 21228 12740
rect 13364 12462 13406 12698
rect 13642 12462 20950 12698
rect 21186 12462 21228 12698
rect 13364 12420 21228 12462
rect 6372 12018 13684 12060
rect 6372 11782 6414 12018
rect 6650 11782 13406 12018
rect 13642 11782 13684 12018
rect 6372 11740 13684 11782
rect 17596 12018 26012 12060
rect 17596 11782 17638 12018
rect 17874 11782 21870 12018
rect 22106 11782 25734 12018
rect 25970 11782 26012 12018
rect 17596 11740 26012 11782
rect 13364 10658 25092 10700
rect 13364 10422 13406 10658
rect 13642 10422 24814 10658
rect 25050 10422 25092 10658
rect 13364 10380 25092 10422
rect 6004 9978 16444 10020
rect 6004 9742 6046 9978
rect 6282 9742 16166 9978
rect 16402 9742 16444 9978
rect 6004 9700 16444 9742
rect 8764 8618 17916 8660
rect 8764 8382 8806 8618
rect 9042 8382 17638 8618
rect 17874 8382 17916 8618
rect 8764 8340 17916 8382
rect 7660 7938 23436 7980
rect 7660 7702 7702 7938
rect 7938 7702 23158 7938
rect 23394 7702 23436 7938
rect 7660 7660 23436 7702
rect 3796 7258 13500 7300
rect 3796 7022 3838 7258
rect 4074 7022 13222 7258
rect 13458 7022 13500 7258
rect 3796 6980 13500 7022
rect 16124 7258 23804 7300
rect 16124 7022 16166 7258
rect 16402 7022 23526 7258
rect 23762 7022 23804 7258
rect 16124 6980 23804 7022
rect 5268 6578 17916 6620
rect 5268 6342 5310 6578
rect 5546 6342 17638 6578
rect 17874 6342 17916 6578
rect 5268 6300 17916 6342
rect 3796 5898 19388 5940
rect 3796 5662 3838 5898
rect 4074 5662 19110 5898
rect 19346 5662 19388 5898
rect 3796 5620 19388 5662
rect 9316 5218 22884 5260
rect 9316 4982 9358 5218
rect 9594 4982 22606 5218
rect 22842 4982 22884 5218
rect 9316 4940 22884 4982
rect 4532 4538 17732 4580
rect 4532 4302 4574 4538
rect 4810 4302 17454 4538
rect 17690 4302 17732 4538
rect 4532 4260 17732 4302
rect 13548 3178 23620 3220
rect 13548 2942 13590 3178
rect 13826 2942 23342 3178
rect 23578 2942 23620 3178
rect 13548 2900 23620 2942
rect 2876 2498 17364 2540
rect 2876 2262 2918 2498
rect 3154 2262 17086 2498
rect 17322 2262 17364 2498
rect 2876 2220 17364 2262
use sky130_fd_sc_hd__fill_2  FILLER_0_7 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1748 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_6__A1 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_4__A1
timestamp 1604681595
transform 1 0 1564 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_4_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_16
timestamp 1604681595
transform 1 0 2576 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_12
timestamp 1604681595
transform 1 0 2208 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11
timestamp 1604681595
transform 1 0 2116 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_6__A0
timestamp 1604681595
transform 1 0 2760 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_4__A0
timestamp 1604681595
transform 1 0 2392 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_20 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2944 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_24 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3312 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23
timestamp 1604681595
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3404 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1604681595
transform 1 0 3588 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_40
timestamp 1604681595
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_36
timestamp 1604681595
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4324 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1604681595
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_53
timestamp 1604681595
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58
timestamp 1604681595
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1604681595
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_4__S
timestamp 1604681595
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_62
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 7176 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 7176 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_5__A1
timestamp 1604681595
transform 1 0 6992 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_89
timestamp 1604681595
transform 1 0 9292 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_85
timestamp 1604681595
transform 1 0 8924 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89
timestamp 1604681595
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1604681595
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 9476 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_5__A0
timestamp 1604681595
transform 1 0 9108 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 9660 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 10028 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_1_112
timestamp 1604681595
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_116
timestamp 1604681595
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1604681595
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1604681595
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_125
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12880 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_1_142
timestamp 1604681595
transform 1 0 14168 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_148
timestamp 1604681595
transform 1 0 14720 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1604681595
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1604681595
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 14904 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_165
timestamp 1604681595
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 15088 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_1_175
timestamp 1604681595
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_171
timestamp 1604681595
transform 1 0 16836 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1604681595
transform 1 0 16652 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1604681595
transform 1 0 16836 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 17020 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _115_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 17020 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_177
timestamp 1604681595
transform 1 0 17388 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_179
timestamp 1604681595
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_182
timestamp 1604681595
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_197
timestamp 1604681595
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_193
timestamp 1604681595
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_196
timestamp 1604681595
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_200
timestamp 1604681595
transform 1 0 19504 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1604681595
transform 1 0 19780 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19596 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1604681595
transform 1 0 19964 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 20608 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1604681595
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_213
timestamp 1604681595
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_210
timestamp 1604681595
transform 1 0 20424 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 20976 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_214
timestamp 1604681595
transform 1 0 20792 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_4_
timestamp 1604681595
transform 1 0 21160 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_227
timestamp 1604681595
transform 1 0 21988 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_227
timestamp 1604681595
transform 1 0 21988 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 22172 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_238
timestamp 1604681595
transform 1 0 23000 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_234
timestamp 1604681595
transform 1 0 22632 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_231
timestamp 1604681595
transform 1 0 22356 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_235
timestamp 1604681595
transform 1 0 22724 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_231
timestamp 1604681595
transform 1 0 22356 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 22540 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 22816 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 22448 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1604681595
transform 1 0 22816 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_244
timestamp 1604681595
transform 1 0 23552 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_240
timestamp 1604681595
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1604681595
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_254
timestamp 1604681595
transform 1 0 24472 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 24656 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_258
timestamp 1604681595
transform 1 0 24840 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_262
timestamp 1604681595
transform 1 0 25208 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_258
timestamp 1604681595
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 25024 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 25208 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_268
timestamp 1604681595
transform 1 0 25760 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_269
timestamp 1604681595
transform 1 0 25852 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 25392 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _031_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 25576 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 26036 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 26312 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 26404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_273
timestamp 1604681595
transform 1 0 26220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_272
timestamp 1604681595
transform 1 0 26128 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_276
timestamp 1604681595
transform 1 0 26496 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1604681595
transform 1 0 2944 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_6_
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_7__A0
timestamp 1604681595
transform 1 0 2392 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_7__S
timestamp 1604681595
transform 1 0 2760 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_12
timestamp 1604681595
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_16
timestamp 1604681595
transform 1 0 2576 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_6__S
timestamp 1604681595
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_23
timestamp 1604681595
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 6532 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 5980 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 6348 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_51
timestamp 1604681595
transform 1 0 5796 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_55
timestamp 1604681595
transform 1 0 6164 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_5_
timestamp 1604681595
transform 1 0 7820 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_5__S
timestamp 1604681595
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_65
timestamp 1604681595
transform 1 0 7084 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_69
timestamp 1604681595
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_82
timestamp 1604681595
transform 1 0 8648 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_3_
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_4__S
timestamp 1604681595
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_88
timestamp 1604681595
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_102
timestamp 1604681595
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1604681595
transform 1 0 11224 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 11040 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_106
timestamp 1604681595
transform 1 0 10856 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_119
timestamp 1604681595
transform 1 0 12052 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_125
timestamp 1604681595
transform 1 0 12604 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12788 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 13984 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1604681595
transform 1 0 13616 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_142
timestamp 1604681595
transform 1 0 14168 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_146
timestamp 1604681595
transform 1 0 14536 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_150
timestamp 1604681595
transform 1 0 14904 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_163
timestamp 1604681595
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16836 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 16652 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_167
timestamp 1604681595
transform 1 0 16468 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_180
timestamp 1604681595
transform 1 0 17664 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_186
timestamp 1604681595
transform 1 0 18216 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1604681595
transform 1 0 18400 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 19872 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19504 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_197
timestamp 1604681595
transform 1 0 19228 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_202
timestamp 1604681595
transform 1 0 19688 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_206
timestamp 1604681595
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 21896 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_210
timestamp 1604681595
transform 1 0 20424 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_224
timestamp 1604681595
transform 1 0 21712 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_228
timestamp 1604681595
transform 1 0 22080 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_1_
timestamp 1604681595
transform 1 0 24012 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 22448 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 23644 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 22264 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_241
timestamp 1604681595
transform 1 0 23276 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_247
timestamp 1604681595
transform 1 0 23828 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 25024 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 25392 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 25760 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_258
timestamp 1604681595
transform 1 0 24840 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_262
timestamp 1604681595
transform 1 0 25208 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_266
timestamp 1604681595
transform 1 0 25576 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_270
timestamp 1604681595
transform 1 0 25944 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 26128 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_274
timestamp 1604681595
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1604681595
transform 1 0 2944 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_7_
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_7__A1
timestamp 1604681595
transform 1 0 2760 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_12
timestamp 1604681595
transform 1 0 2208 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_16
timestamp 1604681595
transform 1 0 2576 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 3956 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3772 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_23
timestamp 1604681595
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_27
timestamp 1604681595
transform 1 0 3588 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 5888 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 6256 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_50
timestamp 1604681595
transform 1 0 5704 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1604681595
transform 1 0 6072 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_58
timestamp 1604681595
transform 1 0 6440 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 7176 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 6992 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_4_
timestamp 1604681595
transform 1 0 9660 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_4__A1
timestamp 1604681595
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_4__A0
timestamp 1604681595
transform 1 0 9108 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 10672 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_85
timestamp 1604681595
transform 1 0 8924 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_89
timestamp 1604681595
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_102
timestamp 1604681595
transform 1 0 10488 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1604681595
transform 1 0 11224 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 11040 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_106
timestamp 1604681595
transform 1 0 10856 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_114
timestamp 1604681595
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_118
timestamp 1604681595
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1604681595
transform 1 0 13984 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_132
timestamp 1604681595
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_136
timestamp 1604681595
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15548 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 15364 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 14996 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_149
timestamp 1604681595
transform 1 0 14812 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_153
timestamp 1604681595
transform 1 0 15180 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1604681595
transform 1 0 16376 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_170
timestamp 1604681595
transform 1 0 16744 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 16560 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_174
timestamp 1604681595
transform 1 0 17112 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 16928 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_179
timestamp 1604681595
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_184
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 18216 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 18400 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 19964 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 19780 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_197
timestamp 1604681595
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_201
timestamp 1604681595
transform 1 0 19596 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1604681595
transform 1 0 21528 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 20976 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 21344 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_214
timestamp 1604681595
transform 1 0 20792 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_218
timestamp 1604681595
transform 1 0 21160 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 22540 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 22908 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_231
timestamp 1604681595
transform 1 0 22356 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_235
timestamp 1604681595
transform 1 0 22724 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_239
timestamp 1604681595
transform 1 0 23092 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1604681595
transform 1 0 25208 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 24656 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1604681595
transform 1 0 25760 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_254
timestamp 1604681595
transform 1 0 24472 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_258
timestamp 1604681595
transform 1 0 24840 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_266
timestamp 1604681595
transform 1 0 25576 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_270
timestamp 1604681595
transform 1 0 25944 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 26128 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_274
timestamp 1604681595
transform 1 0 26312 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 1472 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 2944 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 2484 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_13
timestamp 1604681595
transform 1 0 2300 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_17
timestamp 1604681595
transform 1 0 2668 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 3312 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_22
timestamp 1604681595
transform 1 0 3128 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_26
timestamp 1604681595
transform 1 0 3496 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_41
timestamp 1604681595
transform 1 0 4876 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 5704 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 5152 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_1__A0
timestamp 1604681595
transform 1 0 5520 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 6716 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_46
timestamp 1604681595
transform 1 0 5336 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_59
timestamp 1604681595
transform 1 0 6532 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 7268 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 7084 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 8740 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l5_in_0__A0
timestamp 1604681595
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_63
timestamp 1604681595
transform 1 0 6900 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_76
timestamp 1604681595
transform 1 0 8096 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_81
timestamp 1604681595
transform 1 0 8556 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 9108 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1604681595
transform 1 0 8924 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_89
timestamp 1604681595
transform 1 0 9292 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_102
timestamp 1604681595
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1604681595
transform 1 0 11868 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1604681595
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11684 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_106
timestamp 1604681595
transform 1 0 10856 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_112
timestamp 1604681595
transform 1 0 11408 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13432 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 13248 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12880 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_126
timestamp 1604681595
transform 1 0 12696 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_130
timestamp 1604681595
transform 1 0 13064 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_143
timestamp 1604681595
transform 1 0 14260 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_147
timestamp 1604681595
transform 1 0 14628 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 18032 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17848 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 17480 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_173
timestamp 1604681595
transform 1 0 17020 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_177
timestamp 1604681595
transform 1 0 17388 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_180
timestamp 1604681595
transform 1 0 17664 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19964 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_203
timestamp 1604681595
transform 1 0 19780 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_207
timestamp 1604681595
transform 1 0 20148 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 21896 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_211
timestamp 1604681595
transform 1 0 20516 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_224
timestamp 1604681595
transform 1 0 21712 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_228
timestamp 1604681595
transform 1 0 22080 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 24012 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1604681595
transform 1 0 22448 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 23644 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 22264 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_241
timestamp 1604681595
transform 1 0 23276 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_247
timestamp 1604681595
transform 1 0 23828 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 25024 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 25392 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 25760 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_258
timestamp 1604681595
transform 1 0 24840 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_262
timestamp 1604681595
transform 1 0 25208 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_266
timestamp 1604681595
transform 1 0 25576 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_270
timestamp 1604681595
transform 1 0 25944 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 26128 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_274
timestamp 1604681595
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_4_
timestamp 1604681595
transform 1 0 2944 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 2760 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 2392 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_12
timestamp 1604681595
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_16
timestamp 1604681595
transform 1 0 2576 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_29
timestamp 1604681595
transform 1 0 3772 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_33
timestamp 1604681595
transform 1 0 4140 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_36
timestamp 1604681595
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_40
timestamp 1604681595
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5152 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_1__S
timestamp 1604681595
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_53
timestamp 1604681595
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1604681595
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_2_
timestamp 1604681595
transform 1 0 7544 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_2__S
timestamp 1604681595
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 6992 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 8556 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_66
timestamp 1604681595
transform 1 0 7176 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_79
timestamp 1604681595
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_83
timestamp 1604681595
transform 1 0 8740 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 9108 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10672 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 10488 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l5_in_0__S
timestamp 1604681595
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_96
timestamp 1604681595
transform 1 0 9936 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_100
timestamp 1604681595
transform 1 0 10304 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_113
timestamp 1604681595
transform 1 0 11500 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_118
timestamp 1604681595
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_4_
timestamp 1604681595
transform 1 0 13984 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_132
timestamp 1604681595
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_136
timestamp 1604681595
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15548 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_149
timestamp 1604681595
transform 1 0 14812 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_153
timestamp 1604681595
transform 1 0 15180 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_156
timestamp 1604681595
transform 1 0 15456 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1604681595
transform 1 0 16376 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_170
timestamp 1604681595
transform 1 0 16744 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 16560 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_174
timestamp 1604681595
transform 1 0 17112 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 16928 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_178
timestamp 1604681595
transform 1 0 17480 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17296 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_184
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 18216 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 18768 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 18584 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_188
timestamp 1604681595
transform 1 0 18400 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 21252 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 21068 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20700 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_211
timestamp 1604681595
transform 1 0 20516 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_215
timestamp 1604681595
transform 1 0 20884 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_228
timestamp 1604681595
transform 1 0 22080 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 22264 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 22632 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_232
timestamp 1604681595
transform 1 0 22448 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_236
timestamp 1604681595
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_240
timestamp 1604681595
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 25024 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_254
timestamp 1604681595
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_258
timestamp 1604681595
transform 1 0 24840 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_268
timestamp 1604681595
transform 1 0 25760 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 26312 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_272
timestamp 1604681595
transform 1 0 26128 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_276
timestamp 1604681595
transform 1 0 26496 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_10
timestamp 1604681595
transform 1 0 2024 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_6
timestamp 1604681595
transform 1 0 1656 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 1840 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_16
timestamp 1604681595
transform 1 0 2576 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_12
timestamp 1604681595
transform 1 0 2208 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 2760 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 2392 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1604681595
transform 1 0 2944 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 2392 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1604681595
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_23
timestamp 1604681595
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_37
timestamp 1604681595
transform 1 0 4508 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_33
timestamp 1604681595
transform 1 0 4140 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 4324 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4692 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4232 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4876 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_7_50
timestamp 1604681595
transform 1 0 5704 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_47
timestamp 1604681595
transform 1 0 5428 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_43
timestamp 1604681595
transform 1 0 5060 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_1__A1
timestamp 1604681595
transform 1 0 5612 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 5244 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_1_
timestamp 1604681595
transform 1 0 5796 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1604681595
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_54
timestamp 1604681595
transform 1 0 6072 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_60
timestamp 1604681595
transform 1 0 6624 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_2__A0
timestamp 1604681595
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 7360 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 7360 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 7176 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l5_in_0__A1
timestamp 1604681595
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 7176 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_2__A1
timestamp 1604681595
transform 1 0 8372 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_64
timestamp 1604681595
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_77
timestamp 1604681595
transform 1 0 8188 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_81
timestamp 1604681595
transform 1 0 8556 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_91
timestamp 1604681595
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_87
timestamp 1604681595
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_89
timestamp 1604681595
transform 1 0 9292 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1604681595
transform 1 0 8924 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_4__D
timestamp 1604681595
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 9108 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l5_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_102
timestamp 1604681595
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_4_
timestamp 1604681595
transform 1 0 9844 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_114
timestamp 1604681595
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_114
timestamp 1604681595
transform 1 0 11592 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_110
timestamp 1604681595
transform 1 0 11224 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_106
timestamp 1604681595
transform 1 0 10856 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 11040 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 11408 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_118
timestamp 1604681595
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11776 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11960 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 13984 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 14352 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_137
timestamp 1604681595
transform 1 0 13708 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_142
timestamp 1604681595
transform 1 0 14168 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_142
timestamp 1604681595
transform 1 0 14168 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_150
timestamp 1604681595
transform 1 0 14904 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_146
timestamp 1604681595
transform 1 0 14536 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_150
timestamp 1604681595
transform 1 0 14904 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_146
timestamp 1604681595
transform 1 0 14536 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14720 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 15088 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_2_
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_163
timestamp 1604681595
transform 1 0 16100 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16284 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15272 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_7_173
timestamp 1604681595
transform 1 0 17020 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_174
timestamp 1604681595
transform 1 0 17112 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_167
timestamp 1604681595
transform 1 0 16468 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 17296 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 16652 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1604681595
transform 1 0 16836 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_179
timestamp 1604681595
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_178
timestamp 1604681595
transform 1 0 17480 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 17664 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_4_
timestamp 1604681595
transform 1 0 17848 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_193
timestamp 1604681595
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_191
timestamp 1604681595
transform 1 0 18676 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 18860 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_201
timestamp 1604681595
transform 1 0 19596 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_197
timestamp 1604681595
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_195
timestamp 1604681595
transform 1 0 19044 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 19228 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19412 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_7_205
timestamp 1604681595
transform 1 0 19964 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_205
timestamp 1604681595
transform 1 0 19964 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19780 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 20240 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_215
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1604681595
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_209
timestamp 1604681595
transform 1 0 20332 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 21068 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 20424 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_229
timestamp 1604681595
transform 1 0 22172 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_219
timestamp 1604681595
transform 1 0 21252 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 21528 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 20424 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_7_237
timestamp 1604681595
transform 1 0 22908 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_233
timestamp 1604681595
transform 1 0 22540 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 22356 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_240
timestamp 1604681595
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_247
timestamp 1604681595
transform 1 0 23828 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_241
timestamp 1604681595
transform 1 0 23276 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 23644 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l4_in_0_
timestamp 1604681595
transform 1 0 24012 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_6_258
timestamp 1604681595
transform 1 0 24840 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 25024 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_264
timestamp 1604681595
transform 1 0 25392 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_262
timestamp 1604681595
transform 1 0 25208 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25392 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_266
timestamp 1604681595
transform 1 0 25576 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_4__CLK
timestamp 1604681595
transform 1 0 25576 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_268
timestamp 1604681595
transform 1 0 25760 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 25760 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_270
timestamp 1604681595
transform 1 0 25944 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 25944 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 26128 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 26312 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_274
timestamp 1604681595
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_272
timestamp 1604681595
transform 1 0 26128 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_276
timestamp 1604681595
transform 1 0 26496 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1472 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_27
timestamp 1604681595
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_23
timestamp 1604681595
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_36
timestamp 1604681595
transform 1 0 4416 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4600 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4232 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4784 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6716 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_59
timestamp 1604681595
transform 1 0 6532 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7268 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_7__S
timestamp 1604681595
transform 1 0 8280 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_3__A1
timestamp 1604681595
transform 1 0 8648 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_63
timestamp 1604681595
transform 1 0 6900 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_76
timestamp 1604681595
transform 1 0 8096 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_80
timestamp 1604681595
transform 1 0 8464 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10120 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 9936 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_84
timestamp 1604681595
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_88
timestamp 1604681595
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_93
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12604 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 12052 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_117
timestamp 1604681595
transform 1 0 11868 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_121
timestamp 1604681595
transform 1 0 12236 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1604681595
transform 1 0 14168 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 13616 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_134
timestamp 1604681595
transform 1 0 13432 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1604681595
transform 1 0 13800 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_145
timestamp 1604681595
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16192 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16008 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 15456 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_149
timestamp 1604681595
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_158
timestamp 1604681595
transform 1 0 15640 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1604681595
transform 1 0 17848 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 17664 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17296 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_173
timestamp 1604681595
transform 1 0 17020 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_178
timestamp 1604681595
transform 1 0 17480 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19412 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20148 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 19228 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 18860 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_191
timestamp 1604681595
transform 1 0 18676 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_195
timestamp 1604681595
transform 1 0 19044 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_205
timestamp 1604681595
transform 1 0 19964 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 21896 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20516 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_209
timestamp 1604681595
transform 1 0 20332 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1604681595
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_224
timestamp 1604681595
transform 1 0 21712 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_228
timestamp 1604681595
transform 1 0 22080 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 23276 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 22264 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 22632 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_232
timestamp 1604681595
transform 1 0 22448 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_236
timestamp 1604681595
transform 1 0 22816 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_240
timestamp 1604681595
transform 1 0 23184 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 25208 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25576 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 25944 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_260
timestamp 1604681595
transform 1 0 25024 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_264
timestamp 1604681595
transform 1 0 25392 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_268
timestamp 1604681595
transform 1 0 25760 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_272
timestamp 1604681595
transform 1 0 26128 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 1472 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2484 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_13
timestamp 1604681595
transform 1 0 2300 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_17
timestamp 1604681595
transform 1 0 2668 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 3956 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3772 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_21
timestamp 1604681595
transform 1 0 3036 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_27
timestamp 1604681595
transform 1 0 3588 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_40
timestamp 1604681595
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_44
timestamp 1604681595
transform 1 0 5152 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 5336 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_48
timestamp 1604681595
transform 1 0 5520 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1604681595
transform 1 0 5612 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_53
timestamp 1604681595
transform 1 0 5980 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_62
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_3_
timestamp 1604681595
transform 1 0 7544 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_7__A1
timestamp 1604681595
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_7__A0
timestamp 1604681595
transform 1 0 7360 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6992 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_66
timestamp 1604681595
transform 1 0 7176 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_79
timestamp 1604681595
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_83
timestamp 1604681595
transform 1 0 8740 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9844 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 9108 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 8924 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_90
timestamp 1604681595
transform 1 0 9384 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_3_
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_114
timestamp 1604681595
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_118
timestamp 1604681595
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1604681595
transform 1 0 13984 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_132
timestamp 1604681595
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_136
timestamp 1604681595
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_2_
timestamp 1604681595
transform 1 0 16376 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 15456 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 14996 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_149
timestamp 1604681595
transform 1 0 14812 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_153
timestamp 1604681595
transform 1 0 15180 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_158
timestamp 1604681595
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_162
timestamp 1604681595
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18216 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_175
timestamp 1604681595
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_179
timestamp 1604681595
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_184
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20148 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 19964 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19596 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_195
timestamp 1604681595
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_199
timestamp 1604681595
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_203
timestamp 1604681595
transform 1 0 19780 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1604681595
transform 1 0 21712 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 21528 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 21160 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_216
timestamp 1604681595
transform 1 0 20976 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_220
timestamp 1604681595
transform 1 0 21344 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 23920 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1604681595
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_233
timestamp 1604681595
transform 1 0 22540 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_237
timestamp 1604681595
transform 1 0 22908 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_240
timestamp 1604681595
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_245
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1604681595
transform 1 0 25484 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 24932 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 25300 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_257
timestamp 1604681595
transform 1 0 24748 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_261
timestamp 1604681595
transform 1 0 25116 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_269
timestamp 1604681595
transform 1 0 25852 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 26036 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 26404 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_273
timestamp 1604681595
transform 1 0 26220 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4692 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 4232 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 3312 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_22
timestamp 1604681595
transform 1 0 3128 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_26
timestamp 1604681595
transform 1 0 3496 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_36
timestamp 1604681595
transform 1 0 4416 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6348 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1604681595
transform 1 0 5704 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 6072 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_48
timestamp 1604681595
transform 1 0 5520 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_52
timestamp 1604681595
transform 1 0 5888 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_56
timestamp 1604681595
transform 1 0 6256 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_7_
timestamp 1604681595
transform 1 0 7912 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_3__S
timestamp 1604681595
transform 1 0 7544 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_66
timestamp 1604681595
transform 1 0 7176 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_72
timestamp 1604681595
transform 1 0 7728 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_83
timestamp 1604681595
transform 1 0 8740 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1604681595
transform 1 0 10120 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9844 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_3__A0
timestamp 1604681595
transform 1 0 8924 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_87
timestamp 1604681595
transform 1 0 9108 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_97
timestamp 1604681595
transform 1 0 10028 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1604681595
transform 1 0 11868 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11684 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11316 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_107
timestamp 1604681595
transform 1 0 10948 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_113
timestamp 1604681595
transform 1 0 11500 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 13432 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 12880 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13248 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_126
timestamp 1604681595
transform 1 0 12696 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_130
timestamp 1604681595
transform 1 0 13064 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_143
timestamp 1604681595
transform 1 0 14260 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1604681595
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_147
timestamp 1604681595
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_161
timestamp 1604681595
transform 1 0 15916 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_157
timestamp 1604681595
transform 1 0 15548 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 15732 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 16284 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18216 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_184
timestamp 1604681595
transform 1 0 18032 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18768 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 20148 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 18584 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 19780 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_188
timestamp 1604681595
transform 1 0 18400 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_201
timestamp 1604681595
transform 1 0 19596 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_205
timestamp 1604681595
transform 1 0 19964 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 20516 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_209
timestamp 1604681595
transform 1 0 20332 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_213
timestamp 1604681595
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1604681595
transform 1 0 23368 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 24012 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 22816 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 23184 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_234
timestamp 1604681595
transform 1 0 22632 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_238
timestamp 1604681595
transform 1 0 23000 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_246
timestamp 1604681595
transform 1 0 23736 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 24472 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1604681595
transform 1 0 25484 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 25852 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_251
timestamp 1604681595
transform 1 0 24196 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_263
timestamp 1604681595
transform 1 0 25300 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_267
timestamp 1604681595
transform 1 0 25668 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 26220 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_271
timestamp 1604681595
transform 1 0 26036 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2668 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2116 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_9
timestamp 1604681595
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_13
timestamp 1604681595
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 4232 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 3680 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_26
timestamp 1604681595
transform 1 0 3496 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_30
timestamp 1604681595
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_53
timestamp 1604681595
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1604681595
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_6_
timestamp 1604681595
transform 1 0 7912 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_6__A1
timestamp 1604681595
transform 1 0 7728 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_6__A0
timestamp 1604681595
transform 1 0 7360 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_66
timestamp 1604681595
transform 1 0 7176 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_70
timestamp 1604681595
transform 1 0 7544 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_83
timestamp 1604681595
transform 1 0 8740 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9476 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 9292 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 8924 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_87
timestamp 1604681595
transform 1 0 9108 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_97
timestamp 1604681595
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_101
timestamp 1604681595
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1604681595
transform 1 0 10764 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_114
timestamp 1604681595
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_118
timestamp 1604681595
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 13984 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1604681595
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_132
timestamp 1604681595
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_136
timestamp 1604681595
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 15916 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16284 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_159
timestamp 1604681595
transform 1 0 15732 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_163
timestamp 1604681595
transform 1 0 16100 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16468 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_173
timestamp 1604681595
transform 1 0 17020 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_179
timestamp 1604681595
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19964 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_203
timestamp 1604681595
transform 1 0 19780 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_207
timestamp 1604681595
transform 1 0 20148 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_3_
timestamp 1604681595
transform 1 0 20516 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 20332 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21528 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1604681595
transform 1 0 21896 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_220
timestamp 1604681595
transform 1 0 21344 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_224
timestamp 1604681595
transform 1 0 21712 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_228
timestamp 1604681595
transform 1 0 22080 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1604681595
transform 1 0 22448 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 22264 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_236
timestamp 1604681595
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_240
timestamp 1604681595
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1604681595
transform 1 0 25208 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1604681595
transform 1 0 25760 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 24656 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 25024 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_254
timestamp 1604681595
transform 1 0 24472 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_258
timestamp 1604681595
transform 1 0 24840 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_266
timestamp 1604681595
transform 1 0 25576 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_270
timestamp 1604681595
transform 1 0 25944 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 26128 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_274
timestamp 1604681595
transform 1 0 26312 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 2116 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_6
timestamp 1604681595
transform 1 0 1656 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_10
timestamp 1604681595
transform 1 0 2024 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_13
timestamp 1604681595
transform 1 0 2300 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_4_
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_23
timestamp 1604681595
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_41
timestamp 1604681595
transform 1 0 4876 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 6072 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1604681595
transform 1 0 5796 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 5520 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_46
timestamp 1604681595
transform 1 0 5336 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_50
timestamp 1604681595
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1604681595
transform 1 0 8556 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_6__S
timestamp 1604681595
transform 1 0 8004 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_73
timestamp 1604681595
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_77
timestamp 1604681595
transform 1 0 8188 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_84
timestamp 1604681595
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_88
timestamp 1604681595
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_102
timestamp 1604681595
transform 1 0 10488 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11500 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 10764 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 11132 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_107
timestamp 1604681595
transform 1 0 10948 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_111
timestamp 1604681595
transform 1 0 11316 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1604681595
transform 1 0 14076 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 13800 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_132
timestamp 1604681595
transform 1 0 13248 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_136
timestamp 1604681595
transform 1 0 13616 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_140
timestamp 1604681595
transform 1 0 13984 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_145
timestamp 1604681595
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14628 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_149
timestamp 1604681595
transform 1 0 14812 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 17940 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 17756 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 17204 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_173
timestamp 1604681595
transform 1 0 17020 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_177
timestamp 1604681595
transform 1 0 17388 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 19872 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_202
timestamp 1604681595
transform 1 0 19688 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_206
timestamp 1604681595
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 20424 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21896 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_213
timestamp 1604681595
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_224
timestamp 1604681595
transform 1 0 21712 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_228
timestamp 1604681595
transform 1 0 22080 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24012 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1604681595
transform 1 0 22448 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 23460 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23828 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 22264 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_241
timestamp 1604681595
transform 1 0 23276 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_245
timestamp 1604681595
transform 1 0 23644 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 25024 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25392 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 25760 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_258
timestamp 1604681595
transform 1 0 24840 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_262
timestamp 1604681595
transform 1 0 25208 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_266
timestamp 1604681595
transform 1 0 25576 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_270
timestamp 1604681595
transform 1 0 25944 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 26128 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_274
timestamp 1604681595
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_276
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 1564 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_7
timestamp 1604681595
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_6
timestamp 1604681595
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_1__S
timestamp 1604681595
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_10
timestamp 1604681595
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1604681595
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 2116 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_23
timestamp 1604681595
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_30
timestamp 1604681595
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_38
timestamp 1604681595
transform 1 0 4600 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_34
timestamp 1604681595
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_14_41
timestamp 1604681595
transform 1 0 4876 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_46
timestamp 1604681595
transform 1 0 5336 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 5152 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5612 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_58
timestamp 1604681595
transform 1 0 6440 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1604681595
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_53
timestamp 1604681595
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6624 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_62
timestamp 1604681595
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_66
timestamp 1604681595
transform 1 0 7176 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 7268 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7176 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 7452 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_79
timestamp 1604681595
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_75
timestamp 1604681595
transform 1 0 8004 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_82
timestamp 1604681595
transform 1 0 8648 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_78
timestamp 1604681595
transform 1 0 8280 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 8188 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 8464 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 8740 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9016 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 8832 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_86
timestamp 1604681595
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1604681595
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_102
timestamp 1604681595
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_110
timestamp 1604681595
transform 1 0 11224 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_106
timestamp 1604681595
transform 1 0 10856 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_109
timestamp 1604681595
transform 1 0 11132 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_105
timestamp 1604681595
transform 1 0 10764 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 11040 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 11500 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 10948 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_119
timestamp 1604681595
transform 1 0 12052 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_115
timestamp 1604681595
transform 1 0 11684 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 11500 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_14_132
timestamp 1604681595
transform 1 0 13248 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_132
timestamp 1604681595
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13432 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_140
timestamp 1604681595
transform 1 0 13984 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_136
timestamp 1604681595
transform 1 0 13616 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_136
timestamp 1604681595
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 13800 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1604681595
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13984 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1604681595
transform 1 0 14076 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_145
timestamp 1604681595
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_149
timestamp 1604681595
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_156
timestamp 1604681595
transform 1 0 15456 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_153
timestamp 1604681595
transform 1 0 15180 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_149
timestamp 1604681595
transform 1 0 14812 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1604681595
transform 1 0 16376 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15548 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_13_170
timestamp 1604681595
transform 1 0 16744 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16560 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_173
timestamp 1604681595
transform 1 0 17020 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 17204 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 17112 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_177
timestamp 1604681595
transform 1 0 17388 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_177
timestamp 1604681595
transform 1 0 17388 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 17664 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1604681595
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 17848 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1604681595
transform 1 0 18124 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1604681595
transform 1 0 18584 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 18676 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_188
timestamp 1604681595
transform 1 0 18400 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_192
timestamp 1604681595
transform 1 0 18768 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_189
timestamp 1604681595
transform 1 0 18492 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 18952 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 19044 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_193
timestamp 1604681595
transform 1 0 18860 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 19136 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 19228 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_206
timestamp 1604681595
transform 1 0 20056 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_205
timestamp 1604681595
transform 1 0 19964 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 20148 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 20240 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 20700 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 20516 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_209
timestamp 1604681595
transform 1 0 20332 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_210
timestamp 1604681595
transform 1 0 20424 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_238
timestamp 1604681595
transform 1 0 23000 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_234
timestamp 1604681595
transform 1 0 22632 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_236
timestamp 1604681595
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_232
timestamp 1604681595
transform 1 0 22448 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 22632 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 22816 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_240
timestamp 1604681595
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 23184 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 23368 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_14_251
timestamp 1604681595
transform 1 0 24196 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 24380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_255
timestamp 1604681595
transform 1 0 24564 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 24748 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1604681595
transform 1 0 24932 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_263
timestamp 1604681595
transform 1 0 25300 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_264
timestamp 1604681595
transform 1 0 25392 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_267
timestamp 1604681595
transform 1 0 25668 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_268
timestamp 1604681595
transform 1 0 25760 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 25852 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 25484 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1604681595
transform 1 0 25576 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 25944 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 26312 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 26220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_272
timestamp 1604681595
transform 1 0 26128 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_276
timestamp 1604681595
transform 1 0 26496 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_271
timestamp 1604681595
transform 1 0 26036 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_1_
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_12
timestamp 1604681595
transform 1 0 2208 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_16
timestamp 1604681595
transform 1 0 2576 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 3036 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_15_40
timestamp 1604681595
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_44
timestamp 1604681595
transform 1 0 5152 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1604681595
transform 1 0 5336 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1604681595
transform 1 0 5520 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1604681595
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_52
timestamp 1604681595
transform 1 0 5888 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_71
timestamp 1604681595
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_75
timestamp 1604681595
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_79
timestamp 1604681595
transform 1 0 8372 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_83
timestamp 1604681595
transform 1 0 8740 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9016 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_113
timestamp 1604681595
transform 1 0 11500 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_109
timestamp 1604681595
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_105
timestamp 1604681595
transform 1 0 10764 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_118
timestamp 1604681595
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1604681595
transform 1 0 13984 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_132
timestamp 1604681595
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_136
timestamp 1604681595
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_3_
timestamp 1604681595
transform 1 0 16376 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_149
timestamp 1604681595
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_153
timestamp 1604681595
transform 1 0 15180 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_158
timestamp 1604681595
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_162
timestamp 1604681595
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 18216 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1604681595
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_175
timestamp 1604681595
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_179
timestamp 1604681595
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_184
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1604681595
transform 1 0 18400 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 19504 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 19320 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 18952 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_192
timestamp 1604681595
transform 1 0 18768 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_196
timestamp 1604681595
transform 1 0 19136 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 21068 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 20884 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 20516 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 22080 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_209
timestamp 1604681595
transform 1 0 20332 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_213
timestamp 1604681595
transform 1 0 20700 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_226
timestamp 1604681595
transform 1 0 21896 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_4_
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A
timestamp 1604681595
transform 1 0 22448 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_4__D
timestamp 1604681595
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_230
timestamp 1604681595
transform 1 0 22264 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_234
timestamp 1604681595
transform 1 0 22632 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_240
timestamp 1604681595
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 25576 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_4__CLK
timestamp 1604681595
transform 1 0 25944 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_264
timestamp 1604681595
transform 1 0 25392 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_268
timestamp 1604681595
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 26312 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_272
timestamp 1604681595
transform 1 0 26128 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_276
timestamp 1604681595
transform 1 0 26496 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_6
timestamp 1604681595
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_10
timestamp 1604681595
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_23
timestamp 1604681595
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1604681595
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6532 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 5980 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6348 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_51
timestamp 1604681595
transform 1 0 5796 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_55
timestamp 1604681595
transform 1 0 6164 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1604681595
transform 1 0 8556 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 8372 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 8004 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 7636 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_68
timestamp 1604681595
transform 1 0 7360 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_73
timestamp 1604681595
transform 1 0 7820 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_77
timestamp 1604681595
transform 1 0 8188 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1604681595
transform 1 0 10212 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 9844 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_84
timestamp 1604681595
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_88
timestamp 1604681595
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_97
timestamp 1604681595
transform 1 0 10028 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 11776 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 11224 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 11592 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_108
timestamp 1604681595
transform 1 0 11040 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_112
timestamp 1604681595
transform 1 0 11408 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 13984 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 14352 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_135
timestamp 1604681595
transform 1 0 13524 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1604681595
transform 1 0 13892 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_142
timestamp 1604681595
transform 1 0 14168 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15640 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14720 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 15456 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_146
timestamp 1604681595
transform 1 0 14536 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_150
timestamp 1604681595
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_154
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 18308 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 17572 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_177
timestamp 1604681595
transform 1 0 17388 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_181
timestamp 1604681595
transform 1 0 17756 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_186
timestamp 1604681595
transform 1 0 18216 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 20240 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_206
timestamp 1604681595
transform 1 0 20056 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 21896 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_210
timestamp 1604681595
transform 1 0 20424 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_224
timestamp 1604681595
transform 1 0 21712 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_228
timestamp 1604681595
transform 1 0 22080 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1604681595
transform 1 0 22448 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23644 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 22264 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1604681595
transform 1 0 23000 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 23368 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_236
timestamp 1604681595
transform 1 0 22816 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_240
timestamp 1604681595
transform 1 0 23184 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_244
timestamp 1604681595
transform 1 0 23552 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 25576 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 25944 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_264
timestamp 1604681595
transform 1 0 25392 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_268
timestamp 1604681595
transform 1 0 25760 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_272
timestamp 1604681595
transform 1 0 26128 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_2_
timestamp 1604681595
transform 1 0 2576 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1604681595
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_7
timestamp 1604681595
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_11
timestamp 1604681595
transform 1 0 2116 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 4140 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1604681595
transform 1 0 3956 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_25
timestamp 1604681595
transform 1 0 3404 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_29
timestamp 1604681595
transform 1 0 3772 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_52
timestamp 1604681595
transform 1 0 5888 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1604681595
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 8372 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_71
timestamp 1604681595
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_75
timestamp 1604681595
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 9384 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_88
timestamp 1604681595
transform 1 0 9200 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_92
timestamp 1604681595
transform 1 0 9568 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_97
timestamp 1604681595
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_101
timestamp 1604681595
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12512 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1604681595
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_114
timestamp 1604681595
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_118
timestamp 1604681595
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1604681595
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_143
timestamp 1604681595
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1604681595
transform 1 0 15272 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1604681595
transform 1 0 15088 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_147
timestamp 1604681595
transform 1 0 14628 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_151
timestamp 1604681595
transform 1 0 14996 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_158
timestamp 1604681595
transform 1 0 15640 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_162
timestamp 1604681595
transform 1 0 16008 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_4_
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1604681595
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_179
timestamp 1604681595
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 19964 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19136 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 19780 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_193
timestamp 1604681595
transform 1 0 18860 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_198
timestamp 1604681595
transform 1 0 19320 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_202
timestamp 1604681595
transform 1 0 19688 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 21528 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 20976 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 21344 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_214
timestamp 1604681595
transform 1 0 20792 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_218
timestamp 1604681595
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 22540 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_231
timestamp 1604681595
transform 1 0 22356 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_235
timestamp 1604681595
transform 1 0 22724 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_240
timestamp 1604681595
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1604681595
transform 1 0 25208 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1604681595
transform 1 0 25760 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 24656 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_254
timestamp 1604681595
transform 1 0 24472 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_258
timestamp 1604681595
transform 1 0 24840 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_266
timestamp 1604681595
transform 1 0 25576 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_270
timestamp 1604681595
transform 1 0 25944 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 26128 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_274
timestamp 1604681595
transform 1 0 26312 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_6
timestamp 1604681595
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_10
timestamp 1604681595
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4876 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1604681595
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_36
timestamp 1604681595
transform 1 0 4416 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_40
timestamp 1604681595
transform 1 0 4784 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 5428 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 5244 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_43
timestamp 1604681595
transform 1 0 5060 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 7360 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 7728 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_66
timestamp 1604681595
transform 1 0 7176 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_70
timestamp 1604681595
transform 1 0 7544 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_74
timestamp 1604681595
transform 1 0 7912 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_84
timestamp 1604681595
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_88
timestamp 1604681595
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_98
timestamp 1604681595
transform 1 0 10120 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1604681595
transform 1 0 9844 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_102
timestamp 1604681595
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 10304 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10856 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12604 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12052 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_115
timestamp 1604681595
transform 1 0 11684 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_121
timestamp 1604681595
transform 1 0 12236 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1604681595
transform 1 0 14444 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 16008 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 15824 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 15456 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_149
timestamp 1604681595
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_154
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_158
timestamp 1604681595
transform 1 0 15640 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 18032 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_181
timestamp 1604681595
transform 1 0 17756 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_186
timestamp 1604681595
transform 1 0 18216 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19136 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18952 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 18584 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 20148 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_192
timestamp 1604681595
transform 1 0 18768 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_205
timestamp 1604681595
transform 1 0 19964 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 22080 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_209
timestamp 1604681595
transform 1 0 20332 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_224
timestamp 1604681595
transform 1 0 21712 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1604681595
transform 1 0 22632 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23736 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 22448 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 23184 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 23552 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_230
timestamp 1604681595
transform 1 0 22264 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_238
timestamp 1604681595
transform 1 0 23000 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_242
timestamp 1604681595
transform 1 0 23368 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25668 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_265
timestamp 1604681595
transform 1 0 25484 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_269
timestamp 1604681595
transform 1 0 25852 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 26036 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_273
timestamp 1604681595
transform 1 0 26220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1564 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_30
timestamp 1604681595
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1604681595
transform 1 0 3496 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_22
timestamp 1604681595
transform 1 0 3128 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_28
timestamp 1604681595
transform 1 0 3680 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_24
timestamp 1604681595
transform 1 0 3312 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 3680 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3312 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 3496 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 3956 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_33
timestamp 1604681595
transform 1 0 4140 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4692 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 4508 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_37
timestamp 1604681595
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_36
timestamp 1604681595
transform 1 0 4416 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4692 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4876 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_52
timestamp 1604681595
transform 1 0 5888 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_48
timestamp 1604681595
transform 1 0 5520 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_50
timestamp 1604681595
transform 1 0 5704 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l5_in_0__A1
timestamp 1604681595
transform 1 0 5704 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1604681595
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_54
timestamp 1604681595
transform 1 0 6072 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6072 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 6256 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_19_72
timestamp 1604681595
transform 1 0 7728 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_2_
timestamp 1604681595
transform 1 0 6900 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1604681595
transform 1 0 8648 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_79
timestamp 1604681595
transform 1 0 8372 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_75
timestamp 1604681595
transform 1 0 8004 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_76
timestamp 1604681595
transform 1 0 8096 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8464 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 7912 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 8280 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 8464 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1604681595
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_99
timestamp 1604681595
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_103
timestamp 1604681595
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_86
timestamp 1604681595
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 1604681595
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_112
timestamp 1604681595
transform 1 0 11408 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_114
timestamp 1604681595
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_107
timestamp 1604681595
transform 1 0 10948 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11592 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 10764 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1604681595
transform 1 0 11316 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_116
timestamp 1604681595
transform 1 0 11776 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_118
timestamp 1604681595
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 11960 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1604681595
transform 1 0 12144 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_134
timestamp 1604681595
transform 1 0 13432 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_129
timestamp 1604681595
transform 1 0 12972 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 13248 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1604681595
transform 1 0 13248 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1604681595
transform 1 0 13800 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_141
timestamp 1604681595
transform 1 0 14076 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 13984 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 14260 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 13616 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1604681595
transform 1 0 14168 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_145
timestamp 1604681595
transform 1 0 14444 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_145
timestamp 1604681595
transform 1 0 14444 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1604681595
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 14812 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 14628 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1604681595
transform 1 0 14812 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_162
timestamp 1604681595
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_158
timestamp 1604681595
transform 1 0 15640 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1604681595
transform 1 0 16376 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_20_173
timestamp 1604681595
transform 1 0 17020 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_175
timestamp 1604681595
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17204 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_177
timestamp 1604681595
transform 1 0 17388 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_179
timestamp 1604681595
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 17572 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l4_in_0_
timestamp 1604681595
transform 1 0 17756 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 18308 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1604681595
transform 1 0 18952 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_190
timestamp 1604681595
transform 1 0 18584 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 19136 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 18768 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_206
timestamp 1604681595
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_198
timestamp 1604681595
transform 1 0 19320 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_208
timestamp 1604681595
transform 1 0 20240 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1604681595
transform 1 0 20240 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 19504 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1604681595
transform 1 0 19688 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18492 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_210
timestamp 1604681595
transform 1 0 20424 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_212
timestamp 1604681595
transform 1 0 20608 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1604681595
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 20424 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1604681595
transform 1 0 20792 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 20976 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1604681595
transform 1 0 20976 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_224
timestamp 1604681595
transform 1 0 21712 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_220
timestamp 1604681595
transform 1 0 21344 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_229
timestamp 1604681595
transform 1 0 22172 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1604681595
transform 1 0 21804 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 21896 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 21988 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 21528 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 22080 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_19_236
timestamp 1604681595
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 22356 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1604681595
transform 1 0 22540 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_247
timestamp 1604681595
transform 1 0 23828 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_240
timestamp 1604681595
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l4_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 24012 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_251
timestamp 1604681595
transform 1 0 24196 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_258
timestamp 1604681595
transform 1 0 24840 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_254
timestamp 1604681595
transform 1 0 24472 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 24380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 24656 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_1_
timestamp 1604681595
transform 1 0 24564 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_268
timestamp 1604681595
transform 1 0 25760 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_264
timestamp 1604681595
transform 1 0 25392 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_268
timestamp 1604681595
transform 1 0 25760 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25576 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 25024 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 25944 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 25944 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 26312 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_272
timestamp 1604681595
transform 1 0 26128 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_276
timestamp 1604681595
transform 1 0 26496 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_272
timestamp 1604681595
transform 1 0 26128 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_4_
timestamp 1604681595
transform 1 0 1564 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1604681595
transform 1 0 4048 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1604681595
transform 1 0 3864 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_1__A1
timestamp 1604681595
transform 1 0 3496 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_24
timestamp 1604681595
transform 1 0 3312 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_28
timestamp 1604681595
transform 1 0 3680 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_36
timestamp 1604681595
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_40
timestamp 1604681595
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1604681595
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_53
timestamp 1604681595
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1604681595
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8464 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8280 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_71
timestamp 1604681595
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_75
timestamp 1604681595
transform 1 0 8004 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10028 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 9476 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_89
timestamp 1604681595
transform 1 0 9292 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_93
timestamp 1604681595
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_106
timestamp 1604681595
transform 1 0 10856 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11040 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1604681595
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604681595
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_114
timestamp 1604681595
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_123
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 13064 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12880 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_127
timestamp 1604681595
transform 1 0 12788 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1604681595
transform 1 0 16376 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 16192 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 15824 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15456 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15088 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_149
timestamp 1604681595
transform 1 0 14812 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_154
timestamp 1604681595
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_158
timestamp 1604681595
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_162
timestamp 1604681595
transform 1 0 16008 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_175
timestamp 1604681595
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_179
timestamp 1604681595
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 20240 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_203
timestamp 1604681595
transform 1 0 19780 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_207
timestamp 1604681595
transform 1 0 20148 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1604681595
transform 1 0 20792 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 20608 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 21804 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 22172 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_210
timestamp 1604681595
transform 1 0 20424 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_223
timestamp 1604681595
transform 1 0 21620 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_227
timestamp 1604681595
transform 1 0 21988 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1604681595
transform 1 0 22448 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1604681595
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_231
timestamp 1604681595
transform 1 0 22356 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_236
timestamp 1604681595
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_240
timestamp 1604681595
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 25576 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25944 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_264
timestamp 1604681595
transform 1 0 25392 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_268
timestamp 1604681595
transform 1 0 25760 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 26312 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_272
timestamp 1604681595
transform 1 0 26128 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_276
timestamp 1604681595
transform 1 0 26496 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1604681595
transform 1 0 2944 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l5_in_0_
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l5_in_0__S
timestamp 1604681595
transform 1 0 2392 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_4__D
timestamp 1604681595
transform 1 0 2760 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_12
timestamp 1604681595
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_16
timestamp 1604681595
transform 1 0 2576 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_1__A0
timestamp 1604681595
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_23
timestamp 1604681595
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6532 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6348 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 5980 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_51
timestamp 1604681595
transform 1 0 5796 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_55
timestamp 1604681595
transform 1 0 6164 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1604681595
transform 1 0 8096 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8648 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 7544 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7912 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_68
timestamp 1604681595
transform 1 0 7360 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_72
timestamp 1604681595
transform 1 0 7728 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_80
timestamp 1604681595
transform 1 0 8464 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10396 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 9200 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10028 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_84
timestamp 1604681595
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1604681595
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_99
timestamp 1604681595
transform 1 0 10212 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 12328 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_120
timestamp 1604681595
transform 1 0 12144 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_124
timestamp 1604681595
transform 1 0 12512 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12880 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 13892 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12696 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14260 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_137
timestamp 1604681595
transform 1 0 13708 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1604681595
transform 1 0 14076 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_145
timestamp 1604681595
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_154
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_149
timestamp 1604681595
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1604681595
transform 1 0 15364 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_165
timestamp 1604681595
transform 1 0 16284 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_162
timestamp 1604681595
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_158
timestamp 1604681595
transform 1 0 15640 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 16100 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16376 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_2_
timestamp 1604681595
transform 1 0 17940 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 17664 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_175
timestamp 1604681595
transform 1 0 17204 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_179
timestamp 1604681595
transform 1 0 17572 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_182
timestamp 1604681595
transform 1 0 17848 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1604681595
transform 1 0 19688 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19228 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 20240 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1604681595
transform 1 0 18768 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_196
timestamp 1604681595
transform 1 0 19136 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_199
timestamp 1604681595
transform 1 0 19412 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_206
timestamp 1604681595
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 21252 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21068 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_210
timestamp 1604681595
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_228
timestamp 1604681595
transform 1 0 22080 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1604681595
transform 1 0 22816 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23828 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23644 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23276 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 22448 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_234
timestamp 1604681595
transform 1 0 22632 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_239
timestamp 1604681595
transform 1 0 23092 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_243
timestamp 1604681595
transform 1 0 23460 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 25760 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_266
timestamp 1604681595
transform 1 0 25576 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_270
timestamp 1604681595
transform 1 0 25944 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 26128 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_274
timestamp 1604681595
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 2760 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1472 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 2576 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 2208 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_10
timestamp 1604681595
transform 1 0 2024 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_14
timestamp 1604681595
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 4692 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_37
timestamp 1604681595
transform 1 0 4508 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_41
timestamp 1604681595
transform 1 0 4876 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5244 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 5060 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1604681595
transform 1 0 5796 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1604681595
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8740 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_81
timestamp 1604681595
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9292 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9108 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_85
timestamp 1604681595
transform 1 0 8924 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11224 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_108
timestamp 1604681595
transform 1 0 11040 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_112
timestamp 1604681595
transform 1 0 11408 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_118
timestamp 1604681595
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 13984 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_132
timestamp 1604681595
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_136
timestamp 1604681595
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 16100 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_159
timestamp 1604681595
transform 1 0 15732 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_165
timestamp 1604681595
transform 1 0 16284 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1604681595
transform 1 0 16836 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1604681595
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 16468 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1604681595
transform 1 0 16652 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_175
timestamp 1604681595
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_179
timestamp 1604681595
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19964 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_203
timestamp 1604681595
transform 1 0 19780 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_207
timestamp 1604681595
transform 1 0 20148 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 20976 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 20516 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20332 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_214
timestamp 1604681595
transform 1 0 20792 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 22908 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_235
timestamp 1604681595
transform 1 0 22724 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_239
timestamp 1604681595
transform 1 0 23092 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 24656 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 25024 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_254
timestamp 1604681595
transform 1 0 24472 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_258
timestamp 1604681595
transform 1 0 24840 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_268
timestamp 1604681595
transform 1 0 25760 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 26312 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_272
timestamp 1604681595
transform 1 0 26128 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_276
timestamp 1604681595
transform 1 0 26496 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 2208 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_3__S
timestamp 1604681595
transform 1 0 1564 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_2__S
timestamp 1604681595
transform 1 0 1932 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_7
timestamp 1604681595
transform 1 0 1748 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_11
timestamp 1604681595
transform 1 0 2116 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1604681595
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_25
timestamp 1604681595
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_21
timestamp 1604681595
transform 1 0 3036 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_36
timestamp 1604681595
transform 1 0 4416 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_32
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 4508 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1604681595
transform 1 0 4692 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 6256 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 5704 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 6072 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_48
timestamp 1604681595
transform 1 0 5520 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_52
timestamp 1604681595
transform 1 0 5888 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 8740 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_2__A1
timestamp 1604681595
transform 1 0 8188 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_3__A1
timestamp 1604681595
transform 1 0 8556 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_75
timestamp 1604681595
transform 1 0 8004 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_79
timestamp 1604681595
transform 1 0 8372 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10672 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 10212 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_86
timestamp 1604681595
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1604681595
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_96
timestamp 1604681595
transform 1 0 9936 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_101
timestamp 1604681595
transform 1 0 10396 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 12604 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_123
timestamp 1604681595
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 13156 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 14168 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 12972 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_127
timestamp 1604681595
transform 1 0 12788 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_140
timestamp 1604681595
transform 1 0 13984 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_144
timestamp 1604681595
transform 1 0 14352 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 1604681595
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_148
timestamp 1604681595
transform 1 0 14720 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14904 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 14536 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_162
timestamp 1604681595
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_158
timestamp 1604681595
transform 1 0 15640 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 15824 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 15456 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_3_
timestamp 1604681595
transform 1 0 16100 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_1_
timestamp 1604681595
transform 1 0 17664 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 17480 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 17112 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_172
timestamp 1604681595
transform 1 0 16928 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_176
timestamp 1604681595
transform 1 0 17296 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19044 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 18676 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 20240 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_189
timestamp 1604681595
transform 1 0 18492 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_193
timestamp 1604681595
transform 1 0 18860 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_206
timestamp 1604681595
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 21896 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_210
timestamp 1604681595
transform 1 0 20424 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_224
timestamp 1604681595
transform 1 0 21712 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_228
timestamp 1604681595
transform 1 0 22080 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1604681595
transform 1 0 24012 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1604681595
transform 1 0 22448 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 23644 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 22264 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_241
timestamp 1604681595
transform 1 0 23276 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_247
timestamp 1604681595
transform 1 0 23828 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 25024 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 25392 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 25760 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_258
timestamp 1604681595
transform 1 0 24840 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_262
timestamp 1604681595
transform 1 0 25208 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_266
timestamp 1604681595
transform 1 0 25576 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_270
timestamp 1604681595
transform 1 0 25944 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 26128 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_274
timestamp 1604681595
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_3_
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_12
timestamp 1604681595
transform 1 0 2208 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_18
timestamp 1604681595
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 3128 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4692 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 4140 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4508 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_31
timestamp 1604681595
transform 1 0 3956 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_35
timestamp 1604681595
transform 1 0 4324 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 6256 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 5704 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 6072 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_48
timestamp 1604681595
transform 1 0 5520 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_52
timestamp 1604681595
transform 1 0 5888 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1604681595
transform 1 0 8648 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 7084 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 8464 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8096 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_74
timestamp 1604681595
transform 1 0 7912 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_78
timestamp 1604681595
transform 1 0 8280 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l4_in_0_
timestamp 1604681595
transform 1 0 10212 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9660 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10028 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_91
timestamp 1604681595
transform 1 0 9476 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_95
timestamp 1604681595
transform 1 0 9844 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_3_
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11224 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_108
timestamp 1604681595
transform 1 0 11040 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_112
timestamp 1604681595
transform 1 0 11408 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_118
timestamp 1604681595
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 14352 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 13800 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_132
timestamp 1604681595
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_136
timestamp 1604681595
transform 1 0 13616 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_140
timestamp 1604681595
transform 1 0 13984 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 14536 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_25_165
timestamp 1604681595
transform 1 0 16284 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 17572 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 16468 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1604681595
transform 1 0 17020 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_169
timestamp 1604681595
transform 1 0 16652 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_175
timestamp 1604681595
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 1604681595
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 20148 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_203
timestamp 1604681595
transform 1 0 19780 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l4_in_0_
timestamp 1604681595
transform 1 0 20700 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 20516 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 21712 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_209
timestamp 1604681595
transform 1 0 20332 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1604681595
transform 1 0 21528 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_226
timestamp 1604681595
transform 1 0 21896 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1604681595
transform 1 0 22448 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1604681595
transform 1 0 22264 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_236
timestamp 1604681595
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_240
timestamp 1604681595
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 24656 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 25024 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_254
timestamp 1604681595
transform 1 0 24472 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_258
timestamp 1604681595
transform 1 0 24840 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_268
timestamp 1604681595
transform 1 0 25760 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 26312 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_272
timestamp 1604681595
transform 1 0 26128 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_276
timestamp 1604681595
transform 1 0 26496 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_2_
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_5_
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_16
timestamp 1604681595
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_12
timestamp 1604681595
transform 1 0 2208 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_16
timestamp 1604681595
transform 1 0 2576 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_12
timestamp 1604681595
transform 1 0 2208 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l5_in_0__A0
timestamp 1604681595
transform 1 0 2760 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_7__S
timestamp 1604681595
transform 1 0 2392 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_7__A0
timestamp 1604681595
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_7__A1
timestamp 1604681595
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_20
timestamp 1604681595
transform 1 0 2944 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1604681595
transform 1 0 2944 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_23
timestamp 1604681595
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1604681595
transform 1 0 3128 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_35
timestamp 1604681595
transform 1 0 4324 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_31
timestamp 1604681595
transform 1 0 3956 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 4140 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4508 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4692 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_41
timestamp 1604681595
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_52
timestamp 1604681595
transform 1 0 5888 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_48
timestamp 1604681595
transform 1 0 5520 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_45
timestamp 1604681595
transform 1 0 5244 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 5428 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 5704 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5612 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1604681595
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_62
timestamp 1604681595
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_58
timestamp 1604681595
transform 1 0 6440 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6624 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7176 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 8648 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 6992 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_2__A0
timestamp 1604681595
transform 1 0 8188 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_75
timestamp 1604681595
transform 1 0 8004 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_79
timestamp 1604681595
transform 1 0 8372 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_81
timestamp 1604681595
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_85
timestamp 1604681595
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_91
timestamp 1604681595
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_88
timestamp 1604681595
transform 1 0 9200 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_84
timestamp 1604681595
transform 1 0 8832 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 9292 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 9108 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_3_
timestamp 1604681595
transform 1 0 9292 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_102
timestamp 1604681595
transform 1 0 10488 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_98
timestamp 1604681595
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_102
timestamp 1604681595
transform 1 0 10488 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 10304 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 10672 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_114
timestamp 1604681595
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1604681595
transform 1 0 11224 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_114
timestamp 1604681595
transform 1 0 11592 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_110
timestamp 1604681595
transform 1 0 11224 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_106
timestamp 1604681595
transform 1 0 10856 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 11408 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 11040 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 11408 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1604681595
transform 1 0 10856 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_118
timestamp 1604681595
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 11684 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_27_132
timestamp 1604681595
transform 1 0 13248 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_134
timestamp 1604681595
transform 1 0 13432 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_138
timestamp 1604681595
transform 1 0 13800 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1604681595
transform 1 0 13800 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13616 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13616 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_144
timestamp 1604681595
transform 1 0 14352 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13984 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 14168 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1604681595
transform 1 0 14168 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_145
timestamp 1604681595
transform 1 0 14444 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 14720 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1604681595
transform 1 0 15456 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 14536 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 14628 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_149
timestamp 1604681595
transform 1 0 14812 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_154
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_165
timestamp 1604681595
transform 1 0 16284 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 16836 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 16468 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_169
timestamp 1604681595
transform 1 0 16652 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_167
timestamp 1604681595
transform 1 0 16468 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_171
timestamp 1604681595
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1604681595
transform 1 0 17020 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 17204 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 16928 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_174
timestamp 1604681595
transform 1 0 17112 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_177
timestamp 1604681595
transform 1 0 17388 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_178
timestamp 1604681595
transform 1 0 17480 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_181
timestamp 1604681595
transform 1 0 17756 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 17572 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17940 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_2_
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18124 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1604681595
transform 1 0 19780 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 19044 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1604681595
transform 1 0 19596 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20056 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_204
timestamp 1604681595
transform 1 0 19872 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_208
timestamp 1604681595
transform 1 0 20240 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_193
timestamp 1604681595
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_197
timestamp 1604681595
transform 1 0 19228 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_207
timestamp 1604681595
transform 1 0 20148 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 20884 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 20700 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 20332 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_211
timestamp 1604681595
transform 1 0 20516 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_238
timestamp 1604681595
transform 1 0 23000 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_234
timestamp 1604681595
transform 1 0 22632 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_238
timestamp 1604681595
transform 1 0 23000 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_234
timestamp 1604681595
transform 1 0 22632 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 22816 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 23184 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_3_
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_3_
timestamp 1604681595
transform 1 0 23368 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_254
timestamp 1604681595
transform 1 0 24472 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_255
timestamp 1604681595
transform 1 0 24564 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_251
timestamp 1604681595
transform 1 0 24196 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 24380 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 24656 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_258
timestamp 1604681595
transform 1 0 24840 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 24748 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 25024 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24932 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1604681595
transform 1 0 25208 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_270
timestamp 1604681595
transform 1 0 25944 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_266
timestamp 1604681595
transform 1 0 25576 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_269
timestamp 1604681595
transform 1 0 25852 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_265
timestamp 1604681595
transform 1 0 25484 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25668 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1604681595
transform 1 0 25760 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 26036 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 26128 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_273
timestamp 1604681595
transform 1 0 26220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_274
timestamp 1604681595
transform 1 0 26312 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_7_
timestamp 1604681595
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_5__A1
timestamp 1604681595
transform 1 0 1840 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_5__A0
timestamp 1604681595
transform 1 0 2208 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_6
timestamp 1604681595
transform 1 0 1656 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_10
timestamp 1604681595
transform 1 0 2024 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 4140 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l4_in_1__S
timestamp 1604681595
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_23
timestamp 1604681595
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_27
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6624 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 6072 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6440 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_52
timestamp 1604681595
transform 1 0 5888 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_56
timestamp 1604681595
transform 1 0 6256 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8188 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 7636 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8004 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_69
timestamp 1604681595
transform 1 0 7452 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_73
timestamp 1604681595
transform 1 0 7820 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_83
timestamp 1604681595
transform 1 0 8740 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_2_
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 9292 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 8924 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_87
timestamp 1604681595
transform 1 0 9108 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_91
timestamp 1604681595
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_102
timestamp 1604681595
transform 1 0 10488 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 11224 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1604681595
transform 1 0 11040 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 12420 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_106
timestamp 1604681595
transform 1 0 10856 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_119
timestamp 1604681595
transform 1 0 12052 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_125
timestamp 1604681595
transform 1 0 12604 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 13156 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_129
timestamp 1604681595
transform 1 0 12972 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_133
timestamp 1604681595
transform 1 0 13340 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_145
timestamp 1604681595
transform 1 0 14444 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 16284 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_149
timestamp 1604681595
transform 1 0 14812 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_163
timestamp 1604681595
transform 1 0 16100 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 16928 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 16744 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_167
timestamp 1604681595
transform 1 0 16468 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19504 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 18860 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19228 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20240 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_191
timestamp 1604681595
transform 1 0 18676 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_195
timestamp 1604681595
transform 1 0 19044 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_199
timestamp 1604681595
transform 1 0 19412 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_206
timestamp 1604681595
transform 1 0 20056 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_1_
timestamp 1604681595
transform 1 0 20976 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 21988 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_210
timestamp 1604681595
transform 1 0 20424 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_225
timestamp 1604681595
transform 1 0 21804 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_229
timestamp 1604681595
transform 1 0 22172 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_3_
timestamp 1604681595
transform 1 0 24104 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_2_
timestamp 1604681595
transform 1 0 22540 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 23644 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 22356 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_242
timestamp 1604681595
transform 1 0 23368 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_247
timestamp 1604681595
transform 1 0 23828 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 25116 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 25484 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 25852 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_259
timestamp 1604681595
transform 1 0 24932 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_263
timestamp 1604681595
transform 1 0 25300 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_267
timestamp 1604681595
transform 1 0 25668 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 26220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_271
timestamp 1604681595
transform 1 0 26036 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_3_
timestamp 1604681595
transform 1 0 2024 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_5__S
timestamp 1604681595
transform 1 0 1564 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_7
timestamp 1604681595
transform 1 0 1748 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_19
timestamp 1604681595
transform 1 0 2852 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 3588 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1604681595
transform 1 0 4600 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3404 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_3__S
timestamp 1604681595
transform 1 0 3036 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_23
timestamp 1604681595
transform 1 0 3220 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_36
timestamp 1604681595
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_40
timestamp 1604681595
transform 1 0 4784 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_53
timestamp 1604681595
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1604681595
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_62
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 7728 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1604681595
transform 1 0 7544 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6992 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_66
timestamp 1604681595
transform 1 0 7176 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_4_
timestamp 1604681595
transform 1 0 10488 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 10304 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 9936 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_91
timestamp 1604681595
transform 1 0 9476 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_95
timestamp 1604681595
transform 1 0 9844 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_98
timestamp 1604681595
transform 1 0 10120 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 11500 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_111
timestamp 1604681595
transform 1 0 11316 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_115
timestamp 1604681595
transform 1 0 11684 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_119
timestamp 1604681595
transform 1 0 12052 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13524 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1604681595
transform 1 0 12972 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13340 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_127
timestamp 1604681595
transform 1 0 12788 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_131
timestamp 1604681595
transform 1 0 13156 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_144
timestamp 1604681595
transform 1 0 14352 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 15456 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 15272 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 14904 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14536 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_148
timestamp 1604681595
transform 1 0 14720 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_152
timestamp 1604681595
transform 1 0 15088 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_175
timestamp 1604681595
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_179
timestamp 1604681595
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 19688 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 19504 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_193
timestamp 1604681595
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_197
timestamp 1604681595
transform 1 0 19228 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 22172 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 21988 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 21620 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_221
timestamp 1604681595
transform 1 0 21436 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1604681595
transform 1 0 21804 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 22908 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_235
timestamp 1604681595
transform 1 0 22724 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_239
timestamp 1604681595
transform 1 0 23092 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1604681595
transform 1 0 25208 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 24656 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1604681595
transform 1 0 25760 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 25024 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_254
timestamp 1604681595
transform 1 0 24472 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_258
timestamp 1604681595
transform 1 0 24840 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_266
timestamp 1604681595
transform 1 0 25576 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_270
timestamp 1604681595
transform 1 0 25944 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 26128 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_274
timestamp 1604681595
transform 1 0 26312 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_6__A1
timestamp 1604681595
transform 1 0 2024 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 1656 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_8
timestamp 1604681595
transform 1 0 1840 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_12
timestamp 1604681595
transform 1 0 2208 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_2__S
timestamp 1604681595
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 4600 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_23
timestamp 1604681595
transform 1 0 3220 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1604681595
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_36
timestamp 1604681595
transform 1 0 4416 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_40
timestamp 1604681595
transform 1 0 4784 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6808 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5244 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 5060 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6624 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 6256 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_54
timestamp 1604681595
transform 1 0 6072 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_58
timestamp 1604681595
transform 1 0 6440 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1604681595
transform 1 0 8372 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 7820 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 8188 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_71
timestamp 1604681595
transform 1 0 7636 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_75
timestamp 1604681595
transform 1 0 8004 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_83
timestamp 1604681595
transform 1 0 8740 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 9016 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_88
timestamp 1604681595
transform 1 0 9200 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 12144 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 11592 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11960 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_112
timestamp 1604681595
transform 1 0 11408 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_116
timestamp 1604681595
transform 1 0 11776 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14076 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14444 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_139
timestamp 1604681595
transform 1 0 13892 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_143
timestamp 1604681595
transform 1 0 14260 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 16284 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_147
timestamp 1604681595
transform 1 0 14628 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_163
timestamp 1604681595
transform 1 0 16100 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16836 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 18032 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 16652 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_167
timestamp 1604681595
transform 1 0 16468 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_180
timestamp 1604681595
transform 1 0 17664 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_186
timestamp 1604681595
transform 1 0 18216 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18400 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 20240 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 19596 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_197
timestamp 1604681595
transform 1 0 19228 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_203
timestamp 1604681595
transform 1 0 19780 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_207
timestamp 1604681595
transform 1 0 20148 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 21896 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_210
timestamp 1604681595
transform 1 0 20424 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_224
timestamp 1604681595
transform 1 0 21712 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_228
timestamp 1604681595
transform 1 0 22080 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_2_
timestamp 1604681595
transform 1 0 24012 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l4_in_0_
timestamp 1604681595
transform 1 0 22448 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 23644 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 22264 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_241
timestamp 1604681595
transform 1 0 23276 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_247
timestamp 1604681595
transform 1 0 23828 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_2__A0
timestamp 1604681595
transform 1 0 25024 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_3__A1
timestamp 1604681595
transform 1 0 25392 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25760 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_258
timestamp 1604681595
transform 1 0 24840 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_262
timestamp 1604681595
transform 1 0 25208 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_266
timestamp 1604681595
transform 1 0 25576 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_270
timestamp 1604681595
transform 1 0 25944 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 26128 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_274
timestamp 1604681595
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_276
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_6_
timestamp 1604681595
transform 1 0 2024 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_6__A0
timestamp 1604681595
transform 1 0 1840 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_7
timestamp 1604681595
transform 1 0 1748 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_19
timestamp 1604681595
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_2_
timestamp 1604681595
transform 1 0 3588 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 3036 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 3404 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_23
timestamp 1604681595
transform 1 0 3220 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_36
timestamp 1604681595
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_40
timestamp 1604681595
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 5152 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_53
timestamp 1604681595
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1604681595
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_62
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 7268 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 7084 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 8280 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_2__A1
timestamp 1604681595
transform 1 0 8648 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_76
timestamp 1604681595
transform 1 0 8096 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_80
timestamp 1604681595
transform 1 0 8464 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1604681595
transform 1 0 8832 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9844 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 9660 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 9292 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_87
timestamp 1604681595
transform 1 0 9108 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_91
timestamp 1604681595
transform 1 0 9476 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_114
timestamp 1604681595
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_118
timestamp 1604681595
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12880 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 12696 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15364 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 15180 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 14812 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 16376 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_147
timestamp 1604681595
transform 1 0 14628 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_151
timestamp 1604681595
transform 1 0 14996 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_164
timestamp 1604681595
transform 1 0 16192 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_168
timestamp 1604681595
transform 1 0 16560 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 16744 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1604681595
transform 1 0 16928 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_175
timestamp 1604681595
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_179
timestamp 1604681595
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_184
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 18216 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 18676 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_31_188
timestamp 1604681595
transform 1 0 18400 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1604681595
transform 1 0 21160 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20884 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_210
timestamp 1604681595
transform 1 0 20424 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_214
timestamp 1604681595
transform 1 0 20792 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_217
timestamp 1604681595
transform 1 0 21068 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_227
timestamp 1604681595
transform 1 0 21988 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_2_
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 22448 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 22816 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_2__S
timestamp 1604681595
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_231
timestamp 1604681595
transform 1 0 22356 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_234
timestamp 1604681595
transform 1 0 22632 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_238
timestamp 1604681595
transform 1 0 23000 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604681595
transform 1 0 25208 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1604681595
transform 1 0 25760 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_3__S
timestamp 1604681595
transform 1 0 24656 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_2__A1
timestamp 1604681595
transform 1 0 25024 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_254
timestamp 1604681595
transform 1 0 24472 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_258
timestamp 1604681595
transform 1 0 24840 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_266
timestamp 1604681595
transform 1 0 25576 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_270
timestamp 1604681595
transform 1 0 25944 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_3__A0
timestamp 1604681595
transform 1 0 26128 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_274
timestamp 1604681595
transform 1 0 26312 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 2392 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_4__A0
timestamp 1604681595
transform 1 0 1564 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_6__S
timestamp 1604681595
transform 1 0 2024 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_7
timestamp 1604681595
transform 1 0 1748 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_12
timestamp 1604681595
transform 1 0 2208 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 3404 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_3__A0
timestamp 1604681595
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_23
timestamp 1604681595
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_27
timestamp 1604681595
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6808 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5980 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6348 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_51
timestamp 1604681595
transform 1 0 5796 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_55
timestamp 1604681595
transform 1 0 6164 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_59
timestamp 1604681595
transform 1 0 6532 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 8740 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_81
timestamp 1604681595
transform 1 0 8556 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1604681595
transform 1 0 9936 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_85
timestamp 1604681595
transform 1 0 8924 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_89
timestamp 1604681595
transform 1 0 9292 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1604681595
transform 1 0 11500 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 12512 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 10948 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 11316 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_105
timestamp 1604681595
transform 1 0 10764 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_109
timestamp 1604681595
transform 1 0 11132 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_122
timestamp 1604681595
transform 1 0 12328 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 13064 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12880 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 14076 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_126
timestamp 1604681595
transform 1 0 12696 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_139
timestamp 1604681595
transform 1 0 13892 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_143
timestamp 1604681595
transform 1 0 14260 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15364 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14628 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_149
timestamp 1604681595
transform 1 0 14812 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_154
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 17848 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 17664 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 17296 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_174
timestamp 1604681595
transform 1 0 17112 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_178
timestamp 1604681595
transform 1 0 17480 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 19780 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20240 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_201
timestamp 1604681595
transform 1 0 19596 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_205
timestamp 1604681595
transform 1 0 19964 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 21896 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_210
timestamp 1604681595
transform 1 0 20424 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_224
timestamp 1604681595
transform 1 0 21712 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_228
timestamp 1604681595
transform 1 0 22080 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_3_
timestamp 1604681595
transform 1 0 24012 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_2_
timestamp 1604681595
transform 1 0 22448 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 23644 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 22264 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_241
timestamp 1604681595
transform 1 0 23276 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_247
timestamp 1604681595
transform 1 0 23828 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 25024 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 25392 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25760 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_258
timestamp 1604681595
transform 1 0 24840 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_262
timestamp 1604681595
transform 1 0 25208 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_266
timestamp 1604681595
transform 1 0 25576 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_270
timestamp 1604681595
transform 1 0 25944 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 26128 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_274
timestamp 1604681595
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_7
timestamp 1604681595
transform 1 0 1748 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_4__S
timestamp 1604681595
transform 1 0 1932 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_4__A1
timestamp 1604681595
transform 1 0 1564 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_4_
timestamp 1604681595
transform 1 0 1564 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_34_11
timestamp 1604681595
transform 1 0 2116 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_18
timestamp 1604681595
transform 1 0 2760 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_14
timestamp 1604681595
transform 1 0 2392 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 2576 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 2944 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1604681595
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_23
timestamp 1604681595
transform 1 0 3220 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_31
timestamp 1604681595
transform 1 0 3956 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 3128 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_36
timestamp 1604681595
transform 1 0 4416 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_32
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_35
timestamp 1604681595
transform 1 0 4324 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l4_in_1__A0
timestamp 1604681595
transform 1 0 4600 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 4232 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4508 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4140 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4692 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_4_
timestamp 1604681595
transform 1 0 4784 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_33_48
timestamp 1604681595
transform 1 0 5520 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_4__D
timestamp 1604681595
transform 1 0 5704 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_56
timestamp 1604681595
transform 1 0 6256 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_52
timestamp 1604681595
transform 1 0 5888 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 6072 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_59
timestamp 1604681595
transform 1 0 6532 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 6808 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_71
timestamp 1604681595
transform 1 0 7636 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_68
timestamp 1604681595
transform 1 0 7360 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_64
timestamp 1604681595
transform 1 0 6992 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_70
timestamp 1604681595
transform 1 0 7544 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_66
timestamp 1604681595
transform 1 0 7176 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 7452 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 7360 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 7728 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_74
timestamp 1604681595
transform 1 0 7912 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 7820 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 8096 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 8004 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 8280 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_34_91
timestamp 1604681595
transform 1 0 9476 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_88
timestamp 1604681595
transform 1 0 9200 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_84
timestamp 1604681595
transform 1 0 8832 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_91
timestamp 1604681595
transform 1 0 9476 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_87
timestamp 1604681595
transform 1 0 9108 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 9292 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 9292 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 9660 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_104
timestamp 1604681595
transform 1 0 10672 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 9844 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_34_112
timestamp 1604681595
transform 1 0 11408 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_112
timestamp 1604681595
transform 1 0 11408 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_108
timestamp 1604681595
transform 1 0 11040 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 11224 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 10856 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 11684 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_118
timestamp 1604681595
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_117
timestamp 1604681595
transform 1 0 11868 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12420 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 12052 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_121
timestamp 1604681595
transform 1 0 12236 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_34_125
timestamp 1604681595
transform 1 0 12604 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 12696 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 13432 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 14444 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 13800 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_132
timestamp 1604681595
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_136
timestamp 1604681595
transform 1 0 13616 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_140
timestamp 1604681595
transform 1 0 13984 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_144
timestamp 1604681595
transform 1 0 14352 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_145
timestamp 1604681595
transform 1 0 14444 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_154
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_149
timestamp 1604681595
transform 1 0 14812 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_156
timestamp 1604681595
transform 1 0 15456 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14628 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 15456 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1604681595
transform 1 0 14628 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_158
timestamp 1604681595
transform 1 0 15640 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_160
timestamp 1604681595
transform 1 0 15824 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 15640 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 16008 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1604681595
transform 1 0 16192 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 15824 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_33_173
timestamp 1604681595
transform 1 0 17020 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_186
timestamp 1604681595
transform 1 0 18216 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_183
timestamp 1604681595
transform 1 0 17940 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_179
timestamp 1604681595
transform 1 0 17572 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_177
timestamp 1604681595
transform 1 0 17388 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 18032 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_2_
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1604681595
transform 1 0 18308 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_34_196
timestamp 1604681595
transform 1 0 19136 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_197
timestamp 1604681595
transform 1 0 19228 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_193
timestamp 1604681595
transform 1 0 18860 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_207
timestamp 1604681595
transform 1 0 20148 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_203
timestamp 1604681595
transform 1 0 19780 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_200
timestamp 1604681595
transform 1 0 19504 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 19964 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 19412 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 19596 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1604681595
transform 1 0 19596 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_34_211
timestamp 1604681595
transform 1 0 20516 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_217
timestamp 1604681595
transform 1 0 21068 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_214
timestamp 1604681595
transform 1 0 20792 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_210
timestamp 1604681595
transform 1 0 20424 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 20332 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 20884 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21160 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_228
timestamp 1604681595
transform 1 0 22080 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_224
timestamp 1604681595
transform 1 0 21712 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_227
timestamp 1604681595
transform 1 0 21988 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 21896 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 22172 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_1__A1
timestamp 1604681595
transform 1 0 22540 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 22264 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_231
timestamp 1604681595
transform 1 0 22356 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_232
timestamp 1604681595
transform 1 0 22448 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 22724 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_235
timestamp 1604681595
transform 1 0 22724 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 22908 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_1__A0
timestamp 1604681595
transform 1 0 23092 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_239
timestamp 1604681595
transform 1 0 23092 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_237
timestamp 1604681595
transform 1 0 22908 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_243
timestamp 1604681595
transform 1 0 23460 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_1__S
timestamp 1604681595
transform 1 0 23276 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_1_
timestamp 1604681595
transform 1 0 23276 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1604681595
transform 1 0 24104 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_254
timestamp 1604681595
transform 1 0 24472 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_254
timestamp 1604681595
transform 1 0 24472 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 24656 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 24288 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 24840 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 24840 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_34_267 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 25668 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_268
timestamp 1604681595
transform 1 0 25760 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_260
timestamp 1604681595
transform 1 0 25024 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 25944 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_272
timestamp 1604681595
transform 1 0 26128 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_276
timestamp 1604681595
transform 1 0 26496 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 2668 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 2484 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 2116 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_9
timestamp 1604681595
transform 1 0 1932 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_13
timestamp 1604681595
transform 1 0 2300 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 4232 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 4048 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3680 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_26
timestamp 1604681595
transform 1 0 3496 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_30
timestamp 1604681595
transform 1 0 3864 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_51
timestamp 1604681595
transform 1 0 5796 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_47
timestamp 1604681595
transform 1 0 5428 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_43
timestamp 1604681595
transform 1 0 5060 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l5_in_0__A1
timestamp 1604681595
transform 1 0 5612 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l5_in_0__S
timestamp 1604681595
transform 1 0 5244 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_55
timestamp 1604681595
transform 1 0 6164 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l5_in_0__A0
timestamp 1604681595
transform 1 0 5980 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 8740 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_81
timestamp 1604681595
transform 1 0 8556 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 9292 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A
timestamp 1604681595
transform 1 0 9108 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_85
timestamp 1604681595
transform 1 0 8924 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11224 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_108
timestamp 1604681595
transform 1 0 11040 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_112
timestamp 1604681595
transform 1 0 11408 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_118
timestamp 1604681595
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13616 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13984 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14352 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_132
timestamp 1604681595
transform 1 0 13248 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_138
timestamp 1604681595
transform 1 0 13800 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_142
timestamp 1604681595
transform 1 0 14168 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 14904 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 14720 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_146
timestamp 1604681595
transform 1 0 14536 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 16836 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1604681595
transform 1 0 16652 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_173
timestamp 1604681595
transform 1 0 17020 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_177
timestamp 1604681595
transform 1 0 17388 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_3_
timestamp 1604681595
transform 1 0 19596 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 19412 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 19044 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_193
timestamp 1604681595
transform 1 0 18860 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_197
timestamp 1604681595
transform 1 0 19228 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21160 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 22172 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20976 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_210
timestamp 1604681595
transform 1 0 20424 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_214
timestamp 1604681595
transform 1 0 20792 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_227
timestamp 1604681595
transform 1 0 21988 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l5_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 22540 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l5_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_231
timestamp 1604681595
transform 1 0 22356 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_235
timestamp 1604681595
transform 1 0 22724 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_240
timestamp 1604681595
transform 1 0 23184 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1604681595
transform 1 0 25208 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1604681595
transform 1 0 25760 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 24656 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l5_in_0__A0
timestamp 1604681595
transform 1 0 25024 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_254
timestamp 1604681595
transform 1 0 24472 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_258
timestamp 1604681595
transform 1 0 24840 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_266
timestamp 1604681595
transform 1 0 25576 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_270 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 25944 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_276
timestamp 1604681595
transform 1 0 26496 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1932 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 2668 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1604681595
transform 1 0 1380 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_7
timestamp 1604681595
transform 1 0 1748 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_15
timestamp 1604681595
transform 1 0 2484 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_19
timestamp 1604681595
transform 1 0 2852 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_27
timestamp 1604681595
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_23
timestamp 1604681595
transform 1 0 3220 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3404 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l4_in_1__A1
timestamp 1604681595
transform 1 0 3036 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_36
timestamp 1604681595
transform 1 0 4416 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_32
timestamp 1604681595
transform 1 0 4048 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 4232 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l5_in_0_
timestamp 1604681595
transform 1 0 4692 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6164 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6808 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 5704 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_48
timestamp 1604681595
transform 1 0 5520 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_52
timestamp 1604681595
transform 1 0 5888 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_57
timestamp 1604681595
transform 1 0 6348 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_61
timestamp 1604681595
transform 1 0 6716 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6992 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_36_83
timestamp 1604681595
transform 1 0 8740 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _129_
timestamp 1604681595
transform 1 0 9844 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 9200 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10396 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_87
timestamp 1604681595
transform 1 0 9108 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_90
timestamp 1604681595
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_93
timestamp 1604681595
transform 1 0 9660 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_99
timestamp 1604681595
transform 1 0 10212 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_103
timestamp 1604681595
transform 1 0 10580 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10948 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 10764 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12880 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 13432 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_126
timestamp 1604681595
transform 1 0 12696 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_130
timestamp 1604681595
transform 1 0 13064 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_145
timestamp 1604681595
transform 1 0 14444 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 16284 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 14996 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 14628 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_149
timestamp 1604681595
transform 1 0 14812 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_163
timestamp 1604681595
transform 1 0 16100 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_3_
timestamp 1604681595
transform 1 0 16836 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 18032 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 16652 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_167
timestamp 1604681595
transform 1 0 16468 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_180
timestamp 1604681595
transform 1 0 17664 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_186
timestamp 1604681595
transform 1 0 18216 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18400 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 19596 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 19964 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_197
timestamp 1604681595
transform 1 0 19228 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_203
timestamp 1604681595
transform 1 0 19780 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_207
timestamp 1604681595
transform 1 0 20148 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1604681595
transform 1 0 20884 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 21896 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21344 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 21712 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20608 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_211
timestamp 1604681595
transform 1 0 20516 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_218
timestamp 1604681595
transform 1 0 21160 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_222
timestamp 1604681595
transform 1 0 21528 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1604681595
transform 1 0 23920 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l5_in_0__S
timestamp 1604681595
transform 1 0 23644 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 23276 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 22908 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_235
timestamp 1604681595
transform 1 0 22724 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_239
timestamp 1604681595
transform 1 0 23092 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_243
timestamp 1604681595
transform 1 0 23460 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_247
timestamp 1604681595
transform 1 0 23828 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_257 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 24748 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_269
timestamp 1604681595
transform 1 0 25852 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1604681595
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1604681595
transform 1 0 2484 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1604681595
transform 1 0 1380 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__A
timestamp 1604681595
transform 1 0 1932 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2300 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_7
timestamp 1604681595
transform 1 0 1748 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_11
timestamp 1604681595
transform 1 0 2116 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_19
timestamp 1604681595
transform 1 0 2852 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1604681595
transform 1 0 3588 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1604681595
transform 1 0 4140 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A
timestamp 1604681595
transform 1 0 3036 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4600 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 3404 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_23
timestamp 1604681595
transform 1 0 3220 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_31
timestamp 1604681595
transform 1 0 3956 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_35
timestamp 1604681595
transform 1 0 4324 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_40
timestamp 1604681595
transform 1 0 4784 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4968 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_53
timestamp 1604681595
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1604681595
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_62
timestamp 1604681595
transform 1 0 6808 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7360 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7176 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8372 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8740 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_77
timestamp 1604681595
transform 1 0 8188 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_81
timestamp 1604681595
transform 1 0 8556 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 9200 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 10580 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 10212 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_85
timestamp 1604681595
transform 1 0 8924 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_97
timestamp 1604681595
transform 1 0 10028 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_101
timestamp 1604681595
transform 1 0 10396 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_114
timestamp 1604681595
transform 1 0 11592 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_118
timestamp 1604681595
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1604681595
transform 1 0 14076 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13432 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 13800 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_132
timestamp 1604681595
transform 1 0 13248 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_136
timestamp 1604681595
transform 1 0 13616 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_140
timestamp 1604681595
transform 1 0 13984 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_145
timestamp 1604681595
transform 1 0 14444 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l4_in_0_
timestamp 1604681595
transform 1 0 15180 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 14996 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1604681595
transform 1 0 16284 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 14628 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_149
timestamp 1604681595
transform 1 0 14812 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_162
timestamp 1604681595
transform 1 0 16008 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1604681595
transform 1 0 16836 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 18032 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 16652 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_167
timestamp 1604681595
transform 1 0 16468 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_175
timestamp 1604681595
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_179
timestamp 1604681595
transform 1 0 17572 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 19596 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 19044 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 19412 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_193
timestamp 1604681595
transform 1 0 18860 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_197
timestamp 1604681595
transform 1 0 19228 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21436 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 21068 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 20608 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_210
timestamp 1604681595
transform 1 0 20424 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_214
timestamp 1604681595
transform 1 0 20792 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_219
timestamp 1604681595
transform 1 0 21252 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_234
timestamp 1604681595
transform 1 0 22632 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_230
timestamp 1604681595
transform 1 0 22264 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 23000 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 22448 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_245
timestamp 1604681595
transform 1 0 23644 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_240
timestamp 1604681595
transform 1 0 23184 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 23368 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 23828 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1604681595
transform 1 0 24012 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25024 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_258
timestamp 1604681595
transform 1 0 24840 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_262
timestamp 1604681595
transform 1 0 25208 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_274
timestamp 1604681595
transform 1 0 26312 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2208 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__056__A
timestamp 1604681595
transform 1 0 1564 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_3__A1
timestamp 1604681595
transform 1 0 2024 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_3__A0
timestamp 1604681595
transform 1 0 2944 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1604681595
transform 1 0 1380 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_7
timestamp 1604681595
transform 1 0 1748 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_18
timestamp 1604681595
transform 1 0 2760 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_26
timestamp 1604681595
transform 1 0 3496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_22
timestamp 1604681595
transform 1 0 3128 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_2__A0
timestamp 1604681595
transform 1 0 3588 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_32
timestamp 1604681595
transform 1 0 4048 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1604681595
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 4232 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_36
timestamp 1604681595
transform 1 0 4416 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 4692 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4876 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6164 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5612 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 5980 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_47
timestamp 1604681595
transform 1 0 5428 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_51
timestamp 1604681595
transform 1 0 5796 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7728 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7360 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_64
timestamp 1604681595
transform 1 0 6992 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_70
timestamp 1604681595
transform 1 0 7544 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_81
timestamp 1604681595
transform 1 0 8556 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_93
timestamp 1604681595
transform 1 0 9660 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_91
timestamp 1604681595
transform 1 0 9476 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_87
timestamp 1604681595
transform 1 0 9108 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 8924 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 9292 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_100
timestamp 1604681595
transform 1 0 10304 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_97
timestamp 1604681595
transform 1 0 10028 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 10120 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10488 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10672 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12236 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 11684 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 12052 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_113
timestamp 1604681595
transform 1 0 11500 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_117
timestamp 1604681595
transform 1 0 11868 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13800 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13248 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 13616 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_130
timestamp 1604681595
transform 1 0 13064 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_134
timestamp 1604681595
transform 1 0 13432 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_144
timestamp 1604681595
transform 1 0 14352 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 14536 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 14904 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16284 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_148
timestamp 1604681595
transform 1 0 14720 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_152
timestamp 1604681595
transform 1 0 15088 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_163
timestamp 1604681595
transform 1 0 16100 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1604681595
transform 1 0 16836 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18032 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 16652 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_167
timestamp 1604681595
transform 1 0 16468 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_180
timestamp 1604681595
transform 1 0 17664 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_186
timestamp 1604681595
transform 1 0 18216 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1604681595
transform 1 0 18400 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20148 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 19412 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 19780 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1604681595
transform 1 0 19228 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_201
timestamp 1604681595
transform 1 0 19596 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_205
timestamp 1604681595
transform 1 0 19964 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 21068 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 22080 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_209
timestamp 1604681595
transform 1 0 20332 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_215
timestamp 1604681595
transform 1 0 20884 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_226
timestamp 1604681595
transform 1 0 21896 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1604681595
transform 1 0 23460 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 23276 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 22908 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 22448 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_230
timestamp 1604681595
transform 1 0 22264 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_234
timestamp 1604681595
transform 1 0 22632 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_239
timestamp 1604681595
transform 1 0 23092 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25024 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 24472 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 24840 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_252
timestamp 1604681595
transform 1 0 24288 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_256
timestamp 1604681595
transform 1 0 24656 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_266
timestamp 1604681595
transform 1 0 25576 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604681595
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_274
timestamp 1604681595
transform 1 0 26312 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_276
timestamp 1604681595
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1604681595
transform 1 0 1380 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1604681595
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_7
timestamp 1604681595
transform 1 0 1748 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_7
timestamp 1604681595
transform 1 0 1748 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 1932 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__057__A
timestamp 1604681595
transform 1 0 1932 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_11
timestamp 1604681595
transform 1 0 2116 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_11
timestamp 1604681595
transform 1 0 2116 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 2300 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__058__A
timestamp 1604681595
transform 1 0 2300 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_19
timestamp 1604681595
transform 1 0 2852 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_19
timestamp 1604681595
transform 1 0 2852 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1604681595
transform 1 0 2484 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1604681595
transform 1 0 2484 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_23
timestamp 1604681595
transform 1 0 3220 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_23
timestamp 1604681595
transform 1 0 3220 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3036 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_4__CLK
timestamp 1604681595
transform 1 0 3404 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A
timestamp 1604681595
transform 1 0 3036 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1604681595
transform 1 0 3588 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_36
timestamp 1604681595
transform 1 0 4416 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_32
timestamp 1604681595
transform 1 0 4048 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_35
timestamp 1604681595
transform 1 0 4324 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_31
timestamp 1604681595
transform 1 0 3956 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 4232 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A
timestamp 1604681595
transform 1 0 4140 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_5__S
timestamp 1604681595
transform 1 0 4600 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604681595
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_40
timestamp 1604681595
transform 1 0 4784 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_4__CLK
timestamp 1604681595
transform 1 0 4784 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_46
timestamp 1604681595
transform 1 0 5336 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_42
timestamp 1604681595
transform 1 0 4968 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_5__A1
timestamp 1604681595
transform 1 0 5152 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_5__A0
timestamp 1604681595
transform 1 0 4968 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_5_
timestamp 1604681595
transform 1 0 5152 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _133_
timestamp 1604681595
transform 1 0 6164 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__A
timestamp 1604681595
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 5980 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_53
timestamp 1604681595
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_52
timestamp 1604681595
transform 1 0 5888 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604681595
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__A
timestamp 1604681595
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6716 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1604681595
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_59
timestamp 1604681595
transform 1 0 6532 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_62
timestamp 1604681595
transform 1 0 6808 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_40_67
timestamp 1604681595
transform 1 0 7268 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_63
timestamp 1604681595
transform 1 0 6900 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__A
timestamp 1604681595
transform 1 0 7084 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _131_
timestamp 1604681595
transform 1 0 7084 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_72
timestamp 1604681595
transform 1 0 7728 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_69
timestamp 1604681595
transform 1 0 7452 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7728 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _134_
timestamp 1604681595
transform 1 0 7360 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_76
timestamp 1604681595
transform 1 0 8096 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_74
timestamp 1604681595
transform 1 0 7912 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__A
timestamp 1604681595
transform 1 0 8188 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _127_
timestamp 1604681595
transform 1 0 8188 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_79
timestamp 1604681595
transform 1 0 8372 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_81
timestamp 1604681595
transform 1 0 8556 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _130_
timestamp 1604681595
transform 1 0 8464 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__A
timestamp 1604681595
transform 1 0 8740 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_93
timestamp 1604681595
transform 1 0 9660 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_91
timestamp 1604681595
transform 1 0 9476 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_88
timestamp 1604681595
transform 1 0 9200 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_84
timestamp 1604681595
transform 1 0 8832 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_85
timestamp 1604681595
transform 1 0 8924 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 9292 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 9108 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604681595
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 9292 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_40_97
timestamp 1604681595
transform 1 0 10028 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_102
timestamp 1604681595
transform 1 0 10488 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_98
timestamp 1604681595
transform 1 0 10120 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 9844 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 10304 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1604681595
transform 1 0 10120 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 10672 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_111
timestamp 1604681595
transform 1 0 11316 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_107
timestamp 1604681595
transform 1 0 10948 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_114
timestamp 1604681595
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_106
timestamp 1604681595
transform 1 0 10856 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 11500 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11040 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 11132 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1604681595
transform 1 0 11224 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_118
timestamp 1604681595
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1604681595
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604681595
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 11684 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1604681595
transform 1 0 12420 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_124
timestamp 1604681595
transform 1 0 12512 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_128
timestamp 1604681595
transform 1 0 12880 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_132
timestamp 1604681595
transform 1 0 13248 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 13064 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 12696 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13432 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13248 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_40_141
timestamp 1604681595
transform 1 0 14076 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_140
timestamp 1604681595
transform 1 0 13984 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_136
timestamp 1604681595
transform 1 0 13616 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 14352 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13800 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 14352 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_150
timestamp 1604681595
transform 1 0 14904 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_146
timestamp 1604681595
transform 1 0 14536 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_155
timestamp 1604681595
transform 1 0 15364 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 14720 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604681595
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_3_
timestamp 1604681595
transform 1 0 14536 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_163
timestamp 1604681595
transform 1 0 16100 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_159
timestamp 1604681595
transform 1 0 15732 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16284 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_4__S
timestamp 1604681595
transform 1 0 15916 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 15548 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16100 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_167
timestamp 1604681595
transform 1 0 16468 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_176
timestamp 1604681595
transform 1 0 17296 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_172
timestamp 1604681595
transform 1 0 16928 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16652 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_4__A1
timestamp 1604681595
transform 1 0 17112 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_4_
timestamp 1604681595
transform 1 0 16836 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_186
timestamp 1604681595
transform 1 0 18216 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_180
timestamp 1604681595
transform 1 0 17664 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_180
timestamp 1604681595
transform 1 0 17664 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18032 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_4__A0
timestamp 1604681595
transform 1 0 17480 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604681595
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1604681595
transform 1 0 18952 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_197
timestamp 1604681595
transform 1 0 19228 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_193
timestamp 1604681595
transform 1 0 18860 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19136 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19044 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18400 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_206
timestamp 1604681595
transform 1 0 20056 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_198
timestamp 1604681595
transform 1 0 19320 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_203
timestamp 1604681595
transform 1 0 19780 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 19504 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19596 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19964 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20148 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1604681595
transform 1 0 19688 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1604681595
transform 1 0 20240 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_215
timestamp 1604681595
transform 1 0 20884 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_210
timestamp 1604681595
transform 1 0 20424 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_216
timestamp 1604681595
transform 1 0 20976 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 20608 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_5__A1
timestamp 1604681595
transform 1 0 21160 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604681595
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_5_
timestamp 1604681595
transform 1 0 20976 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_225
timestamp 1604681595
transform 1 0 21804 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_220
timestamp 1604681595
transform 1 0 21344 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_5__A0
timestamp 1604681595
transform 1 0 21528 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_6__A1
timestamp 1604681595
transform 1 0 21988 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 21712 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_229
timestamp 1604681595
transform 1 0 22172 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_237
timestamp 1604681595
transform 1 0 22908 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_233
timestamp 1604681595
transform 1 0 22540 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_237
timestamp 1604681595
transform 1 0 22908 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_233
timestamp 1604681595
transform 1 0 22540 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_5__S
timestamp 1604681595
transform 1 0 22724 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_7__S
timestamp 1604681595
transform 1 0 22724 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_7__A0
timestamp 1604681595
transform 1 0 22356 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_241
timestamp 1604681595
transform 1 0 23276 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 23184 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604681595
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23368 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_40_256
timestamp 1604681595
transform 1 0 24656 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_251
timestamp 1604681595
transform 1 0 24196 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_39_258
timestamp 1604681595
transform 1 0 24840 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_254
timestamp 1604681595
transform 1 0 24472 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 24472 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1604681595
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1604681595
transform 1 0 24932 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_270
timestamp 1604681595
transform 1 0 25944 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_266
timestamp 1604681595
transform 1 0 25576 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_261
timestamp 1604681595
transform 1 0 25116 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1604681595
transform 1 0 25760 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1604681595
transform 1 0 25208 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_263
timestamp 1604681595
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604681595
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 26128 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_274
timestamp 1604681595
transform 1 0 26312 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1604681595
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1604681595
transform 1 0 1380 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1604681595
transform 1 0 2484 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A
timestamp 1604681595
transform 1 0 1932 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__059__A
timestamp 1604681595
transform 1 0 2300 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_7
timestamp 1604681595
transform 1 0 1748 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_11
timestamp 1604681595
transform 1 0 2116 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_19
timestamp 1604681595
transform 1 0 2852 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1604681595
transform 1 0 3036 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_23
timestamp 1604681595
transform 1 0 3220 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_35
timestamp 1604681595
transform 1 0 4324 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604681595
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_47
timestamp 1604681595
transform 1 0 5428 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_59
timestamp 1604681595
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_62
timestamp 1604681595
transform 1 0 6808 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1604681595
transform 1 0 7452 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _132_
timestamp 1604681595
transform 1 0 8556 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1604681595
transform 1 0 8004 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A
timestamp 1604681595
transform 1 0 8372 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 6992 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_66
timestamp 1604681595
transform 1 0 7176 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_73
timestamp 1604681595
transform 1 0 7820 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_77
timestamp 1604681595
transform 1 0 8188 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _128_
timestamp 1604681595
transform 1 0 9660 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 10580 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 10212 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__A
timestamp 1604681595
transform 1 0 9108 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__128__A
timestamp 1604681595
transform 1 0 9476 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_85
timestamp 1604681595
transform 1 0 8924 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_89
timestamp 1604681595
transform 1 0 9292 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_97
timestamp 1604681595
transform 1 0 10028 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_101
timestamp 1604681595
transform 1 0 10396 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1604681595
transform 1 0 10764 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604681595
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1604681595
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1604681595
transform 1 0 12604 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_114
timestamp 1604681595
transform 1 0 11592 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_118
timestamp 1604681595
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_123
timestamp 1604681595
transform 1 0 12420 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13432 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1604681595
transform 1 0 12972 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 14168 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_127
timestamp 1604681595
transform 1 0 12788 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_131
timestamp 1604681595
transform 1 0 13156 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_140
timestamp 1604681595
transform 1 0 13984 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_144
timestamp 1604681595
transform 1 0 14352 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16284 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 14720 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 15732 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 16100 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 14536 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_157
timestamp 1604681595
transform 1 0 15548 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_161
timestamp 1604681595
transform 1 0 15916 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18032 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604681595
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1604681595
transform 1 0 17296 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17664 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_174
timestamp 1604681595
transform 1 0 17112 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_178
timestamp 1604681595
transform 1 0 17480 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_182
timestamp 1604681595
transform 1 0 17848 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1604681595
transform 1 0 19780 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__A
timestamp 1604681595
transform 1 0 18860 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 19228 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_190
timestamp 1604681595
transform 1 0 18584 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_195
timestamp 1604681595
transform 1 0 19044 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_199
timestamp 1604681595
transform 1 0 19412 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_207
timestamp 1604681595
transform 1 0 20148 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1604681595
transform 1 0 20884 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_6_
timestamp 1604681595
transform 1 0 21988 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1604681595
transform 1 0 21436 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A
timestamp 1604681595
transform 1 0 20332 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A
timestamp 1604681595
transform 1 0 20700 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_6__A0
timestamp 1604681595
transform 1 0 21804 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_211
timestamp 1604681595
transform 1 0 20516 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_219
timestamp 1604681595
transform 1 0 21252 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_223
timestamp 1604681595
transform 1 0 21620 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604681595
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_7__A1
timestamp 1604681595
transform 1 0 23000 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_4__A1
timestamp 1604681595
transform 1 0 23920 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_4__A0
timestamp 1604681595
transform 1 0 23368 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_236
timestamp 1604681595
transform 1 0 22816 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_240
timestamp 1604681595
transform 1 0 23184 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_245
timestamp 1604681595
transform 1 0 23644 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_250
timestamp 1604681595
transform 1 0 24104 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 24472 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 24288 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_4__S
timestamp 1604681595
transform 1 0 25484 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_263
timestamp 1604681595
transform 1 0 25300 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_267
timestamp 1604681595
transform 1 0 25668 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_275
timestamp 1604681595
transform 1 0 26404 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1604681595
transform 1 0 1380 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_7
timestamp 1604681595
transform 1 0 1748 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_19
timestamp 1604681595
transform 1 0 2852 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604681595
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1604681595
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604681595
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1604681595
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_56
timestamp 1604681595
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _135_
timestamp 1604681595
transform 1 0 8556 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 7728 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 8372 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_63
timestamp 1604681595
transform 1 0 6900 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_71
timestamp 1604681595
transform 1 0 7636 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_74
timestamp 1604681595
transform 1 0 7912 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_78
timestamp 1604681595
transform 1 0 8280 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1604681595
transform 1 0 8924 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 9108 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_89
timestamp 1604681595
transform 1 0 9292 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 9476 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604681595
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_94
timestamp 1604681595
transform 1 0 9752 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9936 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_98
timestamp 1604681595
transform 1 0 10120 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1604681595
transform 1 0 10304 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_104
timestamp 1604681595
transform 1 0 10672 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1604681595
transform 1 0 11408 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604681595
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1604681595
transform 1 0 10856 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11224 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 12144 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_108
timestamp 1604681595
transform 1 0 11040 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_116
timestamp 1604681595
transform 1 0 11776 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_122
timestamp 1604681595
transform 1 0 12328 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_125
timestamp 1604681595
transform 1 0 12604 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1604681595
transform 1 0 12972 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 14076 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13524 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13892 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 12788 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_133
timestamp 1604681595
transform 1 0 13340 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_137
timestamp 1604681595
transform 1 0 13708 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 15456 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604681595
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 14812 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 15180 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_147
timestamp 1604681595
transform 1 0 14628 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_151
timestamp 1604681595
transform 1 0 14996 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_165
timestamp 1604681595
transform 1 0 16284 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_169
timestamp 1604681595
transform 1 0 16652 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16836 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16468 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_173
timestamp 1604681595
transform 1 0 17020 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1604681595
transform 1 0 17112 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_178
timestamp 1604681595
transform 1 0 17480 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 17664 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_182
timestamp 1604681595
transform 1 0 17848 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 18032 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604681595
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_187
timestamp 1604681595
transform 1 0 18308 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1604681595
transform 1 0 19964 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _126_
timestamp 1604681595
transform 1 0 18860 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 18492 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_191
timestamp 1604681595
transform 1 0 18676 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_197
timestamp 1604681595
transform 1 0 19228 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1604681595
transform 1 0 21252 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604681595
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1604681595
transform 1 0 20884 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_6__S
timestamp 1604681595
transform 1 0 21988 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_209
timestamp 1604681595
transform 1 0 20332 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_218
timestamp 1604681595
transform 1 0 21160 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_223
timestamp 1604681595
transform 1 0 21620 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_229
timestamp 1604681595
transform 1 0 22172 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_4_
timestamp 1604681595
transform 1 0 24012 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_7_
timestamp 1604681595
transform 1 0 22356 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604681595
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_240
timestamp 1604681595
transform 1 0 23184 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 25024 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_258
timestamp 1604681595
transform 1 0 24840 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_262
timestamp 1604681595
transform 1 0 25208 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_274
timestamp 1604681595
transform 1 0 26312 0 -1 25568
box -38 -48 314 592
<< labels >>
rlabel metal2 s 202 0 258 480 6 bottom_left_grid_pin_42_
port 0 nsew default input
rlabel metal2 s 662 0 718 480 6 bottom_left_grid_pin_43_
port 1 nsew default input
rlabel metal2 s 1214 0 1270 480 6 bottom_left_grid_pin_44_
port 2 nsew default input
rlabel metal2 s 1766 0 1822 480 6 bottom_left_grid_pin_45_
port 3 nsew default input
rlabel metal2 s 2318 0 2374 480 6 bottom_left_grid_pin_46_
port 4 nsew default input
rlabel metal2 s 2870 0 2926 480 6 bottom_left_grid_pin_47_
port 5 nsew default input
rlabel metal2 s 3422 0 3478 480 6 bottom_left_grid_pin_48_
port 6 nsew default input
rlabel metal2 s 3974 0 4030 480 6 bottom_left_grid_pin_49_
port 7 nsew default input
rlabel metal2 s 5078 0 5134 480 6 ccff_head
port 8 nsew default input
rlabel metal2 s 5630 0 5686 480 6 ccff_tail
port 9 nsew default tristate
rlabel metal3 s 0 4904 480 5024 6 chanx_left_in[0]
port 10 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[10]
port 11 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[11]
port 12 nsew default input
rlabel metal3 s 0 11840 480 11960 6 chanx_left_in[12]
port 13 nsew default input
rlabel metal3 s 0 12520 480 12640 6 chanx_left_in[13]
port 14 nsew default input
rlabel metal3 s 0 13064 480 13184 6 chanx_left_in[14]
port 15 nsew default input
rlabel metal3 s 0 13608 480 13728 6 chanx_left_in[15]
port 16 nsew default input
rlabel metal3 s 0 14288 480 14408 6 chanx_left_in[16]
port 17 nsew default input
rlabel metal3 s 0 14832 480 14952 6 chanx_left_in[17]
port 18 nsew default input
rlabel metal3 s 0 15376 480 15496 6 chanx_left_in[18]
port 19 nsew default input
rlabel metal3 s 0 15920 480 16040 6 chanx_left_in[19]
port 20 nsew default input
rlabel metal3 s 0 5448 480 5568 6 chanx_left_in[1]
port 21 nsew default input
rlabel metal3 s 0 5992 480 6112 6 chanx_left_in[2]
port 22 nsew default input
rlabel metal3 s 0 6672 480 6792 6 chanx_left_in[3]
port 23 nsew default input
rlabel metal3 s 0 7216 480 7336 6 chanx_left_in[4]
port 24 nsew default input
rlabel metal3 s 0 7760 480 7880 6 chanx_left_in[5]
port 25 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_in[6]
port 26 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[7]
port 27 nsew default input
rlabel metal3 s 0 9528 480 9648 6 chanx_left_in[8]
port 28 nsew default input
rlabel metal3 s 0 10072 480 10192 6 chanx_left_in[9]
port 29 nsew default input
rlabel metal3 s 0 16600 480 16720 6 chanx_left_out[0]
port 30 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 chanx_left_out[10]
port 31 nsew default tristate
rlabel metal3 s 0 22992 480 23112 6 chanx_left_out[11]
port 32 nsew default tristate
rlabel metal3 s 0 23536 480 23656 6 chanx_left_out[12]
port 33 nsew default tristate
rlabel metal3 s 0 24080 480 24200 6 chanx_left_out[13]
port 34 nsew default tristate
rlabel metal3 s 0 24760 480 24880 6 chanx_left_out[14]
port 35 nsew default tristate
rlabel metal3 s 0 25304 480 25424 6 chanx_left_out[15]
port 36 nsew default tristate
rlabel metal3 s 0 25848 480 25968 6 chanx_left_out[16]
port 37 nsew default tristate
rlabel metal3 s 0 26528 480 26648 6 chanx_left_out[17]
port 38 nsew default tristate
rlabel metal3 s 0 27072 480 27192 6 chanx_left_out[18]
port 39 nsew default tristate
rlabel metal3 s 0 27616 480 27736 6 chanx_left_out[19]
port 40 nsew default tristate
rlabel metal3 s 0 17144 480 17264 6 chanx_left_out[1]
port 41 nsew default tristate
rlabel metal3 s 0 17688 480 17808 6 chanx_left_out[2]
port 42 nsew default tristate
rlabel metal3 s 0 18368 480 18488 6 chanx_left_out[3]
port 43 nsew default tristate
rlabel metal3 s 0 18912 480 19032 6 chanx_left_out[4]
port 44 nsew default tristate
rlabel metal3 s 0 19456 480 19576 6 chanx_left_out[5]
port 45 nsew default tristate
rlabel metal3 s 0 20000 480 20120 6 chanx_left_out[6]
port 46 nsew default tristate
rlabel metal3 s 0 20680 480 20800 6 chanx_left_out[7]
port 47 nsew default tristate
rlabel metal3 s 0 21224 480 21344 6 chanx_left_out[8]
port 48 nsew default tristate
rlabel metal3 s 0 21768 480 21888 6 chanx_left_out[9]
port 49 nsew default tristate
rlabel metal3 s 27520 4904 28000 5024 6 chanx_right_in[0]
port 50 nsew default input
rlabel metal3 s 27520 10752 28000 10872 6 chanx_right_in[10]
port 51 nsew default input
rlabel metal3 s 27520 11296 28000 11416 6 chanx_right_in[11]
port 52 nsew default input
rlabel metal3 s 27520 11840 28000 11960 6 chanx_right_in[12]
port 53 nsew default input
rlabel metal3 s 27520 12520 28000 12640 6 chanx_right_in[13]
port 54 nsew default input
rlabel metal3 s 27520 13064 28000 13184 6 chanx_right_in[14]
port 55 nsew default input
rlabel metal3 s 27520 13608 28000 13728 6 chanx_right_in[15]
port 56 nsew default input
rlabel metal3 s 27520 14288 28000 14408 6 chanx_right_in[16]
port 57 nsew default input
rlabel metal3 s 27520 14832 28000 14952 6 chanx_right_in[17]
port 58 nsew default input
rlabel metal3 s 27520 15376 28000 15496 6 chanx_right_in[18]
port 59 nsew default input
rlabel metal3 s 27520 15920 28000 16040 6 chanx_right_in[19]
port 60 nsew default input
rlabel metal3 s 27520 5448 28000 5568 6 chanx_right_in[1]
port 61 nsew default input
rlabel metal3 s 27520 5992 28000 6112 6 chanx_right_in[2]
port 62 nsew default input
rlabel metal3 s 27520 6672 28000 6792 6 chanx_right_in[3]
port 63 nsew default input
rlabel metal3 s 27520 7216 28000 7336 6 chanx_right_in[4]
port 64 nsew default input
rlabel metal3 s 27520 7760 28000 7880 6 chanx_right_in[5]
port 65 nsew default input
rlabel metal3 s 27520 8440 28000 8560 6 chanx_right_in[6]
port 66 nsew default input
rlabel metal3 s 27520 8984 28000 9104 6 chanx_right_in[7]
port 67 nsew default input
rlabel metal3 s 27520 9528 28000 9648 6 chanx_right_in[8]
port 68 nsew default input
rlabel metal3 s 27520 10072 28000 10192 6 chanx_right_in[9]
port 69 nsew default input
rlabel metal3 s 27520 16600 28000 16720 6 chanx_right_out[0]
port 70 nsew default tristate
rlabel metal3 s 27520 22448 28000 22568 6 chanx_right_out[10]
port 71 nsew default tristate
rlabel metal3 s 27520 22992 28000 23112 6 chanx_right_out[11]
port 72 nsew default tristate
rlabel metal3 s 27520 23536 28000 23656 6 chanx_right_out[12]
port 73 nsew default tristate
rlabel metal3 s 27520 24080 28000 24200 6 chanx_right_out[13]
port 74 nsew default tristate
rlabel metal3 s 27520 24760 28000 24880 6 chanx_right_out[14]
port 75 nsew default tristate
rlabel metal3 s 27520 25304 28000 25424 6 chanx_right_out[15]
port 76 nsew default tristate
rlabel metal3 s 27520 25848 28000 25968 6 chanx_right_out[16]
port 77 nsew default tristate
rlabel metal3 s 27520 26528 28000 26648 6 chanx_right_out[17]
port 78 nsew default tristate
rlabel metal3 s 27520 27072 28000 27192 6 chanx_right_out[18]
port 79 nsew default tristate
rlabel metal3 s 27520 27616 28000 27736 6 chanx_right_out[19]
port 80 nsew default tristate
rlabel metal3 s 27520 17144 28000 17264 6 chanx_right_out[1]
port 81 nsew default tristate
rlabel metal3 s 27520 17688 28000 17808 6 chanx_right_out[2]
port 82 nsew default tristate
rlabel metal3 s 27520 18368 28000 18488 6 chanx_right_out[3]
port 83 nsew default tristate
rlabel metal3 s 27520 18912 28000 19032 6 chanx_right_out[4]
port 84 nsew default tristate
rlabel metal3 s 27520 19456 28000 19576 6 chanx_right_out[5]
port 85 nsew default tristate
rlabel metal3 s 27520 20000 28000 20120 6 chanx_right_out[6]
port 86 nsew default tristate
rlabel metal3 s 27520 20680 28000 20800 6 chanx_right_out[7]
port 87 nsew default tristate
rlabel metal3 s 27520 21224 28000 21344 6 chanx_right_out[8]
port 88 nsew default tristate
rlabel metal3 s 27520 21768 28000 21888 6 chanx_right_out[9]
port 89 nsew default tristate
rlabel metal2 s 6182 0 6238 480 6 chany_bottom_in[0]
port 90 nsew default input
rlabel metal2 s 11702 0 11758 480 6 chany_bottom_in[10]
port 91 nsew default input
rlabel metal2 s 12254 0 12310 480 6 chany_bottom_in[11]
port 92 nsew default input
rlabel metal2 s 12806 0 12862 480 6 chany_bottom_in[12]
port 93 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[13]
port 94 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chany_bottom_in[14]
port 95 nsew default input
rlabel metal2 s 14370 0 14426 480 6 chany_bottom_in[15]
port 96 nsew default input
rlabel metal2 s 14922 0 14978 480 6 chany_bottom_in[16]
port 97 nsew default input
rlabel metal2 s 15474 0 15530 480 6 chany_bottom_in[17]
port 98 nsew default input
rlabel metal2 s 16026 0 16082 480 6 chany_bottom_in[18]
port 99 nsew default input
rlabel metal2 s 16578 0 16634 480 6 chany_bottom_in[19]
port 100 nsew default input
rlabel metal2 s 6734 0 6790 480 6 chany_bottom_in[1]
port 101 nsew default input
rlabel metal2 s 7286 0 7342 480 6 chany_bottom_in[2]
port 102 nsew default input
rlabel metal2 s 7838 0 7894 480 6 chany_bottom_in[3]
port 103 nsew default input
rlabel metal2 s 8390 0 8446 480 6 chany_bottom_in[4]
port 104 nsew default input
rlabel metal2 s 8942 0 8998 480 6 chany_bottom_in[5]
port 105 nsew default input
rlabel metal2 s 9494 0 9550 480 6 chany_bottom_in[6]
port 106 nsew default input
rlabel metal2 s 10046 0 10102 480 6 chany_bottom_in[7]
port 107 nsew default input
rlabel metal2 s 10598 0 10654 480 6 chany_bottom_in[8]
port 108 nsew default input
rlabel metal2 s 11150 0 11206 480 6 chany_bottom_in[9]
port 109 nsew default input
rlabel metal2 s 17130 0 17186 480 6 chany_bottom_out[0]
port 110 nsew default tristate
rlabel metal2 s 22650 0 22706 480 6 chany_bottom_out[10]
port 111 nsew default tristate
rlabel metal2 s 23202 0 23258 480 6 chany_bottom_out[11]
port 112 nsew default tristate
rlabel metal2 s 23754 0 23810 480 6 chany_bottom_out[12]
port 113 nsew default tristate
rlabel metal2 s 24306 0 24362 480 6 chany_bottom_out[13]
port 114 nsew default tristate
rlabel metal2 s 24858 0 24914 480 6 chany_bottom_out[14]
port 115 nsew default tristate
rlabel metal2 s 25410 0 25466 480 6 chany_bottom_out[15]
port 116 nsew default tristate
rlabel metal2 s 25962 0 26018 480 6 chany_bottom_out[16]
port 117 nsew default tristate
rlabel metal2 s 26514 0 26570 480 6 chany_bottom_out[17]
port 118 nsew default tristate
rlabel metal2 s 27066 0 27122 480 6 chany_bottom_out[18]
port 119 nsew default tristate
rlabel metal2 s 27618 0 27674 480 6 chany_bottom_out[19]
port 120 nsew default tristate
rlabel metal2 s 17682 0 17738 480 6 chany_bottom_out[1]
port 121 nsew default tristate
rlabel metal2 s 18234 0 18290 480 6 chany_bottom_out[2]
port 122 nsew default tristate
rlabel metal2 s 18786 0 18842 480 6 chany_bottom_out[3]
port 123 nsew default tristate
rlabel metal2 s 19338 0 19394 480 6 chany_bottom_out[4]
port 124 nsew default tristate
rlabel metal2 s 19890 0 19946 480 6 chany_bottom_out[5]
port 125 nsew default tristate
rlabel metal2 s 20442 0 20498 480 6 chany_bottom_out[6]
port 126 nsew default tristate
rlabel metal2 s 20994 0 21050 480 6 chany_bottom_out[7]
port 127 nsew default tristate
rlabel metal2 s 21546 0 21602 480 6 chany_bottom_out[8]
port 128 nsew default tristate
rlabel metal2 s 22098 0 22154 480 6 chany_bottom_out[9]
port 129 nsew default tristate
rlabel metal2 s 4894 27520 4950 28000 6 chany_top_in[0]
port 130 nsew default input
rlabel metal2 s 10782 27520 10838 28000 6 chany_top_in[10]
port 131 nsew default input
rlabel metal2 s 11334 27520 11390 28000 6 chany_top_in[11]
port 132 nsew default input
rlabel metal2 s 11886 27520 11942 28000 6 chany_top_in[12]
port 133 nsew default input
rlabel metal2 s 12530 27520 12586 28000 6 chany_top_in[13]
port 134 nsew default input
rlabel metal2 s 13082 27520 13138 28000 6 chany_top_in[14]
port 135 nsew default input
rlabel metal2 s 13634 27520 13690 28000 6 chany_top_in[15]
port 136 nsew default input
rlabel metal2 s 14278 27520 14334 28000 6 chany_top_in[16]
port 137 nsew default input
rlabel metal2 s 14830 27520 14886 28000 6 chany_top_in[17]
port 138 nsew default input
rlabel metal2 s 15382 27520 15438 28000 6 chany_top_in[18]
port 139 nsew default input
rlabel metal2 s 16026 27520 16082 28000 6 chany_top_in[19]
port 140 nsew default input
rlabel metal2 s 5538 27520 5594 28000 6 chany_top_in[1]
port 141 nsew default input
rlabel metal2 s 6090 27520 6146 28000 6 chany_top_in[2]
port 142 nsew default input
rlabel metal2 s 6642 27520 6698 28000 6 chany_top_in[3]
port 143 nsew default input
rlabel metal2 s 7286 27520 7342 28000 6 chany_top_in[4]
port 144 nsew default input
rlabel metal2 s 7838 27520 7894 28000 6 chany_top_in[5]
port 145 nsew default input
rlabel metal2 s 8390 27520 8446 28000 6 chany_top_in[6]
port 146 nsew default input
rlabel metal2 s 9034 27520 9090 28000 6 chany_top_in[7]
port 147 nsew default input
rlabel metal2 s 9586 27520 9642 28000 6 chany_top_in[8]
port 148 nsew default input
rlabel metal2 s 10138 27520 10194 28000 6 chany_top_in[9]
port 149 nsew default input
rlabel metal2 s 16578 27520 16634 28000 6 chany_top_out[0]
port 150 nsew default tristate
rlabel metal2 s 22374 27520 22430 28000 6 chany_top_out[10]
port 151 nsew default tristate
rlabel metal2 s 23018 27520 23074 28000 6 chany_top_out[11]
port 152 nsew default tristate
rlabel metal2 s 23570 27520 23626 28000 6 chany_top_out[12]
port 153 nsew default tristate
rlabel metal2 s 24122 27520 24178 28000 6 chany_top_out[13]
port 154 nsew default tristate
rlabel metal2 s 24766 27520 24822 28000 6 chany_top_out[14]
port 155 nsew default tristate
rlabel metal2 s 25318 27520 25374 28000 6 chany_top_out[15]
port 156 nsew default tristate
rlabel metal2 s 25870 27520 25926 28000 6 chany_top_out[16]
port 157 nsew default tristate
rlabel metal2 s 26514 27520 26570 28000 6 chany_top_out[17]
port 158 nsew default tristate
rlabel metal2 s 27066 27520 27122 28000 6 chany_top_out[18]
port 159 nsew default tristate
rlabel metal2 s 27618 27520 27674 28000 6 chany_top_out[19]
port 160 nsew default tristate
rlabel metal2 s 17130 27520 17186 28000 6 chany_top_out[1]
port 161 nsew default tristate
rlabel metal2 s 17774 27520 17830 28000 6 chany_top_out[2]
port 162 nsew default tristate
rlabel metal2 s 18326 27520 18382 28000 6 chany_top_out[3]
port 163 nsew default tristate
rlabel metal2 s 18878 27520 18934 28000 6 chany_top_out[4]
port 164 nsew default tristate
rlabel metal2 s 19522 27520 19578 28000 6 chany_top_out[5]
port 165 nsew default tristate
rlabel metal2 s 20074 27520 20130 28000 6 chany_top_out[6]
port 166 nsew default tristate
rlabel metal2 s 20626 27520 20682 28000 6 chany_top_out[7]
port 167 nsew default tristate
rlabel metal2 s 21270 27520 21326 28000 6 chany_top_out[8]
port 168 nsew default tristate
rlabel metal2 s 21822 27520 21878 28000 6 chany_top_out[9]
port 169 nsew default tristate
rlabel metal3 s 0 280 480 400 6 left_bottom_grid_pin_34_
port 170 nsew default input
rlabel metal3 s 0 824 480 944 6 left_bottom_grid_pin_35_
port 171 nsew default input
rlabel metal3 s 0 1368 480 1488 6 left_bottom_grid_pin_36_
port 172 nsew default input
rlabel metal3 s 0 1912 480 2032 6 left_bottom_grid_pin_37_
port 173 nsew default input
rlabel metal3 s 0 2592 480 2712 6 left_bottom_grid_pin_38_
port 174 nsew default input
rlabel metal3 s 0 3136 480 3256 6 left_bottom_grid_pin_39_
port 175 nsew default input
rlabel metal3 s 0 3680 480 3800 6 left_bottom_grid_pin_40_
port 176 nsew default input
rlabel metal3 s 0 4360 480 4480 6 left_bottom_grid_pin_41_
port 177 nsew default input
rlabel metal2 s 4526 0 4582 480 6 prog_clk
port 178 nsew default input
rlabel metal3 s 27520 280 28000 400 6 right_bottom_grid_pin_34_
port 179 nsew default input
rlabel metal3 s 27520 824 28000 944 6 right_bottom_grid_pin_35_
port 180 nsew default input
rlabel metal3 s 27520 1368 28000 1488 6 right_bottom_grid_pin_36_
port 181 nsew default input
rlabel metal3 s 27520 1912 28000 2032 6 right_bottom_grid_pin_37_
port 182 nsew default input
rlabel metal3 s 27520 2592 28000 2712 6 right_bottom_grid_pin_38_
port 183 nsew default input
rlabel metal3 s 27520 3136 28000 3256 6 right_bottom_grid_pin_39_
port 184 nsew default input
rlabel metal3 s 27520 3680 28000 3800 6 right_bottom_grid_pin_40_
port 185 nsew default input
rlabel metal3 s 27520 4360 28000 4480 6 right_bottom_grid_pin_41_
port 186 nsew default input
rlabel metal2 s 294 27520 350 28000 6 top_left_grid_pin_42_
port 187 nsew default input
rlabel metal2 s 846 27520 902 28000 6 top_left_grid_pin_43_
port 188 nsew default input
rlabel metal2 s 1398 27520 1454 28000 6 top_left_grid_pin_44_
port 189 nsew default input
rlabel metal2 s 2042 27520 2098 28000 6 top_left_grid_pin_45_
port 190 nsew default input
rlabel metal2 s 2594 27520 2650 28000 6 top_left_grid_pin_46_
port 191 nsew default input
rlabel metal2 s 3146 27520 3202 28000 6 top_left_grid_pin_47_
port 192 nsew default input
rlabel metal2 s 3790 27520 3846 28000 6 top_left_grid_pin_48_
port 193 nsew default input
rlabel metal2 s 4342 27520 4398 28000 6 top_left_grid_pin_49_
port 194 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 VPWR
port 195 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 VGND
port 196 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
